VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO sky130_osu_ring_oscillator_mpr2aa_8_b0r1
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 0.005 0.01 ;
  SIZE 81.785 BY 8.955 ;
  SYMMETRY X Y R90 ;
  SITE CoreSite ;
  OBS
    LAYER met3 ;
      RECT 73.57 7.04 73.94 7.41 ;
      RECT 73.61 6.72 73.945 7.085 ;
      RECT 73.61 6.72 73.995 7.03 ;
      RECT 73.61 6.72 76.4 7.025 ;
      RECT 76.095 2.85 76.4 7.025 ;
      RECT 76.06 2.85 76.43 3.22 ;
      RECT 75.32 0.815 75.625 4.02 ;
      RECT 75.07 2.975 75.625 3.705 ;
      RECT 75.28 0.815 75.65 1.185 ;
      RECT 71.43 1.85 71.76 2.745 ;
      RECT 70.55 2.015 70.88 2.745 ;
      RECT 71.425 1.85 71.795 2.65 ;
      RECT 74.59 1.85 74.92 2.58 ;
      RECT 74.55 1.735 74.73 2.385 ;
      RECT 70.56 1.85 74.92 2.22 ;
      RECT 71.05 3.535 71.38 3.865 ;
      RECT 69.845 3.55 71.38 3.85 ;
      RECT 69.845 2.43 70.145 3.85 ;
      RECT 69.59 2.415 69.92 2.745 ;
      RECT 57.785 7.04 58.155 7.41 ;
      RECT 57.825 6.72 58.16 7.085 ;
      RECT 57.825 6.72 58.21 7.03 ;
      RECT 57.825 6.72 60.615 7.025 ;
      RECT 60.31 2.85 60.615 7.025 ;
      RECT 60.275 2.85 60.645 3.22 ;
      RECT 59.535 0.815 59.84 4.02 ;
      RECT 59.285 2.975 59.84 3.705 ;
      RECT 59.495 0.815 59.865 1.185 ;
      RECT 55.645 1.85 55.975 2.745 ;
      RECT 54.765 2.015 55.095 2.745 ;
      RECT 55.64 1.85 56.01 2.65 ;
      RECT 58.805 1.85 59.135 2.58 ;
      RECT 58.765 1.735 58.945 2.385 ;
      RECT 54.775 1.85 59.135 2.22 ;
      RECT 55.265 3.535 55.595 3.865 ;
      RECT 54.06 3.55 55.595 3.85 ;
      RECT 54.06 2.43 54.36 3.85 ;
      RECT 53.805 2.415 54.135 2.745 ;
      RECT 42 7.04 42.37 7.41 ;
      RECT 42.04 6.72 42.375 7.085 ;
      RECT 42.04 6.72 42.425 7.03 ;
      RECT 42.04 6.72 44.83 7.025 ;
      RECT 44.525 2.85 44.83 7.025 ;
      RECT 44.49 2.85 44.86 3.22 ;
      RECT 43.75 0.815 44.055 4.02 ;
      RECT 43.5 2.975 44.055 3.705 ;
      RECT 43.71 0.815 44.08 1.185 ;
      RECT 39.86 1.85 40.19 2.745 ;
      RECT 38.98 2.015 39.31 2.745 ;
      RECT 39.855 1.85 40.225 2.65 ;
      RECT 43.02 1.85 43.35 2.58 ;
      RECT 42.98 1.735 43.16 2.385 ;
      RECT 38.99 1.85 43.35 2.22 ;
      RECT 39.48 3.535 39.81 3.865 ;
      RECT 38.275 3.55 39.81 3.85 ;
      RECT 38.275 2.43 38.575 3.85 ;
      RECT 38.02 2.415 38.35 2.745 ;
      RECT 26.225 7.04 26.595 7.41 ;
      RECT 26.265 6.72 26.6 7.085 ;
      RECT 26.265 6.72 26.65 7.03 ;
      RECT 26.265 6.72 29.055 7.025 ;
      RECT 28.75 2.85 29.055 7.025 ;
      RECT 28.715 2.85 29.085 3.22 ;
      RECT 27.975 0.815 28.28 4.02 ;
      RECT 27.725 2.975 28.28 3.705 ;
      RECT 27.935 0.815 28.305 1.185 ;
      RECT 24.085 1.85 24.415 2.745 ;
      RECT 23.205 2.015 23.535 2.745 ;
      RECT 24.08 1.85 24.45 2.65 ;
      RECT 27.245 1.85 27.575 2.58 ;
      RECT 27.205 1.735 27.385 2.385 ;
      RECT 23.215 1.85 27.575 2.22 ;
      RECT 23.705 3.535 24.035 3.865 ;
      RECT 22.5 3.55 24.035 3.85 ;
      RECT 22.5 2.43 22.8 3.85 ;
      RECT 22.245 2.415 22.575 2.745 ;
      RECT 10.445 7.04 10.815 7.41 ;
      RECT 10.485 6.72 10.82 7.085 ;
      RECT 10.485 6.72 10.87 7.03 ;
      RECT 10.485 6.72 13.275 7.025 ;
      RECT 12.97 2.85 13.275 7.025 ;
      RECT 12.935 2.85 13.305 3.22 ;
      RECT 12.195 0.815 12.5 4.02 ;
      RECT 11.945 2.975 12.5 3.705 ;
      RECT 12.155 0.815 12.525 1.185 ;
      RECT 8.305 1.85 8.635 2.745 ;
      RECT 7.425 2.015 7.755 2.745 ;
      RECT 8.3 1.85 8.67 2.65 ;
      RECT 11.465 1.85 11.795 2.58 ;
      RECT 11.425 1.735 11.605 2.385 ;
      RECT 7.435 1.85 11.795 2.22 ;
      RECT 7.925 3.535 8.255 3.865 ;
      RECT 6.72 3.55 8.255 3.85 ;
      RECT 6.72 2.43 7.02 3.85 ;
      RECT 6.465 2.415 6.795 2.745 ;
      RECT 0.055 8.565 0.865 8.945 ;
      RECT -0.005 8.575 0.865 8.88 ;
      RECT 72.99 2.575 73.32 3.305 ;
      RECT 68.87 2.415 69.2 3.145 ;
      RECT 67.87 1.855 68.2 2.585 ;
      RECT 66.43 2.575 66.76 3.305 ;
      RECT 57.205 2.575 57.535 3.305 ;
      RECT 53.085 2.415 53.415 3.145 ;
      RECT 52.085 1.855 52.415 2.585 ;
      RECT 50.645 2.575 50.975 3.305 ;
      RECT 41.42 2.575 41.75 3.305 ;
      RECT 37.3 2.415 37.63 3.145 ;
      RECT 36.3 1.855 36.63 2.585 ;
      RECT 34.86 2.575 35.19 3.305 ;
      RECT 25.645 2.575 25.975 3.305 ;
      RECT 21.525 2.415 21.855 3.145 ;
      RECT 20.525 1.855 20.855 2.585 ;
      RECT 19.085 2.575 19.415 3.305 ;
      RECT 9.865 2.575 10.195 3.305 ;
      RECT 5.745 2.415 6.075 3.145 ;
      RECT 4.745 1.855 5.075 2.585 ;
      RECT 3.305 2.575 3.635 3.305 ;
      RECT 0.64 4.26 1.45 4.64 ;
      RECT 0.585 -0.01 1.395 0.37 ;
    LAYER via2 ;
      RECT 76.145 2.935 76.345 3.135 ;
      RECT 75.365 0.9 75.565 1.1 ;
      RECT 75.135 3.04 75.335 3.24 ;
      RECT 74.655 2.315 74.855 2.515 ;
      RECT 73.655 7.125 73.855 7.325 ;
      RECT 73.055 3.04 73.255 3.24 ;
      RECT 71.495 2.48 71.695 2.68 ;
      RECT 71.115 3.6 71.315 3.8 ;
      RECT 70.615 2.48 70.815 2.68 ;
      RECT 69.655 2.48 69.855 2.68 ;
      RECT 68.935 2.48 69.135 2.68 ;
      RECT 67.935 1.92 68.135 2.12 ;
      RECT 66.495 3.04 66.695 3.24 ;
      RECT 60.36 2.935 60.56 3.135 ;
      RECT 59.58 0.9 59.78 1.1 ;
      RECT 59.35 3.04 59.55 3.24 ;
      RECT 58.87 2.315 59.07 2.515 ;
      RECT 57.87 7.125 58.07 7.325 ;
      RECT 57.27 3.04 57.47 3.24 ;
      RECT 55.71 2.48 55.91 2.68 ;
      RECT 55.33 3.6 55.53 3.8 ;
      RECT 54.83 2.48 55.03 2.68 ;
      RECT 53.87 2.48 54.07 2.68 ;
      RECT 53.15 2.48 53.35 2.68 ;
      RECT 52.15 1.92 52.35 2.12 ;
      RECT 50.71 3.04 50.91 3.24 ;
      RECT 44.575 2.935 44.775 3.135 ;
      RECT 43.795 0.9 43.995 1.1 ;
      RECT 43.565 3.04 43.765 3.24 ;
      RECT 43.085 2.315 43.285 2.515 ;
      RECT 42.085 7.125 42.285 7.325 ;
      RECT 41.485 3.04 41.685 3.24 ;
      RECT 39.925 2.48 40.125 2.68 ;
      RECT 39.545 3.6 39.745 3.8 ;
      RECT 39.045 2.48 39.245 2.68 ;
      RECT 38.085 2.48 38.285 2.68 ;
      RECT 37.365 2.48 37.565 2.68 ;
      RECT 36.365 1.92 36.565 2.12 ;
      RECT 34.925 3.04 35.125 3.24 ;
      RECT 28.8 2.935 29 3.135 ;
      RECT 28.02 0.9 28.22 1.1 ;
      RECT 27.79 3.04 27.99 3.24 ;
      RECT 27.31 2.315 27.51 2.515 ;
      RECT 26.31 7.125 26.51 7.325 ;
      RECT 25.71 3.04 25.91 3.24 ;
      RECT 24.15 2.48 24.35 2.68 ;
      RECT 23.77 3.6 23.97 3.8 ;
      RECT 23.27 2.48 23.47 2.68 ;
      RECT 22.31 2.48 22.51 2.68 ;
      RECT 21.59 2.48 21.79 2.68 ;
      RECT 20.59 1.92 20.79 2.12 ;
      RECT 19.15 3.04 19.35 3.24 ;
      RECT 13.02 2.935 13.22 3.135 ;
      RECT 12.24 0.9 12.44 1.1 ;
      RECT 12.01 3.04 12.21 3.24 ;
      RECT 11.53 2.315 11.73 2.515 ;
      RECT 10.53 7.125 10.73 7.325 ;
      RECT 9.93 3.04 10.13 3.24 ;
      RECT 8.37 2.48 8.57 2.68 ;
      RECT 7.99 3.6 8.19 3.8 ;
      RECT 7.49 2.48 7.69 2.68 ;
      RECT 6.53 2.48 6.73 2.68 ;
      RECT 5.81 2.48 6.01 2.68 ;
      RECT 4.81 1.92 5.01 2.12 ;
      RECT 3.37 3.04 3.57 3.24 ;
      RECT 0.925 4.35 1.125 4.55 ;
      RECT 0.87 0.08 1.07 0.28 ;
      RECT 0.34 8.655 0.54 8.855 ;
    LAYER met2 ;
      RECT 1.24 8.4 81.405 8.57 ;
      RECT 81.235 7.275 81.405 8.57 ;
      RECT 1.24 6.255 1.41 8.57 ;
      RECT 81.205 7.275 81.555 7.625 ;
      RECT 1.175 6.255 1.465 6.605 ;
      RECT 78.045 6.22 78.365 6.545 ;
      RECT 78.075 5.695 78.245 6.545 ;
      RECT 78.075 5.695 78.25 6.045 ;
      RECT 78.075 5.695 79.05 5.87 ;
      RECT 78.875 1.965 79.05 5.87 ;
      RECT 78.82 1.965 79.17 2.315 ;
      RECT 78.845 6.655 79.17 6.98 ;
      RECT 77.73 6.745 79.17 6.915 ;
      RECT 77.73 2.395 77.89 6.915 ;
      RECT 78.045 2.365 78.365 2.685 ;
      RECT 77.73 2.395 78.365 2.565 ;
      RECT 76.995 5.855 77.345 6.205 ;
      RECT 77.065 2.705 77.24 6.205 ;
      RECT 76.99 2.705 77.34 3.055 ;
      RECT 67.815 1.92 68.075 2.18 ;
      RECT 67.87 1.88 68.175 2.16 ;
      RECT 67.87 1.42 68.045 2.18 ;
      RECT 76.385 1.34 76.735 1.69 ;
      RECT 67.87 1.42 76.735 1.595 ;
      RECT 76.06 2.85 76.43 3.22 ;
      RECT 76.145 2.235 76.315 3.22 ;
      RECT 72.165 2.455 72.4 2.715 ;
      RECT 75.31 2.235 75.475 2.495 ;
      RECT 75.215 2.225 75.23 2.495 ;
      RECT 75.31 2.235 76.315 2.415 ;
      RECT 73.815 1.795 73.855 1.935 ;
      RECT 75.23 2.23 75.31 2.495 ;
      RECT 75.175 2.225 75.215 2.461 ;
      RECT 75.161 2.225 75.175 2.461 ;
      RECT 75.075 2.23 75.161 2.463 ;
      RECT 75.03 2.237 75.075 2.465 ;
      RECT 75 2.237 75.03 2.467 ;
      RECT 74.975 2.232 75 2.469 ;
      RECT 74.945 2.228 74.975 2.478 ;
      RECT 74.935 2.225 74.945 2.49 ;
      RECT 74.93 2.225 74.935 2.498 ;
      RECT 74.925 2.225 74.93 2.503 ;
      RECT 74.915 2.224 74.925 2.513 ;
      RECT 74.91 2.223 74.915 2.523 ;
      RECT 74.895 2.222 74.91 2.528 ;
      RECT 74.867 2.219 74.895 2.555 ;
      RECT 74.781 2.211 74.867 2.555 ;
      RECT 74.695 2.2 74.781 2.555 ;
      RECT 74.655 2.185 74.695 2.555 ;
      RECT 74.615 2.159 74.655 2.555 ;
      RECT 74.61 2.141 74.615 2.367 ;
      RECT 74.6 2.137 74.61 2.357 ;
      RECT 74.585 2.127 74.6 2.344 ;
      RECT 74.565 2.111 74.585 2.329 ;
      RECT 74.55 2.096 74.565 2.314 ;
      RECT 74.54 2.085 74.55 2.304 ;
      RECT 74.515 2.069 74.54 2.293 ;
      RECT 74.51 2.056 74.515 2.283 ;
      RECT 74.505 2.052 74.51 2.278 ;
      RECT 74.45 2.038 74.505 2.256 ;
      RECT 74.411 2.019 74.45 2.22 ;
      RECT 74.325 1.993 74.411 2.173 ;
      RECT 74.321 1.975 74.325 2.139 ;
      RECT 74.235 1.956 74.321 2.117 ;
      RECT 74.23 1.938 74.235 2.095 ;
      RECT 74.225 1.936 74.23 2.093 ;
      RECT 74.215 1.935 74.225 2.088 ;
      RECT 74.155 1.922 74.215 2.074 ;
      RECT 74.11 1.9 74.155 2.053 ;
      RECT 74.05 1.877 74.11 2.032 ;
      RECT 73.986 1.852 74.05 2.007 ;
      RECT 73.9 1.822 73.986 1.976 ;
      RECT 73.885 1.802 73.9 1.955 ;
      RECT 73.855 1.797 73.885 1.946 ;
      RECT 73.802 1.795 73.815 1.935 ;
      RECT 73.716 1.795 73.802 1.937 ;
      RECT 73.63 1.795 73.716 1.939 ;
      RECT 73.61 1.795 73.63 1.943 ;
      RECT 73.565 1.797 73.61 1.954 ;
      RECT 73.525 1.807 73.565 1.97 ;
      RECT 73.521 1.816 73.525 1.978 ;
      RECT 73.435 1.836 73.521 1.994 ;
      RECT 73.425 1.855 73.435 2.012 ;
      RECT 73.42 1.857 73.425 2.015 ;
      RECT 73.41 1.861 73.42 2.018 ;
      RECT 73.39 1.866 73.41 2.028 ;
      RECT 73.36 1.876 73.39 2.048 ;
      RECT 73.355 1.883 73.36 2.062 ;
      RECT 73.345 1.887 73.355 2.069 ;
      RECT 73.33 1.895 73.345 2.08 ;
      RECT 73.32 1.905 73.33 2.091 ;
      RECT 73.31 1.912 73.32 2.099 ;
      RECT 73.285 1.925 73.31 2.114 ;
      RECT 73.221 1.961 73.285 2.153 ;
      RECT 73.135 2.024 73.221 2.217 ;
      RECT 73.1 2.075 73.135 2.27 ;
      RECT 73.095 2.092 73.1 2.287 ;
      RECT 73.08 2.101 73.095 2.294 ;
      RECT 73.06 2.116 73.08 2.308 ;
      RECT 73.055 2.127 73.06 2.318 ;
      RECT 73.035 2.14 73.055 2.328 ;
      RECT 73.03 2.15 73.035 2.338 ;
      RECT 73.015 2.155 73.03 2.347 ;
      RECT 73.005 2.165 73.015 2.358 ;
      RECT 72.975 2.182 73.005 2.375 ;
      RECT 72.965 2.2 72.975 2.393 ;
      RECT 72.95 2.211 72.965 2.404 ;
      RECT 72.91 2.235 72.95 2.42 ;
      RECT 72.875 2.269 72.91 2.437 ;
      RECT 72.845 2.292 72.875 2.449 ;
      RECT 72.83 2.302 72.845 2.458 ;
      RECT 72.79 2.312 72.83 2.469 ;
      RECT 72.77 2.323 72.79 2.481 ;
      RECT 72.765 2.327 72.77 2.488 ;
      RECT 72.75 2.331 72.765 2.493 ;
      RECT 72.74 2.336 72.75 2.498 ;
      RECT 72.735 2.339 72.74 2.501 ;
      RECT 72.705 2.345 72.735 2.508 ;
      RECT 72.67 2.355 72.705 2.522 ;
      RECT 72.61 2.37 72.67 2.542 ;
      RECT 72.555 2.39 72.61 2.566 ;
      RECT 72.526 2.405 72.555 2.584 ;
      RECT 72.44 2.425 72.526 2.609 ;
      RECT 72.435 2.44 72.44 2.629 ;
      RECT 72.425 2.443 72.435 2.63 ;
      RECT 72.4 2.45 72.425 2.715 ;
      RECT 75.095 2.943 75.375 3.28 ;
      RECT 75.095 2.953 75.38 3.238 ;
      RECT 75.095 2.962 75.385 3.135 ;
      RECT 75.095 2.977 75.39 3.003 ;
      RECT 75.095 2.805 75.355 3.28 ;
      RECT 65.395 6.655 65.745 7.005 ;
      RECT 74.22 6.61 74.57 6.96 ;
      RECT 65.395 6.685 74.57 6.885 ;
      RECT 72.815 3.685 72.825 3.875 ;
      RECT 71.075 3.56 71.355 3.84 ;
      RECT 74.12 2.5 74.125 2.985 ;
      RECT 74.015 2.5 74.075 2.76 ;
      RECT 74.34 3.47 74.345 3.545 ;
      RECT 74.33 3.337 74.34 3.58 ;
      RECT 74.32 3.172 74.33 3.601 ;
      RECT 74.315 3.042 74.32 3.617 ;
      RECT 74.305 2.932 74.315 3.633 ;
      RECT 74.3 2.831 74.305 3.65 ;
      RECT 74.295 2.813 74.3 3.66 ;
      RECT 74.29 2.795 74.295 3.67 ;
      RECT 74.28 2.77 74.29 3.685 ;
      RECT 74.275 2.75 74.28 3.7 ;
      RECT 74.255 2.5 74.275 3.725 ;
      RECT 74.24 2.5 74.255 3.758 ;
      RECT 74.21 2.5 74.24 3.78 ;
      RECT 74.19 2.5 74.21 3.794 ;
      RECT 74.17 2.5 74.19 3.31 ;
      RECT 74.185 3.377 74.19 3.799 ;
      RECT 74.18 3.407 74.185 3.801 ;
      RECT 74.175 3.42 74.18 3.804 ;
      RECT 74.17 3.43 74.175 3.808 ;
      RECT 74.165 2.5 74.17 3.228 ;
      RECT 74.165 3.44 74.17 3.81 ;
      RECT 74.16 2.5 74.165 3.205 ;
      RECT 74.15 3.462 74.165 3.81 ;
      RECT 74.145 2.5 74.16 3.15 ;
      RECT 74.14 3.487 74.15 3.81 ;
      RECT 74.14 2.5 74.145 3.095 ;
      RECT 74.13 2.5 74.14 3.043 ;
      RECT 74.135 3.5 74.14 3.811 ;
      RECT 74.13 3.512 74.135 3.812 ;
      RECT 74.125 2.5 74.13 3.003 ;
      RECT 74.125 3.525 74.13 3.813 ;
      RECT 74.11 3.54 74.125 3.814 ;
      RECT 74.115 2.5 74.12 2.965 ;
      RECT 74.11 2.5 74.115 2.93 ;
      RECT 74.105 2.5 74.11 2.905 ;
      RECT 74.1 3.567 74.11 3.816 ;
      RECT 74.095 2.5 74.105 2.863 ;
      RECT 74.095 3.585 74.1 3.817 ;
      RECT 74.09 2.5 74.095 2.823 ;
      RECT 74.09 3.592 74.095 3.818 ;
      RECT 74.085 2.5 74.09 2.795 ;
      RECT 74.08 3.61 74.09 3.819 ;
      RECT 74.075 2.5 74.085 2.775 ;
      RECT 74.07 3.63 74.08 3.821 ;
      RECT 74.06 3.647 74.07 3.822 ;
      RECT 74.025 3.67 74.06 3.825 ;
      RECT 73.97 3.688 74.025 3.831 ;
      RECT 73.884 3.696 73.97 3.84 ;
      RECT 73.798 3.707 73.884 3.851 ;
      RECT 73.712 3.717 73.798 3.862 ;
      RECT 73.626 3.727 73.712 3.874 ;
      RECT 73.54 3.737 73.626 3.885 ;
      RECT 73.52 3.743 73.54 3.891 ;
      RECT 73.44 3.745 73.52 3.895 ;
      RECT 73.435 3.744 73.44 3.9 ;
      RECT 73.427 3.743 73.435 3.9 ;
      RECT 73.341 3.739 73.427 3.898 ;
      RECT 73.255 3.731 73.341 3.895 ;
      RECT 73.169 3.722 73.255 3.891 ;
      RECT 73.083 3.714 73.169 3.888 ;
      RECT 72.997 3.706 73.083 3.884 ;
      RECT 72.911 3.697 72.997 3.881 ;
      RECT 72.825 3.689 72.911 3.877 ;
      RECT 72.77 3.682 72.815 3.875 ;
      RECT 72.685 3.675 72.77 3.873 ;
      RECT 72.611 3.667 72.685 3.869 ;
      RECT 72.525 3.659 72.611 3.866 ;
      RECT 72.522 3.655 72.525 3.864 ;
      RECT 72.436 3.651 72.522 3.863 ;
      RECT 72.35 3.643 72.436 3.86 ;
      RECT 72.265 3.638 72.35 3.857 ;
      RECT 72.179 3.635 72.265 3.854 ;
      RECT 72.093 3.633 72.179 3.851 ;
      RECT 72.007 3.63 72.093 3.848 ;
      RECT 71.921 3.627 72.007 3.845 ;
      RECT 71.835 3.624 71.921 3.842 ;
      RECT 71.759 3.622 71.835 3.839 ;
      RECT 71.673 3.619 71.759 3.836 ;
      RECT 71.587 3.616 71.673 3.834 ;
      RECT 71.501 3.614 71.587 3.831 ;
      RECT 71.415 3.611 71.501 3.828 ;
      RECT 71.355 3.602 71.415 3.826 ;
      RECT 73.865 3.22 73.94 3.48 ;
      RECT 73.845 3.2 73.85 3.48 ;
      RECT 73.165 2.985 73.27 3.28 ;
      RECT 67.61 2.96 67.68 3.22 ;
      RECT 73.505 2.835 73.51 3.206 ;
      RECT 73.495 2.89 73.5 3.206 ;
      RECT 73.8 2.06 73.86 2.32 ;
      RECT 73.855 3.215 73.865 3.48 ;
      RECT 73.85 3.205 73.855 3.48 ;
      RECT 73.77 3.152 73.845 3.48 ;
      RECT 73.795 2.06 73.8 2.34 ;
      RECT 73.785 2.06 73.795 2.36 ;
      RECT 73.77 2.06 73.785 2.39 ;
      RECT 73.755 2.06 73.77 2.433 ;
      RECT 73.75 3.095 73.77 3.48 ;
      RECT 73.74 2.06 73.755 2.47 ;
      RECT 73.735 3.075 73.75 3.48 ;
      RECT 73.735 2.06 73.74 2.493 ;
      RECT 73.725 2.06 73.735 2.518 ;
      RECT 73.695 3.042 73.735 3.48 ;
      RECT 73.7 2.06 73.725 2.568 ;
      RECT 73.695 2.06 73.7 2.623 ;
      RECT 73.69 2.06 73.695 2.665 ;
      RECT 73.68 3.005 73.695 3.48 ;
      RECT 73.685 2.06 73.69 2.708 ;
      RECT 73.68 2.06 73.685 2.773 ;
      RECT 73.675 2.06 73.68 2.795 ;
      RECT 73.675 2.993 73.68 3.345 ;
      RECT 73.67 2.06 73.675 2.863 ;
      RECT 73.67 2.985 73.675 3.328 ;
      RECT 73.665 2.06 73.67 2.908 ;
      RECT 73.66 2.967 73.67 3.305 ;
      RECT 73.66 2.06 73.665 2.945 ;
      RECT 73.65 2.06 73.66 3.285 ;
      RECT 73.645 2.06 73.65 3.268 ;
      RECT 73.64 2.06 73.645 3.253 ;
      RECT 73.635 2.06 73.64 3.238 ;
      RECT 73.615 2.06 73.635 3.228 ;
      RECT 73.61 2.06 73.615 3.218 ;
      RECT 73.6 2.06 73.61 3.214 ;
      RECT 73.595 2.337 73.6 3.213 ;
      RECT 73.59 2.36 73.595 3.212 ;
      RECT 73.585 2.39 73.59 3.211 ;
      RECT 73.58 2.417 73.585 3.21 ;
      RECT 73.575 2.445 73.58 3.21 ;
      RECT 73.57 2.472 73.575 3.21 ;
      RECT 73.565 2.492 73.57 3.21 ;
      RECT 73.56 2.52 73.565 3.21 ;
      RECT 73.55 2.562 73.56 3.21 ;
      RECT 73.54 2.607 73.55 3.209 ;
      RECT 73.535 2.66 73.54 3.208 ;
      RECT 73.53 2.692 73.535 3.207 ;
      RECT 73.525 2.712 73.53 3.206 ;
      RECT 73.52 2.75 73.525 3.206 ;
      RECT 73.515 2.772 73.52 3.206 ;
      RECT 73.51 2.797 73.515 3.206 ;
      RECT 73.5 2.862 73.505 3.206 ;
      RECT 73.485 2.922 73.495 3.206 ;
      RECT 73.47 2.932 73.485 3.206 ;
      RECT 73.45 2.942 73.47 3.206 ;
      RECT 73.42 2.947 73.45 3.203 ;
      RECT 73.36 2.957 73.42 3.2 ;
      RECT 73.34 2.966 73.36 3.205 ;
      RECT 73.315 2.972 73.34 3.218 ;
      RECT 73.295 2.977 73.315 3.233 ;
      RECT 73.27 2.982 73.295 3.28 ;
      RECT 73.141 2.984 73.165 3.28 ;
      RECT 73.055 2.979 73.141 3.28 ;
      RECT 73.015 2.976 73.055 3.28 ;
      RECT 72.965 2.978 73.015 3.26 ;
      RECT 72.935 2.982 72.965 3.26 ;
      RECT 72.856 2.992 72.935 3.26 ;
      RECT 72.77 3.007 72.856 3.261 ;
      RECT 72.72 3.017 72.77 3.262 ;
      RECT 72.712 3.02 72.72 3.262 ;
      RECT 72.626 3.022 72.712 3.263 ;
      RECT 72.54 3.026 72.626 3.263 ;
      RECT 72.454 3.03 72.54 3.264 ;
      RECT 72.368 3.033 72.454 3.265 ;
      RECT 72.282 3.037 72.368 3.265 ;
      RECT 72.196 3.041 72.282 3.266 ;
      RECT 72.11 3.044 72.196 3.267 ;
      RECT 72.024 3.048 72.11 3.267 ;
      RECT 71.938 3.052 72.024 3.268 ;
      RECT 71.852 3.056 71.938 3.269 ;
      RECT 71.766 3.059 71.852 3.269 ;
      RECT 71.68 3.063 71.766 3.27 ;
      RECT 71.65 3.065 71.68 3.27 ;
      RECT 71.564 3.068 71.65 3.271 ;
      RECT 71.478 3.072 71.564 3.272 ;
      RECT 71.392 3.076 71.478 3.273 ;
      RECT 71.306 3.079 71.392 3.273 ;
      RECT 71.22 3.083 71.306 3.274 ;
      RECT 71.185 3.088 71.22 3.275 ;
      RECT 71.13 3.098 71.185 3.282 ;
      RECT 71.105 3.11 71.13 3.292 ;
      RECT 71.07 3.123 71.105 3.3 ;
      RECT 71.03 3.14 71.07 3.323 ;
      RECT 71.01 3.153 71.03 3.35 ;
      RECT 70.98 3.165 71.01 3.378 ;
      RECT 70.975 3.173 70.98 3.398 ;
      RECT 70.97 3.176 70.975 3.408 ;
      RECT 70.92 3.188 70.97 3.442 ;
      RECT 70.91 3.203 70.92 3.475 ;
      RECT 70.9 3.209 70.91 3.488 ;
      RECT 70.89 3.216 70.9 3.5 ;
      RECT 70.865 3.229 70.89 3.518 ;
      RECT 70.85 3.244 70.865 3.54 ;
      RECT 70.84 3.252 70.85 3.556 ;
      RECT 70.825 3.261 70.84 3.571 ;
      RECT 70.815 3.271 70.825 3.585 ;
      RECT 70.796 3.284 70.815 3.602 ;
      RECT 70.71 3.329 70.796 3.667 ;
      RECT 70.695 3.374 70.71 3.725 ;
      RECT 70.69 3.383 70.695 3.738 ;
      RECT 70.68 3.39 70.69 3.743 ;
      RECT 70.675 3.395 70.68 3.747 ;
      RECT 70.655 3.405 70.675 3.754 ;
      RECT 70.63 3.425 70.655 3.768 ;
      RECT 70.595 3.45 70.63 3.788 ;
      RECT 70.58 3.473 70.595 3.803 ;
      RECT 70.57 3.483 70.58 3.808 ;
      RECT 70.56 3.491 70.57 3.815 ;
      RECT 70.55 3.5 70.56 3.821 ;
      RECT 70.53 3.512 70.55 3.823 ;
      RECT 70.52 3.525 70.53 3.825 ;
      RECT 70.495 3.54 70.52 3.828 ;
      RECT 70.475 3.557 70.495 3.832 ;
      RECT 70.435 3.585 70.475 3.838 ;
      RECT 70.37 3.632 70.435 3.847 ;
      RECT 70.355 3.665 70.37 3.855 ;
      RECT 70.35 3.672 70.355 3.857 ;
      RECT 70.3 3.697 70.35 3.862 ;
      RECT 70.285 3.721 70.3 3.869 ;
      RECT 70.235 3.726 70.285 3.87 ;
      RECT 70.149 3.73 70.235 3.87 ;
      RECT 70.063 3.73 70.149 3.87 ;
      RECT 69.977 3.73 70.063 3.871 ;
      RECT 69.891 3.73 69.977 3.871 ;
      RECT 69.805 3.73 69.891 3.871 ;
      RECT 69.739 3.73 69.805 3.871 ;
      RECT 69.653 3.73 69.739 3.872 ;
      RECT 69.567 3.73 69.653 3.872 ;
      RECT 69.481 3.731 69.567 3.873 ;
      RECT 69.395 3.731 69.481 3.873 ;
      RECT 69.309 3.731 69.395 3.873 ;
      RECT 69.223 3.731 69.309 3.874 ;
      RECT 69.137 3.731 69.223 3.874 ;
      RECT 69.051 3.732 69.137 3.875 ;
      RECT 68.965 3.732 69.051 3.875 ;
      RECT 68.945 3.732 68.965 3.875 ;
      RECT 68.859 3.732 68.945 3.875 ;
      RECT 68.773 3.732 68.859 3.875 ;
      RECT 68.687 3.733 68.773 3.875 ;
      RECT 68.601 3.733 68.687 3.875 ;
      RECT 68.515 3.733 68.601 3.875 ;
      RECT 68.429 3.734 68.515 3.875 ;
      RECT 68.343 3.734 68.429 3.875 ;
      RECT 68.257 3.734 68.343 3.875 ;
      RECT 68.171 3.734 68.257 3.875 ;
      RECT 68.085 3.735 68.171 3.875 ;
      RECT 68.035 3.732 68.085 3.875 ;
      RECT 68.025 3.73 68.035 3.874 ;
      RECT 68.021 3.73 68.025 3.873 ;
      RECT 67.935 3.725 68.021 3.868 ;
      RECT 67.913 3.718 67.935 3.862 ;
      RECT 67.827 3.709 67.913 3.856 ;
      RECT 67.741 3.696 67.827 3.847 ;
      RECT 67.655 3.682 67.741 3.837 ;
      RECT 67.61 3.672 67.655 3.83 ;
      RECT 67.59 2.96 67.61 3.238 ;
      RECT 67.59 3.665 67.61 3.826 ;
      RECT 67.56 2.96 67.59 3.26 ;
      RECT 67.55 3.632 67.59 3.823 ;
      RECT 67.545 2.96 67.56 3.28 ;
      RECT 67.545 3.597 67.55 3.821 ;
      RECT 67.54 2.96 67.545 3.405 ;
      RECT 67.54 3.557 67.545 3.821 ;
      RECT 67.53 2.96 67.54 3.821 ;
      RECT 67.455 2.96 67.53 3.815 ;
      RECT 67.425 2.96 67.455 3.805 ;
      RECT 67.42 2.96 67.425 3.797 ;
      RECT 67.415 3.002 67.42 3.79 ;
      RECT 67.405 3.071 67.415 3.781 ;
      RECT 67.4 3.141 67.405 3.733 ;
      RECT 67.395 3.205 67.4 3.63 ;
      RECT 67.39 3.24 67.395 3.585 ;
      RECT 67.388 3.277 67.39 3.477 ;
      RECT 67.385 3.285 67.388 3.47 ;
      RECT 67.38 3.35 67.385 3.413 ;
      RECT 71.455 2.44 71.735 2.72 ;
      RECT 71.445 2.44 71.735 2.583 ;
      RECT 71.4 2.305 71.66 2.565 ;
      RECT 71.4 2.42 71.715 2.565 ;
      RECT 71.4 2.39 71.71 2.565 ;
      RECT 71.4 2.377 71.7 2.565 ;
      RECT 71.4 2.367 71.695 2.565 ;
      RECT 67.375 2.35 67.635 2.61 ;
      RECT 71.145 1.9 71.405 2.16 ;
      RECT 71.135 1.925 71.405 2.12 ;
      RECT 71.13 1.925 71.135 2.119 ;
      RECT 71.06 1.92 71.13 2.111 ;
      RECT 70.975 1.907 71.06 2.094 ;
      RECT 70.971 1.899 70.975 2.084 ;
      RECT 70.885 1.892 70.971 2.074 ;
      RECT 70.876 1.884 70.885 2.064 ;
      RECT 70.79 1.877 70.876 2.052 ;
      RECT 70.77 1.868 70.79 2.038 ;
      RECT 70.715 1.863 70.77 2.03 ;
      RECT 70.705 1.857 70.715 2.024 ;
      RECT 70.685 1.855 70.705 2.02 ;
      RECT 70.677 1.854 70.685 2.016 ;
      RECT 70.591 1.846 70.677 2.005 ;
      RECT 70.505 1.832 70.591 1.985 ;
      RECT 70.445 1.82 70.505 1.97 ;
      RECT 70.435 1.815 70.445 1.965 ;
      RECT 70.385 1.815 70.435 1.967 ;
      RECT 70.338 1.817 70.385 1.971 ;
      RECT 70.252 1.824 70.338 1.976 ;
      RECT 70.166 1.832 70.252 1.982 ;
      RECT 70.08 1.841 70.166 1.988 ;
      RECT 70.021 1.847 70.08 1.993 ;
      RECT 69.935 1.852 70.021 1.999 ;
      RECT 69.86 1.857 69.935 2.005 ;
      RECT 69.821 1.859 69.86 2.01 ;
      RECT 69.735 1.856 69.821 2.015 ;
      RECT 69.65 1.854 69.735 2.022 ;
      RECT 69.618 1.853 69.65 2.025 ;
      RECT 69.532 1.852 69.618 2.026 ;
      RECT 69.446 1.851 69.532 2.027 ;
      RECT 69.36 1.85 69.446 2.027 ;
      RECT 69.274 1.849 69.36 2.028 ;
      RECT 69.188 1.848 69.274 2.029 ;
      RECT 69.102 1.847 69.188 2.03 ;
      RECT 69.016 1.846 69.102 2.03 ;
      RECT 68.93 1.845 69.016 2.031 ;
      RECT 68.88 1.845 68.93 2.032 ;
      RECT 68.866 1.846 68.88 2.032 ;
      RECT 68.78 1.853 68.866 2.033 ;
      RECT 68.706 1.864 68.78 2.034 ;
      RECT 68.62 1.873 68.706 2.035 ;
      RECT 68.585 1.88 68.62 2.05 ;
      RECT 68.56 1.883 68.585 2.08 ;
      RECT 68.535 1.892 68.56 2.109 ;
      RECT 68.525 1.903 68.535 2.129 ;
      RECT 68.515 1.911 68.525 2.143 ;
      RECT 68.51 1.917 68.515 2.153 ;
      RECT 68.485 1.934 68.51 2.17 ;
      RECT 68.47 1.956 68.485 2.198 ;
      RECT 68.44 1.982 68.47 2.228 ;
      RECT 68.42 2.011 68.44 2.258 ;
      RECT 68.415 2.026 68.42 2.275 ;
      RECT 68.395 2.041 68.415 2.29 ;
      RECT 68.385 2.059 68.395 2.308 ;
      RECT 68.375 2.07 68.385 2.323 ;
      RECT 68.325 2.102 68.375 2.349 ;
      RECT 68.32 2.132 68.325 2.369 ;
      RECT 68.31 2.145 68.32 2.375 ;
      RECT 68.301 2.155 68.31 2.383 ;
      RECT 68.29 2.166 68.301 2.391 ;
      RECT 68.285 2.176 68.29 2.397 ;
      RECT 68.27 2.197 68.285 2.404 ;
      RECT 68.255 2.227 68.27 2.412 ;
      RECT 68.22 2.257 68.255 2.418 ;
      RECT 68.195 2.275 68.22 2.425 ;
      RECT 68.145 2.283 68.195 2.434 ;
      RECT 68.12 2.288 68.145 2.443 ;
      RECT 68.065 2.294 68.12 2.453 ;
      RECT 68.06 2.299 68.065 2.461 ;
      RECT 68.046 2.302 68.06 2.463 ;
      RECT 67.96 2.314 68.046 2.475 ;
      RECT 67.95 2.326 67.96 2.488 ;
      RECT 67.865 2.339 67.95 2.5 ;
      RECT 67.821 2.356 67.865 2.514 ;
      RECT 67.735 2.373 67.821 2.53 ;
      RECT 67.705 2.387 67.735 2.544 ;
      RECT 67.695 2.392 67.705 2.549 ;
      RECT 67.635 2.395 67.695 2.558 ;
      RECT 70.525 2.665 70.785 2.925 ;
      RECT 70.525 2.665 70.805 2.778 ;
      RECT 70.525 2.665 70.83 2.745 ;
      RECT 70.525 2.665 70.835 2.725 ;
      RECT 70.575 2.44 70.855 2.72 ;
      RECT 70.13 3.175 70.39 3.435 ;
      RECT 70.12 3.032 70.315 3.373 ;
      RECT 70.115 3.14 70.33 3.365 ;
      RECT 70.11 3.19 70.39 3.355 ;
      RECT 70.1 3.267 70.39 3.34 ;
      RECT 70.12 3.115 70.33 3.373 ;
      RECT 70.13 2.99 70.315 3.435 ;
      RECT 70.13 2.885 70.295 3.435 ;
      RECT 70.14 2.872 70.295 3.435 ;
      RECT 70.14 2.83 70.285 3.435 ;
      RECT 70.145 2.755 70.285 3.435 ;
      RECT 70.175 2.405 70.285 3.435 ;
      RECT 70.18 2.135 70.305 2.758 ;
      RECT 70.15 2.71 70.305 2.758 ;
      RECT 70.165 2.512 70.285 3.435 ;
      RECT 70.155 2.622 70.305 2.758 ;
      RECT 70.18 2.135 70.32 2.615 ;
      RECT 70.18 2.135 70.34 2.49 ;
      RECT 70.145 2.135 70.405 2.395 ;
      RECT 69.615 2.44 69.895 2.72 ;
      RECT 69.6 2.44 69.895 2.7 ;
      RECT 67.655 3.305 67.915 3.565 ;
      RECT 69.44 3.16 69.7 3.42 ;
      RECT 69.42 3.18 69.7 3.395 ;
      RECT 69.377 3.18 69.42 3.394 ;
      RECT 69.291 3.181 69.377 3.391 ;
      RECT 69.205 3.182 69.291 3.387 ;
      RECT 69.13 3.184 69.205 3.384 ;
      RECT 69.107 3.185 69.13 3.382 ;
      RECT 69.021 3.186 69.107 3.38 ;
      RECT 68.935 3.187 69.021 3.377 ;
      RECT 68.911 3.188 68.935 3.375 ;
      RECT 68.825 3.19 68.911 3.372 ;
      RECT 68.74 3.192 68.825 3.373 ;
      RECT 68.683 3.193 68.74 3.379 ;
      RECT 68.597 3.195 68.683 3.389 ;
      RECT 68.511 3.198 68.597 3.402 ;
      RECT 68.425 3.2 68.511 3.414 ;
      RECT 68.411 3.201 68.425 3.421 ;
      RECT 68.325 3.202 68.411 3.429 ;
      RECT 68.285 3.204 68.325 3.438 ;
      RECT 68.276 3.205 68.285 3.441 ;
      RECT 68.19 3.213 68.276 3.447 ;
      RECT 68.17 3.222 68.19 3.455 ;
      RECT 68.085 3.237 68.17 3.463 ;
      RECT 68.025 3.26 68.085 3.474 ;
      RECT 68.015 3.272 68.025 3.479 ;
      RECT 67.975 3.282 68.015 3.483 ;
      RECT 67.92 3.299 67.975 3.491 ;
      RECT 67.915 3.309 67.92 3.495 ;
      RECT 68.981 2.44 69.04 2.837 ;
      RECT 68.895 2.44 69.1 2.828 ;
      RECT 68.89 2.47 69.1 2.823 ;
      RECT 68.856 2.47 69.1 2.821 ;
      RECT 68.77 2.47 69.1 2.815 ;
      RECT 68.725 2.47 69.12 2.793 ;
      RECT 68.725 2.47 69.14 2.748 ;
      RECT 68.685 2.47 69.14 2.738 ;
      RECT 68.895 2.44 69.175 2.72 ;
      RECT 68.63 2.44 68.89 2.7 ;
      RECT 66.455 3 66.735 3.28 ;
      RECT 66.425 2.962 66.68 3.265 ;
      RECT 66.42 2.963 66.68 3.263 ;
      RECT 66.415 2.964 66.68 3.257 ;
      RECT 66.41 2.967 66.68 3.25 ;
      RECT 66.405 3 66.735 3.243 ;
      RECT 66.375 2.97 66.68 3.23 ;
      RECT 66.375 2.997 66.7 3.23 ;
      RECT 66.375 2.987 66.695 3.23 ;
      RECT 66.375 2.972 66.69 3.23 ;
      RECT 66.455 2.959 66.67 3.28 ;
      RECT 66.541 2.957 66.67 3.28 ;
      RECT 66.627 2.955 66.655 3.28 ;
      RECT 62.26 6.22 62.58 6.545 ;
      RECT 62.29 5.695 62.46 6.545 ;
      RECT 62.29 5.695 62.465 6.045 ;
      RECT 62.29 5.695 63.265 5.87 ;
      RECT 63.09 1.965 63.265 5.87 ;
      RECT 63.035 1.965 63.385 2.315 ;
      RECT 63.06 6.655 63.385 6.98 ;
      RECT 61.945 6.745 63.385 6.915 ;
      RECT 61.945 2.395 62.105 6.915 ;
      RECT 62.26 2.365 62.58 2.685 ;
      RECT 61.945 2.395 62.58 2.565 ;
      RECT 61.21 5.855 61.56 6.205 ;
      RECT 61.28 2.705 61.455 6.205 ;
      RECT 61.205 2.705 61.555 3.055 ;
      RECT 52.03 1.92 52.29 2.18 ;
      RECT 52.085 1.88 52.39 2.16 ;
      RECT 52.085 1.42 52.26 2.18 ;
      RECT 60.6 1.34 60.95 1.69 ;
      RECT 52.085 1.42 60.95 1.595 ;
      RECT 60.275 2.85 60.645 3.22 ;
      RECT 60.36 2.235 60.53 3.22 ;
      RECT 56.38 2.455 56.615 2.715 ;
      RECT 59.525 2.235 59.69 2.495 ;
      RECT 59.43 2.225 59.445 2.495 ;
      RECT 59.525 2.235 60.53 2.415 ;
      RECT 58.03 1.795 58.07 1.935 ;
      RECT 59.445 2.23 59.525 2.495 ;
      RECT 59.39 2.225 59.43 2.461 ;
      RECT 59.376 2.225 59.39 2.461 ;
      RECT 59.29 2.23 59.376 2.463 ;
      RECT 59.245 2.237 59.29 2.465 ;
      RECT 59.215 2.237 59.245 2.467 ;
      RECT 59.19 2.232 59.215 2.469 ;
      RECT 59.16 2.228 59.19 2.478 ;
      RECT 59.15 2.225 59.16 2.49 ;
      RECT 59.145 2.225 59.15 2.498 ;
      RECT 59.14 2.225 59.145 2.503 ;
      RECT 59.13 2.224 59.14 2.513 ;
      RECT 59.125 2.223 59.13 2.523 ;
      RECT 59.11 2.222 59.125 2.528 ;
      RECT 59.082 2.219 59.11 2.555 ;
      RECT 58.996 2.211 59.082 2.555 ;
      RECT 58.91 2.2 58.996 2.555 ;
      RECT 58.87 2.185 58.91 2.555 ;
      RECT 58.83 2.159 58.87 2.555 ;
      RECT 58.825 2.141 58.83 2.367 ;
      RECT 58.815 2.137 58.825 2.357 ;
      RECT 58.8 2.127 58.815 2.344 ;
      RECT 58.78 2.111 58.8 2.329 ;
      RECT 58.765 2.096 58.78 2.314 ;
      RECT 58.755 2.085 58.765 2.304 ;
      RECT 58.73 2.069 58.755 2.293 ;
      RECT 58.725 2.056 58.73 2.283 ;
      RECT 58.72 2.052 58.725 2.278 ;
      RECT 58.665 2.038 58.72 2.256 ;
      RECT 58.626 2.019 58.665 2.22 ;
      RECT 58.54 1.993 58.626 2.173 ;
      RECT 58.536 1.975 58.54 2.139 ;
      RECT 58.45 1.956 58.536 2.117 ;
      RECT 58.445 1.938 58.45 2.095 ;
      RECT 58.44 1.936 58.445 2.093 ;
      RECT 58.43 1.935 58.44 2.088 ;
      RECT 58.37 1.922 58.43 2.074 ;
      RECT 58.325 1.9 58.37 2.053 ;
      RECT 58.265 1.877 58.325 2.032 ;
      RECT 58.201 1.852 58.265 2.007 ;
      RECT 58.115 1.822 58.201 1.976 ;
      RECT 58.1 1.802 58.115 1.955 ;
      RECT 58.07 1.797 58.1 1.946 ;
      RECT 58.017 1.795 58.03 1.935 ;
      RECT 57.931 1.795 58.017 1.937 ;
      RECT 57.845 1.795 57.931 1.939 ;
      RECT 57.825 1.795 57.845 1.943 ;
      RECT 57.78 1.797 57.825 1.954 ;
      RECT 57.74 1.807 57.78 1.97 ;
      RECT 57.736 1.816 57.74 1.978 ;
      RECT 57.65 1.836 57.736 1.994 ;
      RECT 57.64 1.855 57.65 2.012 ;
      RECT 57.635 1.857 57.64 2.015 ;
      RECT 57.625 1.861 57.635 2.018 ;
      RECT 57.605 1.866 57.625 2.028 ;
      RECT 57.575 1.876 57.605 2.048 ;
      RECT 57.57 1.883 57.575 2.062 ;
      RECT 57.56 1.887 57.57 2.069 ;
      RECT 57.545 1.895 57.56 2.08 ;
      RECT 57.535 1.905 57.545 2.091 ;
      RECT 57.525 1.912 57.535 2.099 ;
      RECT 57.5 1.925 57.525 2.114 ;
      RECT 57.436 1.961 57.5 2.153 ;
      RECT 57.35 2.024 57.436 2.217 ;
      RECT 57.315 2.075 57.35 2.27 ;
      RECT 57.31 2.092 57.315 2.287 ;
      RECT 57.295 2.101 57.31 2.294 ;
      RECT 57.275 2.116 57.295 2.308 ;
      RECT 57.27 2.127 57.275 2.318 ;
      RECT 57.25 2.14 57.27 2.328 ;
      RECT 57.245 2.15 57.25 2.338 ;
      RECT 57.23 2.155 57.245 2.347 ;
      RECT 57.22 2.165 57.23 2.358 ;
      RECT 57.19 2.182 57.22 2.375 ;
      RECT 57.18 2.2 57.19 2.393 ;
      RECT 57.165 2.211 57.18 2.404 ;
      RECT 57.125 2.235 57.165 2.42 ;
      RECT 57.09 2.269 57.125 2.437 ;
      RECT 57.06 2.292 57.09 2.449 ;
      RECT 57.045 2.302 57.06 2.458 ;
      RECT 57.005 2.312 57.045 2.469 ;
      RECT 56.985 2.323 57.005 2.481 ;
      RECT 56.98 2.327 56.985 2.488 ;
      RECT 56.965 2.331 56.98 2.493 ;
      RECT 56.955 2.336 56.965 2.498 ;
      RECT 56.95 2.339 56.955 2.501 ;
      RECT 56.92 2.345 56.95 2.508 ;
      RECT 56.885 2.355 56.92 2.522 ;
      RECT 56.825 2.37 56.885 2.542 ;
      RECT 56.77 2.39 56.825 2.566 ;
      RECT 56.741 2.405 56.77 2.584 ;
      RECT 56.655 2.425 56.741 2.609 ;
      RECT 56.65 2.44 56.655 2.629 ;
      RECT 56.64 2.443 56.65 2.63 ;
      RECT 56.615 2.45 56.64 2.715 ;
      RECT 59.31 2.943 59.59 3.28 ;
      RECT 59.31 2.953 59.595 3.238 ;
      RECT 59.31 2.962 59.6 3.135 ;
      RECT 59.31 2.977 59.605 3.003 ;
      RECT 59.31 2.805 59.57 3.28 ;
      RECT 49.61 6.655 49.96 7.005 ;
      RECT 58.435 6.61 58.785 6.96 ;
      RECT 49.61 6.685 58.785 6.885 ;
      RECT 57.03 3.685 57.04 3.875 ;
      RECT 55.29 3.56 55.57 3.84 ;
      RECT 58.335 2.5 58.34 2.985 ;
      RECT 58.23 2.5 58.29 2.76 ;
      RECT 58.555 3.47 58.56 3.545 ;
      RECT 58.545 3.337 58.555 3.58 ;
      RECT 58.535 3.172 58.545 3.601 ;
      RECT 58.53 3.042 58.535 3.617 ;
      RECT 58.52 2.932 58.53 3.633 ;
      RECT 58.515 2.831 58.52 3.65 ;
      RECT 58.51 2.813 58.515 3.66 ;
      RECT 58.505 2.795 58.51 3.67 ;
      RECT 58.495 2.77 58.505 3.685 ;
      RECT 58.49 2.75 58.495 3.7 ;
      RECT 58.47 2.5 58.49 3.725 ;
      RECT 58.455 2.5 58.47 3.758 ;
      RECT 58.425 2.5 58.455 3.78 ;
      RECT 58.405 2.5 58.425 3.794 ;
      RECT 58.385 2.5 58.405 3.31 ;
      RECT 58.4 3.377 58.405 3.799 ;
      RECT 58.395 3.407 58.4 3.801 ;
      RECT 58.39 3.42 58.395 3.804 ;
      RECT 58.385 3.43 58.39 3.808 ;
      RECT 58.38 2.5 58.385 3.228 ;
      RECT 58.38 3.44 58.385 3.81 ;
      RECT 58.375 2.5 58.38 3.205 ;
      RECT 58.365 3.462 58.38 3.81 ;
      RECT 58.36 2.5 58.375 3.15 ;
      RECT 58.355 3.487 58.365 3.81 ;
      RECT 58.355 2.5 58.36 3.095 ;
      RECT 58.345 2.5 58.355 3.043 ;
      RECT 58.35 3.5 58.355 3.811 ;
      RECT 58.345 3.512 58.35 3.812 ;
      RECT 58.34 2.5 58.345 3.003 ;
      RECT 58.34 3.525 58.345 3.813 ;
      RECT 58.325 3.54 58.34 3.814 ;
      RECT 58.33 2.5 58.335 2.965 ;
      RECT 58.325 2.5 58.33 2.93 ;
      RECT 58.32 2.5 58.325 2.905 ;
      RECT 58.315 3.567 58.325 3.816 ;
      RECT 58.31 2.5 58.32 2.863 ;
      RECT 58.31 3.585 58.315 3.817 ;
      RECT 58.305 2.5 58.31 2.823 ;
      RECT 58.305 3.592 58.31 3.818 ;
      RECT 58.3 2.5 58.305 2.795 ;
      RECT 58.295 3.61 58.305 3.819 ;
      RECT 58.29 2.5 58.3 2.775 ;
      RECT 58.285 3.63 58.295 3.821 ;
      RECT 58.275 3.647 58.285 3.822 ;
      RECT 58.24 3.67 58.275 3.825 ;
      RECT 58.185 3.688 58.24 3.831 ;
      RECT 58.099 3.696 58.185 3.84 ;
      RECT 58.013 3.707 58.099 3.851 ;
      RECT 57.927 3.717 58.013 3.862 ;
      RECT 57.841 3.727 57.927 3.874 ;
      RECT 57.755 3.737 57.841 3.885 ;
      RECT 57.735 3.743 57.755 3.891 ;
      RECT 57.655 3.745 57.735 3.895 ;
      RECT 57.65 3.744 57.655 3.9 ;
      RECT 57.642 3.743 57.65 3.9 ;
      RECT 57.556 3.739 57.642 3.898 ;
      RECT 57.47 3.731 57.556 3.895 ;
      RECT 57.384 3.722 57.47 3.891 ;
      RECT 57.298 3.714 57.384 3.888 ;
      RECT 57.212 3.706 57.298 3.884 ;
      RECT 57.126 3.697 57.212 3.881 ;
      RECT 57.04 3.689 57.126 3.877 ;
      RECT 56.985 3.682 57.03 3.875 ;
      RECT 56.9 3.675 56.985 3.873 ;
      RECT 56.826 3.667 56.9 3.869 ;
      RECT 56.74 3.659 56.826 3.866 ;
      RECT 56.737 3.655 56.74 3.864 ;
      RECT 56.651 3.651 56.737 3.863 ;
      RECT 56.565 3.643 56.651 3.86 ;
      RECT 56.48 3.638 56.565 3.857 ;
      RECT 56.394 3.635 56.48 3.854 ;
      RECT 56.308 3.633 56.394 3.851 ;
      RECT 56.222 3.63 56.308 3.848 ;
      RECT 56.136 3.627 56.222 3.845 ;
      RECT 56.05 3.624 56.136 3.842 ;
      RECT 55.974 3.622 56.05 3.839 ;
      RECT 55.888 3.619 55.974 3.836 ;
      RECT 55.802 3.616 55.888 3.834 ;
      RECT 55.716 3.614 55.802 3.831 ;
      RECT 55.63 3.611 55.716 3.828 ;
      RECT 55.57 3.602 55.63 3.826 ;
      RECT 58.08 3.22 58.155 3.48 ;
      RECT 58.06 3.2 58.065 3.48 ;
      RECT 57.38 2.985 57.485 3.28 ;
      RECT 51.825 2.96 51.895 3.22 ;
      RECT 57.72 2.835 57.725 3.206 ;
      RECT 57.71 2.89 57.715 3.206 ;
      RECT 58.015 2.06 58.075 2.32 ;
      RECT 58.07 3.215 58.08 3.48 ;
      RECT 58.065 3.205 58.07 3.48 ;
      RECT 57.985 3.152 58.06 3.48 ;
      RECT 58.01 2.06 58.015 2.34 ;
      RECT 58 2.06 58.01 2.36 ;
      RECT 57.985 2.06 58 2.39 ;
      RECT 57.97 2.06 57.985 2.433 ;
      RECT 57.965 3.095 57.985 3.48 ;
      RECT 57.955 2.06 57.97 2.47 ;
      RECT 57.95 3.075 57.965 3.48 ;
      RECT 57.95 2.06 57.955 2.493 ;
      RECT 57.94 2.06 57.95 2.518 ;
      RECT 57.91 3.042 57.95 3.48 ;
      RECT 57.915 2.06 57.94 2.568 ;
      RECT 57.91 2.06 57.915 2.623 ;
      RECT 57.905 2.06 57.91 2.665 ;
      RECT 57.895 3.005 57.91 3.48 ;
      RECT 57.9 2.06 57.905 2.708 ;
      RECT 57.895 2.06 57.9 2.773 ;
      RECT 57.89 2.06 57.895 2.795 ;
      RECT 57.89 2.993 57.895 3.345 ;
      RECT 57.885 2.06 57.89 2.863 ;
      RECT 57.885 2.985 57.89 3.328 ;
      RECT 57.88 2.06 57.885 2.908 ;
      RECT 57.875 2.967 57.885 3.305 ;
      RECT 57.875 2.06 57.88 2.945 ;
      RECT 57.865 2.06 57.875 3.285 ;
      RECT 57.86 2.06 57.865 3.268 ;
      RECT 57.855 2.06 57.86 3.253 ;
      RECT 57.85 2.06 57.855 3.238 ;
      RECT 57.83 2.06 57.85 3.228 ;
      RECT 57.825 2.06 57.83 3.218 ;
      RECT 57.815 2.06 57.825 3.214 ;
      RECT 57.81 2.337 57.815 3.213 ;
      RECT 57.805 2.36 57.81 3.212 ;
      RECT 57.8 2.39 57.805 3.211 ;
      RECT 57.795 2.417 57.8 3.21 ;
      RECT 57.79 2.445 57.795 3.21 ;
      RECT 57.785 2.472 57.79 3.21 ;
      RECT 57.78 2.492 57.785 3.21 ;
      RECT 57.775 2.52 57.78 3.21 ;
      RECT 57.765 2.562 57.775 3.21 ;
      RECT 57.755 2.607 57.765 3.209 ;
      RECT 57.75 2.66 57.755 3.208 ;
      RECT 57.745 2.692 57.75 3.207 ;
      RECT 57.74 2.712 57.745 3.206 ;
      RECT 57.735 2.75 57.74 3.206 ;
      RECT 57.73 2.772 57.735 3.206 ;
      RECT 57.725 2.797 57.73 3.206 ;
      RECT 57.715 2.862 57.72 3.206 ;
      RECT 57.7 2.922 57.71 3.206 ;
      RECT 57.685 2.932 57.7 3.206 ;
      RECT 57.665 2.942 57.685 3.206 ;
      RECT 57.635 2.947 57.665 3.203 ;
      RECT 57.575 2.957 57.635 3.2 ;
      RECT 57.555 2.966 57.575 3.205 ;
      RECT 57.53 2.972 57.555 3.218 ;
      RECT 57.51 2.977 57.53 3.233 ;
      RECT 57.485 2.982 57.51 3.28 ;
      RECT 57.356 2.984 57.38 3.28 ;
      RECT 57.27 2.979 57.356 3.28 ;
      RECT 57.23 2.976 57.27 3.28 ;
      RECT 57.18 2.978 57.23 3.26 ;
      RECT 57.15 2.982 57.18 3.26 ;
      RECT 57.071 2.992 57.15 3.26 ;
      RECT 56.985 3.007 57.071 3.261 ;
      RECT 56.935 3.017 56.985 3.262 ;
      RECT 56.927 3.02 56.935 3.262 ;
      RECT 56.841 3.022 56.927 3.263 ;
      RECT 56.755 3.026 56.841 3.263 ;
      RECT 56.669 3.03 56.755 3.264 ;
      RECT 56.583 3.033 56.669 3.265 ;
      RECT 56.497 3.037 56.583 3.265 ;
      RECT 56.411 3.041 56.497 3.266 ;
      RECT 56.325 3.044 56.411 3.267 ;
      RECT 56.239 3.048 56.325 3.267 ;
      RECT 56.153 3.052 56.239 3.268 ;
      RECT 56.067 3.056 56.153 3.269 ;
      RECT 55.981 3.059 56.067 3.269 ;
      RECT 55.895 3.063 55.981 3.27 ;
      RECT 55.865 3.065 55.895 3.27 ;
      RECT 55.779 3.068 55.865 3.271 ;
      RECT 55.693 3.072 55.779 3.272 ;
      RECT 55.607 3.076 55.693 3.273 ;
      RECT 55.521 3.079 55.607 3.273 ;
      RECT 55.435 3.083 55.521 3.274 ;
      RECT 55.4 3.088 55.435 3.275 ;
      RECT 55.345 3.098 55.4 3.282 ;
      RECT 55.32 3.11 55.345 3.292 ;
      RECT 55.285 3.123 55.32 3.3 ;
      RECT 55.245 3.14 55.285 3.323 ;
      RECT 55.225 3.153 55.245 3.35 ;
      RECT 55.195 3.165 55.225 3.378 ;
      RECT 55.19 3.173 55.195 3.398 ;
      RECT 55.185 3.176 55.19 3.408 ;
      RECT 55.135 3.188 55.185 3.442 ;
      RECT 55.125 3.203 55.135 3.475 ;
      RECT 55.115 3.209 55.125 3.488 ;
      RECT 55.105 3.216 55.115 3.5 ;
      RECT 55.08 3.229 55.105 3.518 ;
      RECT 55.065 3.244 55.08 3.54 ;
      RECT 55.055 3.252 55.065 3.556 ;
      RECT 55.04 3.261 55.055 3.571 ;
      RECT 55.03 3.271 55.04 3.585 ;
      RECT 55.011 3.284 55.03 3.602 ;
      RECT 54.925 3.329 55.011 3.667 ;
      RECT 54.91 3.374 54.925 3.725 ;
      RECT 54.905 3.383 54.91 3.738 ;
      RECT 54.895 3.39 54.905 3.743 ;
      RECT 54.89 3.395 54.895 3.747 ;
      RECT 54.87 3.405 54.89 3.754 ;
      RECT 54.845 3.425 54.87 3.768 ;
      RECT 54.81 3.45 54.845 3.788 ;
      RECT 54.795 3.473 54.81 3.803 ;
      RECT 54.785 3.483 54.795 3.808 ;
      RECT 54.775 3.491 54.785 3.815 ;
      RECT 54.765 3.5 54.775 3.821 ;
      RECT 54.745 3.512 54.765 3.823 ;
      RECT 54.735 3.525 54.745 3.825 ;
      RECT 54.71 3.54 54.735 3.828 ;
      RECT 54.69 3.557 54.71 3.832 ;
      RECT 54.65 3.585 54.69 3.838 ;
      RECT 54.585 3.632 54.65 3.847 ;
      RECT 54.57 3.665 54.585 3.855 ;
      RECT 54.565 3.672 54.57 3.857 ;
      RECT 54.515 3.697 54.565 3.862 ;
      RECT 54.5 3.721 54.515 3.869 ;
      RECT 54.45 3.726 54.5 3.87 ;
      RECT 54.364 3.73 54.45 3.87 ;
      RECT 54.278 3.73 54.364 3.87 ;
      RECT 54.192 3.73 54.278 3.871 ;
      RECT 54.106 3.73 54.192 3.871 ;
      RECT 54.02 3.73 54.106 3.871 ;
      RECT 53.954 3.73 54.02 3.871 ;
      RECT 53.868 3.73 53.954 3.872 ;
      RECT 53.782 3.73 53.868 3.872 ;
      RECT 53.696 3.731 53.782 3.873 ;
      RECT 53.61 3.731 53.696 3.873 ;
      RECT 53.524 3.731 53.61 3.873 ;
      RECT 53.438 3.731 53.524 3.874 ;
      RECT 53.352 3.731 53.438 3.874 ;
      RECT 53.266 3.732 53.352 3.875 ;
      RECT 53.18 3.732 53.266 3.875 ;
      RECT 53.16 3.732 53.18 3.875 ;
      RECT 53.074 3.732 53.16 3.875 ;
      RECT 52.988 3.732 53.074 3.875 ;
      RECT 52.902 3.733 52.988 3.875 ;
      RECT 52.816 3.733 52.902 3.875 ;
      RECT 52.73 3.733 52.816 3.875 ;
      RECT 52.644 3.734 52.73 3.875 ;
      RECT 52.558 3.734 52.644 3.875 ;
      RECT 52.472 3.734 52.558 3.875 ;
      RECT 52.386 3.734 52.472 3.875 ;
      RECT 52.3 3.735 52.386 3.875 ;
      RECT 52.25 3.732 52.3 3.875 ;
      RECT 52.24 3.73 52.25 3.874 ;
      RECT 52.236 3.73 52.24 3.873 ;
      RECT 52.15 3.725 52.236 3.868 ;
      RECT 52.128 3.718 52.15 3.862 ;
      RECT 52.042 3.709 52.128 3.856 ;
      RECT 51.956 3.696 52.042 3.847 ;
      RECT 51.87 3.682 51.956 3.837 ;
      RECT 51.825 3.672 51.87 3.83 ;
      RECT 51.805 2.96 51.825 3.238 ;
      RECT 51.805 3.665 51.825 3.826 ;
      RECT 51.775 2.96 51.805 3.26 ;
      RECT 51.765 3.632 51.805 3.823 ;
      RECT 51.76 2.96 51.775 3.28 ;
      RECT 51.76 3.597 51.765 3.821 ;
      RECT 51.755 2.96 51.76 3.405 ;
      RECT 51.755 3.557 51.76 3.821 ;
      RECT 51.745 2.96 51.755 3.821 ;
      RECT 51.67 2.96 51.745 3.815 ;
      RECT 51.64 2.96 51.67 3.805 ;
      RECT 51.635 2.96 51.64 3.797 ;
      RECT 51.63 3.002 51.635 3.79 ;
      RECT 51.62 3.071 51.63 3.781 ;
      RECT 51.615 3.141 51.62 3.733 ;
      RECT 51.61 3.205 51.615 3.63 ;
      RECT 51.605 3.24 51.61 3.585 ;
      RECT 51.603 3.277 51.605 3.477 ;
      RECT 51.6 3.285 51.603 3.47 ;
      RECT 51.595 3.35 51.6 3.413 ;
      RECT 55.67 2.44 55.95 2.72 ;
      RECT 55.66 2.44 55.95 2.583 ;
      RECT 55.615 2.305 55.875 2.565 ;
      RECT 55.615 2.42 55.93 2.565 ;
      RECT 55.615 2.39 55.925 2.565 ;
      RECT 55.615 2.377 55.915 2.565 ;
      RECT 55.615 2.367 55.91 2.565 ;
      RECT 51.59 2.35 51.85 2.61 ;
      RECT 55.36 1.9 55.62 2.16 ;
      RECT 55.35 1.925 55.62 2.12 ;
      RECT 55.345 1.925 55.35 2.119 ;
      RECT 55.275 1.92 55.345 2.111 ;
      RECT 55.19 1.907 55.275 2.094 ;
      RECT 55.186 1.899 55.19 2.084 ;
      RECT 55.1 1.892 55.186 2.074 ;
      RECT 55.091 1.884 55.1 2.064 ;
      RECT 55.005 1.877 55.091 2.052 ;
      RECT 54.985 1.868 55.005 2.038 ;
      RECT 54.93 1.863 54.985 2.03 ;
      RECT 54.92 1.857 54.93 2.024 ;
      RECT 54.9 1.855 54.92 2.02 ;
      RECT 54.892 1.854 54.9 2.016 ;
      RECT 54.806 1.846 54.892 2.005 ;
      RECT 54.72 1.832 54.806 1.985 ;
      RECT 54.66 1.82 54.72 1.97 ;
      RECT 54.65 1.815 54.66 1.965 ;
      RECT 54.6 1.815 54.65 1.967 ;
      RECT 54.553 1.817 54.6 1.971 ;
      RECT 54.467 1.824 54.553 1.976 ;
      RECT 54.381 1.832 54.467 1.982 ;
      RECT 54.295 1.841 54.381 1.988 ;
      RECT 54.236 1.847 54.295 1.993 ;
      RECT 54.15 1.852 54.236 1.999 ;
      RECT 54.075 1.857 54.15 2.005 ;
      RECT 54.036 1.859 54.075 2.01 ;
      RECT 53.95 1.856 54.036 2.015 ;
      RECT 53.865 1.854 53.95 2.022 ;
      RECT 53.833 1.853 53.865 2.025 ;
      RECT 53.747 1.852 53.833 2.026 ;
      RECT 53.661 1.851 53.747 2.027 ;
      RECT 53.575 1.85 53.661 2.027 ;
      RECT 53.489 1.849 53.575 2.028 ;
      RECT 53.403 1.848 53.489 2.029 ;
      RECT 53.317 1.847 53.403 2.03 ;
      RECT 53.231 1.846 53.317 2.03 ;
      RECT 53.145 1.845 53.231 2.031 ;
      RECT 53.095 1.845 53.145 2.032 ;
      RECT 53.081 1.846 53.095 2.032 ;
      RECT 52.995 1.853 53.081 2.033 ;
      RECT 52.921 1.864 52.995 2.034 ;
      RECT 52.835 1.873 52.921 2.035 ;
      RECT 52.8 1.88 52.835 2.05 ;
      RECT 52.775 1.883 52.8 2.08 ;
      RECT 52.75 1.892 52.775 2.109 ;
      RECT 52.74 1.903 52.75 2.129 ;
      RECT 52.73 1.911 52.74 2.143 ;
      RECT 52.725 1.917 52.73 2.153 ;
      RECT 52.7 1.934 52.725 2.17 ;
      RECT 52.685 1.956 52.7 2.198 ;
      RECT 52.655 1.982 52.685 2.228 ;
      RECT 52.635 2.011 52.655 2.258 ;
      RECT 52.63 2.026 52.635 2.275 ;
      RECT 52.61 2.041 52.63 2.29 ;
      RECT 52.6 2.059 52.61 2.308 ;
      RECT 52.59 2.07 52.6 2.323 ;
      RECT 52.54 2.102 52.59 2.349 ;
      RECT 52.535 2.132 52.54 2.369 ;
      RECT 52.525 2.145 52.535 2.375 ;
      RECT 52.516 2.155 52.525 2.383 ;
      RECT 52.505 2.166 52.516 2.391 ;
      RECT 52.5 2.176 52.505 2.397 ;
      RECT 52.485 2.197 52.5 2.404 ;
      RECT 52.47 2.227 52.485 2.412 ;
      RECT 52.435 2.257 52.47 2.418 ;
      RECT 52.41 2.275 52.435 2.425 ;
      RECT 52.36 2.283 52.41 2.434 ;
      RECT 52.335 2.288 52.36 2.443 ;
      RECT 52.28 2.294 52.335 2.453 ;
      RECT 52.275 2.299 52.28 2.461 ;
      RECT 52.261 2.302 52.275 2.463 ;
      RECT 52.175 2.314 52.261 2.475 ;
      RECT 52.165 2.326 52.175 2.488 ;
      RECT 52.08 2.339 52.165 2.5 ;
      RECT 52.036 2.356 52.08 2.514 ;
      RECT 51.95 2.373 52.036 2.53 ;
      RECT 51.92 2.387 51.95 2.544 ;
      RECT 51.91 2.392 51.92 2.549 ;
      RECT 51.85 2.395 51.91 2.558 ;
      RECT 54.74 2.665 55 2.925 ;
      RECT 54.74 2.665 55.02 2.778 ;
      RECT 54.74 2.665 55.045 2.745 ;
      RECT 54.74 2.665 55.05 2.725 ;
      RECT 54.79 2.44 55.07 2.72 ;
      RECT 54.345 3.175 54.605 3.435 ;
      RECT 54.335 3.032 54.53 3.373 ;
      RECT 54.33 3.14 54.545 3.365 ;
      RECT 54.325 3.19 54.605 3.355 ;
      RECT 54.315 3.267 54.605 3.34 ;
      RECT 54.335 3.115 54.545 3.373 ;
      RECT 54.345 2.99 54.53 3.435 ;
      RECT 54.345 2.885 54.51 3.435 ;
      RECT 54.355 2.872 54.51 3.435 ;
      RECT 54.355 2.83 54.5 3.435 ;
      RECT 54.36 2.755 54.5 3.435 ;
      RECT 54.39 2.405 54.5 3.435 ;
      RECT 54.395 2.135 54.52 2.758 ;
      RECT 54.365 2.71 54.52 2.758 ;
      RECT 54.38 2.512 54.5 3.435 ;
      RECT 54.37 2.622 54.52 2.758 ;
      RECT 54.395 2.135 54.535 2.615 ;
      RECT 54.395 2.135 54.555 2.49 ;
      RECT 54.36 2.135 54.62 2.395 ;
      RECT 53.83 2.44 54.11 2.72 ;
      RECT 53.815 2.44 54.11 2.7 ;
      RECT 51.87 3.305 52.13 3.565 ;
      RECT 53.655 3.16 53.915 3.42 ;
      RECT 53.635 3.18 53.915 3.395 ;
      RECT 53.592 3.18 53.635 3.394 ;
      RECT 53.506 3.181 53.592 3.391 ;
      RECT 53.42 3.182 53.506 3.387 ;
      RECT 53.345 3.184 53.42 3.384 ;
      RECT 53.322 3.185 53.345 3.382 ;
      RECT 53.236 3.186 53.322 3.38 ;
      RECT 53.15 3.187 53.236 3.377 ;
      RECT 53.126 3.188 53.15 3.375 ;
      RECT 53.04 3.19 53.126 3.372 ;
      RECT 52.955 3.192 53.04 3.373 ;
      RECT 52.898 3.193 52.955 3.379 ;
      RECT 52.812 3.195 52.898 3.389 ;
      RECT 52.726 3.198 52.812 3.402 ;
      RECT 52.64 3.2 52.726 3.414 ;
      RECT 52.626 3.201 52.64 3.421 ;
      RECT 52.54 3.202 52.626 3.429 ;
      RECT 52.5 3.204 52.54 3.438 ;
      RECT 52.491 3.205 52.5 3.441 ;
      RECT 52.405 3.213 52.491 3.447 ;
      RECT 52.385 3.222 52.405 3.455 ;
      RECT 52.3 3.237 52.385 3.463 ;
      RECT 52.24 3.26 52.3 3.474 ;
      RECT 52.23 3.272 52.24 3.479 ;
      RECT 52.19 3.282 52.23 3.483 ;
      RECT 52.135 3.299 52.19 3.491 ;
      RECT 52.13 3.309 52.135 3.495 ;
      RECT 53.196 2.44 53.255 2.837 ;
      RECT 53.11 2.44 53.315 2.828 ;
      RECT 53.105 2.47 53.315 2.823 ;
      RECT 53.071 2.47 53.315 2.821 ;
      RECT 52.985 2.47 53.315 2.815 ;
      RECT 52.94 2.47 53.335 2.793 ;
      RECT 52.94 2.47 53.355 2.748 ;
      RECT 52.9 2.47 53.355 2.738 ;
      RECT 53.11 2.44 53.39 2.72 ;
      RECT 52.845 2.44 53.105 2.7 ;
      RECT 50.67 3 50.95 3.28 ;
      RECT 50.64 2.962 50.895 3.265 ;
      RECT 50.635 2.963 50.895 3.263 ;
      RECT 50.63 2.964 50.895 3.257 ;
      RECT 50.625 2.967 50.895 3.25 ;
      RECT 50.62 3 50.95 3.243 ;
      RECT 50.59 2.97 50.895 3.23 ;
      RECT 50.59 2.997 50.915 3.23 ;
      RECT 50.59 2.987 50.91 3.23 ;
      RECT 50.59 2.972 50.905 3.23 ;
      RECT 50.67 2.959 50.885 3.28 ;
      RECT 50.756 2.957 50.885 3.28 ;
      RECT 50.842 2.955 50.87 3.28 ;
      RECT 46.475 6.22 46.795 6.545 ;
      RECT 46.505 5.695 46.675 6.545 ;
      RECT 46.505 5.695 46.68 6.045 ;
      RECT 46.505 5.695 47.48 5.87 ;
      RECT 47.305 1.965 47.48 5.87 ;
      RECT 47.25 1.965 47.6 2.315 ;
      RECT 47.275 6.655 47.6 6.98 ;
      RECT 46.16 6.745 47.6 6.915 ;
      RECT 46.16 2.395 46.32 6.915 ;
      RECT 46.475 2.365 46.795 2.685 ;
      RECT 46.16 2.395 46.795 2.565 ;
      RECT 45.425 5.855 45.775 6.205 ;
      RECT 45.495 2.705 45.67 6.205 ;
      RECT 45.42 2.705 45.77 3.055 ;
      RECT 36.245 1.92 36.505 2.18 ;
      RECT 36.3 1.88 36.605 2.16 ;
      RECT 36.3 1.42 36.475 2.18 ;
      RECT 44.815 1.34 45.165 1.69 ;
      RECT 36.3 1.42 45.165 1.595 ;
      RECT 44.49 2.85 44.86 3.22 ;
      RECT 44.575 2.235 44.745 3.22 ;
      RECT 40.595 2.455 40.83 2.715 ;
      RECT 43.74 2.235 43.905 2.495 ;
      RECT 43.645 2.225 43.66 2.495 ;
      RECT 43.74 2.235 44.745 2.415 ;
      RECT 42.245 1.795 42.285 1.935 ;
      RECT 43.66 2.23 43.74 2.495 ;
      RECT 43.605 2.225 43.645 2.461 ;
      RECT 43.591 2.225 43.605 2.461 ;
      RECT 43.505 2.23 43.591 2.463 ;
      RECT 43.46 2.237 43.505 2.465 ;
      RECT 43.43 2.237 43.46 2.467 ;
      RECT 43.405 2.232 43.43 2.469 ;
      RECT 43.375 2.228 43.405 2.478 ;
      RECT 43.365 2.225 43.375 2.49 ;
      RECT 43.36 2.225 43.365 2.498 ;
      RECT 43.355 2.225 43.36 2.503 ;
      RECT 43.345 2.224 43.355 2.513 ;
      RECT 43.34 2.223 43.345 2.523 ;
      RECT 43.325 2.222 43.34 2.528 ;
      RECT 43.297 2.219 43.325 2.555 ;
      RECT 43.211 2.211 43.297 2.555 ;
      RECT 43.125 2.2 43.211 2.555 ;
      RECT 43.085 2.185 43.125 2.555 ;
      RECT 43.045 2.159 43.085 2.555 ;
      RECT 43.04 2.141 43.045 2.367 ;
      RECT 43.03 2.137 43.04 2.357 ;
      RECT 43.015 2.127 43.03 2.344 ;
      RECT 42.995 2.111 43.015 2.329 ;
      RECT 42.98 2.096 42.995 2.314 ;
      RECT 42.97 2.085 42.98 2.304 ;
      RECT 42.945 2.069 42.97 2.293 ;
      RECT 42.94 2.056 42.945 2.283 ;
      RECT 42.935 2.052 42.94 2.278 ;
      RECT 42.88 2.038 42.935 2.256 ;
      RECT 42.841 2.019 42.88 2.22 ;
      RECT 42.755 1.993 42.841 2.173 ;
      RECT 42.751 1.975 42.755 2.139 ;
      RECT 42.665 1.956 42.751 2.117 ;
      RECT 42.66 1.938 42.665 2.095 ;
      RECT 42.655 1.936 42.66 2.093 ;
      RECT 42.645 1.935 42.655 2.088 ;
      RECT 42.585 1.922 42.645 2.074 ;
      RECT 42.54 1.9 42.585 2.053 ;
      RECT 42.48 1.877 42.54 2.032 ;
      RECT 42.416 1.852 42.48 2.007 ;
      RECT 42.33 1.822 42.416 1.976 ;
      RECT 42.315 1.802 42.33 1.955 ;
      RECT 42.285 1.797 42.315 1.946 ;
      RECT 42.232 1.795 42.245 1.935 ;
      RECT 42.146 1.795 42.232 1.937 ;
      RECT 42.06 1.795 42.146 1.939 ;
      RECT 42.04 1.795 42.06 1.943 ;
      RECT 41.995 1.797 42.04 1.954 ;
      RECT 41.955 1.807 41.995 1.97 ;
      RECT 41.951 1.816 41.955 1.978 ;
      RECT 41.865 1.836 41.951 1.994 ;
      RECT 41.855 1.855 41.865 2.012 ;
      RECT 41.85 1.857 41.855 2.015 ;
      RECT 41.84 1.861 41.85 2.018 ;
      RECT 41.82 1.866 41.84 2.028 ;
      RECT 41.79 1.876 41.82 2.048 ;
      RECT 41.785 1.883 41.79 2.062 ;
      RECT 41.775 1.887 41.785 2.069 ;
      RECT 41.76 1.895 41.775 2.08 ;
      RECT 41.75 1.905 41.76 2.091 ;
      RECT 41.74 1.912 41.75 2.099 ;
      RECT 41.715 1.925 41.74 2.114 ;
      RECT 41.651 1.961 41.715 2.153 ;
      RECT 41.565 2.024 41.651 2.217 ;
      RECT 41.53 2.075 41.565 2.27 ;
      RECT 41.525 2.092 41.53 2.287 ;
      RECT 41.51 2.101 41.525 2.294 ;
      RECT 41.49 2.116 41.51 2.308 ;
      RECT 41.485 2.127 41.49 2.318 ;
      RECT 41.465 2.14 41.485 2.328 ;
      RECT 41.46 2.15 41.465 2.338 ;
      RECT 41.445 2.155 41.46 2.347 ;
      RECT 41.435 2.165 41.445 2.358 ;
      RECT 41.405 2.182 41.435 2.375 ;
      RECT 41.395 2.2 41.405 2.393 ;
      RECT 41.38 2.211 41.395 2.404 ;
      RECT 41.34 2.235 41.38 2.42 ;
      RECT 41.305 2.269 41.34 2.437 ;
      RECT 41.275 2.292 41.305 2.449 ;
      RECT 41.26 2.302 41.275 2.458 ;
      RECT 41.22 2.312 41.26 2.469 ;
      RECT 41.2 2.323 41.22 2.481 ;
      RECT 41.195 2.327 41.2 2.488 ;
      RECT 41.18 2.331 41.195 2.493 ;
      RECT 41.17 2.336 41.18 2.498 ;
      RECT 41.165 2.339 41.17 2.501 ;
      RECT 41.135 2.345 41.165 2.508 ;
      RECT 41.1 2.355 41.135 2.522 ;
      RECT 41.04 2.37 41.1 2.542 ;
      RECT 40.985 2.39 41.04 2.566 ;
      RECT 40.956 2.405 40.985 2.584 ;
      RECT 40.87 2.425 40.956 2.609 ;
      RECT 40.865 2.44 40.87 2.629 ;
      RECT 40.855 2.443 40.865 2.63 ;
      RECT 40.83 2.45 40.855 2.715 ;
      RECT 43.525 2.943 43.805 3.28 ;
      RECT 43.525 2.953 43.81 3.238 ;
      RECT 43.525 2.962 43.815 3.135 ;
      RECT 43.525 2.977 43.82 3.003 ;
      RECT 43.525 2.805 43.785 3.28 ;
      RECT 33.88 6.66 34.23 7.01 ;
      RECT 42.705 6.615 43.055 6.965 ;
      RECT 33.88 6.69 43.055 6.89 ;
      RECT 41.245 3.685 41.255 3.875 ;
      RECT 39.505 3.56 39.785 3.84 ;
      RECT 42.55 2.5 42.555 2.985 ;
      RECT 42.445 2.5 42.505 2.76 ;
      RECT 42.77 3.47 42.775 3.545 ;
      RECT 42.76 3.337 42.77 3.58 ;
      RECT 42.75 3.172 42.76 3.601 ;
      RECT 42.745 3.042 42.75 3.617 ;
      RECT 42.735 2.932 42.745 3.633 ;
      RECT 42.73 2.831 42.735 3.65 ;
      RECT 42.725 2.813 42.73 3.66 ;
      RECT 42.72 2.795 42.725 3.67 ;
      RECT 42.71 2.77 42.72 3.685 ;
      RECT 42.705 2.75 42.71 3.7 ;
      RECT 42.685 2.5 42.705 3.725 ;
      RECT 42.67 2.5 42.685 3.758 ;
      RECT 42.64 2.5 42.67 3.78 ;
      RECT 42.62 2.5 42.64 3.794 ;
      RECT 42.6 2.5 42.62 3.31 ;
      RECT 42.615 3.377 42.62 3.799 ;
      RECT 42.61 3.407 42.615 3.801 ;
      RECT 42.605 3.42 42.61 3.804 ;
      RECT 42.6 3.43 42.605 3.808 ;
      RECT 42.595 2.5 42.6 3.228 ;
      RECT 42.595 3.44 42.6 3.81 ;
      RECT 42.59 2.5 42.595 3.205 ;
      RECT 42.58 3.462 42.595 3.81 ;
      RECT 42.575 2.5 42.59 3.15 ;
      RECT 42.57 3.487 42.58 3.81 ;
      RECT 42.57 2.5 42.575 3.095 ;
      RECT 42.56 2.5 42.57 3.043 ;
      RECT 42.565 3.5 42.57 3.811 ;
      RECT 42.56 3.512 42.565 3.812 ;
      RECT 42.555 2.5 42.56 3.003 ;
      RECT 42.555 3.525 42.56 3.813 ;
      RECT 42.54 3.54 42.555 3.814 ;
      RECT 42.545 2.5 42.55 2.965 ;
      RECT 42.54 2.5 42.545 2.93 ;
      RECT 42.535 2.5 42.54 2.905 ;
      RECT 42.53 3.567 42.54 3.816 ;
      RECT 42.525 2.5 42.535 2.863 ;
      RECT 42.525 3.585 42.53 3.817 ;
      RECT 42.52 2.5 42.525 2.823 ;
      RECT 42.52 3.592 42.525 3.818 ;
      RECT 42.515 2.5 42.52 2.795 ;
      RECT 42.51 3.61 42.52 3.819 ;
      RECT 42.505 2.5 42.515 2.775 ;
      RECT 42.5 3.63 42.51 3.821 ;
      RECT 42.49 3.647 42.5 3.822 ;
      RECT 42.455 3.67 42.49 3.825 ;
      RECT 42.4 3.688 42.455 3.831 ;
      RECT 42.314 3.696 42.4 3.84 ;
      RECT 42.228 3.707 42.314 3.851 ;
      RECT 42.142 3.717 42.228 3.862 ;
      RECT 42.056 3.727 42.142 3.874 ;
      RECT 41.97 3.737 42.056 3.885 ;
      RECT 41.95 3.743 41.97 3.891 ;
      RECT 41.87 3.745 41.95 3.895 ;
      RECT 41.865 3.744 41.87 3.9 ;
      RECT 41.857 3.743 41.865 3.9 ;
      RECT 41.771 3.739 41.857 3.898 ;
      RECT 41.685 3.731 41.771 3.895 ;
      RECT 41.599 3.722 41.685 3.891 ;
      RECT 41.513 3.714 41.599 3.888 ;
      RECT 41.427 3.706 41.513 3.884 ;
      RECT 41.341 3.697 41.427 3.881 ;
      RECT 41.255 3.689 41.341 3.877 ;
      RECT 41.2 3.682 41.245 3.875 ;
      RECT 41.115 3.675 41.2 3.873 ;
      RECT 41.041 3.667 41.115 3.869 ;
      RECT 40.955 3.659 41.041 3.866 ;
      RECT 40.952 3.655 40.955 3.864 ;
      RECT 40.866 3.651 40.952 3.863 ;
      RECT 40.78 3.643 40.866 3.86 ;
      RECT 40.695 3.638 40.78 3.857 ;
      RECT 40.609 3.635 40.695 3.854 ;
      RECT 40.523 3.633 40.609 3.851 ;
      RECT 40.437 3.63 40.523 3.848 ;
      RECT 40.351 3.627 40.437 3.845 ;
      RECT 40.265 3.624 40.351 3.842 ;
      RECT 40.189 3.622 40.265 3.839 ;
      RECT 40.103 3.619 40.189 3.836 ;
      RECT 40.017 3.616 40.103 3.834 ;
      RECT 39.931 3.614 40.017 3.831 ;
      RECT 39.845 3.611 39.931 3.828 ;
      RECT 39.785 3.602 39.845 3.826 ;
      RECT 42.295 3.22 42.37 3.48 ;
      RECT 42.275 3.2 42.28 3.48 ;
      RECT 41.595 2.985 41.7 3.28 ;
      RECT 36.04 2.96 36.11 3.22 ;
      RECT 41.935 2.835 41.94 3.206 ;
      RECT 41.925 2.89 41.93 3.206 ;
      RECT 42.23 2.06 42.29 2.32 ;
      RECT 42.285 3.215 42.295 3.48 ;
      RECT 42.28 3.205 42.285 3.48 ;
      RECT 42.2 3.152 42.275 3.48 ;
      RECT 42.225 2.06 42.23 2.34 ;
      RECT 42.215 2.06 42.225 2.36 ;
      RECT 42.2 2.06 42.215 2.39 ;
      RECT 42.185 2.06 42.2 2.433 ;
      RECT 42.18 3.095 42.2 3.48 ;
      RECT 42.17 2.06 42.185 2.47 ;
      RECT 42.165 3.075 42.18 3.48 ;
      RECT 42.165 2.06 42.17 2.493 ;
      RECT 42.155 2.06 42.165 2.518 ;
      RECT 42.125 3.042 42.165 3.48 ;
      RECT 42.13 2.06 42.155 2.568 ;
      RECT 42.125 2.06 42.13 2.623 ;
      RECT 42.12 2.06 42.125 2.665 ;
      RECT 42.11 3.005 42.125 3.48 ;
      RECT 42.115 2.06 42.12 2.708 ;
      RECT 42.11 2.06 42.115 2.773 ;
      RECT 42.105 2.06 42.11 2.795 ;
      RECT 42.105 2.993 42.11 3.345 ;
      RECT 42.1 2.06 42.105 2.863 ;
      RECT 42.1 2.985 42.105 3.328 ;
      RECT 42.095 2.06 42.1 2.908 ;
      RECT 42.09 2.967 42.1 3.305 ;
      RECT 42.09 2.06 42.095 2.945 ;
      RECT 42.08 2.06 42.09 3.285 ;
      RECT 42.075 2.06 42.08 3.268 ;
      RECT 42.07 2.06 42.075 3.253 ;
      RECT 42.065 2.06 42.07 3.238 ;
      RECT 42.045 2.06 42.065 3.228 ;
      RECT 42.04 2.06 42.045 3.218 ;
      RECT 42.03 2.06 42.04 3.214 ;
      RECT 42.025 2.337 42.03 3.213 ;
      RECT 42.02 2.36 42.025 3.212 ;
      RECT 42.015 2.39 42.02 3.211 ;
      RECT 42.01 2.417 42.015 3.21 ;
      RECT 42.005 2.445 42.01 3.21 ;
      RECT 42 2.472 42.005 3.21 ;
      RECT 41.995 2.492 42 3.21 ;
      RECT 41.99 2.52 41.995 3.21 ;
      RECT 41.98 2.562 41.99 3.21 ;
      RECT 41.97 2.607 41.98 3.209 ;
      RECT 41.965 2.66 41.97 3.208 ;
      RECT 41.96 2.692 41.965 3.207 ;
      RECT 41.955 2.712 41.96 3.206 ;
      RECT 41.95 2.75 41.955 3.206 ;
      RECT 41.945 2.772 41.95 3.206 ;
      RECT 41.94 2.797 41.945 3.206 ;
      RECT 41.93 2.862 41.935 3.206 ;
      RECT 41.915 2.922 41.925 3.206 ;
      RECT 41.9 2.932 41.915 3.206 ;
      RECT 41.88 2.942 41.9 3.206 ;
      RECT 41.85 2.947 41.88 3.203 ;
      RECT 41.79 2.957 41.85 3.2 ;
      RECT 41.77 2.966 41.79 3.205 ;
      RECT 41.745 2.972 41.77 3.218 ;
      RECT 41.725 2.977 41.745 3.233 ;
      RECT 41.7 2.982 41.725 3.28 ;
      RECT 41.571 2.984 41.595 3.28 ;
      RECT 41.485 2.979 41.571 3.28 ;
      RECT 41.445 2.976 41.485 3.28 ;
      RECT 41.395 2.978 41.445 3.26 ;
      RECT 41.365 2.982 41.395 3.26 ;
      RECT 41.286 2.992 41.365 3.26 ;
      RECT 41.2 3.007 41.286 3.261 ;
      RECT 41.15 3.017 41.2 3.262 ;
      RECT 41.142 3.02 41.15 3.262 ;
      RECT 41.056 3.022 41.142 3.263 ;
      RECT 40.97 3.026 41.056 3.263 ;
      RECT 40.884 3.03 40.97 3.264 ;
      RECT 40.798 3.033 40.884 3.265 ;
      RECT 40.712 3.037 40.798 3.265 ;
      RECT 40.626 3.041 40.712 3.266 ;
      RECT 40.54 3.044 40.626 3.267 ;
      RECT 40.454 3.048 40.54 3.267 ;
      RECT 40.368 3.052 40.454 3.268 ;
      RECT 40.282 3.056 40.368 3.269 ;
      RECT 40.196 3.059 40.282 3.269 ;
      RECT 40.11 3.063 40.196 3.27 ;
      RECT 40.08 3.065 40.11 3.27 ;
      RECT 39.994 3.068 40.08 3.271 ;
      RECT 39.908 3.072 39.994 3.272 ;
      RECT 39.822 3.076 39.908 3.273 ;
      RECT 39.736 3.079 39.822 3.273 ;
      RECT 39.65 3.083 39.736 3.274 ;
      RECT 39.615 3.088 39.65 3.275 ;
      RECT 39.56 3.098 39.615 3.282 ;
      RECT 39.535 3.11 39.56 3.292 ;
      RECT 39.5 3.123 39.535 3.3 ;
      RECT 39.46 3.14 39.5 3.323 ;
      RECT 39.44 3.153 39.46 3.35 ;
      RECT 39.41 3.165 39.44 3.378 ;
      RECT 39.405 3.173 39.41 3.398 ;
      RECT 39.4 3.176 39.405 3.408 ;
      RECT 39.35 3.188 39.4 3.442 ;
      RECT 39.34 3.203 39.35 3.475 ;
      RECT 39.33 3.209 39.34 3.488 ;
      RECT 39.32 3.216 39.33 3.5 ;
      RECT 39.295 3.229 39.32 3.518 ;
      RECT 39.28 3.244 39.295 3.54 ;
      RECT 39.27 3.252 39.28 3.556 ;
      RECT 39.255 3.261 39.27 3.571 ;
      RECT 39.245 3.271 39.255 3.585 ;
      RECT 39.226 3.284 39.245 3.602 ;
      RECT 39.14 3.329 39.226 3.667 ;
      RECT 39.125 3.374 39.14 3.725 ;
      RECT 39.12 3.383 39.125 3.738 ;
      RECT 39.11 3.39 39.12 3.743 ;
      RECT 39.105 3.395 39.11 3.747 ;
      RECT 39.085 3.405 39.105 3.754 ;
      RECT 39.06 3.425 39.085 3.768 ;
      RECT 39.025 3.45 39.06 3.788 ;
      RECT 39.01 3.473 39.025 3.803 ;
      RECT 39 3.483 39.01 3.808 ;
      RECT 38.99 3.491 39 3.815 ;
      RECT 38.98 3.5 38.99 3.821 ;
      RECT 38.96 3.512 38.98 3.823 ;
      RECT 38.95 3.525 38.96 3.825 ;
      RECT 38.925 3.54 38.95 3.828 ;
      RECT 38.905 3.557 38.925 3.832 ;
      RECT 38.865 3.585 38.905 3.838 ;
      RECT 38.8 3.632 38.865 3.847 ;
      RECT 38.785 3.665 38.8 3.855 ;
      RECT 38.78 3.672 38.785 3.857 ;
      RECT 38.73 3.697 38.78 3.862 ;
      RECT 38.715 3.721 38.73 3.869 ;
      RECT 38.665 3.726 38.715 3.87 ;
      RECT 38.579 3.73 38.665 3.87 ;
      RECT 38.493 3.73 38.579 3.87 ;
      RECT 38.407 3.73 38.493 3.871 ;
      RECT 38.321 3.73 38.407 3.871 ;
      RECT 38.235 3.73 38.321 3.871 ;
      RECT 38.169 3.73 38.235 3.871 ;
      RECT 38.083 3.73 38.169 3.872 ;
      RECT 37.997 3.73 38.083 3.872 ;
      RECT 37.911 3.731 37.997 3.873 ;
      RECT 37.825 3.731 37.911 3.873 ;
      RECT 37.739 3.731 37.825 3.873 ;
      RECT 37.653 3.731 37.739 3.874 ;
      RECT 37.567 3.731 37.653 3.874 ;
      RECT 37.481 3.732 37.567 3.875 ;
      RECT 37.395 3.732 37.481 3.875 ;
      RECT 37.375 3.732 37.395 3.875 ;
      RECT 37.289 3.732 37.375 3.875 ;
      RECT 37.203 3.732 37.289 3.875 ;
      RECT 37.117 3.733 37.203 3.875 ;
      RECT 37.031 3.733 37.117 3.875 ;
      RECT 36.945 3.733 37.031 3.875 ;
      RECT 36.859 3.734 36.945 3.875 ;
      RECT 36.773 3.734 36.859 3.875 ;
      RECT 36.687 3.734 36.773 3.875 ;
      RECT 36.601 3.734 36.687 3.875 ;
      RECT 36.515 3.735 36.601 3.875 ;
      RECT 36.465 3.732 36.515 3.875 ;
      RECT 36.455 3.73 36.465 3.874 ;
      RECT 36.451 3.73 36.455 3.873 ;
      RECT 36.365 3.725 36.451 3.868 ;
      RECT 36.343 3.718 36.365 3.862 ;
      RECT 36.257 3.709 36.343 3.856 ;
      RECT 36.171 3.696 36.257 3.847 ;
      RECT 36.085 3.682 36.171 3.837 ;
      RECT 36.04 3.672 36.085 3.83 ;
      RECT 36.02 2.96 36.04 3.238 ;
      RECT 36.02 3.665 36.04 3.826 ;
      RECT 35.99 2.96 36.02 3.26 ;
      RECT 35.98 3.632 36.02 3.823 ;
      RECT 35.975 2.96 35.99 3.28 ;
      RECT 35.975 3.597 35.98 3.821 ;
      RECT 35.97 2.96 35.975 3.405 ;
      RECT 35.97 3.557 35.975 3.821 ;
      RECT 35.96 2.96 35.97 3.821 ;
      RECT 35.885 2.96 35.96 3.815 ;
      RECT 35.855 2.96 35.885 3.805 ;
      RECT 35.85 2.96 35.855 3.797 ;
      RECT 35.845 3.002 35.85 3.79 ;
      RECT 35.835 3.071 35.845 3.781 ;
      RECT 35.83 3.141 35.835 3.733 ;
      RECT 35.825 3.205 35.83 3.63 ;
      RECT 35.82 3.24 35.825 3.585 ;
      RECT 35.818 3.277 35.82 3.477 ;
      RECT 35.815 3.285 35.818 3.47 ;
      RECT 35.81 3.35 35.815 3.413 ;
      RECT 39.885 2.44 40.165 2.72 ;
      RECT 39.875 2.44 40.165 2.583 ;
      RECT 39.83 2.305 40.09 2.565 ;
      RECT 39.83 2.42 40.145 2.565 ;
      RECT 39.83 2.39 40.14 2.565 ;
      RECT 39.83 2.377 40.13 2.565 ;
      RECT 39.83 2.367 40.125 2.565 ;
      RECT 35.805 2.35 36.065 2.61 ;
      RECT 39.575 1.9 39.835 2.16 ;
      RECT 39.565 1.925 39.835 2.12 ;
      RECT 39.56 1.925 39.565 2.119 ;
      RECT 39.49 1.92 39.56 2.111 ;
      RECT 39.405 1.907 39.49 2.094 ;
      RECT 39.401 1.899 39.405 2.084 ;
      RECT 39.315 1.892 39.401 2.074 ;
      RECT 39.306 1.884 39.315 2.064 ;
      RECT 39.22 1.877 39.306 2.052 ;
      RECT 39.2 1.868 39.22 2.038 ;
      RECT 39.145 1.863 39.2 2.03 ;
      RECT 39.135 1.857 39.145 2.024 ;
      RECT 39.115 1.855 39.135 2.02 ;
      RECT 39.107 1.854 39.115 2.016 ;
      RECT 39.021 1.846 39.107 2.005 ;
      RECT 38.935 1.832 39.021 1.985 ;
      RECT 38.875 1.82 38.935 1.97 ;
      RECT 38.865 1.815 38.875 1.965 ;
      RECT 38.815 1.815 38.865 1.967 ;
      RECT 38.768 1.817 38.815 1.971 ;
      RECT 38.682 1.824 38.768 1.976 ;
      RECT 38.596 1.832 38.682 1.982 ;
      RECT 38.51 1.841 38.596 1.988 ;
      RECT 38.451 1.847 38.51 1.993 ;
      RECT 38.365 1.852 38.451 1.999 ;
      RECT 38.29 1.857 38.365 2.005 ;
      RECT 38.251 1.859 38.29 2.01 ;
      RECT 38.165 1.856 38.251 2.015 ;
      RECT 38.08 1.854 38.165 2.022 ;
      RECT 38.048 1.853 38.08 2.025 ;
      RECT 37.962 1.852 38.048 2.026 ;
      RECT 37.876 1.851 37.962 2.027 ;
      RECT 37.79 1.85 37.876 2.027 ;
      RECT 37.704 1.849 37.79 2.028 ;
      RECT 37.618 1.848 37.704 2.029 ;
      RECT 37.532 1.847 37.618 2.03 ;
      RECT 37.446 1.846 37.532 2.03 ;
      RECT 37.36 1.845 37.446 2.031 ;
      RECT 37.31 1.845 37.36 2.032 ;
      RECT 37.296 1.846 37.31 2.032 ;
      RECT 37.21 1.853 37.296 2.033 ;
      RECT 37.136 1.864 37.21 2.034 ;
      RECT 37.05 1.873 37.136 2.035 ;
      RECT 37.015 1.88 37.05 2.05 ;
      RECT 36.99 1.883 37.015 2.08 ;
      RECT 36.965 1.892 36.99 2.109 ;
      RECT 36.955 1.903 36.965 2.129 ;
      RECT 36.945 1.911 36.955 2.143 ;
      RECT 36.94 1.917 36.945 2.153 ;
      RECT 36.915 1.934 36.94 2.17 ;
      RECT 36.9 1.956 36.915 2.198 ;
      RECT 36.87 1.982 36.9 2.228 ;
      RECT 36.85 2.011 36.87 2.258 ;
      RECT 36.845 2.026 36.85 2.275 ;
      RECT 36.825 2.041 36.845 2.29 ;
      RECT 36.815 2.059 36.825 2.308 ;
      RECT 36.805 2.07 36.815 2.323 ;
      RECT 36.755 2.102 36.805 2.349 ;
      RECT 36.75 2.132 36.755 2.369 ;
      RECT 36.74 2.145 36.75 2.375 ;
      RECT 36.731 2.155 36.74 2.383 ;
      RECT 36.72 2.166 36.731 2.391 ;
      RECT 36.715 2.176 36.72 2.397 ;
      RECT 36.7 2.197 36.715 2.404 ;
      RECT 36.685 2.227 36.7 2.412 ;
      RECT 36.65 2.257 36.685 2.418 ;
      RECT 36.625 2.275 36.65 2.425 ;
      RECT 36.575 2.283 36.625 2.434 ;
      RECT 36.55 2.288 36.575 2.443 ;
      RECT 36.495 2.294 36.55 2.453 ;
      RECT 36.49 2.299 36.495 2.461 ;
      RECT 36.476 2.302 36.49 2.463 ;
      RECT 36.39 2.314 36.476 2.475 ;
      RECT 36.38 2.326 36.39 2.488 ;
      RECT 36.295 2.339 36.38 2.5 ;
      RECT 36.251 2.356 36.295 2.514 ;
      RECT 36.165 2.373 36.251 2.53 ;
      RECT 36.135 2.387 36.165 2.544 ;
      RECT 36.125 2.392 36.135 2.549 ;
      RECT 36.065 2.395 36.125 2.558 ;
      RECT 38.955 2.665 39.215 2.925 ;
      RECT 38.955 2.665 39.235 2.778 ;
      RECT 38.955 2.665 39.26 2.745 ;
      RECT 38.955 2.665 39.265 2.725 ;
      RECT 39.005 2.44 39.285 2.72 ;
      RECT 38.56 3.175 38.82 3.435 ;
      RECT 38.55 3.032 38.745 3.373 ;
      RECT 38.545 3.14 38.76 3.365 ;
      RECT 38.54 3.19 38.82 3.355 ;
      RECT 38.53 3.267 38.82 3.34 ;
      RECT 38.55 3.115 38.76 3.373 ;
      RECT 38.56 2.99 38.745 3.435 ;
      RECT 38.56 2.885 38.725 3.435 ;
      RECT 38.57 2.872 38.725 3.435 ;
      RECT 38.57 2.83 38.715 3.435 ;
      RECT 38.575 2.755 38.715 3.435 ;
      RECT 38.605 2.405 38.715 3.435 ;
      RECT 38.61 2.135 38.735 2.758 ;
      RECT 38.58 2.71 38.735 2.758 ;
      RECT 38.595 2.512 38.715 3.435 ;
      RECT 38.585 2.622 38.735 2.758 ;
      RECT 38.61 2.135 38.75 2.615 ;
      RECT 38.61 2.135 38.77 2.49 ;
      RECT 38.575 2.135 38.835 2.395 ;
      RECT 38.045 2.44 38.325 2.72 ;
      RECT 38.03 2.44 38.325 2.7 ;
      RECT 36.085 3.305 36.345 3.565 ;
      RECT 37.87 3.16 38.13 3.42 ;
      RECT 37.85 3.18 38.13 3.395 ;
      RECT 37.807 3.18 37.85 3.394 ;
      RECT 37.721 3.181 37.807 3.391 ;
      RECT 37.635 3.182 37.721 3.387 ;
      RECT 37.56 3.184 37.635 3.384 ;
      RECT 37.537 3.185 37.56 3.382 ;
      RECT 37.451 3.186 37.537 3.38 ;
      RECT 37.365 3.187 37.451 3.377 ;
      RECT 37.341 3.188 37.365 3.375 ;
      RECT 37.255 3.19 37.341 3.372 ;
      RECT 37.17 3.192 37.255 3.373 ;
      RECT 37.113 3.193 37.17 3.379 ;
      RECT 37.027 3.195 37.113 3.389 ;
      RECT 36.941 3.198 37.027 3.402 ;
      RECT 36.855 3.2 36.941 3.414 ;
      RECT 36.841 3.201 36.855 3.421 ;
      RECT 36.755 3.202 36.841 3.429 ;
      RECT 36.715 3.204 36.755 3.438 ;
      RECT 36.706 3.205 36.715 3.441 ;
      RECT 36.62 3.213 36.706 3.447 ;
      RECT 36.6 3.222 36.62 3.455 ;
      RECT 36.515 3.237 36.6 3.463 ;
      RECT 36.455 3.26 36.515 3.474 ;
      RECT 36.445 3.272 36.455 3.479 ;
      RECT 36.405 3.282 36.445 3.483 ;
      RECT 36.35 3.299 36.405 3.491 ;
      RECT 36.345 3.309 36.35 3.495 ;
      RECT 37.411 2.44 37.47 2.837 ;
      RECT 37.325 2.44 37.53 2.828 ;
      RECT 37.32 2.47 37.53 2.823 ;
      RECT 37.286 2.47 37.53 2.821 ;
      RECT 37.2 2.47 37.53 2.815 ;
      RECT 37.155 2.47 37.55 2.793 ;
      RECT 37.155 2.47 37.57 2.748 ;
      RECT 37.115 2.47 37.57 2.738 ;
      RECT 37.325 2.44 37.605 2.72 ;
      RECT 37.06 2.44 37.32 2.7 ;
      RECT 34.885 3 35.165 3.28 ;
      RECT 34.855 2.962 35.11 3.265 ;
      RECT 34.85 2.963 35.11 3.263 ;
      RECT 34.845 2.964 35.11 3.257 ;
      RECT 34.84 2.967 35.11 3.25 ;
      RECT 34.835 3 35.165 3.243 ;
      RECT 34.805 2.97 35.11 3.23 ;
      RECT 34.805 2.997 35.13 3.23 ;
      RECT 34.805 2.987 35.125 3.23 ;
      RECT 34.805 2.972 35.12 3.23 ;
      RECT 34.885 2.959 35.1 3.28 ;
      RECT 34.971 2.957 35.1 3.28 ;
      RECT 35.057 2.955 35.085 3.28 ;
      RECT 30.7 6.22 31.02 6.545 ;
      RECT 30.73 5.695 30.9 6.545 ;
      RECT 30.73 5.695 30.905 6.045 ;
      RECT 30.73 5.695 31.705 5.87 ;
      RECT 31.53 1.965 31.705 5.87 ;
      RECT 31.475 1.965 31.825 2.315 ;
      RECT 31.5 6.655 31.825 6.98 ;
      RECT 30.385 6.745 31.825 6.915 ;
      RECT 30.385 2.395 30.545 6.915 ;
      RECT 30.7 2.365 31.02 2.685 ;
      RECT 30.385 2.395 31.02 2.565 ;
      RECT 29.65 5.855 30 6.205 ;
      RECT 29.72 2.705 29.895 6.205 ;
      RECT 29.645 2.705 29.995 3.055 ;
      RECT 20.47 1.92 20.73 2.18 ;
      RECT 20.525 1.88 20.83 2.16 ;
      RECT 20.525 1.42 20.7 2.18 ;
      RECT 29.04 1.34 29.39 1.69 ;
      RECT 20.525 1.42 29.39 1.595 ;
      RECT 28.715 2.85 29.085 3.22 ;
      RECT 28.8 2.235 28.97 3.22 ;
      RECT 24.82 2.455 25.055 2.715 ;
      RECT 27.965 2.235 28.13 2.495 ;
      RECT 27.87 2.225 27.885 2.495 ;
      RECT 27.965 2.235 28.97 2.415 ;
      RECT 26.47 1.795 26.51 1.935 ;
      RECT 27.885 2.23 27.965 2.495 ;
      RECT 27.83 2.225 27.87 2.461 ;
      RECT 27.816 2.225 27.83 2.461 ;
      RECT 27.73 2.23 27.816 2.463 ;
      RECT 27.685 2.237 27.73 2.465 ;
      RECT 27.655 2.237 27.685 2.467 ;
      RECT 27.63 2.232 27.655 2.469 ;
      RECT 27.6 2.228 27.63 2.478 ;
      RECT 27.59 2.225 27.6 2.49 ;
      RECT 27.585 2.225 27.59 2.498 ;
      RECT 27.58 2.225 27.585 2.503 ;
      RECT 27.57 2.224 27.58 2.513 ;
      RECT 27.565 2.223 27.57 2.523 ;
      RECT 27.55 2.222 27.565 2.528 ;
      RECT 27.522 2.219 27.55 2.555 ;
      RECT 27.436 2.211 27.522 2.555 ;
      RECT 27.35 2.2 27.436 2.555 ;
      RECT 27.31 2.185 27.35 2.555 ;
      RECT 27.27 2.159 27.31 2.555 ;
      RECT 27.265 2.141 27.27 2.367 ;
      RECT 27.255 2.137 27.265 2.357 ;
      RECT 27.24 2.127 27.255 2.344 ;
      RECT 27.22 2.111 27.24 2.329 ;
      RECT 27.205 2.096 27.22 2.314 ;
      RECT 27.195 2.085 27.205 2.304 ;
      RECT 27.17 2.069 27.195 2.293 ;
      RECT 27.165 2.056 27.17 2.283 ;
      RECT 27.16 2.052 27.165 2.278 ;
      RECT 27.105 2.038 27.16 2.256 ;
      RECT 27.066 2.019 27.105 2.22 ;
      RECT 26.98 1.993 27.066 2.173 ;
      RECT 26.976 1.975 26.98 2.139 ;
      RECT 26.89 1.956 26.976 2.117 ;
      RECT 26.885 1.938 26.89 2.095 ;
      RECT 26.88 1.936 26.885 2.093 ;
      RECT 26.87 1.935 26.88 2.088 ;
      RECT 26.81 1.922 26.87 2.074 ;
      RECT 26.765 1.9 26.81 2.053 ;
      RECT 26.705 1.877 26.765 2.032 ;
      RECT 26.641 1.852 26.705 2.007 ;
      RECT 26.555 1.822 26.641 1.976 ;
      RECT 26.54 1.802 26.555 1.955 ;
      RECT 26.51 1.797 26.54 1.946 ;
      RECT 26.457 1.795 26.47 1.935 ;
      RECT 26.371 1.795 26.457 1.937 ;
      RECT 26.285 1.795 26.371 1.939 ;
      RECT 26.265 1.795 26.285 1.943 ;
      RECT 26.22 1.797 26.265 1.954 ;
      RECT 26.18 1.807 26.22 1.97 ;
      RECT 26.176 1.816 26.18 1.978 ;
      RECT 26.09 1.836 26.176 1.994 ;
      RECT 26.08 1.855 26.09 2.012 ;
      RECT 26.075 1.857 26.08 2.015 ;
      RECT 26.065 1.861 26.075 2.018 ;
      RECT 26.045 1.866 26.065 2.028 ;
      RECT 26.015 1.876 26.045 2.048 ;
      RECT 26.01 1.883 26.015 2.062 ;
      RECT 26 1.887 26.01 2.069 ;
      RECT 25.985 1.895 26 2.08 ;
      RECT 25.975 1.905 25.985 2.091 ;
      RECT 25.965 1.912 25.975 2.099 ;
      RECT 25.94 1.925 25.965 2.114 ;
      RECT 25.876 1.961 25.94 2.153 ;
      RECT 25.79 2.024 25.876 2.217 ;
      RECT 25.755 2.075 25.79 2.27 ;
      RECT 25.75 2.092 25.755 2.287 ;
      RECT 25.735 2.101 25.75 2.294 ;
      RECT 25.715 2.116 25.735 2.308 ;
      RECT 25.71 2.127 25.715 2.318 ;
      RECT 25.69 2.14 25.71 2.328 ;
      RECT 25.685 2.15 25.69 2.338 ;
      RECT 25.67 2.155 25.685 2.347 ;
      RECT 25.66 2.165 25.67 2.358 ;
      RECT 25.63 2.182 25.66 2.375 ;
      RECT 25.62 2.2 25.63 2.393 ;
      RECT 25.605 2.211 25.62 2.404 ;
      RECT 25.565 2.235 25.605 2.42 ;
      RECT 25.53 2.269 25.565 2.437 ;
      RECT 25.5 2.292 25.53 2.449 ;
      RECT 25.485 2.302 25.5 2.458 ;
      RECT 25.445 2.312 25.485 2.469 ;
      RECT 25.425 2.323 25.445 2.481 ;
      RECT 25.42 2.327 25.425 2.488 ;
      RECT 25.405 2.331 25.42 2.493 ;
      RECT 25.395 2.336 25.405 2.498 ;
      RECT 25.39 2.339 25.395 2.501 ;
      RECT 25.36 2.345 25.39 2.508 ;
      RECT 25.325 2.355 25.36 2.522 ;
      RECT 25.265 2.37 25.325 2.542 ;
      RECT 25.21 2.39 25.265 2.566 ;
      RECT 25.181 2.405 25.21 2.584 ;
      RECT 25.095 2.425 25.181 2.609 ;
      RECT 25.09 2.44 25.095 2.629 ;
      RECT 25.08 2.443 25.09 2.63 ;
      RECT 25.055 2.45 25.08 2.715 ;
      RECT 27.75 2.943 28.03 3.28 ;
      RECT 27.75 2.953 28.035 3.238 ;
      RECT 27.75 2.962 28.04 3.135 ;
      RECT 27.75 2.977 28.045 3.003 ;
      RECT 27.75 2.805 28.01 3.28 ;
      RECT 18.1 6.655 18.45 7.005 ;
      RECT 26.925 6.61 27.275 6.96 ;
      RECT 18.1 6.685 27.275 6.885 ;
      RECT 25.47 3.685 25.48 3.875 ;
      RECT 23.73 3.56 24.01 3.84 ;
      RECT 26.775 2.5 26.78 2.985 ;
      RECT 26.67 2.5 26.73 2.76 ;
      RECT 26.995 3.47 27 3.545 ;
      RECT 26.985 3.337 26.995 3.58 ;
      RECT 26.975 3.172 26.985 3.601 ;
      RECT 26.97 3.042 26.975 3.617 ;
      RECT 26.96 2.932 26.97 3.633 ;
      RECT 26.955 2.831 26.96 3.65 ;
      RECT 26.95 2.813 26.955 3.66 ;
      RECT 26.945 2.795 26.95 3.67 ;
      RECT 26.935 2.77 26.945 3.685 ;
      RECT 26.93 2.75 26.935 3.7 ;
      RECT 26.91 2.5 26.93 3.725 ;
      RECT 26.895 2.5 26.91 3.758 ;
      RECT 26.865 2.5 26.895 3.78 ;
      RECT 26.845 2.5 26.865 3.794 ;
      RECT 26.825 2.5 26.845 3.31 ;
      RECT 26.84 3.377 26.845 3.799 ;
      RECT 26.835 3.407 26.84 3.801 ;
      RECT 26.83 3.42 26.835 3.804 ;
      RECT 26.825 3.43 26.83 3.808 ;
      RECT 26.82 2.5 26.825 3.228 ;
      RECT 26.82 3.44 26.825 3.81 ;
      RECT 26.815 2.5 26.82 3.205 ;
      RECT 26.805 3.462 26.82 3.81 ;
      RECT 26.8 2.5 26.815 3.15 ;
      RECT 26.795 3.487 26.805 3.81 ;
      RECT 26.795 2.5 26.8 3.095 ;
      RECT 26.785 2.5 26.795 3.043 ;
      RECT 26.79 3.5 26.795 3.811 ;
      RECT 26.785 3.512 26.79 3.812 ;
      RECT 26.78 2.5 26.785 3.003 ;
      RECT 26.78 3.525 26.785 3.813 ;
      RECT 26.765 3.54 26.78 3.814 ;
      RECT 26.77 2.5 26.775 2.965 ;
      RECT 26.765 2.5 26.77 2.93 ;
      RECT 26.76 2.5 26.765 2.905 ;
      RECT 26.755 3.567 26.765 3.816 ;
      RECT 26.75 2.5 26.76 2.863 ;
      RECT 26.75 3.585 26.755 3.817 ;
      RECT 26.745 2.5 26.75 2.823 ;
      RECT 26.745 3.592 26.75 3.818 ;
      RECT 26.74 2.5 26.745 2.795 ;
      RECT 26.735 3.61 26.745 3.819 ;
      RECT 26.73 2.5 26.74 2.775 ;
      RECT 26.725 3.63 26.735 3.821 ;
      RECT 26.715 3.647 26.725 3.822 ;
      RECT 26.68 3.67 26.715 3.825 ;
      RECT 26.625 3.688 26.68 3.831 ;
      RECT 26.539 3.696 26.625 3.84 ;
      RECT 26.453 3.707 26.539 3.851 ;
      RECT 26.367 3.717 26.453 3.862 ;
      RECT 26.281 3.727 26.367 3.874 ;
      RECT 26.195 3.737 26.281 3.885 ;
      RECT 26.175 3.743 26.195 3.891 ;
      RECT 26.095 3.745 26.175 3.895 ;
      RECT 26.09 3.744 26.095 3.9 ;
      RECT 26.082 3.743 26.09 3.9 ;
      RECT 25.996 3.739 26.082 3.898 ;
      RECT 25.91 3.731 25.996 3.895 ;
      RECT 25.824 3.722 25.91 3.891 ;
      RECT 25.738 3.714 25.824 3.888 ;
      RECT 25.652 3.706 25.738 3.884 ;
      RECT 25.566 3.697 25.652 3.881 ;
      RECT 25.48 3.689 25.566 3.877 ;
      RECT 25.425 3.682 25.47 3.875 ;
      RECT 25.34 3.675 25.425 3.873 ;
      RECT 25.266 3.667 25.34 3.869 ;
      RECT 25.18 3.659 25.266 3.866 ;
      RECT 25.177 3.655 25.18 3.864 ;
      RECT 25.091 3.651 25.177 3.863 ;
      RECT 25.005 3.643 25.091 3.86 ;
      RECT 24.92 3.638 25.005 3.857 ;
      RECT 24.834 3.635 24.92 3.854 ;
      RECT 24.748 3.633 24.834 3.851 ;
      RECT 24.662 3.63 24.748 3.848 ;
      RECT 24.576 3.627 24.662 3.845 ;
      RECT 24.49 3.624 24.576 3.842 ;
      RECT 24.414 3.622 24.49 3.839 ;
      RECT 24.328 3.619 24.414 3.836 ;
      RECT 24.242 3.616 24.328 3.834 ;
      RECT 24.156 3.614 24.242 3.831 ;
      RECT 24.07 3.611 24.156 3.828 ;
      RECT 24.01 3.602 24.07 3.826 ;
      RECT 26.52 3.22 26.595 3.48 ;
      RECT 26.5 3.2 26.505 3.48 ;
      RECT 25.82 2.985 25.925 3.28 ;
      RECT 20.265 2.96 20.335 3.22 ;
      RECT 26.16 2.835 26.165 3.206 ;
      RECT 26.15 2.89 26.155 3.206 ;
      RECT 26.455 2.06 26.515 2.32 ;
      RECT 26.51 3.215 26.52 3.48 ;
      RECT 26.505 3.205 26.51 3.48 ;
      RECT 26.425 3.152 26.5 3.48 ;
      RECT 26.45 2.06 26.455 2.34 ;
      RECT 26.44 2.06 26.45 2.36 ;
      RECT 26.425 2.06 26.44 2.39 ;
      RECT 26.41 2.06 26.425 2.433 ;
      RECT 26.405 3.095 26.425 3.48 ;
      RECT 26.395 2.06 26.41 2.47 ;
      RECT 26.39 3.075 26.405 3.48 ;
      RECT 26.39 2.06 26.395 2.493 ;
      RECT 26.38 2.06 26.39 2.518 ;
      RECT 26.35 3.042 26.39 3.48 ;
      RECT 26.355 2.06 26.38 2.568 ;
      RECT 26.35 2.06 26.355 2.623 ;
      RECT 26.345 2.06 26.35 2.665 ;
      RECT 26.335 3.005 26.35 3.48 ;
      RECT 26.34 2.06 26.345 2.708 ;
      RECT 26.335 2.06 26.34 2.773 ;
      RECT 26.33 2.06 26.335 2.795 ;
      RECT 26.33 2.993 26.335 3.345 ;
      RECT 26.325 2.06 26.33 2.863 ;
      RECT 26.325 2.985 26.33 3.328 ;
      RECT 26.32 2.06 26.325 2.908 ;
      RECT 26.315 2.967 26.325 3.305 ;
      RECT 26.315 2.06 26.32 2.945 ;
      RECT 26.305 2.06 26.315 3.285 ;
      RECT 26.3 2.06 26.305 3.268 ;
      RECT 26.295 2.06 26.3 3.253 ;
      RECT 26.29 2.06 26.295 3.238 ;
      RECT 26.27 2.06 26.29 3.228 ;
      RECT 26.265 2.06 26.27 3.218 ;
      RECT 26.255 2.06 26.265 3.214 ;
      RECT 26.25 2.337 26.255 3.213 ;
      RECT 26.245 2.36 26.25 3.212 ;
      RECT 26.24 2.39 26.245 3.211 ;
      RECT 26.235 2.417 26.24 3.21 ;
      RECT 26.23 2.445 26.235 3.21 ;
      RECT 26.225 2.472 26.23 3.21 ;
      RECT 26.22 2.492 26.225 3.21 ;
      RECT 26.215 2.52 26.22 3.21 ;
      RECT 26.205 2.562 26.215 3.21 ;
      RECT 26.195 2.607 26.205 3.209 ;
      RECT 26.19 2.66 26.195 3.208 ;
      RECT 26.185 2.692 26.19 3.207 ;
      RECT 26.18 2.712 26.185 3.206 ;
      RECT 26.175 2.75 26.18 3.206 ;
      RECT 26.17 2.772 26.175 3.206 ;
      RECT 26.165 2.797 26.17 3.206 ;
      RECT 26.155 2.862 26.16 3.206 ;
      RECT 26.14 2.922 26.15 3.206 ;
      RECT 26.125 2.932 26.14 3.206 ;
      RECT 26.105 2.942 26.125 3.206 ;
      RECT 26.075 2.947 26.105 3.203 ;
      RECT 26.015 2.957 26.075 3.2 ;
      RECT 25.995 2.966 26.015 3.205 ;
      RECT 25.97 2.972 25.995 3.218 ;
      RECT 25.95 2.977 25.97 3.233 ;
      RECT 25.925 2.982 25.95 3.28 ;
      RECT 25.796 2.984 25.82 3.28 ;
      RECT 25.71 2.979 25.796 3.28 ;
      RECT 25.67 2.976 25.71 3.28 ;
      RECT 25.62 2.978 25.67 3.26 ;
      RECT 25.59 2.982 25.62 3.26 ;
      RECT 25.511 2.992 25.59 3.26 ;
      RECT 25.425 3.007 25.511 3.261 ;
      RECT 25.375 3.017 25.425 3.262 ;
      RECT 25.367 3.02 25.375 3.262 ;
      RECT 25.281 3.022 25.367 3.263 ;
      RECT 25.195 3.026 25.281 3.263 ;
      RECT 25.109 3.03 25.195 3.264 ;
      RECT 25.023 3.033 25.109 3.265 ;
      RECT 24.937 3.037 25.023 3.265 ;
      RECT 24.851 3.041 24.937 3.266 ;
      RECT 24.765 3.044 24.851 3.267 ;
      RECT 24.679 3.048 24.765 3.267 ;
      RECT 24.593 3.052 24.679 3.268 ;
      RECT 24.507 3.056 24.593 3.269 ;
      RECT 24.421 3.059 24.507 3.269 ;
      RECT 24.335 3.063 24.421 3.27 ;
      RECT 24.305 3.065 24.335 3.27 ;
      RECT 24.219 3.068 24.305 3.271 ;
      RECT 24.133 3.072 24.219 3.272 ;
      RECT 24.047 3.076 24.133 3.273 ;
      RECT 23.961 3.079 24.047 3.273 ;
      RECT 23.875 3.083 23.961 3.274 ;
      RECT 23.84 3.088 23.875 3.275 ;
      RECT 23.785 3.098 23.84 3.282 ;
      RECT 23.76 3.11 23.785 3.292 ;
      RECT 23.725 3.123 23.76 3.3 ;
      RECT 23.685 3.14 23.725 3.323 ;
      RECT 23.665 3.153 23.685 3.35 ;
      RECT 23.635 3.165 23.665 3.378 ;
      RECT 23.63 3.173 23.635 3.398 ;
      RECT 23.625 3.176 23.63 3.408 ;
      RECT 23.575 3.188 23.625 3.442 ;
      RECT 23.565 3.203 23.575 3.475 ;
      RECT 23.555 3.209 23.565 3.488 ;
      RECT 23.545 3.216 23.555 3.5 ;
      RECT 23.52 3.229 23.545 3.518 ;
      RECT 23.505 3.244 23.52 3.54 ;
      RECT 23.495 3.252 23.505 3.556 ;
      RECT 23.48 3.261 23.495 3.571 ;
      RECT 23.47 3.271 23.48 3.585 ;
      RECT 23.451 3.284 23.47 3.602 ;
      RECT 23.365 3.329 23.451 3.667 ;
      RECT 23.35 3.374 23.365 3.725 ;
      RECT 23.345 3.383 23.35 3.738 ;
      RECT 23.335 3.39 23.345 3.743 ;
      RECT 23.33 3.395 23.335 3.747 ;
      RECT 23.31 3.405 23.33 3.754 ;
      RECT 23.285 3.425 23.31 3.768 ;
      RECT 23.25 3.45 23.285 3.788 ;
      RECT 23.235 3.473 23.25 3.803 ;
      RECT 23.225 3.483 23.235 3.808 ;
      RECT 23.215 3.491 23.225 3.815 ;
      RECT 23.205 3.5 23.215 3.821 ;
      RECT 23.185 3.512 23.205 3.823 ;
      RECT 23.175 3.525 23.185 3.825 ;
      RECT 23.15 3.54 23.175 3.828 ;
      RECT 23.13 3.557 23.15 3.832 ;
      RECT 23.09 3.585 23.13 3.838 ;
      RECT 23.025 3.632 23.09 3.847 ;
      RECT 23.01 3.665 23.025 3.855 ;
      RECT 23.005 3.672 23.01 3.857 ;
      RECT 22.955 3.697 23.005 3.862 ;
      RECT 22.94 3.721 22.955 3.869 ;
      RECT 22.89 3.726 22.94 3.87 ;
      RECT 22.804 3.73 22.89 3.87 ;
      RECT 22.718 3.73 22.804 3.87 ;
      RECT 22.632 3.73 22.718 3.871 ;
      RECT 22.546 3.73 22.632 3.871 ;
      RECT 22.46 3.73 22.546 3.871 ;
      RECT 22.394 3.73 22.46 3.871 ;
      RECT 22.308 3.73 22.394 3.872 ;
      RECT 22.222 3.73 22.308 3.872 ;
      RECT 22.136 3.731 22.222 3.873 ;
      RECT 22.05 3.731 22.136 3.873 ;
      RECT 21.964 3.731 22.05 3.873 ;
      RECT 21.878 3.731 21.964 3.874 ;
      RECT 21.792 3.731 21.878 3.874 ;
      RECT 21.706 3.732 21.792 3.875 ;
      RECT 21.62 3.732 21.706 3.875 ;
      RECT 21.6 3.732 21.62 3.875 ;
      RECT 21.514 3.732 21.6 3.875 ;
      RECT 21.428 3.732 21.514 3.875 ;
      RECT 21.342 3.733 21.428 3.875 ;
      RECT 21.256 3.733 21.342 3.875 ;
      RECT 21.17 3.733 21.256 3.875 ;
      RECT 21.084 3.734 21.17 3.875 ;
      RECT 20.998 3.734 21.084 3.875 ;
      RECT 20.912 3.734 20.998 3.875 ;
      RECT 20.826 3.734 20.912 3.875 ;
      RECT 20.74 3.735 20.826 3.875 ;
      RECT 20.69 3.732 20.74 3.875 ;
      RECT 20.68 3.73 20.69 3.874 ;
      RECT 20.676 3.73 20.68 3.873 ;
      RECT 20.59 3.725 20.676 3.868 ;
      RECT 20.568 3.718 20.59 3.862 ;
      RECT 20.482 3.709 20.568 3.856 ;
      RECT 20.396 3.696 20.482 3.847 ;
      RECT 20.31 3.682 20.396 3.837 ;
      RECT 20.265 3.672 20.31 3.83 ;
      RECT 20.245 2.96 20.265 3.238 ;
      RECT 20.245 3.665 20.265 3.826 ;
      RECT 20.215 2.96 20.245 3.26 ;
      RECT 20.205 3.632 20.245 3.823 ;
      RECT 20.2 2.96 20.215 3.28 ;
      RECT 20.2 3.597 20.205 3.821 ;
      RECT 20.195 2.96 20.2 3.405 ;
      RECT 20.195 3.557 20.2 3.821 ;
      RECT 20.185 2.96 20.195 3.821 ;
      RECT 20.11 2.96 20.185 3.815 ;
      RECT 20.08 2.96 20.11 3.805 ;
      RECT 20.075 2.96 20.08 3.797 ;
      RECT 20.07 3.002 20.075 3.79 ;
      RECT 20.06 3.071 20.07 3.781 ;
      RECT 20.055 3.141 20.06 3.733 ;
      RECT 20.05 3.205 20.055 3.63 ;
      RECT 20.045 3.24 20.05 3.585 ;
      RECT 20.043 3.277 20.045 3.477 ;
      RECT 20.04 3.285 20.043 3.47 ;
      RECT 20.035 3.35 20.04 3.413 ;
      RECT 24.11 2.44 24.39 2.72 ;
      RECT 24.1 2.44 24.39 2.583 ;
      RECT 24.055 2.305 24.315 2.565 ;
      RECT 24.055 2.42 24.37 2.565 ;
      RECT 24.055 2.39 24.365 2.565 ;
      RECT 24.055 2.377 24.355 2.565 ;
      RECT 24.055 2.367 24.35 2.565 ;
      RECT 20.03 2.35 20.29 2.61 ;
      RECT 23.8 1.9 24.06 2.16 ;
      RECT 23.79 1.925 24.06 2.12 ;
      RECT 23.785 1.925 23.79 2.119 ;
      RECT 23.715 1.92 23.785 2.111 ;
      RECT 23.63 1.907 23.715 2.094 ;
      RECT 23.626 1.899 23.63 2.084 ;
      RECT 23.54 1.892 23.626 2.074 ;
      RECT 23.531 1.884 23.54 2.064 ;
      RECT 23.445 1.877 23.531 2.052 ;
      RECT 23.425 1.868 23.445 2.038 ;
      RECT 23.37 1.863 23.425 2.03 ;
      RECT 23.36 1.857 23.37 2.024 ;
      RECT 23.34 1.855 23.36 2.02 ;
      RECT 23.332 1.854 23.34 2.016 ;
      RECT 23.246 1.846 23.332 2.005 ;
      RECT 23.16 1.832 23.246 1.985 ;
      RECT 23.1 1.82 23.16 1.97 ;
      RECT 23.09 1.815 23.1 1.965 ;
      RECT 23.04 1.815 23.09 1.967 ;
      RECT 22.993 1.817 23.04 1.971 ;
      RECT 22.907 1.824 22.993 1.976 ;
      RECT 22.821 1.832 22.907 1.982 ;
      RECT 22.735 1.841 22.821 1.988 ;
      RECT 22.676 1.847 22.735 1.993 ;
      RECT 22.59 1.852 22.676 1.999 ;
      RECT 22.515 1.857 22.59 2.005 ;
      RECT 22.476 1.859 22.515 2.01 ;
      RECT 22.39 1.856 22.476 2.015 ;
      RECT 22.305 1.854 22.39 2.022 ;
      RECT 22.273 1.853 22.305 2.025 ;
      RECT 22.187 1.852 22.273 2.026 ;
      RECT 22.101 1.851 22.187 2.027 ;
      RECT 22.015 1.85 22.101 2.027 ;
      RECT 21.929 1.849 22.015 2.028 ;
      RECT 21.843 1.848 21.929 2.029 ;
      RECT 21.757 1.847 21.843 2.03 ;
      RECT 21.671 1.846 21.757 2.03 ;
      RECT 21.585 1.845 21.671 2.031 ;
      RECT 21.535 1.845 21.585 2.032 ;
      RECT 21.521 1.846 21.535 2.032 ;
      RECT 21.435 1.853 21.521 2.033 ;
      RECT 21.361 1.864 21.435 2.034 ;
      RECT 21.275 1.873 21.361 2.035 ;
      RECT 21.24 1.88 21.275 2.05 ;
      RECT 21.215 1.883 21.24 2.08 ;
      RECT 21.19 1.892 21.215 2.109 ;
      RECT 21.18 1.903 21.19 2.129 ;
      RECT 21.17 1.911 21.18 2.143 ;
      RECT 21.165 1.917 21.17 2.153 ;
      RECT 21.14 1.934 21.165 2.17 ;
      RECT 21.125 1.956 21.14 2.198 ;
      RECT 21.095 1.982 21.125 2.228 ;
      RECT 21.075 2.011 21.095 2.258 ;
      RECT 21.07 2.026 21.075 2.275 ;
      RECT 21.05 2.041 21.07 2.29 ;
      RECT 21.04 2.059 21.05 2.308 ;
      RECT 21.03 2.07 21.04 2.323 ;
      RECT 20.98 2.102 21.03 2.349 ;
      RECT 20.975 2.132 20.98 2.369 ;
      RECT 20.965 2.145 20.975 2.375 ;
      RECT 20.956 2.155 20.965 2.383 ;
      RECT 20.945 2.166 20.956 2.391 ;
      RECT 20.94 2.176 20.945 2.397 ;
      RECT 20.925 2.197 20.94 2.404 ;
      RECT 20.91 2.227 20.925 2.412 ;
      RECT 20.875 2.257 20.91 2.418 ;
      RECT 20.85 2.275 20.875 2.425 ;
      RECT 20.8 2.283 20.85 2.434 ;
      RECT 20.775 2.288 20.8 2.443 ;
      RECT 20.72 2.294 20.775 2.453 ;
      RECT 20.715 2.299 20.72 2.461 ;
      RECT 20.701 2.302 20.715 2.463 ;
      RECT 20.615 2.314 20.701 2.475 ;
      RECT 20.605 2.326 20.615 2.488 ;
      RECT 20.52 2.339 20.605 2.5 ;
      RECT 20.476 2.356 20.52 2.514 ;
      RECT 20.39 2.373 20.476 2.53 ;
      RECT 20.36 2.387 20.39 2.544 ;
      RECT 20.35 2.392 20.36 2.549 ;
      RECT 20.29 2.395 20.35 2.558 ;
      RECT 23.18 2.665 23.44 2.925 ;
      RECT 23.18 2.665 23.46 2.778 ;
      RECT 23.18 2.665 23.485 2.745 ;
      RECT 23.18 2.665 23.49 2.725 ;
      RECT 23.23 2.44 23.51 2.72 ;
      RECT 22.785 3.175 23.045 3.435 ;
      RECT 22.775 3.032 22.97 3.373 ;
      RECT 22.77 3.14 22.985 3.365 ;
      RECT 22.765 3.19 23.045 3.355 ;
      RECT 22.755 3.267 23.045 3.34 ;
      RECT 22.775 3.115 22.985 3.373 ;
      RECT 22.785 2.99 22.97 3.435 ;
      RECT 22.785 2.885 22.95 3.435 ;
      RECT 22.795 2.872 22.95 3.435 ;
      RECT 22.795 2.83 22.94 3.435 ;
      RECT 22.8 2.755 22.94 3.435 ;
      RECT 22.83 2.405 22.94 3.435 ;
      RECT 22.835 2.135 22.96 2.758 ;
      RECT 22.805 2.71 22.96 2.758 ;
      RECT 22.82 2.512 22.94 3.435 ;
      RECT 22.81 2.622 22.96 2.758 ;
      RECT 22.835 2.135 22.975 2.615 ;
      RECT 22.835 2.135 22.995 2.49 ;
      RECT 22.8 2.135 23.06 2.395 ;
      RECT 22.27 2.44 22.55 2.72 ;
      RECT 22.255 2.44 22.55 2.7 ;
      RECT 20.31 3.305 20.57 3.565 ;
      RECT 22.095 3.16 22.355 3.42 ;
      RECT 22.075 3.18 22.355 3.395 ;
      RECT 22.032 3.18 22.075 3.394 ;
      RECT 21.946 3.181 22.032 3.391 ;
      RECT 21.86 3.182 21.946 3.387 ;
      RECT 21.785 3.184 21.86 3.384 ;
      RECT 21.762 3.185 21.785 3.382 ;
      RECT 21.676 3.186 21.762 3.38 ;
      RECT 21.59 3.187 21.676 3.377 ;
      RECT 21.566 3.188 21.59 3.375 ;
      RECT 21.48 3.19 21.566 3.372 ;
      RECT 21.395 3.192 21.48 3.373 ;
      RECT 21.338 3.193 21.395 3.379 ;
      RECT 21.252 3.195 21.338 3.389 ;
      RECT 21.166 3.198 21.252 3.402 ;
      RECT 21.08 3.2 21.166 3.414 ;
      RECT 21.066 3.201 21.08 3.421 ;
      RECT 20.98 3.202 21.066 3.429 ;
      RECT 20.94 3.204 20.98 3.438 ;
      RECT 20.931 3.205 20.94 3.441 ;
      RECT 20.845 3.213 20.931 3.447 ;
      RECT 20.825 3.222 20.845 3.455 ;
      RECT 20.74 3.237 20.825 3.463 ;
      RECT 20.68 3.26 20.74 3.474 ;
      RECT 20.67 3.272 20.68 3.479 ;
      RECT 20.63 3.282 20.67 3.483 ;
      RECT 20.575 3.299 20.63 3.491 ;
      RECT 20.57 3.309 20.575 3.495 ;
      RECT 21.636 2.44 21.695 2.837 ;
      RECT 21.55 2.44 21.755 2.828 ;
      RECT 21.545 2.47 21.755 2.823 ;
      RECT 21.511 2.47 21.755 2.821 ;
      RECT 21.425 2.47 21.755 2.815 ;
      RECT 21.38 2.47 21.775 2.793 ;
      RECT 21.38 2.47 21.795 2.748 ;
      RECT 21.34 2.47 21.795 2.738 ;
      RECT 21.55 2.44 21.83 2.72 ;
      RECT 21.285 2.44 21.545 2.7 ;
      RECT 19.11 3 19.39 3.28 ;
      RECT 19.08 2.962 19.335 3.265 ;
      RECT 19.075 2.963 19.335 3.263 ;
      RECT 19.07 2.964 19.335 3.257 ;
      RECT 19.065 2.967 19.335 3.25 ;
      RECT 19.06 3 19.39 3.243 ;
      RECT 19.03 2.97 19.335 3.23 ;
      RECT 19.03 2.997 19.355 3.23 ;
      RECT 19.03 2.987 19.35 3.23 ;
      RECT 19.03 2.972 19.345 3.23 ;
      RECT 19.11 2.959 19.325 3.28 ;
      RECT 19.196 2.957 19.325 3.28 ;
      RECT 19.282 2.955 19.31 3.28 ;
      RECT 14.92 6.22 15.24 6.545 ;
      RECT 14.95 5.695 15.12 6.545 ;
      RECT 14.95 5.695 15.125 6.045 ;
      RECT 14.95 5.695 15.925 5.87 ;
      RECT 15.75 1.965 15.925 5.87 ;
      RECT 15.695 1.965 16.045 2.315 ;
      RECT 15.72 6.655 16.045 6.98 ;
      RECT 14.605 6.745 16.045 6.915 ;
      RECT 14.605 2.395 14.765 6.915 ;
      RECT 14.92 2.365 15.24 2.685 ;
      RECT 14.605 2.395 15.24 2.565 ;
      RECT 13.87 5.855 14.22 6.205 ;
      RECT 13.94 2.705 14.115 6.205 ;
      RECT 13.865 2.705 14.215 3.055 ;
      RECT 4.69 1.92 4.95 2.18 ;
      RECT 4.745 1.88 5.05 2.16 ;
      RECT 4.745 1.42 4.92 2.18 ;
      RECT 13.26 1.34 13.61 1.69 ;
      RECT 4.745 1.42 13.61 1.595 ;
      RECT 12.935 2.85 13.305 3.22 ;
      RECT 13.02 2.235 13.19 3.22 ;
      RECT 9.04 2.455 9.275 2.715 ;
      RECT 12.185 2.235 12.35 2.495 ;
      RECT 12.09 2.225 12.105 2.495 ;
      RECT 12.185 2.235 13.19 2.415 ;
      RECT 10.69 1.795 10.73 1.935 ;
      RECT 12.105 2.23 12.185 2.495 ;
      RECT 12.05 2.225 12.09 2.461 ;
      RECT 12.036 2.225 12.05 2.461 ;
      RECT 11.95 2.23 12.036 2.463 ;
      RECT 11.905 2.237 11.95 2.465 ;
      RECT 11.875 2.237 11.905 2.467 ;
      RECT 11.85 2.232 11.875 2.469 ;
      RECT 11.82 2.228 11.85 2.478 ;
      RECT 11.81 2.225 11.82 2.49 ;
      RECT 11.805 2.225 11.81 2.498 ;
      RECT 11.8 2.225 11.805 2.503 ;
      RECT 11.79 2.224 11.8 2.513 ;
      RECT 11.785 2.223 11.79 2.523 ;
      RECT 11.77 2.222 11.785 2.528 ;
      RECT 11.742 2.219 11.77 2.555 ;
      RECT 11.656 2.211 11.742 2.555 ;
      RECT 11.57 2.2 11.656 2.555 ;
      RECT 11.53 2.185 11.57 2.555 ;
      RECT 11.49 2.159 11.53 2.555 ;
      RECT 11.485 2.141 11.49 2.367 ;
      RECT 11.475 2.137 11.485 2.357 ;
      RECT 11.46 2.127 11.475 2.344 ;
      RECT 11.44 2.111 11.46 2.329 ;
      RECT 11.425 2.096 11.44 2.314 ;
      RECT 11.415 2.085 11.425 2.304 ;
      RECT 11.39 2.069 11.415 2.293 ;
      RECT 11.385 2.056 11.39 2.283 ;
      RECT 11.38 2.052 11.385 2.278 ;
      RECT 11.325 2.038 11.38 2.256 ;
      RECT 11.286 2.019 11.325 2.22 ;
      RECT 11.2 1.993 11.286 2.173 ;
      RECT 11.196 1.975 11.2 2.139 ;
      RECT 11.11 1.956 11.196 2.117 ;
      RECT 11.105 1.938 11.11 2.095 ;
      RECT 11.1 1.936 11.105 2.093 ;
      RECT 11.09 1.935 11.1 2.088 ;
      RECT 11.03 1.922 11.09 2.074 ;
      RECT 10.985 1.9 11.03 2.053 ;
      RECT 10.925 1.877 10.985 2.032 ;
      RECT 10.861 1.852 10.925 2.007 ;
      RECT 10.775 1.822 10.861 1.976 ;
      RECT 10.76 1.802 10.775 1.955 ;
      RECT 10.73 1.797 10.76 1.946 ;
      RECT 10.677 1.795 10.69 1.935 ;
      RECT 10.591 1.795 10.677 1.937 ;
      RECT 10.505 1.795 10.591 1.939 ;
      RECT 10.485 1.795 10.505 1.943 ;
      RECT 10.44 1.797 10.485 1.954 ;
      RECT 10.4 1.807 10.44 1.97 ;
      RECT 10.396 1.816 10.4 1.978 ;
      RECT 10.31 1.836 10.396 1.994 ;
      RECT 10.3 1.855 10.31 2.012 ;
      RECT 10.295 1.857 10.3 2.015 ;
      RECT 10.285 1.861 10.295 2.018 ;
      RECT 10.265 1.866 10.285 2.028 ;
      RECT 10.235 1.876 10.265 2.048 ;
      RECT 10.23 1.883 10.235 2.062 ;
      RECT 10.22 1.887 10.23 2.069 ;
      RECT 10.205 1.895 10.22 2.08 ;
      RECT 10.195 1.905 10.205 2.091 ;
      RECT 10.185 1.912 10.195 2.099 ;
      RECT 10.16 1.925 10.185 2.114 ;
      RECT 10.096 1.961 10.16 2.153 ;
      RECT 10.01 2.024 10.096 2.217 ;
      RECT 9.975 2.075 10.01 2.27 ;
      RECT 9.97 2.092 9.975 2.287 ;
      RECT 9.955 2.101 9.97 2.294 ;
      RECT 9.935 2.116 9.955 2.308 ;
      RECT 9.93 2.127 9.935 2.318 ;
      RECT 9.91 2.14 9.93 2.328 ;
      RECT 9.905 2.15 9.91 2.338 ;
      RECT 9.89 2.155 9.905 2.347 ;
      RECT 9.88 2.165 9.89 2.358 ;
      RECT 9.85 2.182 9.88 2.375 ;
      RECT 9.84 2.2 9.85 2.393 ;
      RECT 9.825 2.211 9.84 2.404 ;
      RECT 9.785 2.235 9.825 2.42 ;
      RECT 9.75 2.269 9.785 2.437 ;
      RECT 9.72 2.292 9.75 2.449 ;
      RECT 9.705 2.302 9.72 2.458 ;
      RECT 9.665 2.312 9.705 2.469 ;
      RECT 9.645 2.323 9.665 2.481 ;
      RECT 9.64 2.327 9.645 2.488 ;
      RECT 9.625 2.331 9.64 2.493 ;
      RECT 9.615 2.336 9.625 2.498 ;
      RECT 9.61 2.339 9.615 2.501 ;
      RECT 9.58 2.345 9.61 2.508 ;
      RECT 9.545 2.355 9.58 2.522 ;
      RECT 9.485 2.37 9.545 2.542 ;
      RECT 9.43 2.39 9.485 2.566 ;
      RECT 9.401 2.405 9.43 2.584 ;
      RECT 9.315 2.425 9.401 2.609 ;
      RECT 9.31 2.44 9.315 2.629 ;
      RECT 9.3 2.443 9.31 2.63 ;
      RECT 9.275 2.45 9.3 2.715 ;
      RECT 11.97 2.943 12.25 3.28 ;
      RECT 11.97 2.953 12.255 3.238 ;
      RECT 11.97 2.962 12.26 3.135 ;
      RECT 11.97 2.977 12.265 3.003 ;
      RECT 11.97 2.805 12.23 3.28 ;
      RECT 1.55 6.995 1.84 7.345 ;
      RECT 1.55 7.085 2.955 7.255 ;
      RECT 2.785 6.685 2.955 7.255 ;
      RECT 11.115 6.605 11.465 6.955 ;
      RECT 2.785 6.685 11.465 6.855 ;
      RECT 9.69 3.685 9.7 3.875 ;
      RECT 7.95 3.56 8.23 3.84 ;
      RECT 10.995 2.5 11 2.985 ;
      RECT 10.89 2.5 10.95 2.76 ;
      RECT 11.215 3.47 11.22 3.545 ;
      RECT 11.205 3.337 11.215 3.58 ;
      RECT 11.195 3.172 11.205 3.601 ;
      RECT 11.19 3.042 11.195 3.617 ;
      RECT 11.18 2.932 11.19 3.633 ;
      RECT 11.175 2.831 11.18 3.65 ;
      RECT 11.17 2.813 11.175 3.66 ;
      RECT 11.165 2.795 11.17 3.67 ;
      RECT 11.155 2.77 11.165 3.685 ;
      RECT 11.15 2.75 11.155 3.7 ;
      RECT 11.13 2.5 11.15 3.725 ;
      RECT 11.115 2.5 11.13 3.758 ;
      RECT 11.085 2.5 11.115 3.78 ;
      RECT 11.065 2.5 11.085 3.794 ;
      RECT 11.045 2.5 11.065 3.31 ;
      RECT 11.06 3.377 11.065 3.799 ;
      RECT 11.055 3.407 11.06 3.801 ;
      RECT 11.05 3.42 11.055 3.804 ;
      RECT 11.045 3.43 11.05 3.808 ;
      RECT 11.04 2.5 11.045 3.228 ;
      RECT 11.04 3.44 11.045 3.81 ;
      RECT 11.035 2.5 11.04 3.205 ;
      RECT 11.025 3.462 11.04 3.81 ;
      RECT 11.02 2.5 11.035 3.15 ;
      RECT 11.015 3.487 11.025 3.81 ;
      RECT 11.015 2.5 11.02 3.095 ;
      RECT 11.005 2.5 11.015 3.043 ;
      RECT 11.01 3.5 11.015 3.811 ;
      RECT 11.005 3.512 11.01 3.812 ;
      RECT 11 2.5 11.005 3.003 ;
      RECT 11 3.525 11.005 3.813 ;
      RECT 10.985 3.54 11 3.814 ;
      RECT 10.99 2.5 10.995 2.965 ;
      RECT 10.985 2.5 10.99 2.93 ;
      RECT 10.98 2.5 10.985 2.905 ;
      RECT 10.975 3.567 10.985 3.816 ;
      RECT 10.97 2.5 10.98 2.863 ;
      RECT 10.97 3.585 10.975 3.817 ;
      RECT 10.965 2.5 10.97 2.823 ;
      RECT 10.965 3.592 10.97 3.818 ;
      RECT 10.96 2.5 10.965 2.795 ;
      RECT 10.955 3.61 10.965 3.819 ;
      RECT 10.95 2.5 10.96 2.775 ;
      RECT 10.945 3.63 10.955 3.821 ;
      RECT 10.935 3.647 10.945 3.822 ;
      RECT 10.9 3.67 10.935 3.825 ;
      RECT 10.845 3.688 10.9 3.831 ;
      RECT 10.759 3.696 10.845 3.84 ;
      RECT 10.673 3.707 10.759 3.851 ;
      RECT 10.587 3.717 10.673 3.862 ;
      RECT 10.501 3.727 10.587 3.874 ;
      RECT 10.415 3.737 10.501 3.885 ;
      RECT 10.395 3.743 10.415 3.891 ;
      RECT 10.315 3.745 10.395 3.895 ;
      RECT 10.31 3.744 10.315 3.9 ;
      RECT 10.302 3.743 10.31 3.9 ;
      RECT 10.216 3.739 10.302 3.898 ;
      RECT 10.13 3.731 10.216 3.895 ;
      RECT 10.044 3.722 10.13 3.891 ;
      RECT 9.958 3.714 10.044 3.888 ;
      RECT 9.872 3.706 9.958 3.884 ;
      RECT 9.786 3.697 9.872 3.881 ;
      RECT 9.7 3.689 9.786 3.877 ;
      RECT 9.645 3.682 9.69 3.875 ;
      RECT 9.56 3.675 9.645 3.873 ;
      RECT 9.486 3.667 9.56 3.869 ;
      RECT 9.4 3.659 9.486 3.866 ;
      RECT 9.397 3.655 9.4 3.864 ;
      RECT 9.311 3.651 9.397 3.863 ;
      RECT 9.225 3.643 9.311 3.86 ;
      RECT 9.14 3.638 9.225 3.857 ;
      RECT 9.054 3.635 9.14 3.854 ;
      RECT 8.968 3.633 9.054 3.851 ;
      RECT 8.882 3.63 8.968 3.848 ;
      RECT 8.796 3.627 8.882 3.845 ;
      RECT 8.71 3.624 8.796 3.842 ;
      RECT 8.634 3.622 8.71 3.839 ;
      RECT 8.548 3.619 8.634 3.836 ;
      RECT 8.462 3.616 8.548 3.834 ;
      RECT 8.376 3.614 8.462 3.831 ;
      RECT 8.29 3.611 8.376 3.828 ;
      RECT 8.23 3.602 8.29 3.826 ;
      RECT 10.74 3.22 10.815 3.48 ;
      RECT 10.72 3.2 10.725 3.48 ;
      RECT 10.04 2.985 10.145 3.28 ;
      RECT 4.485 2.96 4.555 3.22 ;
      RECT 10.38 2.835 10.385 3.206 ;
      RECT 10.37 2.89 10.375 3.206 ;
      RECT 10.675 2.06 10.735 2.32 ;
      RECT 10.73 3.215 10.74 3.48 ;
      RECT 10.725 3.205 10.73 3.48 ;
      RECT 10.645 3.152 10.72 3.48 ;
      RECT 10.67 2.06 10.675 2.34 ;
      RECT 10.66 2.06 10.67 2.36 ;
      RECT 10.645 2.06 10.66 2.39 ;
      RECT 10.63 2.06 10.645 2.433 ;
      RECT 10.625 3.095 10.645 3.48 ;
      RECT 10.615 2.06 10.63 2.47 ;
      RECT 10.61 3.075 10.625 3.48 ;
      RECT 10.61 2.06 10.615 2.493 ;
      RECT 10.6 2.06 10.61 2.518 ;
      RECT 10.57 3.042 10.61 3.48 ;
      RECT 10.575 2.06 10.6 2.568 ;
      RECT 10.57 2.06 10.575 2.623 ;
      RECT 10.565 2.06 10.57 2.665 ;
      RECT 10.555 3.005 10.57 3.48 ;
      RECT 10.56 2.06 10.565 2.708 ;
      RECT 10.555 2.06 10.56 2.773 ;
      RECT 10.55 2.06 10.555 2.795 ;
      RECT 10.55 2.993 10.555 3.345 ;
      RECT 10.545 2.06 10.55 2.863 ;
      RECT 10.545 2.985 10.55 3.328 ;
      RECT 10.54 2.06 10.545 2.908 ;
      RECT 10.535 2.967 10.545 3.305 ;
      RECT 10.535 2.06 10.54 2.945 ;
      RECT 10.525 2.06 10.535 3.285 ;
      RECT 10.52 2.06 10.525 3.268 ;
      RECT 10.515 2.06 10.52 3.253 ;
      RECT 10.51 2.06 10.515 3.238 ;
      RECT 10.49 2.06 10.51 3.228 ;
      RECT 10.485 2.06 10.49 3.218 ;
      RECT 10.475 2.06 10.485 3.214 ;
      RECT 10.47 2.337 10.475 3.213 ;
      RECT 10.465 2.36 10.47 3.212 ;
      RECT 10.46 2.39 10.465 3.211 ;
      RECT 10.455 2.417 10.46 3.21 ;
      RECT 10.45 2.445 10.455 3.21 ;
      RECT 10.445 2.472 10.45 3.21 ;
      RECT 10.44 2.492 10.445 3.21 ;
      RECT 10.435 2.52 10.44 3.21 ;
      RECT 10.425 2.562 10.435 3.21 ;
      RECT 10.415 2.607 10.425 3.209 ;
      RECT 10.41 2.66 10.415 3.208 ;
      RECT 10.405 2.692 10.41 3.207 ;
      RECT 10.4 2.712 10.405 3.206 ;
      RECT 10.395 2.75 10.4 3.206 ;
      RECT 10.39 2.772 10.395 3.206 ;
      RECT 10.385 2.797 10.39 3.206 ;
      RECT 10.375 2.862 10.38 3.206 ;
      RECT 10.36 2.922 10.37 3.206 ;
      RECT 10.345 2.932 10.36 3.206 ;
      RECT 10.325 2.942 10.345 3.206 ;
      RECT 10.295 2.947 10.325 3.203 ;
      RECT 10.235 2.957 10.295 3.2 ;
      RECT 10.215 2.966 10.235 3.205 ;
      RECT 10.19 2.972 10.215 3.218 ;
      RECT 10.17 2.977 10.19 3.233 ;
      RECT 10.145 2.982 10.17 3.28 ;
      RECT 10.016 2.984 10.04 3.28 ;
      RECT 9.93 2.979 10.016 3.28 ;
      RECT 9.89 2.976 9.93 3.28 ;
      RECT 9.84 2.978 9.89 3.26 ;
      RECT 9.81 2.982 9.84 3.26 ;
      RECT 9.731 2.992 9.81 3.26 ;
      RECT 9.645 3.007 9.731 3.261 ;
      RECT 9.595 3.017 9.645 3.262 ;
      RECT 9.587 3.02 9.595 3.262 ;
      RECT 9.501 3.022 9.587 3.263 ;
      RECT 9.415 3.026 9.501 3.263 ;
      RECT 9.329 3.03 9.415 3.264 ;
      RECT 9.243 3.033 9.329 3.265 ;
      RECT 9.157 3.037 9.243 3.265 ;
      RECT 9.071 3.041 9.157 3.266 ;
      RECT 8.985 3.044 9.071 3.267 ;
      RECT 8.899 3.048 8.985 3.267 ;
      RECT 8.813 3.052 8.899 3.268 ;
      RECT 8.727 3.056 8.813 3.269 ;
      RECT 8.641 3.059 8.727 3.269 ;
      RECT 8.555 3.063 8.641 3.27 ;
      RECT 8.525 3.065 8.555 3.27 ;
      RECT 8.439 3.068 8.525 3.271 ;
      RECT 8.353 3.072 8.439 3.272 ;
      RECT 8.267 3.076 8.353 3.273 ;
      RECT 8.181 3.079 8.267 3.273 ;
      RECT 8.095 3.083 8.181 3.274 ;
      RECT 8.06 3.088 8.095 3.275 ;
      RECT 8.005 3.098 8.06 3.282 ;
      RECT 7.98 3.11 8.005 3.292 ;
      RECT 7.945 3.123 7.98 3.3 ;
      RECT 7.905 3.14 7.945 3.323 ;
      RECT 7.885 3.153 7.905 3.35 ;
      RECT 7.855 3.165 7.885 3.378 ;
      RECT 7.85 3.173 7.855 3.398 ;
      RECT 7.845 3.176 7.85 3.408 ;
      RECT 7.795 3.188 7.845 3.442 ;
      RECT 7.785 3.203 7.795 3.475 ;
      RECT 7.775 3.209 7.785 3.488 ;
      RECT 7.765 3.216 7.775 3.5 ;
      RECT 7.74 3.229 7.765 3.518 ;
      RECT 7.725 3.244 7.74 3.54 ;
      RECT 7.715 3.252 7.725 3.556 ;
      RECT 7.7 3.261 7.715 3.571 ;
      RECT 7.69 3.271 7.7 3.585 ;
      RECT 7.671 3.284 7.69 3.602 ;
      RECT 7.585 3.329 7.671 3.667 ;
      RECT 7.57 3.374 7.585 3.725 ;
      RECT 7.565 3.383 7.57 3.738 ;
      RECT 7.555 3.39 7.565 3.743 ;
      RECT 7.55 3.395 7.555 3.747 ;
      RECT 7.53 3.405 7.55 3.754 ;
      RECT 7.505 3.425 7.53 3.768 ;
      RECT 7.47 3.45 7.505 3.788 ;
      RECT 7.455 3.473 7.47 3.803 ;
      RECT 7.445 3.483 7.455 3.808 ;
      RECT 7.435 3.491 7.445 3.815 ;
      RECT 7.425 3.5 7.435 3.821 ;
      RECT 7.405 3.512 7.425 3.823 ;
      RECT 7.395 3.525 7.405 3.825 ;
      RECT 7.37 3.54 7.395 3.828 ;
      RECT 7.35 3.557 7.37 3.832 ;
      RECT 7.31 3.585 7.35 3.838 ;
      RECT 7.245 3.632 7.31 3.847 ;
      RECT 7.23 3.665 7.245 3.855 ;
      RECT 7.225 3.672 7.23 3.857 ;
      RECT 7.175 3.697 7.225 3.862 ;
      RECT 7.16 3.721 7.175 3.869 ;
      RECT 7.11 3.726 7.16 3.87 ;
      RECT 7.024 3.73 7.11 3.87 ;
      RECT 6.938 3.73 7.024 3.87 ;
      RECT 6.852 3.73 6.938 3.871 ;
      RECT 6.766 3.73 6.852 3.871 ;
      RECT 6.68 3.73 6.766 3.871 ;
      RECT 6.614 3.73 6.68 3.871 ;
      RECT 6.528 3.73 6.614 3.872 ;
      RECT 6.442 3.73 6.528 3.872 ;
      RECT 6.356 3.731 6.442 3.873 ;
      RECT 6.27 3.731 6.356 3.873 ;
      RECT 6.184 3.731 6.27 3.873 ;
      RECT 6.098 3.731 6.184 3.874 ;
      RECT 6.012 3.731 6.098 3.874 ;
      RECT 5.926 3.732 6.012 3.875 ;
      RECT 5.84 3.732 5.926 3.875 ;
      RECT 5.82 3.732 5.84 3.875 ;
      RECT 5.734 3.732 5.82 3.875 ;
      RECT 5.648 3.732 5.734 3.875 ;
      RECT 5.562 3.733 5.648 3.875 ;
      RECT 5.476 3.733 5.562 3.875 ;
      RECT 5.39 3.733 5.476 3.875 ;
      RECT 5.304 3.734 5.39 3.875 ;
      RECT 5.218 3.734 5.304 3.875 ;
      RECT 5.132 3.734 5.218 3.875 ;
      RECT 5.046 3.734 5.132 3.875 ;
      RECT 4.96 3.735 5.046 3.875 ;
      RECT 4.91 3.732 4.96 3.875 ;
      RECT 4.9 3.73 4.91 3.874 ;
      RECT 4.896 3.73 4.9 3.873 ;
      RECT 4.81 3.725 4.896 3.868 ;
      RECT 4.788 3.718 4.81 3.862 ;
      RECT 4.702 3.709 4.788 3.856 ;
      RECT 4.616 3.696 4.702 3.847 ;
      RECT 4.53 3.682 4.616 3.837 ;
      RECT 4.485 3.672 4.53 3.83 ;
      RECT 4.465 2.96 4.485 3.238 ;
      RECT 4.465 3.665 4.485 3.826 ;
      RECT 4.435 2.96 4.465 3.26 ;
      RECT 4.425 3.632 4.465 3.823 ;
      RECT 4.42 2.96 4.435 3.28 ;
      RECT 4.42 3.597 4.425 3.821 ;
      RECT 4.415 2.96 4.42 3.405 ;
      RECT 4.415 3.557 4.42 3.821 ;
      RECT 4.405 2.96 4.415 3.821 ;
      RECT 4.33 2.96 4.405 3.815 ;
      RECT 4.3 2.96 4.33 3.805 ;
      RECT 4.295 2.96 4.3 3.797 ;
      RECT 4.29 3.002 4.295 3.79 ;
      RECT 4.28 3.071 4.29 3.781 ;
      RECT 4.275 3.141 4.28 3.733 ;
      RECT 4.27 3.205 4.275 3.63 ;
      RECT 4.265 3.24 4.27 3.585 ;
      RECT 4.263 3.277 4.265 3.477 ;
      RECT 4.26 3.285 4.263 3.47 ;
      RECT 4.255 3.35 4.26 3.413 ;
      RECT 8.33 2.44 8.61 2.72 ;
      RECT 8.32 2.44 8.61 2.583 ;
      RECT 8.275 2.305 8.535 2.565 ;
      RECT 8.275 2.42 8.59 2.565 ;
      RECT 8.275 2.39 8.585 2.565 ;
      RECT 8.275 2.377 8.575 2.565 ;
      RECT 8.275 2.367 8.57 2.565 ;
      RECT 4.25 2.35 4.51 2.61 ;
      RECT 8.02 1.9 8.28 2.16 ;
      RECT 8.01 1.925 8.28 2.12 ;
      RECT 8.005 1.925 8.01 2.119 ;
      RECT 7.935 1.92 8.005 2.111 ;
      RECT 7.85 1.907 7.935 2.094 ;
      RECT 7.846 1.899 7.85 2.084 ;
      RECT 7.76 1.892 7.846 2.074 ;
      RECT 7.751 1.884 7.76 2.064 ;
      RECT 7.665 1.877 7.751 2.052 ;
      RECT 7.645 1.868 7.665 2.038 ;
      RECT 7.59 1.863 7.645 2.03 ;
      RECT 7.58 1.857 7.59 2.024 ;
      RECT 7.56 1.855 7.58 2.02 ;
      RECT 7.552 1.854 7.56 2.016 ;
      RECT 7.466 1.846 7.552 2.005 ;
      RECT 7.38 1.832 7.466 1.985 ;
      RECT 7.32 1.82 7.38 1.97 ;
      RECT 7.31 1.815 7.32 1.965 ;
      RECT 7.26 1.815 7.31 1.967 ;
      RECT 7.213 1.817 7.26 1.971 ;
      RECT 7.127 1.824 7.213 1.976 ;
      RECT 7.041 1.832 7.127 1.982 ;
      RECT 6.955 1.841 7.041 1.988 ;
      RECT 6.896 1.847 6.955 1.993 ;
      RECT 6.81 1.852 6.896 1.999 ;
      RECT 6.735 1.857 6.81 2.005 ;
      RECT 6.696 1.859 6.735 2.01 ;
      RECT 6.61 1.856 6.696 2.015 ;
      RECT 6.525 1.854 6.61 2.022 ;
      RECT 6.493 1.853 6.525 2.025 ;
      RECT 6.407 1.852 6.493 2.026 ;
      RECT 6.321 1.851 6.407 2.027 ;
      RECT 6.235 1.85 6.321 2.027 ;
      RECT 6.149 1.849 6.235 2.028 ;
      RECT 6.063 1.848 6.149 2.029 ;
      RECT 5.977 1.847 6.063 2.03 ;
      RECT 5.891 1.846 5.977 2.03 ;
      RECT 5.805 1.845 5.891 2.031 ;
      RECT 5.755 1.845 5.805 2.032 ;
      RECT 5.741 1.846 5.755 2.032 ;
      RECT 5.655 1.853 5.741 2.033 ;
      RECT 5.581 1.864 5.655 2.034 ;
      RECT 5.495 1.873 5.581 2.035 ;
      RECT 5.46 1.88 5.495 2.05 ;
      RECT 5.435 1.883 5.46 2.08 ;
      RECT 5.41 1.892 5.435 2.109 ;
      RECT 5.4 1.903 5.41 2.129 ;
      RECT 5.39 1.911 5.4 2.143 ;
      RECT 5.385 1.917 5.39 2.153 ;
      RECT 5.36 1.934 5.385 2.17 ;
      RECT 5.345 1.956 5.36 2.198 ;
      RECT 5.315 1.982 5.345 2.228 ;
      RECT 5.295 2.011 5.315 2.258 ;
      RECT 5.29 2.026 5.295 2.275 ;
      RECT 5.27 2.041 5.29 2.29 ;
      RECT 5.26 2.059 5.27 2.308 ;
      RECT 5.25 2.07 5.26 2.323 ;
      RECT 5.2 2.102 5.25 2.349 ;
      RECT 5.195 2.132 5.2 2.369 ;
      RECT 5.185 2.145 5.195 2.375 ;
      RECT 5.176 2.155 5.185 2.383 ;
      RECT 5.165 2.166 5.176 2.391 ;
      RECT 5.16 2.176 5.165 2.397 ;
      RECT 5.145 2.197 5.16 2.404 ;
      RECT 5.13 2.227 5.145 2.412 ;
      RECT 5.095 2.257 5.13 2.418 ;
      RECT 5.07 2.275 5.095 2.425 ;
      RECT 5.02 2.283 5.07 2.434 ;
      RECT 4.995 2.288 5.02 2.443 ;
      RECT 4.94 2.294 4.995 2.453 ;
      RECT 4.935 2.299 4.94 2.461 ;
      RECT 4.921 2.302 4.935 2.463 ;
      RECT 4.835 2.314 4.921 2.475 ;
      RECT 4.825 2.326 4.835 2.488 ;
      RECT 4.74 2.339 4.825 2.5 ;
      RECT 4.696 2.356 4.74 2.514 ;
      RECT 4.61 2.373 4.696 2.53 ;
      RECT 4.58 2.387 4.61 2.544 ;
      RECT 4.57 2.392 4.58 2.549 ;
      RECT 4.51 2.395 4.57 2.558 ;
      RECT 7.4 2.665 7.66 2.925 ;
      RECT 7.4 2.665 7.68 2.778 ;
      RECT 7.4 2.665 7.705 2.745 ;
      RECT 7.4 2.665 7.71 2.725 ;
      RECT 7.45 2.44 7.73 2.72 ;
      RECT 7.005 3.175 7.265 3.435 ;
      RECT 6.995 3.032 7.19 3.373 ;
      RECT 6.99 3.14 7.205 3.365 ;
      RECT 6.985 3.19 7.265 3.355 ;
      RECT 6.975 3.267 7.265 3.34 ;
      RECT 6.995 3.115 7.205 3.373 ;
      RECT 7.005 2.99 7.19 3.435 ;
      RECT 7.005 2.885 7.17 3.435 ;
      RECT 7.015 2.872 7.17 3.435 ;
      RECT 7.015 2.83 7.16 3.435 ;
      RECT 7.02 2.755 7.16 3.435 ;
      RECT 7.05 2.405 7.16 3.435 ;
      RECT 7.055 2.135 7.18 2.758 ;
      RECT 7.025 2.71 7.18 2.758 ;
      RECT 7.04 2.512 7.16 3.435 ;
      RECT 7.03 2.622 7.18 2.758 ;
      RECT 7.055 2.135 7.195 2.615 ;
      RECT 7.055 2.135 7.215 2.49 ;
      RECT 7.02 2.135 7.28 2.395 ;
      RECT 6.49 2.44 6.77 2.72 ;
      RECT 6.475 2.44 6.77 2.7 ;
      RECT 4.53 3.305 4.79 3.565 ;
      RECT 6.315 3.16 6.575 3.42 ;
      RECT 6.295 3.18 6.575 3.395 ;
      RECT 6.252 3.18 6.295 3.394 ;
      RECT 6.166 3.181 6.252 3.391 ;
      RECT 6.08 3.182 6.166 3.387 ;
      RECT 6.005 3.184 6.08 3.384 ;
      RECT 5.982 3.185 6.005 3.382 ;
      RECT 5.896 3.186 5.982 3.38 ;
      RECT 5.81 3.187 5.896 3.377 ;
      RECT 5.786 3.188 5.81 3.375 ;
      RECT 5.7 3.19 5.786 3.372 ;
      RECT 5.615 3.192 5.7 3.373 ;
      RECT 5.558 3.193 5.615 3.379 ;
      RECT 5.472 3.195 5.558 3.389 ;
      RECT 5.386 3.198 5.472 3.402 ;
      RECT 5.3 3.2 5.386 3.414 ;
      RECT 5.286 3.201 5.3 3.421 ;
      RECT 5.2 3.202 5.286 3.429 ;
      RECT 5.16 3.204 5.2 3.438 ;
      RECT 5.151 3.205 5.16 3.441 ;
      RECT 5.065 3.213 5.151 3.447 ;
      RECT 5.045 3.222 5.065 3.455 ;
      RECT 4.96 3.237 5.045 3.463 ;
      RECT 4.9 3.26 4.96 3.474 ;
      RECT 4.89 3.272 4.9 3.479 ;
      RECT 4.85 3.282 4.89 3.483 ;
      RECT 4.795 3.299 4.85 3.491 ;
      RECT 4.79 3.309 4.795 3.495 ;
      RECT 5.856 2.44 5.915 2.837 ;
      RECT 5.77 2.44 5.975 2.828 ;
      RECT 5.765 2.47 5.975 2.823 ;
      RECT 5.731 2.47 5.975 2.821 ;
      RECT 5.645 2.47 5.975 2.815 ;
      RECT 5.6 2.47 5.995 2.793 ;
      RECT 5.6 2.47 6.015 2.748 ;
      RECT 5.56 2.47 6.015 2.738 ;
      RECT 5.77 2.44 6.05 2.72 ;
      RECT 5.505 2.44 5.765 2.7 ;
      RECT 3.33 3 3.61 3.28 ;
      RECT 3.3 2.962 3.555 3.265 ;
      RECT 3.295 2.963 3.555 3.263 ;
      RECT 3.29 2.964 3.555 3.257 ;
      RECT 3.285 2.967 3.555 3.25 ;
      RECT 3.28 3 3.61 3.243 ;
      RECT 3.25 2.97 3.555 3.23 ;
      RECT 3.25 2.997 3.575 3.23 ;
      RECT 3.25 2.987 3.57 3.23 ;
      RECT 3.25 2.972 3.565 3.23 ;
      RECT 3.33 2.959 3.545 3.28 ;
      RECT 3.416 2.957 3.545 3.28 ;
      RECT 3.502 2.955 3.53 3.28 ;
      RECT 75.28 0.815 75.65 1.185 ;
      RECT 73.57 7.04 73.94 7.41 ;
      RECT 59.495 0.815 59.865 1.185 ;
      RECT 57.785 7.04 58.155 7.41 ;
      RECT 43.71 0.815 44.08 1.185 ;
      RECT 42 7.04 42.37 7.41 ;
      RECT 27.935 0.815 28.305 1.185 ;
      RECT 26.225 7.04 26.595 7.41 ;
      RECT 12.155 0.815 12.525 1.185 ;
      RECT 10.445 7.04 10.815 7.41 ;
      RECT 0.835 4.26 1.215 4.64 ;
      RECT 0.78 -0.01 1.16 0.37 ;
      RECT 0.25 8.565 0.63 8.945 ;
    LAYER via1 ;
      RECT 81.305 7.375 81.455 7.525 ;
      RECT 78.935 6.74 79.085 6.89 ;
      RECT 78.92 2.065 79.07 2.215 ;
      RECT 78.13 2.45 78.28 2.6 ;
      RECT 78.13 6.325 78.28 6.475 ;
      RECT 77.095 5.955 77.245 6.105 ;
      RECT 77.09 2.805 77.24 2.955 ;
      RECT 76.485 1.44 76.635 1.59 ;
      RECT 76.17 2.96 76.32 3.11 ;
      RECT 75.39 0.925 75.54 1.075 ;
      RECT 75.27 2.29 75.42 2.44 ;
      RECT 75.15 2.86 75.3 3.01 ;
      RECT 74.32 6.71 74.47 6.86 ;
      RECT 74.07 2.555 74.22 2.705 ;
      RECT 73.735 3.275 73.885 3.425 ;
      RECT 73.68 7.15 73.83 7.3 ;
      RECT 73.655 2.115 73.805 2.265 ;
      RECT 72.22 2.51 72.37 2.66 ;
      RECT 71.455 2.36 71.605 2.51 ;
      RECT 71.2 1.955 71.35 2.105 ;
      RECT 70.58 2.72 70.73 2.87 ;
      RECT 70.2 2.19 70.35 2.34 ;
      RECT 70.185 3.23 70.335 3.38 ;
      RECT 69.655 2.495 69.805 2.645 ;
      RECT 69.495 3.215 69.645 3.365 ;
      RECT 68.685 2.495 68.835 2.645 ;
      RECT 67.87 1.975 68.02 2.125 ;
      RECT 67.71 3.36 67.86 3.51 ;
      RECT 67.475 3.015 67.625 3.165 ;
      RECT 67.43 2.405 67.58 2.555 ;
      RECT 66.43 3.025 66.58 3.175 ;
      RECT 65.495 6.755 65.645 6.905 ;
      RECT 63.15 6.74 63.3 6.89 ;
      RECT 63.135 2.065 63.285 2.215 ;
      RECT 62.345 2.45 62.495 2.6 ;
      RECT 62.345 6.325 62.495 6.475 ;
      RECT 61.31 5.955 61.46 6.105 ;
      RECT 61.305 2.805 61.455 2.955 ;
      RECT 60.7 1.44 60.85 1.59 ;
      RECT 60.385 2.96 60.535 3.11 ;
      RECT 59.605 0.925 59.755 1.075 ;
      RECT 59.485 2.29 59.635 2.44 ;
      RECT 59.365 2.86 59.515 3.01 ;
      RECT 58.535 6.71 58.685 6.86 ;
      RECT 58.285 2.555 58.435 2.705 ;
      RECT 57.95 3.275 58.1 3.425 ;
      RECT 57.895 7.15 58.045 7.3 ;
      RECT 57.87 2.115 58.02 2.265 ;
      RECT 56.435 2.51 56.585 2.66 ;
      RECT 55.67 2.36 55.82 2.51 ;
      RECT 55.415 1.955 55.565 2.105 ;
      RECT 54.795 2.72 54.945 2.87 ;
      RECT 54.415 2.19 54.565 2.34 ;
      RECT 54.4 3.23 54.55 3.38 ;
      RECT 53.87 2.495 54.02 2.645 ;
      RECT 53.71 3.215 53.86 3.365 ;
      RECT 52.9 2.495 53.05 2.645 ;
      RECT 52.085 1.975 52.235 2.125 ;
      RECT 51.925 3.36 52.075 3.51 ;
      RECT 51.69 3.015 51.84 3.165 ;
      RECT 51.645 2.405 51.795 2.555 ;
      RECT 50.645 3.025 50.795 3.175 ;
      RECT 49.71 6.755 49.86 6.905 ;
      RECT 47.365 6.74 47.515 6.89 ;
      RECT 47.35 2.065 47.5 2.215 ;
      RECT 46.56 2.45 46.71 2.6 ;
      RECT 46.56 6.325 46.71 6.475 ;
      RECT 45.525 5.955 45.675 6.105 ;
      RECT 45.52 2.805 45.67 2.955 ;
      RECT 44.915 1.44 45.065 1.59 ;
      RECT 44.6 2.96 44.75 3.11 ;
      RECT 43.82 0.925 43.97 1.075 ;
      RECT 43.7 2.29 43.85 2.44 ;
      RECT 43.58 2.86 43.73 3.01 ;
      RECT 42.805 6.715 42.955 6.865 ;
      RECT 42.5 2.555 42.65 2.705 ;
      RECT 42.165 3.275 42.315 3.425 ;
      RECT 42.11 7.15 42.26 7.3 ;
      RECT 42.085 2.115 42.235 2.265 ;
      RECT 40.65 2.51 40.8 2.66 ;
      RECT 39.885 2.36 40.035 2.51 ;
      RECT 39.63 1.955 39.78 2.105 ;
      RECT 39.01 2.72 39.16 2.87 ;
      RECT 38.63 2.19 38.78 2.34 ;
      RECT 38.615 3.23 38.765 3.38 ;
      RECT 38.085 2.495 38.235 2.645 ;
      RECT 37.925 3.215 38.075 3.365 ;
      RECT 37.115 2.495 37.265 2.645 ;
      RECT 36.3 1.975 36.45 2.125 ;
      RECT 36.14 3.36 36.29 3.51 ;
      RECT 35.905 3.015 36.055 3.165 ;
      RECT 35.86 2.405 36.01 2.555 ;
      RECT 34.86 3.025 35.01 3.175 ;
      RECT 33.98 6.76 34.13 6.91 ;
      RECT 31.59 6.74 31.74 6.89 ;
      RECT 31.575 2.065 31.725 2.215 ;
      RECT 30.785 2.45 30.935 2.6 ;
      RECT 30.785 6.325 30.935 6.475 ;
      RECT 29.75 5.955 29.9 6.105 ;
      RECT 29.745 2.805 29.895 2.955 ;
      RECT 29.14 1.44 29.29 1.59 ;
      RECT 28.825 2.96 28.975 3.11 ;
      RECT 28.045 0.925 28.195 1.075 ;
      RECT 27.925 2.29 28.075 2.44 ;
      RECT 27.805 2.86 27.955 3.01 ;
      RECT 27.025 6.71 27.175 6.86 ;
      RECT 26.725 2.555 26.875 2.705 ;
      RECT 26.39 3.275 26.54 3.425 ;
      RECT 26.335 7.15 26.485 7.3 ;
      RECT 26.31 2.115 26.46 2.265 ;
      RECT 24.875 2.51 25.025 2.66 ;
      RECT 24.11 2.36 24.26 2.51 ;
      RECT 23.855 1.955 24.005 2.105 ;
      RECT 23.235 2.72 23.385 2.87 ;
      RECT 22.855 2.19 23.005 2.34 ;
      RECT 22.84 3.23 22.99 3.38 ;
      RECT 22.31 2.495 22.46 2.645 ;
      RECT 22.15 3.215 22.3 3.365 ;
      RECT 21.34 2.495 21.49 2.645 ;
      RECT 20.525 1.975 20.675 2.125 ;
      RECT 20.365 3.36 20.515 3.51 ;
      RECT 20.13 3.015 20.28 3.165 ;
      RECT 20.085 2.405 20.235 2.555 ;
      RECT 19.085 3.025 19.235 3.175 ;
      RECT 18.2 6.755 18.35 6.905 ;
      RECT 15.81 6.74 15.96 6.89 ;
      RECT 15.795 2.065 15.945 2.215 ;
      RECT 15.005 2.45 15.155 2.6 ;
      RECT 15.005 6.325 15.155 6.475 ;
      RECT 13.97 5.955 14.12 6.105 ;
      RECT 13.965 2.805 14.115 2.955 ;
      RECT 13.36 1.44 13.51 1.59 ;
      RECT 13.045 2.96 13.195 3.11 ;
      RECT 12.265 0.925 12.415 1.075 ;
      RECT 12.145 2.29 12.295 2.44 ;
      RECT 12.025 2.86 12.175 3.01 ;
      RECT 11.215 6.705 11.365 6.855 ;
      RECT 10.945 2.555 11.095 2.705 ;
      RECT 10.61 3.275 10.76 3.425 ;
      RECT 10.555 7.15 10.705 7.3 ;
      RECT 10.53 2.115 10.68 2.265 ;
      RECT 9.095 2.51 9.245 2.66 ;
      RECT 8.33 2.36 8.48 2.51 ;
      RECT 8.075 1.955 8.225 2.105 ;
      RECT 7.455 2.72 7.605 2.87 ;
      RECT 7.075 2.19 7.225 2.34 ;
      RECT 7.06 3.23 7.21 3.38 ;
      RECT 6.53 2.495 6.68 2.645 ;
      RECT 6.37 3.215 6.52 3.365 ;
      RECT 5.56 2.495 5.71 2.645 ;
      RECT 4.745 1.975 4.895 2.125 ;
      RECT 4.585 3.36 4.735 3.51 ;
      RECT 4.35 3.015 4.5 3.165 ;
      RECT 4.305 2.405 4.455 2.555 ;
      RECT 3.305 3.025 3.455 3.175 ;
      RECT 1.62 7.095 1.77 7.245 ;
      RECT 1.245 6.355 1.395 6.505 ;
      RECT 0.95 4.365 1.1 4.515 ;
      RECT 0.895 0.105 1.045 0.255 ;
      RECT 0.365 8.67 0.515 8.82 ;
    LAYER met1 ;
      RECT -0.005 8.575 81.78 8.88 ;
      RECT 72.865 6.315 73.035 8.88 ;
      RECT 57.08 6.315 57.25 8.88 ;
      RECT 41.295 6.315 41.465 8.88 ;
      RECT 25.52 6.315 25.69 8.88 ;
      RECT 9.74 6.315 9.91 8.88 ;
      RECT 73.235 6.285 73.525 6.515 ;
      RECT 57.45 6.285 57.74 6.515 ;
      RECT 41.665 6.285 41.955 6.515 ;
      RECT 25.89 6.285 26.18 6.515 ;
      RECT 10.11 6.285 10.4 6.515 ;
      RECT 72.865 6.315 73.525 6.485 ;
      RECT 57.08 6.315 57.74 6.485 ;
      RECT 41.295 6.315 41.955 6.485 ;
      RECT 25.52 6.315 26.18 6.485 ;
      RECT 9.74 6.315 10.4 6.485 ;
      RECT 66.18 1.26 75.84 1.74 ;
      RECT 50.395 1.26 60.055 1.74 ;
      RECT 34.61 1.26 44.27 1.74 ;
      RECT 18.835 1.26 28.495 1.74 ;
      RECT 3.055 1.26 12.715 1.74 ;
      RECT 66.18 1.26 75.895 1.59 ;
      RECT 50.395 1.26 60.11 1.59 ;
      RECT 34.61 1.26 44.325 1.59 ;
      RECT 18.835 1.26 28.55 1.59 ;
      RECT 3.055 1.26 12.77 1.59 ;
      RECT 66.295 0 76.01 1.585 ;
      RECT 50.51 0 60.225 1.585 ;
      RECT 34.725 0 44.44 1.585 ;
      RECT 18.95 0 28.665 1.585 ;
      RECT 3.17 0 12.885 1.585 ;
      RECT 0.795 0 1.145 0.325 ;
      RECT 0 0 81.775 0.305 ;
      RECT 0 4.135 81.775 4.745 ;
      RECT 66.18 3.98 75.84 4.745 ;
      RECT 50.395 3.98 60.055 4.745 ;
      RECT 34.61 3.98 44.27 4.745 ;
      RECT 18.835 3.98 28.495 4.745 ;
      RECT 3.055 3.98 12.715 4.745 ;
      RECT 81.175 7.765 81.465 7.995 ;
      RECT 81.235 6.285 81.405 7.995 ;
      RECT 81.205 7.275 81.555 7.625 ;
      RECT 81.175 6.285 81.465 6.515 ;
      RECT 81.175 2.365 81.465 2.595 ;
      RECT 81.235 0.885 81.405 2.595 ;
      RECT 81.175 0.885 81.465 1.115 ;
      RECT 80.765 2.735 81.095 2.965 ;
      RECT 80.765 2.765 81.265 2.935 ;
      RECT 80.765 2.395 80.955 2.965 ;
      RECT 80.185 2.365 80.475 2.595 ;
      RECT 80.185 2.395 80.955 2.565 ;
      RECT 80.245 0.885 80.415 2.595 ;
      RECT 80.185 0.885 80.475 1.115 ;
      RECT 80.185 7.765 80.475 7.995 ;
      RECT 80.245 6.285 80.415 7.995 ;
      RECT 80.185 6.285 80.475 6.515 ;
      RECT 80.185 6.325 81.035 6.485 ;
      RECT 80.865 5.915 81.035 6.485 ;
      RECT 80.185 6.32 80.575 6.485 ;
      RECT 80.805 5.915 81.095 6.145 ;
      RECT 80.805 5.945 81.265 6.115 ;
      RECT 79.815 2.735 80.105 2.965 ;
      RECT 79.815 2.765 80.275 2.935 ;
      RECT 79.875 1.655 80.04 2.965 ;
      RECT 78.39 1.625 78.68 1.855 ;
      RECT 78.39 1.655 80.04 1.825 ;
      RECT 78.45 0.885 78.62 1.855 ;
      RECT 78.39 0.885 78.68 1.115 ;
      RECT 78.39 7.765 78.68 7.995 ;
      RECT 78.45 7.025 78.62 7.995 ;
      RECT 78.45 7.12 80.04 7.29 ;
      RECT 79.87 5.915 80.04 7.29 ;
      RECT 78.39 7.025 78.68 7.255 ;
      RECT 79.815 5.915 80.105 6.145 ;
      RECT 79.815 5.945 80.275 6.115 ;
      RECT 78.82 1.965 79.17 2.315 ;
      RECT 76.485 2.025 79.17 2.195 ;
      RECT 76.485 1.34 76.655 2.195 ;
      RECT 76.385 1.34 76.735 1.69 ;
      RECT 78.845 6.655 79.17 6.98 ;
      RECT 74.22 6.61 74.57 6.96 ;
      RECT 78.82 6.655 79.17 6.885 ;
      RECT 74.04 6.655 74.57 6.885 ;
      RECT 73.87 6.685 79.17 6.855 ;
      RECT 78.045 2.365 78.365 2.685 ;
      RECT 78.015 2.365 78.365 2.595 ;
      RECT 77.845 2.395 78.365 2.565 ;
      RECT 78.045 6.255 78.365 6.545 ;
      RECT 78.015 6.285 78.365 6.515 ;
      RECT 77.845 6.315 78.365 6.485 ;
      RECT 76.99 2.705 77.34 3.055 ;
      RECT 76.99 2.765 77.48 2.935 ;
      RECT 76.995 5.855 77.345 6.205 ;
      RECT 72.24 5.915 72.53 6.145 ;
      RECT 72.24 5.945 77.48 6.115 ;
      RECT 74.68 2.465 74.865 2.675 ;
      RECT 74.67 2.47 74.88 2.668 ;
      RECT 74.67 2.47 74.966 2.645 ;
      RECT 74.67 2.47 75.025 2.62 ;
      RECT 74.67 2.47 75.08 2.6 ;
      RECT 74.67 2.47 75.09 2.588 ;
      RECT 74.67 2.47 75.285 2.527 ;
      RECT 74.67 2.47 75.315 2.51 ;
      RECT 74.67 2.47 75.335 2.5 ;
      RECT 75.215 2.235 75.475 2.495 ;
      RECT 75.2 2.325 75.215 2.542 ;
      RECT 74.735 2.457 75.475 2.495 ;
      RECT 75.186 2.336 75.2 2.548 ;
      RECT 74.775 2.45 75.475 2.495 ;
      RECT 75.1 2.376 75.186 2.567 ;
      RECT 75.025 2.437 75.475 2.495 ;
      RECT 75.095 2.412 75.1 2.584 ;
      RECT 75.08 2.422 75.475 2.495 ;
      RECT 75.09 2.417 75.095 2.586 ;
      RECT 75.385 2.922 75.39 3.014 ;
      RECT 75.38 2.9 75.385 3.031 ;
      RECT 75.375 2.89 75.38 3.043 ;
      RECT 75.365 2.881 75.375 3.053 ;
      RECT 75.36 2.876 75.365 3.061 ;
      RECT 75.355 2.735 75.36 3.064 ;
      RECT 75.321 2.735 75.355 3.075 ;
      RECT 75.235 2.735 75.321 3.11 ;
      RECT 75.155 2.735 75.235 3.158 ;
      RECT 75.126 2.735 75.155 3.182 ;
      RECT 75.04 2.735 75.126 3.188 ;
      RECT 75.035 2.919 75.04 3.193 ;
      RECT 75 2.93 75.035 3.196 ;
      RECT 74.975 2.945 75 3.2 ;
      RECT 74.961 2.954 74.975 3.202 ;
      RECT 74.875 2.981 74.961 3.208 ;
      RECT 74.81 3.022 74.875 3.217 ;
      RECT 74.795 3.042 74.81 3.222 ;
      RECT 74.765 3.052 74.795 3.225 ;
      RECT 74.76 3.062 74.765 3.228 ;
      RECT 74.73 3.067 74.76 3.23 ;
      RECT 74.71 3.072 74.73 3.234 ;
      RECT 74.625 3.075 74.71 3.241 ;
      RECT 74.61 3.072 74.625 3.247 ;
      RECT 74.6 3.069 74.61 3.249 ;
      RECT 74.58 3.066 74.6 3.251 ;
      RECT 74.56 3.062 74.58 3.252 ;
      RECT 74.545 3.058 74.56 3.254 ;
      RECT 74.535 3.055 74.545 3.255 ;
      RECT 74.495 3.049 74.535 3.253 ;
      RECT 74.485 3.044 74.495 3.251 ;
      RECT 74.47 3.041 74.485 3.247 ;
      RECT 74.445 3.036 74.47 3.24 ;
      RECT 74.395 3.027 74.445 3.228 ;
      RECT 74.325 3.013 74.395 3.21 ;
      RECT 74.267 2.998 74.325 3.192 ;
      RECT 74.181 2.981 74.267 3.172 ;
      RECT 74.095 2.96 74.181 3.147 ;
      RECT 74.045 2.945 74.095 3.128 ;
      RECT 74.041 2.939 74.045 3.12 ;
      RECT 73.955 2.929 74.041 3.107 ;
      RECT 73.92 2.914 73.955 3.09 ;
      RECT 73.905 2.907 73.92 3.083 ;
      RECT 73.845 2.895 73.905 3.071 ;
      RECT 73.825 2.882 73.845 3.059 ;
      RECT 73.785 2.873 73.825 3.051 ;
      RECT 73.78 2.865 73.785 3.044 ;
      RECT 73.7 2.855 73.78 3.03 ;
      RECT 73.685 2.842 73.7 3.015 ;
      RECT 73.68 2.84 73.685 3.013 ;
      RECT 73.601 2.828 73.68 3 ;
      RECT 73.515 2.803 73.601 2.975 ;
      RECT 73.5 2.772 73.515 2.96 ;
      RECT 73.485 2.747 73.5 2.956 ;
      RECT 73.47 2.74 73.485 2.952 ;
      RECT 73.295 2.745 73.3 2.948 ;
      RECT 73.29 2.75 73.295 2.943 ;
      RECT 73.3 2.74 73.47 2.95 ;
      RECT 74.015 2.5 74.12 2.76 ;
      RECT 74.83 2.025 74.835 2.25 ;
      RECT 74.96 2.025 75.015 2.235 ;
      RECT 75.015 2.03 75.025 2.228 ;
      RECT 74.921 2.025 74.96 2.238 ;
      RECT 74.835 2.025 74.921 2.245 ;
      RECT 74.815 2.03 74.83 2.251 ;
      RECT 74.805 2.07 74.815 2.253 ;
      RECT 74.775 2.08 74.805 2.255 ;
      RECT 74.77 2.085 74.775 2.257 ;
      RECT 74.745 2.09 74.77 2.259 ;
      RECT 74.73 2.095 74.745 2.261 ;
      RECT 74.715 2.097 74.73 2.263 ;
      RECT 74.71 2.102 74.715 2.265 ;
      RECT 74.66 2.11 74.71 2.268 ;
      RECT 74.635 2.119 74.66 2.273 ;
      RECT 74.625 2.126 74.635 2.278 ;
      RECT 74.62 2.129 74.625 2.282 ;
      RECT 74.6 2.132 74.62 2.291 ;
      RECT 74.57 2.14 74.6 2.311 ;
      RECT 74.541 2.153 74.57 2.333 ;
      RECT 74.455 2.187 74.541 2.377 ;
      RECT 74.45 2.213 74.455 2.415 ;
      RECT 74.445 2.217 74.45 2.424 ;
      RECT 74.41 2.23 74.445 2.457 ;
      RECT 74.4 2.244 74.41 2.495 ;
      RECT 74.395 2.248 74.4 2.508 ;
      RECT 74.39 2.252 74.395 2.513 ;
      RECT 74.38 2.26 74.39 2.525 ;
      RECT 74.375 2.267 74.38 2.54 ;
      RECT 74.35 2.28 74.375 2.565 ;
      RECT 74.31 2.309 74.35 2.62 ;
      RECT 74.295 2.334 74.31 2.675 ;
      RECT 74.285 2.345 74.295 2.698 ;
      RECT 74.28 2.352 74.285 2.71 ;
      RECT 74.275 2.356 74.28 2.718 ;
      RECT 74.22 2.384 74.275 2.76 ;
      RECT 74.2 2.42 74.22 2.76 ;
      RECT 74.185 2.435 74.2 2.76 ;
      RECT 74.13 2.467 74.185 2.76 ;
      RECT 74.12 2.497 74.13 2.76 ;
      RECT 73.73 2.112 73.915 2.35 ;
      RECT 73.715 2.114 73.925 2.345 ;
      RECT 73.6 2.06 73.86 2.32 ;
      RECT 73.595 2.097 73.86 2.274 ;
      RECT 73.59 2.107 73.86 2.271 ;
      RECT 73.585 2.147 73.925 2.265 ;
      RECT 73.58 2.18 73.925 2.255 ;
      RECT 73.59 2.122 73.94 2.193 ;
      RECT 73.887 3.22 73.9 3.75 ;
      RECT 73.801 3.22 73.9 3.749 ;
      RECT 73.801 3.22 73.905 3.748 ;
      RECT 73.715 3.22 73.905 3.746 ;
      RECT 73.71 3.22 73.905 3.743 ;
      RECT 73.71 3.22 73.915 3.741 ;
      RECT 73.705 3.512 73.915 3.738 ;
      RECT 73.705 3.522 73.92 3.735 ;
      RECT 73.705 3.59 73.925 3.731 ;
      RECT 73.695 3.595 73.925 3.73 ;
      RECT 73.695 3.687 73.93 3.727 ;
      RECT 73.68 3.22 73.94 3.48 ;
      RECT 73.61 7.765 73.9 7.995 ;
      RECT 73.67 7.025 73.84 7.995 ;
      RECT 73.585 7.055 73.925 7.4 ;
      RECT 73.61 7.025 73.9 7.4 ;
      RECT 72.91 2.21 72.955 3.745 ;
      RECT 73.11 2.21 73.14 2.425 ;
      RECT 71.485 1.95 71.605 2.16 ;
      RECT 71.145 1.9 71.405 2.16 ;
      RECT 71.145 1.945 71.44 2.15 ;
      RECT 73.15 2.226 73.155 2.28 ;
      RECT 73.145 2.219 73.15 2.413 ;
      RECT 73.14 2.213 73.145 2.42 ;
      RECT 73.095 2.21 73.11 2.433 ;
      RECT 73.09 2.21 73.095 2.455 ;
      RECT 73.085 2.21 73.09 2.503 ;
      RECT 73.08 2.21 73.085 2.523 ;
      RECT 73.07 2.21 73.08 2.63 ;
      RECT 73.065 2.21 73.07 2.693 ;
      RECT 73.06 2.21 73.065 2.75 ;
      RECT 73.055 2.21 73.06 2.758 ;
      RECT 73.04 2.21 73.055 2.865 ;
      RECT 73.03 2.21 73.04 3 ;
      RECT 73.02 2.21 73.03 3.11 ;
      RECT 73.01 2.21 73.02 3.167 ;
      RECT 73.005 2.21 73.01 3.207 ;
      RECT 73 2.21 73.005 3.243 ;
      RECT 72.99 2.21 73 3.283 ;
      RECT 72.985 2.21 72.99 3.325 ;
      RECT 72.965 2.21 72.985 3.39 ;
      RECT 72.97 3.535 72.975 3.715 ;
      RECT 72.965 3.517 72.97 3.723 ;
      RECT 72.96 2.21 72.965 3.453 ;
      RECT 72.96 3.497 72.965 3.73 ;
      RECT 72.955 2.21 72.96 3.74 ;
      RECT 72.9 2.21 72.91 2.51 ;
      RECT 72.905 2.757 72.91 3.745 ;
      RECT 72.9 2.822 72.905 3.745 ;
      RECT 72.895 2.211 72.9 2.5 ;
      RECT 72.89 2.887 72.9 3.745 ;
      RECT 72.885 2.212 72.895 2.49 ;
      RECT 72.875 3 72.89 3.745 ;
      RECT 72.88 2.213 72.885 2.48 ;
      RECT 72.86 2.214 72.88 2.458 ;
      RECT 72.865 3.097 72.875 3.745 ;
      RECT 72.86 3.172 72.865 3.745 ;
      RECT 72.85 2.213 72.86 2.435 ;
      RECT 72.855 3.215 72.86 3.745 ;
      RECT 72.85 3.242 72.855 3.745 ;
      RECT 72.84 2.211 72.85 2.423 ;
      RECT 72.845 3.285 72.85 3.745 ;
      RECT 72.84 3.312 72.845 3.745 ;
      RECT 72.83 2.21 72.84 2.41 ;
      RECT 72.835 3.327 72.84 3.745 ;
      RECT 72.795 3.385 72.835 3.745 ;
      RECT 72.825 2.209 72.83 2.395 ;
      RECT 72.82 2.207 72.825 2.388 ;
      RECT 72.81 2.204 72.82 2.378 ;
      RECT 72.805 2.201 72.81 2.363 ;
      RECT 72.79 2.197 72.805 2.356 ;
      RECT 72.785 3.44 72.795 3.745 ;
      RECT 72.785 2.194 72.79 2.351 ;
      RECT 72.77 2.19 72.785 2.345 ;
      RECT 72.78 3.457 72.785 3.745 ;
      RECT 72.77 3.52 72.78 3.745 ;
      RECT 72.69 2.175 72.77 2.325 ;
      RECT 72.765 3.527 72.77 3.74 ;
      RECT 72.76 3.535 72.765 3.73 ;
      RECT 72.68 2.161 72.69 2.309 ;
      RECT 72.665 2.157 72.68 2.307 ;
      RECT 72.655 2.152 72.665 2.303 ;
      RECT 72.63 2.145 72.655 2.295 ;
      RECT 72.625 2.14 72.63 2.29 ;
      RECT 72.615 2.14 72.625 2.288 ;
      RECT 72.605 2.138 72.615 2.286 ;
      RECT 72.575 2.13 72.605 2.28 ;
      RECT 72.56 2.122 72.575 2.273 ;
      RECT 72.54 2.117 72.56 2.266 ;
      RECT 72.535 2.113 72.54 2.261 ;
      RECT 72.505 2.106 72.535 2.255 ;
      RECT 72.48 2.097 72.505 2.245 ;
      RECT 72.45 2.09 72.48 2.237 ;
      RECT 72.425 2.08 72.45 2.228 ;
      RECT 72.41 2.072 72.425 2.222 ;
      RECT 72.385 2.067 72.41 2.217 ;
      RECT 72.375 2.063 72.385 2.212 ;
      RECT 72.355 2.058 72.375 2.207 ;
      RECT 72.32 2.053 72.355 2.2 ;
      RECT 72.26 2.048 72.32 2.193 ;
      RECT 72.247 2.044 72.26 2.191 ;
      RECT 72.161 2.039 72.247 2.188 ;
      RECT 72.075 2.029 72.161 2.184 ;
      RECT 72.034 2.022 72.075 2.181 ;
      RECT 71.948 2.015 72.034 2.178 ;
      RECT 71.862 2.005 71.948 2.174 ;
      RECT 71.776 1.995 71.862 2.169 ;
      RECT 71.69 1.985 71.776 2.165 ;
      RECT 71.68 1.97 71.69 2.163 ;
      RECT 71.67 1.955 71.68 2.163 ;
      RECT 71.605 1.95 71.67 2.162 ;
      RECT 71.44 1.947 71.485 2.155 ;
      RECT 72.685 2.852 72.69 3.043 ;
      RECT 72.68 2.847 72.685 3.05 ;
      RECT 72.666 2.845 72.68 3.056 ;
      RECT 72.58 2.845 72.666 3.058 ;
      RECT 72.576 2.845 72.58 3.061 ;
      RECT 72.49 2.845 72.576 3.079 ;
      RECT 72.48 2.85 72.49 3.098 ;
      RECT 72.47 2.905 72.48 3.102 ;
      RECT 72.445 2.92 72.47 3.109 ;
      RECT 72.405 2.94 72.445 3.122 ;
      RECT 72.4 2.952 72.405 3.132 ;
      RECT 72.385 2.958 72.4 3.137 ;
      RECT 72.38 2.963 72.385 3.141 ;
      RECT 72.36 2.97 72.38 3.146 ;
      RECT 72.29 2.995 72.36 3.163 ;
      RECT 72.25 3.023 72.29 3.183 ;
      RECT 72.245 3.033 72.25 3.191 ;
      RECT 72.225 3.04 72.245 3.193 ;
      RECT 72.22 3.047 72.225 3.196 ;
      RECT 72.19 3.055 72.22 3.199 ;
      RECT 72.185 3.06 72.19 3.203 ;
      RECT 72.111 3.064 72.185 3.211 ;
      RECT 72.025 3.073 72.111 3.227 ;
      RECT 72.021 3.078 72.025 3.236 ;
      RECT 71.935 3.083 72.021 3.246 ;
      RECT 71.895 3.091 71.935 3.258 ;
      RECT 71.845 3.097 71.895 3.265 ;
      RECT 71.76 3.106 71.845 3.28 ;
      RECT 71.685 3.117 71.76 3.298 ;
      RECT 71.65 3.124 71.685 3.308 ;
      RECT 71.575 3.132 71.65 3.313 ;
      RECT 71.52 3.141 71.575 3.313 ;
      RECT 71.495 3.146 71.52 3.311 ;
      RECT 71.485 3.149 71.495 3.309 ;
      RECT 71.45 3.151 71.485 3.307 ;
      RECT 71.42 3.153 71.45 3.303 ;
      RECT 71.375 3.152 71.42 3.299 ;
      RECT 71.355 3.147 71.375 3.296 ;
      RECT 71.305 3.132 71.355 3.293 ;
      RECT 71.295 3.117 71.305 3.288 ;
      RECT 71.245 3.102 71.295 3.278 ;
      RECT 71.195 3.077 71.245 3.258 ;
      RECT 71.185 3.062 71.195 3.24 ;
      RECT 71.18 3.06 71.185 3.234 ;
      RECT 71.16 3.055 71.18 3.229 ;
      RECT 71.155 3.047 71.16 3.223 ;
      RECT 71.14 3.041 71.155 3.216 ;
      RECT 71.135 3.036 71.14 3.208 ;
      RECT 71.115 3.031 71.135 3.2 ;
      RECT 71.1 3.024 71.115 3.193 ;
      RECT 71.085 3.018 71.1 3.184 ;
      RECT 71.08 3.012 71.085 3.177 ;
      RECT 71.035 2.987 71.08 3.163 ;
      RECT 71.02 2.957 71.035 3.145 ;
      RECT 71.005 2.94 71.02 3.136 ;
      RECT 70.98 2.92 71.005 3.124 ;
      RECT 70.94 2.89 70.98 3.104 ;
      RECT 70.93 2.86 70.94 3.089 ;
      RECT 70.915 2.85 70.93 3.082 ;
      RECT 70.86 2.815 70.915 3.061 ;
      RECT 70.845 2.778 70.86 3.04 ;
      RECT 70.835 2.765 70.845 3.032 ;
      RECT 70.785 2.735 70.835 3.014 ;
      RECT 70.77 2.665 70.785 2.995 ;
      RECT 70.725 2.665 70.77 2.978 ;
      RECT 70.7 2.665 70.725 2.96 ;
      RECT 70.69 2.665 70.7 2.953 ;
      RECT 70.611 2.665 70.69 2.946 ;
      RECT 70.525 2.665 70.611 2.938 ;
      RECT 70.51 2.697 70.525 2.933 ;
      RECT 70.435 2.707 70.51 2.929 ;
      RECT 70.415 2.717 70.435 2.924 ;
      RECT 70.39 2.717 70.415 2.921 ;
      RECT 70.38 2.707 70.39 2.92 ;
      RECT 70.37 2.68 70.38 2.919 ;
      RECT 70.33 2.675 70.37 2.917 ;
      RECT 70.285 2.675 70.33 2.913 ;
      RECT 70.26 2.675 70.285 2.908 ;
      RECT 70.21 2.675 70.26 2.895 ;
      RECT 70.17 2.68 70.18 2.88 ;
      RECT 70.18 2.675 70.21 2.885 ;
      RECT 72.165 2.455 72.425 2.715 ;
      RECT 72.16 2.477 72.425 2.673 ;
      RECT 71.4 2.305 71.62 2.67 ;
      RECT 71.382 2.392 71.62 2.669 ;
      RECT 71.365 2.397 71.62 2.666 ;
      RECT 71.365 2.397 71.64 2.665 ;
      RECT 71.335 2.407 71.64 2.663 ;
      RECT 71.33 2.422 71.64 2.659 ;
      RECT 71.33 2.422 71.645 2.658 ;
      RECT 71.325 2.48 71.645 2.656 ;
      RECT 71.325 2.48 71.655 2.653 ;
      RECT 71.32 2.545 71.655 2.648 ;
      RECT 71.4 2.305 71.66 2.565 ;
      RECT 70.145 2.135 70.405 2.395 ;
      RECT 70.145 2.178 70.491 2.369 ;
      RECT 70.145 2.178 70.535 2.368 ;
      RECT 70.145 2.178 70.555 2.366 ;
      RECT 70.145 2.178 70.655 2.365 ;
      RECT 70.145 2.178 70.675 2.363 ;
      RECT 70.145 2.178 70.685 2.358 ;
      RECT 70.555 2.145 70.745 2.355 ;
      RECT 70.555 2.147 70.75 2.353 ;
      RECT 70.545 2.152 70.755 2.345 ;
      RECT 70.491 2.176 70.755 2.345 ;
      RECT 70.535 2.17 70.545 2.367 ;
      RECT 70.545 2.15 70.75 2.353 ;
      RECT 69.5 3.21 69.705 3.44 ;
      RECT 69.44 3.16 69.495 3.42 ;
      RECT 69.5 3.16 69.7 3.44 ;
      RECT 70.47 3.475 70.475 3.502 ;
      RECT 70.46 3.385 70.47 3.507 ;
      RECT 70.455 3.307 70.46 3.513 ;
      RECT 70.445 3.297 70.455 3.52 ;
      RECT 70.44 3.287 70.445 3.526 ;
      RECT 70.43 3.282 70.44 3.528 ;
      RECT 70.415 3.274 70.43 3.536 ;
      RECT 70.4 3.265 70.415 3.548 ;
      RECT 70.39 3.257 70.4 3.558 ;
      RECT 70.355 3.175 70.39 3.576 ;
      RECT 70.32 3.175 70.355 3.595 ;
      RECT 70.305 3.175 70.32 3.603 ;
      RECT 70.25 3.175 70.305 3.603 ;
      RECT 70.216 3.175 70.25 3.594 ;
      RECT 70.13 3.175 70.216 3.57 ;
      RECT 70.12 3.235 70.13 3.552 ;
      RECT 70.08 3.237 70.12 3.543 ;
      RECT 70.075 3.239 70.08 3.533 ;
      RECT 70.055 3.241 70.075 3.528 ;
      RECT 70.045 3.244 70.055 3.523 ;
      RECT 70.035 3.245 70.045 3.518 ;
      RECT 70.011 3.246 70.035 3.51 ;
      RECT 69.925 3.251 70.011 3.488 ;
      RECT 69.87 3.25 69.925 3.461 ;
      RECT 69.855 3.243 69.87 3.448 ;
      RECT 69.82 3.238 69.855 3.444 ;
      RECT 69.765 3.23 69.82 3.443 ;
      RECT 69.705 3.217 69.765 3.441 ;
      RECT 69.495 3.16 69.5 3.428 ;
      RECT 69.57 2.53 69.755 2.74 ;
      RECT 69.56 2.535 69.77 2.733 ;
      RECT 69.6 2.44 69.86 2.7 ;
      RECT 69.555 2.597 69.86 2.623 ;
      RECT 68.9 2.39 68.905 3.19 ;
      RECT 68.845 2.44 68.875 3.19 ;
      RECT 68.835 2.44 68.84 2.75 ;
      RECT 68.82 2.44 68.825 2.745 ;
      RECT 68.365 2.485 68.38 2.7 ;
      RECT 68.295 2.485 68.38 2.695 ;
      RECT 69.56 2.065 69.63 2.275 ;
      RECT 69.63 2.072 69.64 2.27 ;
      RECT 69.526 2.065 69.56 2.282 ;
      RECT 69.44 2.065 69.526 2.306 ;
      RECT 69.43 2.07 69.44 2.325 ;
      RECT 69.425 2.082 69.43 2.328 ;
      RECT 69.41 2.097 69.425 2.332 ;
      RECT 69.405 2.115 69.41 2.336 ;
      RECT 69.365 2.125 69.405 2.345 ;
      RECT 69.35 2.132 69.365 2.357 ;
      RECT 69.335 2.137 69.35 2.362 ;
      RECT 69.32 2.14 69.335 2.367 ;
      RECT 69.31 2.142 69.32 2.371 ;
      RECT 69.275 2.149 69.31 2.379 ;
      RECT 69.24 2.157 69.275 2.393 ;
      RECT 69.23 2.163 69.24 2.402 ;
      RECT 69.225 2.165 69.23 2.404 ;
      RECT 69.205 2.168 69.225 2.41 ;
      RECT 69.175 2.175 69.205 2.421 ;
      RECT 69.165 2.181 69.175 2.428 ;
      RECT 69.14 2.184 69.165 2.435 ;
      RECT 69.13 2.188 69.14 2.443 ;
      RECT 69.125 2.189 69.13 2.465 ;
      RECT 69.12 2.19 69.125 2.48 ;
      RECT 69.115 2.191 69.12 2.495 ;
      RECT 69.11 2.192 69.115 2.51 ;
      RECT 69.105 2.193 69.11 2.54 ;
      RECT 69.095 2.195 69.105 2.573 ;
      RECT 69.08 2.199 69.095 2.62 ;
      RECT 69.07 2.202 69.08 2.665 ;
      RECT 69.065 2.205 69.07 2.693 ;
      RECT 69.055 2.207 69.065 2.72 ;
      RECT 69.05 2.21 69.055 2.755 ;
      RECT 69.02 2.215 69.05 2.813 ;
      RECT 69.015 2.22 69.02 2.898 ;
      RECT 69.01 2.222 69.015 2.933 ;
      RECT 69.005 2.224 69.01 3.015 ;
      RECT 69 2.226 69.005 3.103 ;
      RECT 68.99 2.228 69 3.185 ;
      RECT 68.975 2.242 68.99 3.19 ;
      RECT 68.94 2.287 68.975 3.19 ;
      RECT 68.93 2.327 68.94 3.19 ;
      RECT 68.915 2.355 68.93 3.19 ;
      RECT 68.91 2.372 68.915 3.19 ;
      RECT 68.905 2.38 68.91 3.19 ;
      RECT 68.895 2.395 68.9 3.19 ;
      RECT 68.89 2.402 68.895 3.19 ;
      RECT 68.88 2.422 68.89 3.19 ;
      RECT 68.875 2.435 68.88 3.19 ;
      RECT 68.84 2.44 68.845 2.775 ;
      RECT 68.825 2.83 68.845 3.19 ;
      RECT 68.825 2.44 68.835 2.748 ;
      RECT 68.82 2.87 68.825 3.19 ;
      RECT 68.77 2.44 68.82 2.743 ;
      RECT 68.815 2.907 68.82 3.19 ;
      RECT 68.805 2.93 68.815 3.19 ;
      RECT 68.8 2.975 68.805 3.19 ;
      RECT 68.79 2.985 68.8 3.183 ;
      RECT 68.716 2.44 68.77 2.737 ;
      RECT 68.63 2.44 68.716 2.73 ;
      RECT 68.581 2.487 68.63 2.723 ;
      RECT 68.495 2.495 68.581 2.716 ;
      RECT 68.48 2.492 68.495 2.711 ;
      RECT 68.466 2.485 68.48 2.71 ;
      RECT 68.38 2.485 68.466 2.705 ;
      RECT 68.285 2.49 68.295 2.69 ;
      RECT 67.875 1.92 67.89 2.32 ;
      RECT 68.07 1.92 68.075 2.18 ;
      RECT 67.815 1.92 67.86 2.18 ;
      RECT 68.27 3.225 68.275 3.43 ;
      RECT 68.265 3.215 68.27 3.435 ;
      RECT 68.26 3.202 68.265 3.44 ;
      RECT 68.255 3.182 68.26 3.44 ;
      RECT 68.23 3.135 68.255 3.44 ;
      RECT 68.195 3.05 68.23 3.44 ;
      RECT 68.19 2.987 68.195 3.44 ;
      RECT 68.185 2.972 68.19 3.44 ;
      RECT 68.17 2.932 68.185 3.44 ;
      RECT 68.165 2.907 68.17 3.44 ;
      RECT 68.155 2.89 68.165 3.44 ;
      RECT 68.12 2.812 68.155 3.44 ;
      RECT 68.115 2.755 68.12 3.44 ;
      RECT 68.11 2.742 68.115 3.44 ;
      RECT 68.1 2.72 68.11 3.44 ;
      RECT 68.09 2.685 68.1 3.44 ;
      RECT 68.08 2.655 68.09 3.44 ;
      RECT 68.07 2.57 68.08 3.083 ;
      RECT 68.077 3.215 68.08 3.44 ;
      RECT 68.075 3.225 68.077 3.44 ;
      RECT 68.065 3.235 68.075 3.435 ;
      RECT 68.06 1.92 68.07 2.315 ;
      RECT 68.065 2.447 68.07 3.058 ;
      RECT 68.06 2.345 68.065 3.041 ;
      RECT 68.05 1.92 68.06 3.017 ;
      RECT 68.045 1.92 68.05 2.988 ;
      RECT 68.04 1.92 68.045 2.978 ;
      RECT 68.02 1.92 68.04 2.94 ;
      RECT 68.015 1.92 68.02 2.898 ;
      RECT 68.01 1.92 68.015 2.878 ;
      RECT 67.98 1.92 68.01 2.828 ;
      RECT 67.97 1.92 67.98 2.775 ;
      RECT 67.965 1.92 67.97 2.748 ;
      RECT 67.96 1.92 67.965 2.733 ;
      RECT 67.95 1.92 67.96 2.71 ;
      RECT 67.94 1.92 67.95 2.685 ;
      RECT 67.935 1.92 67.94 2.625 ;
      RECT 67.925 1.92 67.935 2.563 ;
      RECT 67.92 1.92 67.925 2.483 ;
      RECT 67.915 1.92 67.92 2.448 ;
      RECT 67.91 1.92 67.915 2.423 ;
      RECT 67.905 1.92 67.91 2.408 ;
      RECT 67.9 1.92 67.905 2.378 ;
      RECT 67.895 1.92 67.9 2.355 ;
      RECT 67.89 1.92 67.895 2.328 ;
      RECT 67.86 1.92 67.875 2.315 ;
      RECT 67.015 3.455 67.2 3.665 ;
      RECT 67.005 3.46 67.215 3.658 ;
      RECT 67.005 3.46 67.235 3.63 ;
      RECT 67.005 3.46 67.25 3.609 ;
      RECT 67.005 3.46 67.265 3.607 ;
      RECT 67.005 3.46 67.275 3.606 ;
      RECT 67.005 3.46 67.305 3.603 ;
      RECT 67.655 3.305 67.915 3.565 ;
      RECT 67.615 3.352 67.915 3.548 ;
      RECT 67.606 3.36 67.615 3.551 ;
      RECT 67.2 3.453 67.915 3.548 ;
      RECT 67.52 3.378 67.606 3.558 ;
      RECT 67.215 3.45 67.915 3.548 ;
      RECT 67.461 3.4 67.52 3.57 ;
      RECT 67.235 3.446 67.915 3.548 ;
      RECT 67.375 3.412 67.461 3.581 ;
      RECT 67.25 3.442 67.915 3.548 ;
      RECT 67.32 3.425 67.375 3.593 ;
      RECT 67.265 3.44 67.915 3.548 ;
      RECT 67.305 3.431 67.32 3.599 ;
      RECT 67.275 3.436 67.915 3.548 ;
      RECT 67.42 2.96 67.68 3.22 ;
      RECT 67.42 2.98 67.79 3.19 ;
      RECT 67.42 2.985 67.8 3.185 ;
      RECT 67.611 2.399 67.69 2.63 ;
      RECT 67.525 2.402 67.74 2.625 ;
      RECT 67.52 2.402 67.74 2.62 ;
      RECT 67.52 2.407 67.75 2.618 ;
      RECT 67.495 2.407 67.75 2.615 ;
      RECT 67.495 2.415 67.76 2.613 ;
      RECT 67.375 2.35 67.635 2.61 ;
      RECT 67.375 2.397 67.685 2.61 ;
      RECT 66.63 2.97 66.635 3.23 ;
      RECT 66.46 2.74 66.465 3.23 ;
      RECT 66.345 2.98 66.35 3.205 ;
      RECT 67.055 2.075 67.06 2.285 ;
      RECT 67.06 2.08 67.075 2.28 ;
      RECT 66.995 2.075 67.055 2.293 ;
      RECT 66.98 2.075 66.995 2.303 ;
      RECT 66.93 2.075 66.98 2.32 ;
      RECT 66.91 2.075 66.93 2.343 ;
      RECT 66.895 2.075 66.91 2.355 ;
      RECT 66.875 2.075 66.895 2.365 ;
      RECT 66.865 2.08 66.875 2.374 ;
      RECT 66.86 2.09 66.865 2.379 ;
      RECT 66.855 2.102 66.86 2.383 ;
      RECT 66.845 2.125 66.855 2.388 ;
      RECT 66.84 2.14 66.845 2.392 ;
      RECT 66.835 2.157 66.84 2.395 ;
      RECT 66.83 2.165 66.835 2.398 ;
      RECT 66.82 2.17 66.83 2.402 ;
      RECT 66.815 2.177 66.82 2.407 ;
      RECT 66.805 2.182 66.815 2.411 ;
      RECT 66.78 2.194 66.805 2.422 ;
      RECT 66.76 2.211 66.78 2.438 ;
      RECT 66.735 2.228 66.76 2.46 ;
      RECT 66.7 2.251 66.735 2.518 ;
      RECT 66.68 2.273 66.7 2.58 ;
      RECT 66.675 2.283 66.68 2.615 ;
      RECT 66.665 2.29 66.675 2.653 ;
      RECT 66.66 2.297 66.665 2.673 ;
      RECT 66.655 2.308 66.66 2.71 ;
      RECT 66.65 2.316 66.655 2.775 ;
      RECT 66.64 2.327 66.65 2.828 ;
      RECT 66.635 2.345 66.64 2.898 ;
      RECT 66.63 2.355 66.635 2.935 ;
      RECT 66.625 2.365 66.63 3.23 ;
      RECT 66.62 2.377 66.625 3.23 ;
      RECT 66.615 2.387 66.62 3.23 ;
      RECT 66.605 2.397 66.615 3.23 ;
      RECT 66.595 2.42 66.605 3.23 ;
      RECT 66.58 2.455 66.595 3.23 ;
      RECT 66.54 2.517 66.58 3.23 ;
      RECT 66.535 2.57 66.54 3.23 ;
      RECT 66.51 2.605 66.535 3.23 ;
      RECT 66.495 2.65 66.51 3.23 ;
      RECT 66.49 2.672 66.495 3.23 ;
      RECT 66.48 2.685 66.49 3.23 ;
      RECT 66.47 2.71 66.48 3.23 ;
      RECT 66.465 2.732 66.47 3.23 ;
      RECT 66.44 2.77 66.46 3.23 ;
      RECT 66.4 2.827 66.44 3.23 ;
      RECT 66.395 2.877 66.4 3.23 ;
      RECT 66.39 2.895 66.395 3.23 ;
      RECT 66.385 2.907 66.39 3.23 ;
      RECT 66.375 2.925 66.385 3.23 ;
      RECT 66.365 2.945 66.375 3.205 ;
      RECT 66.36 2.962 66.365 3.205 ;
      RECT 66.35 2.975 66.36 3.205 ;
      RECT 66.32 2.985 66.345 3.205 ;
      RECT 66.31 2.992 66.32 3.205 ;
      RECT 66.295 3.002 66.31 3.2 ;
      RECT 65.39 7.765 65.68 7.995 ;
      RECT 65.45 6.285 65.62 7.995 ;
      RECT 65.395 6.655 65.745 7.005 ;
      RECT 65.39 6.285 65.68 6.515 ;
      RECT 65.39 2.365 65.68 2.595 ;
      RECT 65.45 0.885 65.62 2.595 ;
      RECT 65.39 0.885 65.68 1.115 ;
      RECT 64.98 2.735 65.31 2.965 ;
      RECT 64.98 2.765 65.48 2.935 ;
      RECT 64.98 2.395 65.17 2.965 ;
      RECT 64.4 2.365 64.69 2.595 ;
      RECT 64.4 2.395 65.17 2.565 ;
      RECT 64.46 0.885 64.63 2.595 ;
      RECT 64.4 0.885 64.69 1.115 ;
      RECT 64.4 7.765 64.69 7.995 ;
      RECT 64.46 6.285 64.63 7.995 ;
      RECT 64.4 6.285 64.69 6.515 ;
      RECT 64.4 6.325 65.25 6.485 ;
      RECT 65.08 5.915 65.25 6.485 ;
      RECT 64.4 6.32 64.79 6.485 ;
      RECT 65.02 5.915 65.31 6.145 ;
      RECT 65.02 5.945 65.48 6.115 ;
      RECT 64.03 2.735 64.32 2.965 ;
      RECT 64.03 2.765 64.49 2.935 ;
      RECT 64.09 1.655 64.255 2.965 ;
      RECT 62.605 1.625 62.895 1.855 ;
      RECT 62.605 1.655 64.255 1.825 ;
      RECT 62.665 0.885 62.835 1.855 ;
      RECT 62.605 0.885 62.895 1.115 ;
      RECT 62.605 7.765 62.895 7.995 ;
      RECT 62.665 7.025 62.835 7.995 ;
      RECT 62.665 7.12 64.255 7.29 ;
      RECT 64.085 5.915 64.255 7.29 ;
      RECT 62.605 7.025 62.895 7.255 ;
      RECT 64.03 5.915 64.32 6.145 ;
      RECT 64.03 5.945 64.49 6.115 ;
      RECT 63.035 1.965 63.385 2.315 ;
      RECT 60.7 2.025 63.385 2.195 ;
      RECT 60.7 1.34 60.87 2.195 ;
      RECT 60.6 1.34 60.95 1.69 ;
      RECT 63.06 6.655 63.385 6.98 ;
      RECT 58.435 6.61 58.785 6.96 ;
      RECT 63.035 6.655 63.385 6.885 ;
      RECT 58.255 6.655 58.785 6.885 ;
      RECT 58.085 6.685 63.385 6.855 ;
      RECT 62.26 2.365 62.58 2.685 ;
      RECT 62.23 2.365 62.58 2.595 ;
      RECT 62.06 2.395 62.58 2.565 ;
      RECT 62.26 6.255 62.58 6.545 ;
      RECT 62.23 6.285 62.58 6.515 ;
      RECT 62.06 6.315 62.58 6.485 ;
      RECT 61.205 2.705 61.555 3.055 ;
      RECT 61.205 2.765 61.695 2.935 ;
      RECT 61.21 5.855 61.56 6.205 ;
      RECT 56.455 5.915 56.745 6.145 ;
      RECT 56.455 5.945 61.695 6.115 ;
      RECT 58.895 2.465 59.08 2.675 ;
      RECT 58.885 2.47 59.095 2.668 ;
      RECT 58.885 2.47 59.181 2.645 ;
      RECT 58.885 2.47 59.24 2.62 ;
      RECT 58.885 2.47 59.295 2.6 ;
      RECT 58.885 2.47 59.305 2.588 ;
      RECT 58.885 2.47 59.5 2.527 ;
      RECT 58.885 2.47 59.53 2.51 ;
      RECT 58.885 2.47 59.55 2.5 ;
      RECT 59.43 2.235 59.69 2.495 ;
      RECT 59.415 2.325 59.43 2.542 ;
      RECT 58.95 2.457 59.69 2.495 ;
      RECT 59.401 2.336 59.415 2.548 ;
      RECT 58.99 2.45 59.69 2.495 ;
      RECT 59.315 2.376 59.401 2.567 ;
      RECT 59.24 2.437 59.69 2.495 ;
      RECT 59.31 2.412 59.315 2.584 ;
      RECT 59.295 2.422 59.69 2.495 ;
      RECT 59.305 2.417 59.31 2.586 ;
      RECT 59.6 2.922 59.605 3.014 ;
      RECT 59.595 2.9 59.6 3.031 ;
      RECT 59.59 2.89 59.595 3.043 ;
      RECT 59.58 2.881 59.59 3.053 ;
      RECT 59.575 2.876 59.58 3.061 ;
      RECT 59.57 2.735 59.575 3.064 ;
      RECT 59.536 2.735 59.57 3.075 ;
      RECT 59.45 2.735 59.536 3.11 ;
      RECT 59.37 2.735 59.45 3.158 ;
      RECT 59.341 2.735 59.37 3.182 ;
      RECT 59.255 2.735 59.341 3.188 ;
      RECT 59.25 2.919 59.255 3.193 ;
      RECT 59.215 2.93 59.25 3.196 ;
      RECT 59.19 2.945 59.215 3.2 ;
      RECT 59.176 2.954 59.19 3.202 ;
      RECT 59.09 2.981 59.176 3.208 ;
      RECT 59.025 3.022 59.09 3.217 ;
      RECT 59.01 3.042 59.025 3.222 ;
      RECT 58.98 3.052 59.01 3.225 ;
      RECT 58.975 3.062 58.98 3.228 ;
      RECT 58.945 3.067 58.975 3.23 ;
      RECT 58.925 3.072 58.945 3.234 ;
      RECT 58.84 3.075 58.925 3.241 ;
      RECT 58.825 3.072 58.84 3.247 ;
      RECT 58.815 3.069 58.825 3.249 ;
      RECT 58.795 3.066 58.815 3.251 ;
      RECT 58.775 3.062 58.795 3.252 ;
      RECT 58.76 3.058 58.775 3.254 ;
      RECT 58.75 3.055 58.76 3.255 ;
      RECT 58.71 3.049 58.75 3.253 ;
      RECT 58.7 3.044 58.71 3.251 ;
      RECT 58.685 3.041 58.7 3.247 ;
      RECT 58.66 3.036 58.685 3.24 ;
      RECT 58.61 3.027 58.66 3.228 ;
      RECT 58.54 3.013 58.61 3.21 ;
      RECT 58.482 2.998 58.54 3.192 ;
      RECT 58.396 2.981 58.482 3.172 ;
      RECT 58.31 2.96 58.396 3.147 ;
      RECT 58.26 2.945 58.31 3.128 ;
      RECT 58.256 2.939 58.26 3.12 ;
      RECT 58.17 2.929 58.256 3.107 ;
      RECT 58.135 2.914 58.17 3.09 ;
      RECT 58.12 2.907 58.135 3.083 ;
      RECT 58.06 2.895 58.12 3.071 ;
      RECT 58.04 2.882 58.06 3.059 ;
      RECT 58 2.873 58.04 3.051 ;
      RECT 57.995 2.865 58 3.044 ;
      RECT 57.915 2.855 57.995 3.03 ;
      RECT 57.9 2.842 57.915 3.015 ;
      RECT 57.895 2.84 57.9 3.013 ;
      RECT 57.816 2.828 57.895 3 ;
      RECT 57.73 2.803 57.816 2.975 ;
      RECT 57.715 2.772 57.73 2.96 ;
      RECT 57.7 2.747 57.715 2.956 ;
      RECT 57.685 2.74 57.7 2.952 ;
      RECT 57.51 2.745 57.515 2.948 ;
      RECT 57.505 2.75 57.51 2.943 ;
      RECT 57.515 2.74 57.685 2.95 ;
      RECT 58.23 2.5 58.335 2.76 ;
      RECT 59.045 2.025 59.05 2.25 ;
      RECT 59.175 2.025 59.23 2.235 ;
      RECT 59.23 2.03 59.24 2.228 ;
      RECT 59.136 2.025 59.175 2.238 ;
      RECT 59.05 2.025 59.136 2.245 ;
      RECT 59.03 2.03 59.045 2.251 ;
      RECT 59.02 2.07 59.03 2.253 ;
      RECT 58.99 2.08 59.02 2.255 ;
      RECT 58.985 2.085 58.99 2.257 ;
      RECT 58.96 2.09 58.985 2.259 ;
      RECT 58.945 2.095 58.96 2.261 ;
      RECT 58.93 2.097 58.945 2.263 ;
      RECT 58.925 2.102 58.93 2.265 ;
      RECT 58.875 2.11 58.925 2.268 ;
      RECT 58.85 2.119 58.875 2.273 ;
      RECT 58.84 2.126 58.85 2.278 ;
      RECT 58.835 2.129 58.84 2.282 ;
      RECT 58.815 2.132 58.835 2.291 ;
      RECT 58.785 2.14 58.815 2.311 ;
      RECT 58.756 2.153 58.785 2.333 ;
      RECT 58.67 2.187 58.756 2.377 ;
      RECT 58.665 2.213 58.67 2.415 ;
      RECT 58.66 2.217 58.665 2.424 ;
      RECT 58.625 2.23 58.66 2.457 ;
      RECT 58.615 2.244 58.625 2.495 ;
      RECT 58.61 2.248 58.615 2.508 ;
      RECT 58.605 2.252 58.61 2.513 ;
      RECT 58.595 2.26 58.605 2.525 ;
      RECT 58.59 2.267 58.595 2.54 ;
      RECT 58.565 2.28 58.59 2.565 ;
      RECT 58.525 2.309 58.565 2.62 ;
      RECT 58.51 2.334 58.525 2.675 ;
      RECT 58.5 2.345 58.51 2.698 ;
      RECT 58.495 2.352 58.5 2.71 ;
      RECT 58.49 2.356 58.495 2.718 ;
      RECT 58.435 2.384 58.49 2.76 ;
      RECT 58.415 2.42 58.435 2.76 ;
      RECT 58.4 2.435 58.415 2.76 ;
      RECT 58.345 2.467 58.4 2.76 ;
      RECT 58.335 2.497 58.345 2.76 ;
      RECT 57.945 2.112 58.13 2.35 ;
      RECT 57.93 2.114 58.14 2.345 ;
      RECT 57.815 2.06 58.075 2.32 ;
      RECT 57.81 2.097 58.075 2.274 ;
      RECT 57.805 2.107 58.075 2.271 ;
      RECT 57.8 2.147 58.14 2.265 ;
      RECT 57.795 2.18 58.14 2.255 ;
      RECT 57.805 2.122 58.155 2.193 ;
      RECT 58.102 3.22 58.115 3.75 ;
      RECT 58.016 3.22 58.115 3.749 ;
      RECT 58.016 3.22 58.12 3.748 ;
      RECT 57.93 3.22 58.12 3.746 ;
      RECT 57.925 3.22 58.12 3.743 ;
      RECT 57.925 3.22 58.13 3.741 ;
      RECT 57.92 3.512 58.13 3.738 ;
      RECT 57.92 3.522 58.135 3.735 ;
      RECT 57.92 3.59 58.14 3.731 ;
      RECT 57.91 3.595 58.14 3.73 ;
      RECT 57.91 3.687 58.145 3.727 ;
      RECT 57.895 3.22 58.155 3.48 ;
      RECT 57.825 7.765 58.115 7.995 ;
      RECT 57.885 7.025 58.055 7.995 ;
      RECT 57.8 7.055 58.14 7.4 ;
      RECT 57.825 7.025 58.115 7.4 ;
      RECT 57.125 2.21 57.17 3.745 ;
      RECT 57.325 2.21 57.355 2.425 ;
      RECT 55.7 1.95 55.82 2.16 ;
      RECT 55.36 1.9 55.62 2.16 ;
      RECT 55.36 1.945 55.655 2.15 ;
      RECT 57.365 2.226 57.37 2.28 ;
      RECT 57.36 2.219 57.365 2.413 ;
      RECT 57.355 2.213 57.36 2.42 ;
      RECT 57.31 2.21 57.325 2.433 ;
      RECT 57.305 2.21 57.31 2.455 ;
      RECT 57.3 2.21 57.305 2.503 ;
      RECT 57.295 2.21 57.3 2.523 ;
      RECT 57.285 2.21 57.295 2.63 ;
      RECT 57.28 2.21 57.285 2.693 ;
      RECT 57.275 2.21 57.28 2.75 ;
      RECT 57.27 2.21 57.275 2.758 ;
      RECT 57.255 2.21 57.27 2.865 ;
      RECT 57.245 2.21 57.255 3 ;
      RECT 57.235 2.21 57.245 3.11 ;
      RECT 57.225 2.21 57.235 3.167 ;
      RECT 57.22 2.21 57.225 3.207 ;
      RECT 57.215 2.21 57.22 3.243 ;
      RECT 57.205 2.21 57.215 3.283 ;
      RECT 57.2 2.21 57.205 3.325 ;
      RECT 57.18 2.21 57.2 3.39 ;
      RECT 57.185 3.535 57.19 3.715 ;
      RECT 57.18 3.517 57.185 3.723 ;
      RECT 57.175 2.21 57.18 3.453 ;
      RECT 57.175 3.497 57.18 3.73 ;
      RECT 57.17 2.21 57.175 3.74 ;
      RECT 57.115 2.21 57.125 2.51 ;
      RECT 57.12 2.757 57.125 3.745 ;
      RECT 57.115 2.822 57.12 3.745 ;
      RECT 57.11 2.211 57.115 2.5 ;
      RECT 57.105 2.887 57.115 3.745 ;
      RECT 57.1 2.212 57.11 2.49 ;
      RECT 57.09 3 57.105 3.745 ;
      RECT 57.095 2.213 57.1 2.48 ;
      RECT 57.075 2.214 57.095 2.458 ;
      RECT 57.08 3.097 57.09 3.745 ;
      RECT 57.075 3.172 57.08 3.745 ;
      RECT 57.065 2.213 57.075 2.435 ;
      RECT 57.07 3.215 57.075 3.745 ;
      RECT 57.065 3.242 57.07 3.745 ;
      RECT 57.055 2.211 57.065 2.423 ;
      RECT 57.06 3.285 57.065 3.745 ;
      RECT 57.055 3.312 57.06 3.745 ;
      RECT 57.045 2.21 57.055 2.41 ;
      RECT 57.05 3.327 57.055 3.745 ;
      RECT 57.01 3.385 57.05 3.745 ;
      RECT 57.04 2.209 57.045 2.395 ;
      RECT 57.035 2.207 57.04 2.388 ;
      RECT 57.025 2.204 57.035 2.378 ;
      RECT 57.02 2.201 57.025 2.363 ;
      RECT 57.005 2.197 57.02 2.356 ;
      RECT 57 3.44 57.01 3.745 ;
      RECT 57 2.194 57.005 2.351 ;
      RECT 56.985 2.19 57 2.345 ;
      RECT 56.995 3.457 57 3.745 ;
      RECT 56.985 3.52 56.995 3.745 ;
      RECT 56.905 2.175 56.985 2.325 ;
      RECT 56.98 3.527 56.985 3.74 ;
      RECT 56.975 3.535 56.98 3.73 ;
      RECT 56.895 2.161 56.905 2.309 ;
      RECT 56.88 2.157 56.895 2.307 ;
      RECT 56.87 2.152 56.88 2.303 ;
      RECT 56.845 2.145 56.87 2.295 ;
      RECT 56.84 2.14 56.845 2.29 ;
      RECT 56.83 2.14 56.84 2.288 ;
      RECT 56.82 2.138 56.83 2.286 ;
      RECT 56.79 2.13 56.82 2.28 ;
      RECT 56.775 2.122 56.79 2.273 ;
      RECT 56.755 2.117 56.775 2.266 ;
      RECT 56.75 2.113 56.755 2.261 ;
      RECT 56.72 2.106 56.75 2.255 ;
      RECT 56.695 2.097 56.72 2.245 ;
      RECT 56.665 2.09 56.695 2.237 ;
      RECT 56.64 2.08 56.665 2.228 ;
      RECT 56.625 2.072 56.64 2.222 ;
      RECT 56.6 2.067 56.625 2.217 ;
      RECT 56.59 2.063 56.6 2.212 ;
      RECT 56.57 2.058 56.59 2.207 ;
      RECT 56.535 2.053 56.57 2.2 ;
      RECT 56.475 2.048 56.535 2.193 ;
      RECT 56.462 2.044 56.475 2.191 ;
      RECT 56.376 2.039 56.462 2.188 ;
      RECT 56.29 2.029 56.376 2.184 ;
      RECT 56.249 2.022 56.29 2.181 ;
      RECT 56.163 2.015 56.249 2.178 ;
      RECT 56.077 2.005 56.163 2.174 ;
      RECT 55.991 1.995 56.077 2.169 ;
      RECT 55.905 1.985 55.991 2.165 ;
      RECT 55.895 1.97 55.905 2.163 ;
      RECT 55.885 1.955 55.895 2.163 ;
      RECT 55.82 1.95 55.885 2.162 ;
      RECT 55.655 1.947 55.7 2.155 ;
      RECT 56.9 2.852 56.905 3.043 ;
      RECT 56.895 2.847 56.9 3.05 ;
      RECT 56.881 2.845 56.895 3.056 ;
      RECT 56.795 2.845 56.881 3.058 ;
      RECT 56.791 2.845 56.795 3.061 ;
      RECT 56.705 2.845 56.791 3.079 ;
      RECT 56.695 2.85 56.705 3.098 ;
      RECT 56.685 2.905 56.695 3.102 ;
      RECT 56.66 2.92 56.685 3.109 ;
      RECT 56.62 2.94 56.66 3.122 ;
      RECT 56.615 2.952 56.62 3.132 ;
      RECT 56.6 2.958 56.615 3.137 ;
      RECT 56.595 2.963 56.6 3.141 ;
      RECT 56.575 2.97 56.595 3.146 ;
      RECT 56.505 2.995 56.575 3.163 ;
      RECT 56.465 3.023 56.505 3.183 ;
      RECT 56.46 3.033 56.465 3.191 ;
      RECT 56.44 3.04 56.46 3.193 ;
      RECT 56.435 3.047 56.44 3.196 ;
      RECT 56.405 3.055 56.435 3.199 ;
      RECT 56.4 3.06 56.405 3.203 ;
      RECT 56.326 3.064 56.4 3.211 ;
      RECT 56.24 3.073 56.326 3.227 ;
      RECT 56.236 3.078 56.24 3.236 ;
      RECT 56.15 3.083 56.236 3.246 ;
      RECT 56.11 3.091 56.15 3.258 ;
      RECT 56.06 3.097 56.11 3.265 ;
      RECT 55.975 3.106 56.06 3.28 ;
      RECT 55.9 3.117 55.975 3.298 ;
      RECT 55.865 3.124 55.9 3.308 ;
      RECT 55.79 3.132 55.865 3.313 ;
      RECT 55.735 3.141 55.79 3.313 ;
      RECT 55.71 3.146 55.735 3.311 ;
      RECT 55.7 3.149 55.71 3.309 ;
      RECT 55.665 3.151 55.7 3.307 ;
      RECT 55.635 3.153 55.665 3.303 ;
      RECT 55.59 3.152 55.635 3.299 ;
      RECT 55.57 3.147 55.59 3.296 ;
      RECT 55.52 3.132 55.57 3.293 ;
      RECT 55.51 3.117 55.52 3.288 ;
      RECT 55.46 3.102 55.51 3.278 ;
      RECT 55.41 3.077 55.46 3.258 ;
      RECT 55.4 3.062 55.41 3.24 ;
      RECT 55.395 3.06 55.4 3.234 ;
      RECT 55.375 3.055 55.395 3.229 ;
      RECT 55.37 3.047 55.375 3.223 ;
      RECT 55.355 3.041 55.37 3.216 ;
      RECT 55.35 3.036 55.355 3.208 ;
      RECT 55.33 3.031 55.35 3.2 ;
      RECT 55.315 3.024 55.33 3.193 ;
      RECT 55.3 3.018 55.315 3.184 ;
      RECT 55.295 3.012 55.3 3.177 ;
      RECT 55.25 2.987 55.295 3.163 ;
      RECT 55.235 2.957 55.25 3.145 ;
      RECT 55.22 2.94 55.235 3.136 ;
      RECT 55.195 2.92 55.22 3.124 ;
      RECT 55.155 2.89 55.195 3.104 ;
      RECT 55.145 2.86 55.155 3.089 ;
      RECT 55.13 2.85 55.145 3.082 ;
      RECT 55.075 2.815 55.13 3.061 ;
      RECT 55.06 2.778 55.075 3.04 ;
      RECT 55.05 2.765 55.06 3.032 ;
      RECT 55 2.735 55.05 3.014 ;
      RECT 54.985 2.665 55 2.995 ;
      RECT 54.94 2.665 54.985 2.978 ;
      RECT 54.915 2.665 54.94 2.96 ;
      RECT 54.905 2.665 54.915 2.953 ;
      RECT 54.826 2.665 54.905 2.946 ;
      RECT 54.74 2.665 54.826 2.938 ;
      RECT 54.725 2.697 54.74 2.933 ;
      RECT 54.65 2.707 54.725 2.929 ;
      RECT 54.63 2.717 54.65 2.924 ;
      RECT 54.605 2.717 54.63 2.921 ;
      RECT 54.595 2.707 54.605 2.92 ;
      RECT 54.585 2.68 54.595 2.919 ;
      RECT 54.545 2.675 54.585 2.917 ;
      RECT 54.5 2.675 54.545 2.913 ;
      RECT 54.475 2.675 54.5 2.908 ;
      RECT 54.425 2.675 54.475 2.895 ;
      RECT 54.385 2.68 54.395 2.88 ;
      RECT 54.395 2.675 54.425 2.885 ;
      RECT 56.38 2.455 56.64 2.715 ;
      RECT 56.375 2.477 56.64 2.673 ;
      RECT 55.615 2.305 55.835 2.67 ;
      RECT 55.597 2.392 55.835 2.669 ;
      RECT 55.58 2.397 55.835 2.666 ;
      RECT 55.58 2.397 55.855 2.665 ;
      RECT 55.55 2.407 55.855 2.663 ;
      RECT 55.545 2.422 55.855 2.659 ;
      RECT 55.545 2.422 55.86 2.658 ;
      RECT 55.54 2.48 55.86 2.656 ;
      RECT 55.54 2.48 55.87 2.653 ;
      RECT 55.535 2.545 55.87 2.648 ;
      RECT 55.615 2.305 55.875 2.565 ;
      RECT 54.36 2.135 54.62 2.395 ;
      RECT 54.36 2.178 54.706 2.369 ;
      RECT 54.36 2.178 54.75 2.368 ;
      RECT 54.36 2.178 54.77 2.366 ;
      RECT 54.36 2.178 54.87 2.365 ;
      RECT 54.36 2.178 54.89 2.363 ;
      RECT 54.36 2.178 54.9 2.358 ;
      RECT 54.77 2.145 54.96 2.355 ;
      RECT 54.77 2.147 54.965 2.353 ;
      RECT 54.76 2.152 54.97 2.345 ;
      RECT 54.706 2.176 54.97 2.345 ;
      RECT 54.75 2.17 54.76 2.367 ;
      RECT 54.76 2.15 54.965 2.353 ;
      RECT 53.715 3.21 53.92 3.44 ;
      RECT 53.655 3.16 53.71 3.42 ;
      RECT 53.715 3.16 53.915 3.44 ;
      RECT 54.685 3.475 54.69 3.502 ;
      RECT 54.675 3.385 54.685 3.507 ;
      RECT 54.67 3.307 54.675 3.513 ;
      RECT 54.66 3.297 54.67 3.52 ;
      RECT 54.655 3.287 54.66 3.526 ;
      RECT 54.645 3.282 54.655 3.528 ;
      RECT 54.63 3.274 54.645 3.536 ;
      RECT 54.615 3.265 54.63 3.548 ;
      RECT 54.605 3.257 54.615 3.558 ;
      RECT 54.57 3.175 54.605 3.576 ;
      RECT 54.535 3.175 54.57 3.595 ;
      RECT 54.52 3.175 54.535 3.603 ;
      RECT 54.465 3.175 54.52 3.603 ;
      RECT 54.431 3.175 54.465 3.594 ;
      RECT 54.345 3.175 54.431 3.57 ;
      RECT 54.335 3.235 54.345 3.552 ;
      RECT 54.295 3.237 54.335 3.543 ;
      RECT 54.29 3.239 54.295 3.533 ;
      RECT 54.27 3.241 54.29 3.528 ;
      RECT 54.26 3.244 54.27 3.523 ;
      RECT 54.25 3.245 54.26 3.518 ;
      RECT 54.226 3.246 54.25 3.51 ;
      RECT 54.14 3.251 54.226 3.488 ;
      RECT 54.085 3.25 54.14 3.461 ;
      RECT 54.07 3.243 54.085 3.448 ;
      RECT 54.035 3.238 54.07 3.444 ;
      RECT 53.98 3.23 54.035 3.443 ;
      RECT 53.92 3.217 53.98 3.441 ;
      RECT 53.71 3.16 53.715 3.428 ;
      RECT 53.785 2.53 53.97 2.74 ;
      RECT 53.775 2.535 53.985 2.733 ;
      RECT 53.815 2.44 54.075 2.7 ;
      RECT 53.77 2.597 54.075 2.623 ;
      RECT 53.115 2.39 53.12 3.19 ;
      RECT 53.06 2.44 53.09 3.19 ;
      RECT 53.05 2.44 53.055 2.75 ;
      RECT 53.035 2.44 53.04 2.745 ;
      RECT 52.58 2.485 52.595 2.7 ;
      RECT 52.51 2.485 52.595 2.695 ;
      RECT 53.775 2.065 53.845 2.275 ;
      RECT 53.845 2.072 53.855 2.27 ;
      RECT 53.741 2.065 53.775 2.282 ;
      RECT 53.655 2.065 53.741 2.306 ;
      RECT 53.645 2.07 53.655 2.325 ;
      RECT 53.64 2.082 53.645 2.328 ;
      RECT 53.625 2.097 53.64 2.332 ;
      RECT 53.62 2.115 53.625 2.336 ;
      RECT 53.58 2.125 53.62 2.345 ;
      RECT 53.565 2.132 53.58 2.357 ;
      RECT 53.55 2.137 53.565 2.362 ;
      RECT 53.535 2.14 53.55 2.367 ;
      RECT 53.525 2.142 53.535 2.371 ;
      RECT 53.49 2.149 53.525 2.379 ;
      RECT 53.455 2.157 53.49 2.393 ;
      RECT 53.445 2.163 53.455 2.402 ;
      RECT 53.44 2.165 53.445 2.404 ;
      RECT 53.42 2.168 53.44 2.41 ;
      RECT 53.39 2.175 53.42 2.421 ;
      RECT 53.38 2.181 53.39 2.428 ;
      RECT 53.355 2.184 53.38 2.435 ;
      RECT 53.345 2.188 53.355 2.443 ;
      RECT 53.34 2.189 53.345 2.465 ;
      RECT 53.335 2.19 53.34 2.48 ;
      RECT 53.33 2.191 53.335 2.495 ;
      RECT 53.325 2.192 53.33 2.51 ;
      RECT 53.32 2.193 53.325 2.54 ;
      RECT 53.31 2.195 53.32 2.573 ;
      RECT 53.295 2.199 53.31 2.62 ;
      RECT 53.285 2.202 53.295 2.665 ;
      RECT 53.28 2.205 53.285 2.693 ;
      RECT 53.27 2.207 53.28 2.72 ;
      RECT 53.265 2.21 53.27 2.755 ;
      RECT 53.235 2.215 53.265 2.813 ;
      RECT 53.23 2.22 53.235 2.898 ;
      RECT 53.225 2.222 53.23 2.933 ;
      RECT 53.22 2.224 53.225 3.015 ;
      RECT 53.215 2.226 53.22 3.103 ;
      RECT 53.205 2.228 53.215 3.185 ;
      RECT 53.19 2.242 53.205 3.19 ;
      RECT 53.155 2.287 53.19 3.19 ;
      RECT 53.145 2.327 53.155 3.19 ;
      RECT 53.13 2.355 53.145 3.19 ;
      RECT 53.125 2.372 53.13 3.19 ;
      RECT 53.12 2.38 53.125 3.19 ;
      RECT 53.11 2.395 53.115 3.19 ;
      RECT 53.105 2.402 53.11 3.19 ;
      RECT 53.095 2.422 53.105 3.19 ;
      RECT 53.09 2.435 53.095 3.19 ;
      RECT 53.055 2.44 53.06 2.775 ;
      RECT 53.04 2.83 53.06 3.19 ;
      RECT 53.04 2.44 53.05 2.748 ;
      RECT 53.035 2.87 53.04 3.19 ;
      RECT 52.985 2.44 53.035 2.743 ;
      RECT 53.03 2.907 53.035 3.19 ;
      RECT 53.02 2.93 53.03 3.19 ;
      RECT 53.015 2.975 53.02 3.19 ;
      RECT 53.005 2.985 53.015 3.183 ;
      RECT 52.931 2.44 52.985 2.737 ;
      RECT 52.845 2.44 52.931 2.73 ;
      RECT 52.796 2.487 52.845 2.723 ;
      RECT 52.71 2.495 52.796 2.716 ;
      RECT 52.695 2.492 52.71 2.711 ;
      RECT 52.681 2.485 52.695 2.71 ;
      RECT 52.595 2.485 52.681 2.705 ;
      RECT 52.5 2.49 52.51 2.69 ;
      RECT 52.09 1.92 52.105 2.32 ;
      RECT 52.285 1.92 52.29 2.18 ;
      RECT 52.03 1.92 52.075 2.18 ;
      RECT 52.485 3.225 52.49 3.43 ;
      RECT 52.48 3.215 52.485 3.435 ;
      RECT 52.475 3.202 52.48 3.44 ;
      RECT 52.47 3.182 52.475 3.44 ;
      RECT 52.445 3.135 52.47 3.44 ;
      RECT 52.41 3.05 52.445 3.44 ;
      RECT 52.405 2.987 52.41 3.44 ;
      RECT 52.4 2.972 52.405 3.44 ;
      RECT 52.385 2.932 52.4 3.44 ;
      RECT 52.38 2.907 52.385 3.44 ;
      RECT 52.37 2.89 52.38 3.44 ;
      RECT 52.335 2.812 52.37 3.44 ;
      RECT 52.33 2.755 52.335 3.44 ;
      RECT 52.325 2.742 52.33 3.44 ;
      RECT 52.315 2.72 52.325 3.44 ;
      RECT 52.305 2.685 52.315 3.44 ;
      RECT 52.295 2.655 52.305 3.44 ;
      RECT 52.285 2.57 52.295 3.083 ;
      RECT 52.292 3.215 52.295 3.44 ;
      RECT 52.29 3.225 52.292 3.44 ;
      RECT 52.28 3.235 52.29 3.435 ;
      RECT 52.275 1.92 52.285 2.315 ;
      RECT 52.28 2.447 52.285 3.058 ;
      RECT 52.275 2.345 52.28 3.041 ;
      RECT 52.265 1.92 52.275 3.017 ;
      RECT 52.26 1.92 52.265 2.988 ;
      RECT 52.255 1.92 52.26 2.978 ;
      RECT 52.235 1.92 52.255 2.94 ;
      RECT 52.23 1.92 52.235 2.898 ;
      RECT 52.225 1.92 52.23 2.878 ;
      RECT 52.195 1.92 52.225 2.828 ;
      RECT 52.185 1.92 52.195 2.775 ;
      RECT 52.18 1.92 52.185 2.748 ;
      RECT 52.175 1.92 52.18 2.733 ;
      RECT 52.165 1.92 52.175 2.71 ;
      RECT 52.155 1.92 52.165 2.685 ;
      RECT 52.15 1.92 52.155 2.625 ;
      RECT 52.14 1.92 52.15 2.563 ;
      RECT 52.135 1.92 52.14 2.483 ;
      RECT 52.13 1.92 52.135 2.448 ;
      RECT 52.125 1.92 52.13 2.423 ;
      RECT 52.12 1.92 52.125 2.408 ;
      RECT 52.115 1.92 52.12 2.378 ;
      RECT 52.11 1.92 52.115 2.355 ;
      RECT 52.105 1.92 52.11 2.328 ;
      RECT 52.075 1.92 52.09 2.315 ;
      RECT 51.23 3.455 51.415 3.665 ;
      RECT 51.22 3.46 51.43 3.658 ;
      RECT 51.22 3.46 51.45 3.63 ;
      RECT 51.22 3.46 51.465 3.609 ;
      RECT 51.22 3.46 51.48 3.607 ;
      RECT 51.22 3.46 51.49 3.606 ;
      RECT 51.22 3.46 51.52 3.603 ;
      RECT 51.87 3.305 52.13 3.565 ;
      RECT 51.83 3.352 52.13 3.548 ;
      RECT 51.821 3.36 51.83 3.551 ;
      RECT 51.415 3.453 52.13 3.548 ;
      RECT 51.735 3.378 51.821 3.558 ;
      RECT 51.43 3.45 52.13 3.548 ;
      RECT 51.676 3.4 51.735 3.57 ;
      RECT 51.45 3.446 52.13 3.548 ;
      RECT 51.59 3.412 51.676 3.581 ;
      RECT 51.465 3.442 52.13 3.548 ;
      RECT 51.535 3.425 51.59 3.593 ;
      RECT 51.48 3.44 52.13 3.548 ;
      RECT 51.52 3.431 51.535 3.599 ;
      RECT 51.49 3.436 52.13 3.548 ;
      RECT 51.635 2.96 51.895 3.22 ;
      RECT 51.635 2.98 52.005 3.19 ;
      RECT 51.635 2.985 52.015 3.185 ;
      RECT 51.826 2.399 51.905 2.63 ;
      RECT 51.74 2.402 51.955 2.625 ;
      RECT 51.735 2.402 51.955 2.62 ;
      RECT 51.735 2.407 51.965 2.618 ;
      RECT 51.71 2.407 51.965 2.615 ;
      RECT 51.71 2.415 51.975 2.613 ;
      RECT 51.59 2.35 51.85 2.61 ;
      RECT 51.59 2.397 51.9 2.61 ;
      RECT 50.845 2.97 50.85 3.23 ;
      RECT 50.675 2.74 50.68 3.23 ;
      RECT 50.56 2.98 50.565 3.205 ;
      RECT 51.27 2.075 51.275 2.285 ;
      RECT 51.275 2.08 51.29 2.28 ;
      RECT 51.21 2.075 51.27 2.293 ;
      RECT 51.195 2.075 51.21 2.303 ;
      RECT 51.145 2.075 51.195 2.32 ;
      RECT 51.125 2.075 51.145 2.343 ;
      RECT 51.11 2.075 51.125 2.355 ;
      RECT 51.09 2.075 51.11 2.365 ;
      RECT 51.08 2.08 51.09 2.374 ;
      RECT 51.075 2.09 51.08 2.379 ;
      RECT 51.07 2.102 51.075 2.383 ;
      RECT 51.06 2.125 51.07 2.388 ;
      RECT 51.055 2.14 51.06 2.392 ;
      RECT 51.05 2.157 51.055 2.395 ;
      RECT 51.045 2.165 51.05 2.398 ;
      RECT 51.035 2.17 51.045 2.402 ;
      RECT 51.03 2.177 51.035 2.407 ;
      RECT 51.02 2.182 51.03 2.411 ;
      RECT 50.995 2.194 51.02 2.422 ;
      RECT 50.975 2.211 50.995 2.438 ;
      RECT 50.95 2.228 50.975 2.46 ;
      RECT 50.915 2.251 50.95 2.518 ;
      RECT 50.895 2.273 50.915 2.58 ;
      RECT 50.89 2.283 50.895 2.615 ;
      RECT 50.88 2.29 50.89 2.653 ;
      RECT 50.875 2.297 50.88 2.673 ;
      RECT 50.87 2.308 50.875 2.71 ;
      RECT 50.865 2.316 50.87 2.775 ;
      RECT 50.855 2.327 50.865 2.828 ;
      RECT 50.85 2.345 50.855 2.898 ;
      RECT 50.845 2.355 50.85 2.935 ;
      RECT 50.84 2.365 50.845 3.23 ;
      RECT 50.835 2.377 50.84 3.23 ;
      RECT 50.83 2.387 50.835 3.23 ;
      RECT 50.82 2.397 50.83 3.23 ;
      RECT 50.81 2.42 50.82 3.23 ;
      RECT 50.795 2.455 50.81 3.23 ;
      RECT 50.755 2.517 50.795 3.23 ;
      RECT 50.75 2.57 50.755 3.23 ;
      RECT 50.725 2.605 50.75 3.23 ;
      RECT 50.71 2.65 50.725 3.23 ;
      RECT 50.705 2.672 50.71 3.23 ;
      RECT 50.695 2.685 50.705 3.23 ;
      RECT 50.685 2.71 50.695 3.23 ;
      RECT 50.68 2.732 50.685 3.23 ;
      RECT 50.655 2.77 50.675 3.23 ;
      RECT 50.615 2.827 50.655 3.23 ;
      RECT 50.61 2.877 50.615 3.23 ;
      RECT 50.605 2.895 50.61 3.23 ;
      RECT 50.6 2.907 50.605 3.23 ;
      RECT 50.59 2.925 50.6 3.23 ;
      RECT 50.58 2.945 50.59 3.205 ;
      RECT 50.575 2.962 50.58 3.205 ;
      RECT 50.565 2.975 50.575 3.205 ;
      RECT 50.535 2.985 50.56 3.205 ;
      RECT 50.525 2.992 50.535 3.205 ;
      RECT 50.51 3.002 50.525 3.2 ;
      RECT 49.605 7.765 49.895 7.995 ;
      RECT 49.665 6.285 49.835 7.995 ;
      RECT 49.61 6.655 49.96 7.005 ;
      RECT 49.605 6.285 49.895 6.515 ;
      RECT 49.605 2.365 49.895 2.595 ;
      RECT 49.665 0.885 49.835 2.595 ;
      RECT 49.605 0.885 49.895 1.115 ;
      RECT 49.195 2.735 49.525 2.965 ;
      RECT 49.195 2.765 49.695 2.935 ;
      RECT 49.195 2.395 49.385 2.965 ;
      RECT 48.615 2.365 48.905 2.595 ;
      RECT 48.615 2.395 49.385 2.565 ;
      RECT 48.675 0.885 48.845 2.595 ;
      RECT 48.615 0.885 48.905 1.115 ;
      RECT 48.615 7.765 48.905 7.995 ;
      RECT 48.675 6.285 48.845 7.995 ;
      RECT 48.615 6.285 48.905 6.515 ;
      RECT 48.615 6.325 49.465 6.485 ;
      RECT 49.295 5.915 49.465 6.485 ;
      RECT 48.615 6.32 49.005 6.485 ;
      RECT 49.235 5.915 49.525 6.145 ;
      RECT 49.235 5.945 49.695 6.115 ;
      RECT 48.245 2.735 48.535 2.965 ;
      RECT 48.245 2.765 48.705 2.935 ;
      RECT 48.305 1.655 48.47 2.965 ;
      RECT 46.82 1.625 47.11 1.855 ;
      RECT 46.82 1.655 48.47 1.825 ;
      RECT 46.88 0.885 47.05 1.855 ;
      RECT 46.82 0.885 47.11 1.115 ;
      RECT 46.82 7.765 47.11 7.995 ;
      RECT 46.88 7.025 47.05 7.995 ;
      RECT 46.88 7.12 48.47 7.29 ;
      RECT 48.3 5.915 48.47 7.29 ;
      RECT 46.82 7.025 47.11 7.255 ;
      RECT 48.245 5.915 48.535 6.145 ;
      RECT 48.245 5.945 48.705 6.115 ;
      RECT 47.25 1.965 47.6 2.315 ;
      RECT 44.915 2.025 47.6 2.195 ;
      RECT 44.915 1.34 45.085 2.195 ;
      RECT 44.815 1.34 45.165 1.69 ;
      RECT 47.275 6.655 47.6 6.98 ;
      RECT 42.705 6.615 43.055 6.965 ;
      RECT 47.25 6.655 47.6 6.885 ;
      RECT 42.47 6.655 43.055 6.885 ;
      RECT 42.3 6.685 47.6 6.855 ;
      RECT 46.475 2.365 46.795 2.685 ;
      RECT 46.445 2.365 46.795 2.595 ;
      RECT 46.275 2.395 46.795 2.565 ;
      RECT 46.475 6.255 46.795 6.545 ;
      RECT 46.445 6.285 46.795 6.515 ;
      RECT 46.275 6.315 46.795 6.485 ;
      RECT 45.42 2.705 45.77 3.055 ;
      RECT 45.42 2.765 45.91 2.935 ;
      RECT 45.425 5.855 45.775 6.205 ;
      RECT 40.67 5.915 40.96 6.145 ;
      RECT 40.67 5.945 45.91 6.115 ;
      RECT 43.11 2.465 43.295 2.675 ;
      RECT 43.1 2.47 43.31 2.668 ;
      RECT 43.1 2.47 43.396 2.645 ;
      RECT 43.1 2.47 43.455 2.62 ;
      RECT 43.1 2.47 43.51 2.6 ;
      RECT 43.1 2.47 43.52 2.588 ;
      RECT 43.1 2.47 43.715 2.527 ;
      RECT 43.1 2.47 43.745 2.51 ;
      RECT 43.1 2.47 43.765 2.5 ;
      RECT 43.645 2.235 43.905 2.495 ;
      RECT 43.63 2.325 43.645 2.542 ;
      RECT 43.165 2.457 43.905 2.495 ;
      RECT 43.616 2.336 43.63 2.548 ;
      RECT 43.205 2.45 43.905 2.495 ;
      RECT 43.53 2.376 43.616 2.567 ;
      RECT 43.455 2.437 43.905 2.495 ;
      RECT 43.525 2.412 43.53 2.584 ;
      RECT 43.51 2.422 43.905 2.495 ;
      RECT 43.52 2.417 43.525 2.586 ;
      RECT 43.815 2.922 43.82 3.014 ;
      RECT 43.81 2.9 43.815 3.031 ;
      RECT 43.805 2.89 43.81 3.043 ;
      RECT 43.795 2.881 43.805 3.053 ;
      RECT 43.79 2.876 43.795 3.061 ;
      RECT 43.785 2.735 43.79 3.064 ;
      RECT 43.751 2.735 43.785 3.075 ;
      RECT 43.665 2.735 43.751 3.11 ;
      RECT 43.585 2.735 43.665 3.158 ;
      RECT 43.556 2.735 43.585 3.182 ;
      RECT 43.47 2.735 43.556 3.188 ;
      RECT 43.465 2.919 43.47 3.193 ;
      RECT 43.43 2.93 43.465 3.196 ;
      RECT 43.405 2.945 43.43 3.2 ;
      RECT 43.391 2.954 43.405 3.202 ;
      RECT 43.305 2.981 43.391 3.208 ;
      RECT 43.24 3.022 43.305 3.217 ;
      RECT 43.225 3.042 43.24 3.222 ;
      RECT 43.195 3.052 43.225 3.225 ;
      RECT 43.19 3.062 43.195 3.228 ;
      RECT 43.16 3.067 43.19 3.23 ;
      RECT 43.14 3.072 43.16 3.234 ;
      RECT 43.055 3.075 43.14 3.241 ;
      RECT 43.04 3.072 43.055 3.247 ;
      RECT 43.03 3.069 43.04 3.249 ;
      RECT 43.01 3.066 43.03 3.251 ;
      RECT 42.99 3.062 43.01 3.252 ;
      RECT 42.975 3.058 42.99 3.254 ;
      RECT 42.965 3.055 42.975 3.255 ;
      RECT 42.925 3.049 42.965 3.253 ;
      RECT 42.915 3.044 42.925 3.251 ;
      RECT 42.9 3.041 42.915 3.247 ;
      RECT 42.875 3.036 42.9 3.24 ;
      RECT 42.825 3.027 42.875 3.228 ;
      RECT 42.755 3.013 42.825 3.21 ;
      RECT 42.697 2.998 42.755 3.192 ;
      RECT 42.611 2.981 42.697 3.172 ;
      RECT 42.525 2.96 42.611 3.147 ;
      RECT 42.475 2.945 42.525 3.128 ;
      RECT 42.471 2.939 42.475 3.12 ;
      RECT 42.385 2.929 42.471 3.107 ;
      RECT 42.35 2.914 42.385 3.09 ;
      RECT 42.335 2.907 42.35 3.083 ;
      RECT 42.275 2.895 42.335 3.071 ;
      RECT 42.255 2.882 42.275 3.059 ;
      RECT 42.215 2.873 42.255 3.051 ;
      RECT 42.21 2.865 42.215 3.044 ;
      RECT 42.13 2.855 42.21 3.03 ;
      RECT 42.115 2.842 42.13 3.015 ;
      RECT 42.11 2.84 42.115 3.013 ;
      RECT 42.031 2.828 42.11 3 ;
      RECT 41.945 2.803 42.031 2.975 ;
      RECT 41.93 2.772 41.945 2.96 ;
      RECT 41.915 2.747 41.93 2.956 ;
      RECT 41.9 2.74 41.915 2.952 ;
      RECT 41.725 2.745 41.73 2.948 ;
      RECT 41.72 2.75 41.725 2.943 ;
      RECT 41.73 2.74 41.9 2.95 ;
      RECT 42.445 2.5 42.55 2.76 ;
      RECT 43.26 2.025 43.265 2.25 ;
      RECT 43.39 2.025 43.445 2.235 ;
      RECT 43.445 2.03 43.455 2.228 ;
      RECT 43.351 2.025 43.39 2.238 ;
      RECT 43.265 2.025 43.351 2.245 ;
      RECT 43.245 2.03 43.26 2.251 ;
      RECT 43.235 2.07 43.245 2.253 ;
      RECT 43.205 2.08 43.235 2.255 ;
      RECT 43.2 2.085 43.205 2.257 ;
      RECT 43.175 2.09 43.2 2.259 ;
      RECT 43.16 2.095 43.175 2.261 ;
      RECT 43.145 2.097 43.16 2.263 ;
      RECT 43.14 2.102 43.145 2.265 ;
      RECT 43.09 2.11 43.14 2.268 ;
      RECT 43.065 2.119 43.09 2.273 ;
      RECT 43.055 2.126 43.065 2.278 ;
      RECT 43.05 2.129 43.055 2.282 ;
      RECT 43.03 2.132 43.05 2.291 ;
      RECT 43 2.14 43.03 2.311 ;
      RECT 42.971 2.153 43 2.333 ;
      RECT 42.885 2.187 42.971 2.377 ;
      RECT 42.88 2.213 42.885 2.415 ;
      RECT 42.875 2.217 42.88 2.424 ;
      RECT 42.84 2.23 42.875 2.457 ;
      RECT 42.83 2.244 42.84 2.495 ;
      RECT 42.825 2.248 42.83 2.508 ;
      RECT 42.82 2.252 42.825 2.513 ;
      RECT 42.81 2.26 42.82 2.525 ;
      RECT 42.805 2.267 42.81 2.54 ;
      RECT 42.78 2.28 42.805 2.565 ;
      RECT 42.74 2.309 42.78 2.62 ;
      RECT 42.725 2.334 42.74 2.675 ;
      RECT 42.715 2.345 42.725 2.698 ;
      RECT 42.71 2.352 42.715 2.71 ;
      RECT 42.705 2.356 42.71 2.718 ;
      RECT 42.65 2.384 42.705 2.76 ;
      RECT 42.63 2.42 42.65 2.76 ;
      RECT 42.615 2.435 42.63 2.76 ;
      RECT 42.56 2.467 42.615 2.76 ;
      RECT 42.55 2.497 42.56 2.76 ;
      RECT 42.16 2.112 42.345 2.35 ;
      RECT 42.145 2.114 42.355 2.345 ;
      RECT 42.03 2.06 42.29 2.32 ;
      RECT 42.025 2.097 42.29 2.274 ;
      RECT 42.02 2.107 42.29 2.271 ;
      RECT 42.015 2.147 42.355 2.265 ;
      RECT 42.01 2.18 42.355 2.255 ;
      RECT 42.02 2.122 42.37 2.193 ;
      RECT 42.317 3.22 42.33 3.75 ;
      RECT 42.231 3.22 42.33 3.749 ;
      RECT 42.231 3.22 42.335 3.748 ;
      RECT 42.145 3.22 42.335 3.746 ;
      RECT 42.14 3.22 42.335 3.743 ;
      RECT 42.14 3.22 42.345 3.741 ;
      RECT 42.135 3.512 42.345 3.738 ;
      RECT 42.135 3.522 42.35 3.735 ;
      RECT 42.135 3.59 42.355 3.731 ;
      RECT 42.125 3.595 42.355 3.73 ;
      RECT 42.125 3.687 42.36 3.727 ;
      RECT 42.11 3.22 42.37 3.48 ;
      RECT 42.04 7.765 42.33 7.995 ;
      RECT 42.1 7.025 42.27 7.995 ;
      RECT 42.015 7.055 42.355 7.4 ;
      RECT 42.04 7.025 42.33 7.4 ;
      RECT 41.34 2.21 41.385 3.745 ;
      RECT 41.54 2.21 41.57 2.425 ;
      RECT 39.915 1.95 40.035 2.16 ;
      RECT 39.575 1.9 39.835 2.16 ;
      RECT 39.575 1.945 39.87 2.15 ;
      RECT 41.58 2.226 41.585 2.28 ;
      RECT 41.575 2.219 41.58 2.413 ;
      RECT 41.57 2.213 41.575 2.42 ;
      RECT 41.525 2.21 41.54 2.433 ;
      RECT 41.52 2.21 41.525 2.455 ;
      RECT 41.515 2.21 41.52 2.503 ;
      RECT 41.51 2.21 41.515 2.523 ;
      RECT 41.5 2.21 41.51 2.63 ;
      RECT 41.495 2.21 41.5 2.693 ;
      RECT 41.49 2.21 41.495 2.75 ;
      RECT 41.485 2.21 41.49 2.758 ;
      RECT 41.47 2.21 41.485 2.865 ;
      RECT 41.46 2.21 41.47 3 ;
      RECT 41.45 2.21 41.46 3.11 ;
      RECT 41.44 2.21 41.45 3.167 ;
      RECT 41.435 2.21 41.44 3.207 ;
      RECT 41.43 2.21 41.435 3.243 ;
      RECT 41.42 2.21 41.43 3.283 ;
      RECT 41.415 2.21 41.42 3.325 ;
      RECT 41.395 2.21 41.415 3.39 ;
      RECT 41.4 3.535 41.405 3.715 ;
      RECT 41.395 3.517 41.4 3.723 ;
      RECT 41.39 2.21 41.395 3.453 ;
      RECT 41.39 3.497 41.395 3.73 ;
      RECT 41.385 2.21 41.39 3.74 ;
      RECT 41.33 2.21 41.34 2.51 ;
      RECT 41.335 2.757 41.34 3.745 ;
      RECT 41.33 2.822 41.335 3.745 ;
      RECT 41.325 2.211 41.33 2.5 ;
      RECT 41.32 2.887 41.33 3.745 ;
      RECT 41.315 2.212 41.325 2.49 ;
      RECT 41.305 3 41.32 3.745 ;
      RECT 41.31 2.213 41.315 2.48 ;
      RECT 41.29 2.214 41.31 2.458 ;
      RECT 41.295 3.097 41.305 3.745 ;
      RECT 41.29 3.172 41.295 3.745 ;
      RECT 41.28 2.213 41.29 2.435 ;
      RECT 41.285 3.215 41.29 3.745 ;
      RECT 41.28 3.242 41.285 3.745 ;
      RECT 41.27 2.211 41.28 2.423 ;
      RECT 41.275 3.285 41.28 3.745 ;
      RECT 41.27 3.312 41.275 3.745 ;
      RECT 41.26 2.21 41.27 2.41 ;
      RECT 41.265 3.327 41.27 3.745 ;
      RECT 41.225 3.385 41.265 3.745 ;
      RECT 41.255 2.209 41.26 2.395 ;
      RECT 41.25 2.207 41.255 2.388 ;
      RECT 41.24 2.204 41.25 2.378 ;
      RECT 41.235 2.201 41.24 2.363 ;
      RECT 41.22 2.197 41.235 2.356 ;
      RECT 41.215 3.44 41.225 3.745 ;
      RECT 41.215 2.194 41.22 2.351 ;
      RECT 41.2 2.19 41.215 2.345 ;
      RECT 41.21 3.457 41.215 3.745 ;
      RECT 41.2 3.52 41.21 3.745 ;
      RECT 41.12 2.175 41.2 2.325 ;
      RECT 41.195 3.527 41.2 3.74 ;
      RECT 41.19 3.535 41.195 3.73 ;
      RECT 41.11 2.161 41.12 2.309 ;
      RECT 41.095 2.157 41.11 2.307 ;
      RECT 41.085 2.152 41.095 2.303 ;
      RECT 41.06 2.145 41.085 2.295 ;
      RECT 41.055 2.14 41.06 2.29 ;
      RECT 41.045 2.14 41.055 2.288 ;
      RECT 41.035 2.138 41.045 2.286 ;
      RECT 41.005 2.13 41.035 2.28 ;
      RECT 40.99 2.122 41.005 2.273 ;
      RECT 40.97 2.117 40.99 2.266 ;
      RECT 40.965 2.113 40.97 2.261 ;
      RECT 40.935 2.106 40.965 2.255 ;
      RECT 40.91 2.097 40.935 2.245 ;
      RECT 40.88 2.09 40.91 2.237 ;
      RECT 40.855 2.08 40.88 2.228 ;
      RECT 40.84 2.072 40.855 2.222 ;
      RECT 40.815 2.067 40.84 2.217 ;
      RECT 40.805 2.063 40.815 2.212 ;
      RECT 40.785 2.058 40.805 2.207 ;
      RECT 40.75 2.053 40.785 2.2 ;
      RECT 40.69 2.048 40.75 2.193 ;
      RECT 40.677 2.044 40.69 2.191 ;
      RECT 40.591 2.039 40.677 2.188 ;
      RECT 40.505 2.029 40.591 2.184 ;
      RECT 40.464 2.022 40.505 2.181 ;
      RECT 40.378 2.015 40.464 2.178 ;
      RECT 40.292 2.005 40.378 2.174 ;
      RECT 40.206 1.995 40.292 2.169 ;
      RECT 40.12 1.985 40.206 2.165 ;
      RECT 40.11 1.97 40.12 2.163 ;
      RECT 40.1 1.955 40.11 2.163 ;
      RECT 40.035 1.95 40.1 2.162 ;
      RECT 39.87 1.947 39.915 2.155 ;
      RECT 41.115 2.852 41.12 3.043 ;
      RECT 41.11 2.847 41.115 3.05 ;
      RECT 41.096 2.845 41.11 3.056 ;
      RECT 41.01 2.845 41.096 3.058 ;
      RECT 41.006 2.845 41.01 3.061 ;
      RECT 40.92 2.845 41.006 3.079 ;
      RECT 40.91 2.85 40.92 3.098 ;
      RECT 40.9 2.905 40.91 3.102 ;
      RECT 40.875 2.92 40.9 3.109 ;
      RECT 40.835 2.94 40.875 3.122 ;
      RECT 40.83 2.952 40.835 3.132 ;
      RECT 40.815 2.958 40.83 3.137 ;
      RECT 40.81 2.963 40.815 3.141 ;
      RECT 40.79 2.97 40.81 3.146 ;
      RECT 40.72 2.995 40.79 3.163 ;
      RECT 40.68 3.023 40.72 3.183 ;
      RECT 40.675 3.033 40.68 3.191 ;
      RECT 40.655 3.04 40.675 3.193 ;
      RECT 40.65 3.047 40.655 3.196 ;
      RECT 40.62 3.055 40.65 3.199 ;
      RECT 40.615 3.06 40.62 3.203 ;
      RECT 40.541 3.064 40.615 3.211 ;
      RECT 40.455 3.073 40.541 3.227 ;
      RECT 40.451 3.078 40.455 3.236 ;
      RECT 40.365 3.083 40.451 3.246 ;
      RECT 40.325 3.091 40.365 3.258 ;
      RECT 40.275 3.097 40.325 3.265 ;
      RECT 40.19 3.106 40.275 3.28 ;
      RECT 40.115 3.117 40.19 3.298 ;
      RECT 40.08 3.124 40.115 3.308 ;
      RECT 40.005 3.132 40.08 3.313 ;
      RECT 39.95 3.141 40.005 3.313 ;
      RECT 39.925 3.146 39.95 3.311 ;
      RECT 39.915 3.149 39.925 3.309 ;
      RECT 39.88 3.151 39.915 3.307 ;
      RECT 39.85 3.153 39.88 3.303 ;
      RECT 39.805 3.152 39.85 3.299 ;
      RECT 39.785 3.147 39.805 3.296 ;
      RECT 39.735 3.132 39.785 3.293 ;
      RECT 39.725 3.117 39.735 3.288 ;
      RECT 39.675 3.102 39.725 3.278 ;
      RECT 39.625 3.077 39.675 3.258 ;
      RECT 39.615 3.062 39.625 3.24 ;
      RECT 39.61 3.06 39.615 3.234 ;
      RECT 39.59 3.055 39.61 3.229 ;
      RECT 39.585 3.047 39.59 3.223 ;
      RECT 39.57 3.041 39.585 3.216 ;
      RECT 39.565 3.036 39.57 3.208 ;
      RECT 39.545 3.031 39.565 3.2 ;
      RECT 39.53 3.024 39.545 3.193 ;
      RECT 39.515 3.018 39.53 3.184 ;
      RECT 39.51 3.012 39.515 3.177 ;
      RECT 39.465 2.987 39.51 3.163 ;
      RECT 39.45 2.957 39.465 3.145 ;
      RECT 39.435 2.94 39.45 3.136 ;
      RECT 39.41 2.92 39.435 3.124 ;
      RECT 39.37 2.89 39.41 3.104 ;
      RECT 39.36 2.86 39.37 3.089 ;
      RECT 39.345 2.85 39.36 3.082 ;
      RECT 39.29 2.815 39.345 3.061 ;
      RECT 39.275 2.778 39.29 3.04 ;
      RECT 39.265 2.765 39.275 3.032 ;
      RECT 39.215 2.735 39.265 3.014 ;
      RECT 39.2 2.665 39.215 2.995 ;
      RECT 39.155 2.665 39.2 2.978 ;
      RECT 39.13 2.665 39.155 2.96 ;
      RECT 39.12 2.665 39.13 2.953 ;
      RECT 39.041 2.665 39.12 2.946 ;
      RECT 38.955 2.665 39.041 2.938 ;
      RECT 38.94 2.697 38.955 2.933 ;
      RECT 38.865 2.707 38.94 2.929 ;
      RECT 38.845 2.717 38.865 2.924 ;
      RECT 38.82 2.717 38.845 2.921 ;
      RECT 38.81 2.707 38.82 2.92 ;
      RECT 38.8 2.68 38.81 2.919 ;
      RECT 38.76 2.675 38.8 2.917 ;
      RECT 38.715 2.675 38.76 2.913 ;
      RECT 38.69 2.675 38.715 2.908 ;
      RECT 38.64 2.675 38.69 2.895 ;
      RECT 38.6 2.68 38.61 2.88 ;
      RECT 38.61 2.675 38.64 2.885 ;
      RECT 40.595 2.455 40.855 2.715 ;
      RECT 40.59 2.477 40.855 2.673 ;
      RECT 39.83 2.305 40.05 2.67 ;
      RECT 39.812 2.392 40.05 2.669 ;
      RECT 39.795 2.397 40.05 2.666 ;
      RECT 39.795 2.397 40.07 2.665 ;
      RECT 39.765 2.407 40.07 2.663 ;
      RECT 39.76 2.422 40.07 2.659 ;
      RECT 39.76 2.422 40.075 2.658 ;
      RECT 39.755 2.48 40.075 2.656 ;
      RECT 39.755 2.48 40.085 2.653 ;
      RECT 39.75 2.545 40.085 2.648 ;
      RECT 39.83 2.305 40.09 2.565 ;
      RECT 38.575 2.135 38.835 2.395 ;
      RECT 38.575 2.178 38.921 2.369 ;
      RECT 38.575 2.178 38.965 2.368 ;
      RECT 38.575 2.178 38.985 2.366 ;
      RECT 38.575 2.178 39.085 2.365 ;
      RECT 38.575 2.178 39.105 2.363 ;
      RECT 38.575 2.178 39.115 2.358 ;
      RECT 38.985 2.145 39.175 2.355 ;
      RECT 38.985 2.147 39.18 2.353 ;
      RECT 38.975 2.152 39.185 2.345 ;
      RECT 38.921 2.176 39.185 2.345 ;
      RECT 38.965 2.17 38.975 2.367 ;
      RECT 38.975 2.15 39.18 2.353 ;
      RECT 37.93 3.21 38.135 3.44 ;
      RECT 37.87 3.16 37.925 3.42 ;
      RECT 37.93 3.16 38.13 3.44 ;
      RECT 38.9 3.475 38.905 3.502 ;
      RECT 38.89 3.385 38.9 3.507 ;
      RECT 38.885 3.307 38.89 3.513 ;
      RECT 38.875 3.297 38.885 3.52 ;
      RECT 38.87 3.287 38.875 3.526 ;
      RECT 38.86 3.282 38.87 3.528 ;
      RECT 38.845 3.274 38.86 3.536 ;
      RECT 38.83 3.265 38.845 3.548 ;
      RECT 38.82 3.257 38.83 3.558 ;
      RECT 38.785 3.175 38.82 3.576 ;
      RECT 38.75 3.175 38.785 3.595 ;
      RECT 38.735 3.175 38.75 3.603 ;
      RECT 38.68 3.175 38.735 3.603 ;
      RECT 38.646 3.175 38.68 3.594 ;
      RECT 38.56 3.175 38.646 3.57 ;
      RECT 38.55 3.235 38.56 3.552 ;
      RECT 38.51 3.237 38.55 3.543 ;
      RECT 38.505 3.239 38.51 3.533 ;
      RECT 38.485 3.241 38.505 3.528 ;
      RECT 38.475 3.244 38.485 3.523 ;
      RECT 38.465 3.245 38.475 3.518 ;
      RECT 38.441 3.246 38.465 3.51 ;
      RECT 38.355 3.251 38.441 3.488 ;
      RECT 38.3 3.25 38.355 3.461 ;
      RECT 38.285 3.243 38.3 3.448 ;
      RECT 38.25 3.238 38.285 3.444 ;
      RECT 38.195 3.23 38.25 3.443 ;
      RECT 38.135 3.217 38.195 3.441 ;
      RECT 37.925 3.16 37.93 3.428 ;
      RECT 38 2.53 38.185 2.74 ;
      RECT 37.99 2.535 38.2 2.733 ;
      RECT 38.03 2.44 38.29 2.7 ;
      RECT 37.985 2.597 38.29 2.623 ;
      RECT 37.33 2.39 37.335 3.19 ;
      RECT 37.275 2.44 37.305 3.19 ;
      RECT 37.265 2.44 37.27 2.75 ;
      RECT 37.25 2.44 37.255 2.745 ;
      RECT 36.795 2.485 36.81 2.7 ;
      RECT 36.725 2.485 36.81 2.695 ;
      RECT 37.99 2.065 38.06 2.275 ;
      RECT 38.06 2.072 38.07 2.27 ;
      RECT 37.956 2.065 37.99 2.282 ;
      RECT 37.87 2.065 37.956 2.306 ;
      RECT 37.86 2.07 37.87 2.325 ;
      RECT 37.855 2.082 37.86 2.328 ;
      RECT 37.84 2.097 37.855 2.332 ;
      RECT 37.835 2.115 37.84 2.336 ;
      RECT 37.795 2.125 37.835 2.345 ;
      RECT 37.78 2.132 37.795 2.357 ;
      RECT 37.765 2.137 37.78 2.362 ;
      RECT 37.75 2.14 37.765 2.367 ;
      RECT 37.74 2.142 37.75 2.371 ;
      RECT 37.705 2.149 37.74 2.379 ;
      RECT 37.67 2.157 37.705 2.393 ;
      RECT 37.66 2.163 37.67 2.402 ;
      RECT 37.655 2.165 37.66 2.404 ;
      RECT 37.635 2.168 37.655 2.41 ;
      RECT 37.605 2.175 37.635 2.421 ;
      RECT 37.595 2.181 37.605 2.428 ;
      RECT 37.57 2.184 37.595 2.435 ;
      RECT 37.56 2.188 37.57 2.443 ;
      RECT 37.555 2.189 37.56 2.465 ;
      RECT 37.55 2.19 37.555 2.48 ;
      RECT 37.545 2.191 37.55 2.495 ;
      RECT 37.54 2.192 37.545 2.51 ;
      RECT 37.535 2.193 37.54 2.54 ;
      RECT 37.525 2.195 37.535 2.573 ;
      RECT 37.51 2.199 37.525 2.62 ;
      RECT 37.5 2.202 37.51 2.665 ;
      RECT 37.495 2.205 37.5 2.693 ;
      RECT 37.485 2.207 37.495 2.72 ;
      RECT 37.48 2.21 37.485 2.755 ;
      RECT 37.45 2.215 37.48 2.813 ;
      RECT 37.445 2.22 37.45 2.898 ;
      RECT 37.44 2.222 37.445 2.933 ;
      RECT 37.435 2.224 37.44 3.015 ;
      RECT 37.43 2.226 37.435 3.103 ;
      RECT 37.42 2.228 37.43 3.185 ;
      RECT 37.405 2.242 37.42 3.19 ;
      RECT 37.37 2.287 37.405 3.19 ;
      RECT 37.36 2.327 37.37 3.19 ;
      RECT 37.345 2.355 37.36 3.19 ;
      RECT 37.34 2.372 37.345 3.19 ;
      RECT 37.335 2.38 37.34 3.19 ;
      RECT 37.325 2.395 37.33 3.19 ;
      RECT 37.32 2.402 37.325 3.19 ;
      RECT 37.31 2.422 37.32 3.19 ;
      RECT 37.305 2.435 37.31 3.19 ;
      RECT 37.27 2.44 37.275 2.775 ;
      RECT 37.255 2.83 37.275 3.19 ;
      RECT 37.255 2.44 37.265 2.748 ;
      RECT 37.25 2.87 37.255 3.19 ;
      RECT 37.2 2.44 37.25 2.743 ;
      RECT 37.245 2.907 37.25 3.19 ;
      RECT 37.235 2.93 37.245 3.19 ;
      RECT 37.23 2.975 37.235 3.19 ;
      RECT 37.22 2.985 37.23 3.183 ;
      RECT 37.146 2.44 37.2 2.737 ;
      RECT 37.06 2.44 37.146 2.73 ;
      RECT 37.011 2.487 37.06 2.723 ;
      RECT 36.925 2.495 37.011 2.716 ;
      RECT 36.91 2.492 36.925 2.711 ;
      RECT 36.896 2.485 36.91 2.71 ;
      RECT 36.81 2.485 36.896 2.705 ;
      RECT 36.715 2.49 36.725 2.69 ;
      RECT 36.305 1.92 36.32 2.32 ;
      RECT 36.5 1.92 36.505 2.18 ;
      RECT 36.245 1.92 36.29 2.18 ;
      RECT 36.7 3.225 36.705 3.43 ;
      RECT 36.695 3.215 36.7 3.435 ;
      RECT 36.69 3.202 36.695 3.44 ;
      RECT 36.685 3.182 36.69 3.44 ;
      RECT 36.66 3.135 36.685 3.44 ;
      RECT 36.625 3.05 36.66 3.44 ;
      RECT 36.62 2.987 36.625 3.44 ;
      RECT 36.615 2.972 36.62 3.44 ;
      RECT 36.6 2.932 36.615 3.44 ;
      RECT 36.595 2.907 36.6 3.44 ;
      RECT 36.585 2.89 36.595 3.44 ;
      RECT 36.55 2.812 36.585 3.44 ;
      RECT 36.545 2.755 36.55 3.44 ;
      RECT 36.54 2.742 36.545 3.44 ;
      RECT 36.53 2.72 36.54 3.44 ;
      RECT 36.52 2.685 36.53 3.44 ;
      RECT 36.51 2.655 36.52 3.44 ;
      RECT 36.5 2.57 36.51 3.083 ;
      RECT 36.507 3.215 36.51 3.44 ;
      RECT 36.505 3.225 36.507 3.44 ;
      RECT 36.495 3.235 36.505 3.435 ;
      RECT 36.49 1.92 36.5 2.315 ;
      RECT 36.495 2.447 36.5 3.058 ;
      RECT 36.49 2.345 36.495 3.041 ;
      RECT 36.48 1.92 36.49 3.017 ;
      RECT 36.475 1.92 36.48 2.988 ;
      RECT 36.47 1.92 36.475 2.978 ;
      RECT 36.45 1.92 36.47 2.94 ;
      RECT 36.445 1.92 36.45 2.898 ;
      RECT 36.44 1.92 36.445 2.878 ;
      RECT 36.41 1.92 36.44 2.828 ;
      RECT 36.4 1.92 36.41 2.775 ;
      RECT 36.395 1.92 36.4 2.748 ;
      RECT 36.39 1.92 36.395 2.733 ;
      RECT 36.38 1.92 36.39 2.71 ;
      RECT 36.37 1.92 36.38 2.685 ;
      RECT 36.365 1.92 36.37 2.625 ;
      RECT 36.355 1.92 36.365 2.563 ;
      RECT 36.35 1.92 36.355 2.483 ;
      RECT 36.345 1.92 36.35 2.448 ;
      RECT 36.34 1.92 36.345 2.423 ;
      RECT 36.335 1.92 36.34 2.408 ;
      RECT 36.33 1.92 36.335 2.378 ;
      RECT 36.325 1.92 36.33 2.355 ;
      RECT 36.32 1.92 36.325 2.328 ;
      RECT 36.29 1.92 36.305 2.315 ;
      RECT 35.445 3.455 35.63 3.665 ;
      RECT 35.435 3.46 35.645 3.658 ;
      RECT 35.435 3.46 35.665 3.63 ;
      RECT 35.435 3.46 35.68 3.609 ;
      RECT 35.435 3.46 35.695 3.607 ;
      RECT 35.435 3.46 35.705 3.606 ;
      RECT 35.435 3.46 35.735 3.603 ;
      RECT 36.085 3.305 36.345 3.565 ;
      RECT 36.045 3.352 36.345 3.548 ;
      RECT 36.036 3.36 36.045 3.551 ;
      RECT 35.63 3.453 36.345 3.548 ;
      RECT 35.95 3.378 36.036 3.558 ;
      RECT 35.645 3.45 36.345 3.548 ;
      RECT 35.891 3.4 35.95 3.57 ;
      RECT 35.665 3.446 36.345 3.548 ;
      RECT 35.805 3.412 35.891 3.581 ;
      RECT 35.68 3.442 36.345 3.548 ;
      RECT 35.75 3.425 35.805 3.593 ;
      RECT 35.695 3.44 36.345 3.548 ;
      RECT 35.735 3.431 35.75 3.599 ;
      RECT 35.705 3.436 36.345 3.548 ;
      RECT 35.85 2.96 36.11 3.22 ;
      RECT 35.85 2.98 36.22 3.19 ;
      RECT 35.85 2.985 36.23 3.185 ;
      RECT 36.041 2.399 36.12 2.63 ;
      RECT 35.955 2.402 36.17 2.625 ;
      RECT 35.95 2.402 36.17 2.62 ;
      RECT 35.95 2.407 36.18 2.618 ;
      RECT 35.925 2.407 36.18 2.615 ;
      RECT 35.925 2.415 36.19 2.613 ;
      RECT 35.805 2.35 36.065 2.61 ;
      RECT 35.805 2.397 36.115 2.61 ;
      RECT 35.06 2.97 35.065 3.23 ;
      RECT 34.89 2.74 34.895 3.23 ;
      RECT 34.775 2.98 34.78 3.205 ;
      RECT 35.485 2.075 35.49 2.285 ;
      RECT 35.49 2.08 35.505 2.28 ;
      RECT 35.425 2.075 35.485 2.293 ;
      RECT 35.41 2.075 35.425 2.303 ;
      RECT 35.36 2.075 35.41 2.32 ;
      RECT 35.34 2.075 35.36 2.343 ;
      RECT 35.325 2.075 35.34 2.355 ;
      RECT 35.305 2.075 35.325 2.365 ;
      RECT 35.295 2.08 35.305 2.374 ;
      RECT 35.29 2.09 35.295 2.379 ;
      RECT 35.285 2.102 35.29 2.383 ;
      RECT 35.275 2.125 35.285 2.388 ;
      RECT 35.27 2.14 35.275 2.392 ;
      RECT 35.265 2.157 35.27 2.395 ;
      RECT 35.26 2.165 35.265 2.398 ;
      RECT 35.25 2.17 35.26 2.402 ;
      RECT 35.245 2.177 35.25 2.407 ;
      RECT 35.235 2.182 35.245 2.411 ;
      RECT 35.21 2.194 35.235 2.422 ;
      RECT 35.19 2.211 35.21 2.438 ;
      RECT 35.165 2.228 35.19 2.46 ;
      RECT 35.13 2.251 35.165 2.518 ;
      RECT 35.11 2.273 35.13 2.58 ;
      RECT 35.105 2.283 35.11 2.615 ;
      RECT 35.095 2.29 35.105 2.653 ;
      RECT 35.09 2.297 35.095 2.673 ;
      RECT 35.085 2.308 35.09 2.71 ;
      RECT 35.08 2.316 35.085 2.775 ;
      RECT 35.07 2.327 35.08 2.828 ;
      RECT 35.065 2.345 35.07 2.898 ;
      RECT 35.06 2.355 35.065 2.935 ;
      RECT 35.055 2.365 35.06 3.23 ;
      RECT 35.05 2.377 35.055 3.23 ;
      RECT 35.045 2.387 35.05 3.23 ;
      RECT 35.035 2.397 35.045 3.23 ;
      RECT 35.025 2.42 35.035 3.23 ;
      RECT 35.01 2.455 35.025 3.23 ;
      RECT 34.97 2.517 35.01 3.23 ;
      RECT 34.965 2.57 34.97 3.23 ;
      RECT 34.94 2.605 34.965 3.23 ;
      RECT 34.925 2.65 34.94 3.23 ;
      RECT 34.92 2.672 34.925 3.23 ;
      RECT 34.91 2.685 34.92 3.23 ;
      RECT 34.9 2.71 34.91 3.23 ;
      RECT 34.895 2.732 34.9 3.23 ;
      RECT 34.87 2.77 34.89 3.23 ;
      RECT 34.83 2.827 34.87 3.23 ;
      RECT 34.825 2.877 34.83 3.23 ;
      RECT 34.82 2.895 34.825 3.23 ;
      RECT 34.815 2.907 34.82 3.23 ;
      RECT 34.805 2.925 34.815 3.23 ;
      RECT 34.795 2.945 34.805 3.205 ;
      RECT 34.79 2.962 34.795 3.205 ;
      RECT 34.78 2.975 34.79 3.205 ;
      RECT 34.75 2.985 34.775 3.205 ;
      RECT 34.74 2.992 34.75 3.205 ;
      RECT 34.725 3.002 34.74 3.2 ;
      RECT 33.83 7.765 34.12 7.995 ;
      RECT 33.89 6.285 34.06 7.995 ;
      RECT 33.875 6.66 34.23 7.015 ;
      RECT 33.83 6.285 34.12 6.515 ;
      RECT 33.83 2.365 34.12 2.595 ;
      RECT 33.89 0.885 34.06 2.595 ;
      RECT 33.83 0.885 34.12 1.115 ;
      RECT 33.42 2.735 33.75 2.965 ;
      RECT 33.42 2.765 33.92 2.935 ;
      RECT 33.42 2.395 33.61 2.965 ;
      RECT 32.84 2.365 33.13 2.595 ;
      RECT 32.84 2.395 33.61 2.565 ;
      RECT 32.9 0.885 33.07 2.595 ;
      RECT 32.84 0.885 33.13 1.115 ;
      RECT 32.84 7.765 33.13 7.995 ;
      RECT 32.9 6.285 33.07 7.995 ;
      RECT 32.84 6.285 33.13 6.515 ;
      RECT 32.84 6.325 33.69 6.485 ;
      RECT 33.52 5.915 33.69 6.485 ;
      RECT 32.84 6.32 33.23 6.485 ;
      RECT 33.46 5.915 33.75 6.145 ;
      RECT 33.46 5.945 33.92 6.115 ;
      RECT 32.47 2.735 32.76 2.965 ;
      RECT 32.47 2.765 32.93 2.935 ;
      RECT 32.53 1.655 32.695 2.965 ;
      RECT 31.045 1.625 31.335 1.855 ;
      RECT 31.045 1.655 32.695 1.825 ;
      RECT 31.105 0.885 31.275 1.855 ;
      RECT 31.045 0.885 31.335 1.115 ;
      RECT 31.045 7.765 31.335 7.995 ;
      RECT 31.105 7.025 31.275 7.995 ;
      RECT 31.105 7.12 32.695 7.29 ;
      RECT 32.525 5.915 32.695 7.29 ;
      RECT 31.045 7.025 31.335 7.255 ;
      RECT 32.47 5.915 32.76 6.145 ;
      RECT 32.47 5.945 32.93 6.115 ;
      RECT 31.475 1.965 31.825 2.315 ;
      RECT 29.14 2.025 31.825 2.195 ;
      RECT 29.14 1.34 29.31 2.195 ;
      RECT 29.04 1.34 29.39 1.69 ;
      RECT 31.5 6.655 31.825 6.98 ;
      RECT 26.925 6.61 27.275 6.96 ;
      RECT 31.475 6.655 31.825 6.885 ;
      RECT 26.695 6.655 27.275 6.885 ;
      RECT 26.525 6.685 31.825 6.855 ;
      RECT 30.7 2.365 31.02 2.685 ;
      RECT 30.67 2.365 31.02 2.595 ;
      RECT 30.5 2.395 31.02 2.565 ;
      RECT 30.7 6.255 31.02 6.545 ;
      RECT 30.67 6.285 31.02 6.515 ;
      RECT 30.5 6.315 31.02 6.485 ;
      RECT 29.645 2.705 29.995 3.055 ;
      RECT 29.645 2.765 30.135 2.935 ;
      RECT 29.65 5.855 30 6.205 ;
      RECT 24.895 5.915 25.185 6.145 ;
      RECT 24.895 5.945 30.135 6.115 ;
      RECT 27.335 2.465 27.52 2.675 ;
      RECT 27.325 2.47 27.535 2.668 ;
      RECT 27.325 2.47 27.621 2.645 ;
      RECT 27.325 2.47 27.68 2.62 ;
      RECT 27.325 2.47 27.735 2.6 ;
      RECT 27.325 2.47 27.745 2.588 ;
      RECT 27.325 2.47 27.94 2.527 ;
      RECT 27.325 2.47 27.97 2.51 ;
      RECT 27.325 2.47 27.99 2.5 ;
      RECT 27.87 2.235 28.13 2.495 ;
      RECT 27.855 2.325 27.87 2.542 ;
      RECT 27.39 2.457 28.13 2.495 ;
      RECT 27.841 2.336 27.855 2.548 ;
      RECT 27.43 2.45 28.13 2.495 ;
      RECT 27.755 2.376 27.841 2.567 ;
      RECT 27.68 2.437 28.13 2.495 ;
      RECT 27.75 2.412 27.755 2.584 ;
      RECT 27.735 2.422 28.13 2.495 ;
      RECT 27.745 2.417 27.75 2.586 ;
      RECT 28.04 2.922 28.045 3.014 ;
      RECT 28.035 2.9 28.04 3.031 ;
      RECT 28.03 2.89 28.035 3.043 ;
      RECT 28.02 2.881 28.03 3.053 ;
      RECT 28.015 2.876 28.02 3.061 ;
      RECT 28.01 2.735 28.015 3.064 ;
      RECT 27.976 2.735 28.01 3.075 ;
      RECT 27.89 2.735 27.976 3.11 ;
      RECT 27.81 2.735 27.89 3.158 ;
      RECT 27.781 2.735 27.81 3.182 ;
      RECT 27.695 2.735 27.781 3.188 ;
      RECT 27.69 2.919 27.695 3.193 ;
      RECT 27.655 2.93 27.69 3.196 ;
      RECT 27.63 2.945 27.655 3.2 ;
      RECT 27.616 2.954 27.63 3.202 ;
      RECT 27.53 2.981 27.616 3.208 ;
      RECT 27.465 3.022 27.53 3.217 ;
      RECT 27.45 3.042 27.465 3.222 ;
      RECT 27.42 3.052 27.45 3.225 ;
      RECT 27.415 3.062 27.42 3.228 ;
      RECT 27.385 3.067 27.415 3.23 ;
      RECT 27.365 3.072 27.385 3.234 ;
      RECT 27.28 3.075 27.365 3.241 ;
      RECT 27.265 3.072 27.28 3.247 ;
      RECT 27.255 3.069 27.265 3.249 ;
      RECT 27.235 3.066 27.255 3.251 ;
      RECT 27.215 3.062 27.235 3.252 ;
      RECT 27.2 3.058 27.215 3.254 ;
      RECT 27.19 3.055 27.2 3.255 ;
      RECT 27.15 3.049 27.19 3.253 ;
      RECT 27.14 3.044 27.15 3.251 ;
      RECT 27.125 3.041 27.14 3.247 ;
      RECT 27.1 3.036 27.125 3.24 ;
      RECT 27.05 3.027 27.1 3.228 ;
      RECT 26.98 3.013 27.05 3.21 ;
      RECT 26.922 2.998 26.98 3.192 ;
      RECT 26.836 2.981 26.922 3.172 ;
      RECT 26.75 2.96 26.836 3.147 ;
      RECT 26.7 2.945 26.75 3.128 ;
      RECT 26.696 2.939 26.7 3.12 ;
      RECT 26.61 2.929 26.696 3.107 ;
      RECT 26.575 2.914 26.61 3.09 ;
      RECT 26.56 2.907 26.575 3.083 ;
      RECT 26.5 2.895 26.56 3.071 ;
      RECT 26.48 2.882 26.5 3.059 ;
      RECT 26.44 2.873 26.48 3.051 ;
      RECT 26.435 2.865 26.44 3.044 ;
      RECT 26.355 2.855 26.435 3.03 ;
      RECT 26.34 2.842 26.355 3.015 ;
      RECT 26.335 2.84 26.34 3.013 ;
      RECT 26.256 2.828 26.335 3 ;
      RECT 26.17 2.803 26.256 2.975 ;
      RECT 26.155 2.772 26.17 2.96 ;
      RECT 26.14 2.747 26.155 2.956 ;
      RECT 26.125 2.74 26.14 2.952 ;
      RECT 25.95 2.745 25.955 2.948 ;
      RECT 25.945 2.75 25.95 2.943 ;
      RECT 25.955 2.74 26.125 2.95 ;
      RECT 26.67 2.5 26.775 2.76 ;
      RECT 27.485 2.025 27.49 2.25 ;
      RECT 27.615 2.025 27.67 2.235 ;
      RECT 27.67 2.03 27.68 2.228 ;
      RECT 27.576 2.025 27.615 2.238 ;
      RECT 27.49 2.025 27.576 2.245 ;
      RECT 27.47 2.03 27.485 2.251 ;
      RECT 27.46 2.07 27.47 2.253 ;
      RECT 27.43 2.08 27.46 2.255 ;
      RECT 27.425 2.085 27.43 2.257 ;
      RECT 27.4 2.09 27.425 2.259 ;
      RECT 27.385 2.095 27.4 2.261 ;
      RECT 27.37 2.097 27.385 2.263 ;
      RECT 27.365 2.102 27.37 2.265 ;
      RECT 27.315 2.11 27.365 2.268 ;
      RECT 27.29 2.119 27.315 2.273 ;
      RECT 27.28 2.126 27.29 2.278 ;
      RECT 27.275 2.129 27.28 2.282 ;
      RECT 27.255 2.132 27.275 2.291 ;
      RECT 27.225 2.14 27.255 2.311 ;
      RECT 27.196 2.153 27.225 2.333 ;
      RECT 27.11 2.187 27.196 2.377 ;
      RECT 27.105 2.213 27.11 2.415 ;
      RECT 27.1 2.217 27.105 2.424 ;
      RECT 27.065 2.23 27.1 2.457 ;
      RECT 27.055 2.244 27.065 2.495 ;
      RECT 27.05 2.248 27.055 2.508 ;
      RECT 27.045 2.252 27.05 2.513 ;
      RECT 27.035 2.26 27.045 2.525 ;
      RECT 27.03 2.267 27.035 2.54 ;
      RECT 27.005 2.28 27.03 2.565 ;
      RECT 26.965 2.309 27.005 2.62 ;
      RECT 26.95 2.334 26.965 2.675 ;
      RECT 26.94 2.345 26.95 2.698 ;
      RECT 26.935 2.352 26.94 2.71 ;
      RECT 26.93 2.356 26.935 2.718 ;
      RECT 26.875 2.384 26.93 2.76 ;
      RECT 26.855 2.42 26.875 2.76 ;
      RECT 26.84 2.435 26.855 2.76 ;
      RECT 26.785 2.467 26.84 2.76 ;
      RECT 26.775 2.497 26.785 2.76 ;
      RECT 26.385 2.112 26.57 2.35 ;
      RECT 26.37 2.114 26.58 2.345 ;
      RECT 26.255 2.06 26.515 2.32 ;
      RECT 26.25 2.097 26.515 2.274 ;
      RECT 26.245 2.107 26.515 2.271 ;
      RECT 26.24 2.147 26.58 2.265 ;
      RECT 26.235 2.18 26.58 2.255 ;
      RECT 26.245 2.122 26.595 2.193 ;
      RECT 26.542 3.22 26.555 3.75 ;
      RECT 26.456 3.22 26.555 3.749 ;
      RECT 26.456 3.22 26.56 3.748 ;
      RECT 26.37 3.22 26.56 3.746 ;
      RECT 26.365 3.22 26.56 3.743 ;
      RECT 26.365 3.22 26.57 3.741 ;
      RECT 26.36 3.512 26.57 3.738 ;
      RECT 26.36 3.522 26.575 3.735 ;
      RECT 26.36 3.59 26.58 3.731 ;
      RECT 26.35 3.595 26.58 3.73 ;
      RECT 26.35 3.687 26.585 3.727 ;
      RECT 26.335 3.22 26.595 3.48 ;
      RECT 26.265 7.765 26.555 7.995 ;
      RECT 26.325 7.025 26.495 7.995 ;
      RECT 26.24 7.055 26.58 7.4 ;
      RECT 26.265 7.025 26.555 7.4 ;
      RECT 25.565 2.21 25.61 3.745 ;
      RECT 25.765 2.21 25.795 2.425 ;
      RECT 24.14 1.95 24.26 2.16 ;
      RECT 23.8 1.9 24.06 2.16 ;
      RECT 23.8 1.945 24.095 2.15 ;
      RECT 25.805 2.226 25.81 2.28 ;
      RECT 25.8 2.219 25.805 2.413 ;
      RECT 25.795 2.213 25.8 2.42 ;
      RECT 25.75 2.21 25.765 2.433 ;
      RECT 25.745 2.21 25.75 2.455 ;
      RECT 25.74 2.21 25.745 2.503 ;
      RECT 25.735 2.21 25.74 2.523 ;
      RECT 25.725 2.21 25.735 2.63 ;
      RECT 25.72 2.21 25.725 2.693 ;
      RECT 25.715 2.21 25.72 2.75 ;
      RECT 25.71 2.21 25.715 2.758 ;
      RECT 25.695 2.21 25.71 2.865 ;
      RECT 25.685 2.21 25.695 3 ;
      RECT 25.675 2.21 25.685 3.11 ;
      RECT 25.665 2.21 25.675 3.167 ;
      RECT 25.66 2.21 25.665 3.207 ;
      RECT 25.655 2.21 25.66 3.243 ;
      RECT 25.645 2.21 25.655 3.283 ;
      RECT 25.64 2.21 25.645 3.325 ;
      RECT 25.62 2.21 25.64 3.39 ;
      RECT 25.625 3.535 25.63 3.715 ;
      RECT 25.62 3.517 25.625 3.723 ;
      RECT 25.615 2.21 25.62 3.453 ;
      RECT 25.615 3.497 25.62 3.73 ;
      RECT 25.61 2.21 25.615 3.74 ;
      RECT 25.555 2.21 25.565 2.51 ;
      RECT 25.56 2.757 25.565 3.745 ;
      RECT 25.555 2.822 25.56 3.745 ;
      RECT 25.55 2.211 25.555 2.5 ;
      RECT 25.545 2.887 25.555 3.745 ;
      RECT 25.54 2.212 25.55 2.49 ;
      RECT 25.53 3 25.545 3.745 ;
      RECT 25.535 2.213 25.54 2.48 ;
      RECT 25.515 2.214 25.535 2.458 ;
      RECT 25.52 3.097 25.53 3.745 ;
      RECT 25.515 3.172 25.52 3.745 ;
      RECT 25.505 2.213 25.515 2.435 ;
      RECT 25.51 3.215 25.515 3.745 ;
      RECT 25.505 3.242 25.51 3.745 ;
      RECT 25.495 2.211 25.505 2.423 ;
      RECT 25.5 3.285 25.505 3.745 ;
      RECT 25.495 3.312 25.5 3.745 ;
      RECT 25.485 2.21 25.495 2.41 ;
      RECT 25.49 3.327 25.495 3.745 ;
      RECT 25.45 3.385 25.49 3.745 ;
      RECT 25.48 2.209 25.485 2.395 ;
      RECT 25.475 2.207 25.48 2.388 ;
      RECT 25.465 2.204 25.475 2.378 ;
      RECT 25.46 2.201 25.465 2.363 ;
      RECT 25.445 2.197 25.46 2.356 ;
      RECT 25.44 3.44 25.45 3.745 ;
      RECT 25.44 2.194 25.445 2.351 ;
      RECT 25.425 2.19 25.44 2.345 ;
      RECT 25.435 3.457 25.44 3.745 ;
      RECT 25.425 3.52 25.435 3.745 ;
      RECT 25.345 2.175 25.425 2.325 ;
      RECT 25.42 3.527 25.425 3.74 ;
      RECT 25.415 3.535 25.42 3.73 ;
      RECT 25.335 2.161 25.345 2.309 ;
      RECT 25.32 2.157 25.335 2.307 ;
      RECT 25.31 2.152 25.32 2.303 ;
      RECT 25.285 2.145 25.31 2.295 ;
      RECT 25.28 2.14 25.285 2.29 ;
      RECT 25.27 2.14 25.28 2.288 ;
      RECT 25.26 2.138 25.27 2.286 ;
      RECT 25.23 2.13 25.26 2.28 ;
      RECT 25.215 2.122 25.23 2.273 ;
      RECT 25.195 2.117 25.215 2.266 ;
      RECT 25.19 2.113 25.195 2.261 ;
      RECT 25.16 2.106 25.19 2.255 ;
      RECT 25.135 2.097 25.16 2.245 ;
      RECT 25.105 2.09 25.135 2.237 ;
      RECT 25.08 2.08 25.105 2.228 ;
      RECT 25.065 2.072 25.08 2.222 ;
      RECT 25.04 2.067 25.065 2.217 ;
      RECT 25.03 2.063 25.04 2.212 ;
      RECT 25.01 2.058 25.03 2.207 ;
      RECT 24.975 2.053 25.01 2.2 ;
      RECT 24.915 2.048 24.975 2.193 ;
      RECT 24.902 2.044 24.915 2.191 ;
      RECT 24.816 2.039 24.902 2.188 ;
      RECT 24.73 2.029 24.816 2.184 ;
      RECT 24.689 2.022 24.73 2.181 ;
      RECT 24.603 2.015 24.689 2.178 ;
      RECT 24.517 2.005 24.603 2.174 ;
      RECT 24.431 1.995 24.517 2.169 ;
      RECT 24.345 1.985 24.431 2.165 ;
      RECT 24.335 1.97 24.345 2.163 ;
      RECT 24.325 1.955 24.335 2.163 ;
      RECT 24.26 1.95 24.325 2.162 ;
      RECT 24.095 1.947 24.14 2.155 ;
      RECT 25.34 2.852 25.345 3.043 ;
      RECT 25.335 2.847 25.34 3.05 ;
      RECT 25.321 2.845 25.335 3.056 ;
      RECT 25.235 2.845 25.321 3.058 ;
      RECT 25.231 2.845 25.235 3.061 ;
      RECT 25.145 2.845 25.231 3.079 ;
      RECT 25.135 2.85 25.145 3.098 ;
      RECT 25.125 2.905 25.135 3.102 ;
      RECT 25.1 2.92 25.125 3.109 ;
      RECT 25.06 2.94 25.1 3.122 ;
      RECT 25.055 2.952 25.06 3.132 ;
      RECT 25.04 2.958 25.055 3.137 ;
      RECT 25.035 2.963 25.04 3.141 ;
      RECT 25.015 2.97 25.035 3.146 ;
      RECT 24.945 2.995 25.015 3.163 ;
      RECT 24.905 3.023 24.945 3.183 ;
      RECT 24.9 3.033 24.905 3.191 ;
      RECT 24.88 3.04 24.9 3.193 ;
      RECT 24.875 3.047 24.88 3.196 ;
      RECT 24.845 3.055 24.875 3.199 ;
      RECT 24.84 3.06 24.845 3.203 ;
      RECT 24.766 3.064 24.84 3.211 ;
      RECT 24.68 3.073 24.766 3.227 ;
      RECT 24.676 3.078 24.68 3.236 ;
      RECT 24.59 3.083 24.676 3.246 ;
      RECT 24.55 3.091 24.59 3.258 ;
      RECT 24.5 3.097 24.55 3.265 ;
      RECT 24.415 3.106 24.5 3.28 ;
      RECT 24.34 3.117 24.415 3.298 ;
      RECT 24.305 3.124 24.34 3.308 ;
      RECT 24.23 3.132 24.305 3.313 ;
      RECT 24.175 3.141 24.23 3.313 ;
      RECT 24.15 3.146 24.175 3.311 ;
      RECT 24.14 3.149 24.15 3.309 ;
      RECT 24.105 3.151 24.14 3.307 ;
      RECT 24.075 3.153 24.105 3.303 ;
      RECT 24.03 3.152 24.075 3.299 ;
      RECT 24.01 3.147 24.03 3.296 ;
      RECT 23.96 3.132 24.01 3.293 ;
      RECT 23.95 3.117 23.96 3.288 ;
      RECT 23.9 3.102 23.95 3.278 ;
      RECT 23.85 3.077 23.9 3.258 ;
      RECT 23.84 3.062 23.85 3.24 ;
      RECT 23.835 3.06 23.84 3.234 ;
      RECT 23.815 3.055 23.835 3.229 ;
      RECT 23.81 3.047 23.815 3.223 ;
      RECT 23.795 3.041 23.81 3.216 ;
      RECT 23.79 3.036 23.795 3.208 ;
      RECT 23.77 3.031 23.79 3.2 ;
      RECT 23.755 3.024 23.77 3.193 ;
      RECT 23.74 3.018 23.755 3.184 ;
      RECT 23.735 3.012 23.74 3.177 ;
      RECT 23.69 2.987 23.735 3.163 ;
      RECT 23.675 2.957 23.69 3.145 ;
      RECT 23.66 2.94 23.675 3.136 ;
      RECT 23.635 2.92 23.66 3.124 ;
      RECT 23.595 2.89 23.635 3.104 ;
      RECT 23.585 2.86 23.595 3.089 ;
      RECT 23.57 2.85 23.585 3.082 ;
      RECT 23.515 2.815 23.57 3.061 ;
      RECT 23.5 2.778 23.515 3.04 ;
      RECT 23.49 2.765 23.5 3.032 ;
      RECT 23.44 2.735 23.49 3.014 ;
      RECT 23.425 2.665 23.44 2.995 ;
      RECT 23.38 2.665 23.425 2.978 ;
      RECT 23.355 2.665 23.38 2.96 ;
      RECT 23.345 2.665 23.355 2.953 ;
      RECT 23.266 2.665 23.345 2.946 ;
      RECT 23.18 2.665 23.266 2.938 ;
      RECT 23.165 2.697 23.18 2.933 ;
      RECT 23.09 2.707 23.165 2.929 ;
      RECT 23.07 2.717 23.09 2.924 ;
      RECT 23.045 2.717 23.07 2.921 ;
      RECT 23.035 2.707 23.045 2.92 ;
      RECT 23.025 2.68 23.035 2.919 ;
      RECT 22.985 2.675 23.025 2.917 ;
      RECT 22.94 2.675 22.985 2.913 ;
      RECT 22.915 2.675 22.94 2.908 ;
      RECT 22.865 2.675 22.915 2.895 ;
      RECT 22.825 2.68 22.835 2.88 ;
      RECT 22.835 2.675 22.865 2.885 ;
      RECT 24.82 2.455 25.08 2.715 ;
      RECT 24.815 2.477 25.08 2.673 ;
      RECT 24.055 2.305 24.275 2.67 ;
      RECT 24.037 2.392 24.275 2.669 ;
      RECT 24.02 2.397 24.275 2.666 ;
      RECT 24.02 2.397 24.295 2.665 ;
      RECT 23.99 2.407 24.295 2.663 ;
      RECT 23.985 2.422 24.295 2.659 ;
      RECT 23.985 2.422 24.3 2.658 ;
      RECT 23.98 2.48 24.3 2.656 ;
      RECT 23.98 2.48 24.31 2.653 ;
      RECT 23.975 2.545 24.31 2.648 ;
      RECT 24.055 2.305 24.315 2.565 ;
      RECT 22.8 2.135 23.06 2.395 ;
      RECT 22.8 2.178 23.146 2.369 ;
      RECT 22.8 2.178 23.19 2.368 ;
      RECT 22.8 2.178 23.21 2.366 ;
      RECT 22.8 2.178 23.31 2.365 ;
      RECT 22.8 2.178 23.33 2.363 ;
      RECT 22.8 2.178 23.34 2.358 ;
      RECT 23.21 2.145 23.4 2.355 ;
      RECT 23.21 2.147 23.405 2.353 ;
      RECT 23.2 2.152 23.41 2.345 ;
      RECT 23.146 2.176 23.41 2.345 ;
      RECT 23.19 2.17 23.2 2.367 ;
      RECT 23.2 2.15 23.405 2.353 ;
      RECT 22.155 3.21 22.36 3.44 ;
      RECT 22.095 3.16 22.15 3.42 ;
      RECT 22.155 3.16 22.355 3.44 ;
      RECT 23.125 3.475 23.13 3.502 ;
      RECT 23.115 3.385 23.125 3.507 ;
      RECT 23.11 3.307 23.115 3.513 ;
      RECT 23.1 3.297 23.11 3.52 ;
      RECT 23.095 3.287 23.1 3.526 ;
      RECT 23.085 3.282 23.095 3.528 ;
      RECT 23.07 3.274 23.085 3.536 ;
      RECT 23.055 3.265 23.07 3.548 ;
      RECT 23.045 3.257 23.055 3.558 ;
      RECT 23.01 3.175 23.045 3.576 ;
      RECT 22.975 3.175 23.01 3.595 ;
      RECT 22.96 3.175 22.975 3.603 ;
      RECT 22.905 3.175 22.96 3.603 ;
      RECT 22.871 3.175 22.905 3.594 ;
      RECT 22.785 3.175 22.871 3.57 ;
      RECT 22.775 3.235 22.785 3.552 ;
      RECT 22.735 3.237 22.775 3.543 ;
      RECT 22.73 3.239 22.735 3.533 ;
      RECT 22.71 3.241 22.73 3.528 ;
      RECT 22.7 3.244 22.71 3.523 ;
      RECT 22.69 3.245 22.7 3.518 ;
      RECT 22.666 3.246 22.69 3.51 ;
      RECT 22.58 3.251 22.666 3.488 ;
      RECT 22.525 3.25 22.58 3.461 ;
      RECT 22.51 3.243 22.525 3.448 ;
      RECT 22.475 3.238 22.51 3.444 ;
      RECT 22.42 3.23 22.475 3.443 ;
      RECT 22.36 3.217 22.42 3.441 ;
      RECT 22.15 3.16 22.155 3.428 ;
      RECT 22.225 2.53 22.41 2.74 ;
      RECT 22.215 2.535 22.425 2.733 ;
      RECT 22.255 2.44 22.515 2.7 ;
      RECT 22.21 2.597 22.515 2.623 ;
      RECT 21.555 2.39 21.56 3.19 ;
      RECT 21.5 2.44 21.53 3.19 ;
      RECT 21.49 2.44 21.495 2.75 ;
      RECT 21.475 2.44 21.48 2.745 ;
      RECT 21.02 2.485 21.035 2.7 ;
      RECT 20.95 2.485 21.035 2.695 ;
      RECT 22.215 2.065 22.285 2.275 ;
      RECT 22.285 2.072 22.295 2.27 ;
      RECT 22.181 2.065 22.215 2.282 ;
      RECT 22.095 2.065 22.181 2.306 ;
      RECT 22.085 2.07 22.095 2.325 ;
      RECT 22.08 2.082 22.085 2.328 ;
      RECT 22.065 2.097 22.08 2.332 ;
      RECT 22.06 2.115 22.065 2.336 ;
      RECT 22.02 2.125 22.06 2.345 ;
      RECT 22.005 2.132 22.02 2.357 ;
      RECT 21.99 2.137 22.005 2.362 ;
      RECT 21.975 2.14 21.99 2.367 ;
      RECT 21.965 2.142 21.975 2.371 ;
      RECT 21.93 2.149 21.965 2.379 ;
      RECT 21.895 2.157 21.93 2.393 ;
      RECT 21.885 2.163 21.895 2.402 ;
      RECT 21.88 2.165 21.885 2.404 ;
      RECT 21.86 2.168 21.88 2.41 ;
      RECT 21.83 2.175 21.86 2.421 ;
      RECT 21.82 2.181 21.83 2.428 ;
      RECT 21.795 2.184 21.82 2.435 ;
      RECT 21.785 2.188 21.795 2.443 ;
      RECT 21.78 2.189 21.785 2.465 ;
      RECT 21.775 2.19 21.78 2.48 ;
      RECT 21.77 2.191 21.775 2.495 ;
      RECT 21.765 2.192 21.77 2.51 ;
      RECT 21.76 2.193 21.765 2.54 ;
      RECT 21.75 2.195 21.76 2.573 ;
      RECT 21.735 2.199 21.75 2.62 ;
      RECT 21.725 2.202 21.735 2.665 ;
      RECT 21.72 2.205 21.725 2.693 ;
      RECT 21.71 2.207 21.72 2.72 ;
      RECT 21.705 2.21 21.71 2.755 ;
      RECT 21.675 2.215 21.705 2.813 ;
      RECT 21.67 2.22 21.675 2.898 ;
      RECT 21.665 2.222 21.67 2.933 ;
      RECT 21.66 2.224 21.665 3.015 ;
      RECT 21.655 2.226 21.66 3.103 ;
      RECT 21.645 2.228 21.655 3.185 ;
      RECT 21.63 2.242 21.645 3.19 ;
      RECT 21.595 2.287 21.63 3.19 ;
      RECT 21.585 2.327 21.595 3.19 ;
      RECT 21.57 2.355 21.585 3.19 ;
      RECT 21.565 2.372 21.57 3.19 ;
      RECT 21.56 2.38 21.565 3.19 ;
      RECT 21.55 2.395 21.555 3.19 ;
      RECT 21.545 2.402 21.55 3.19 ;
      RECT 21.535 2.422 21.545 3.19 ;
      RECT 21.53 2.435 21.535 3.19 ;
      RECT 21.495 2.44 21.5 2.775 ;
      RECT 21.48 2.83 21.5 3.19 ;
      RECT 21.48 2.44 21.49 2.748 ;
      RECT 21.475 2.87 21.48 3.19 ;
      RECT 21.425 2.44 21.475 2.743 ;
      RECT 21.47 2.907 21.475 3.19 ;
      RECT 21.46 2.93 21.47 3.19 ;
      RECT 21.455 2.975 21.46 3.19 ;
      RECT 21.445 2.985 21.455 3.183 ;
      RECT 21.371 2.44 21.425 2.737 ;
      RECT 21.285 2.44 21.371 2.73 ;
      RECT 21.236 2.487 21.285 2.723 ;
      RECT 21.15 2.495 21.236 2.716 ;
      RECT 21.135 2.492 21.15 2.711 ;
      RECT 21.121 2.485 21.135 2.71 ;
      RECT 21.035 2.485 21.121 2.705 ;
      RECT 20.94 2.49 20.95 2.69 ;
      RECT 20.53 1.92 20.545 2.32 ;
      RECT 20.725 1.92 20.73 2.18 ;
      RECT 20.47 1.92 20.515 2.18 ;
      RECT 20.925 3.225 20.93 3.43 ;
      RECT 20.92 3.215 20.925 3.435 ;
      RECT 20.915 3.202 20.92 3.44 ;
      RECT 20.91 3.182 20.915 3.44 ;
      RECT 20.885 3.135 20.91 3.44 ;
      RECT 20.85 3.05 20.885 3.44 ;
      RECT 20.845 2.987 20.85 3.44 ;
      RECT 20.84 2.972 20.845 3.44 ;
      RECT 20.825 2.932 20.84 3.44 ;
      RECT 20.82 2.907 20.825 3.44 ;
      RECT 20.81 2.89 20.82 3.44 ;
      RECT 20.775 2.812 20.81 3.44 ;
      RECT 20.77 2.755 20.775 3.44 ;
      RECT 20.765 2.742 20.77 3.44 ;
      RECT 20.755 2.72 20.765 3.44 ;
      RECT 20.745 2.685 20.755 3.44 ;
      RECT 20.735 2.655 20.745 3.44 ;
      RECT 20.725 2.57 20.735 3.083 ;
      RECT 20.732 3.215 20.735 3.44 ;
      RECT 20.73 3.225 20.732 3.44 ;
      RECT 20.72 3.235 20.73 3.435 ;
      RECT 20.715 1.92 20.725 2.315 ;
      RECT 20.72 2.447 20.725 3.058 ;
      RECT 20.715 2.345 20.72 3.041 ;
      RECT 20.705 1.92 20.715 3.017 ;
      RECT 20.7 1.92 20.705 2.988 ;
      RECT 20.695 1.92 20.7 2.978 ;
      RECT 20.675 1.92 20.695 2.94 ;
      RECT 20.67 1.92 20.675 2.898 ;
      RECT 20.665 1.92 20.67 2.878 ;
      RECT 20.635 1.92 20.665 2.828 ;
      RECT 20.625 1.92 20.635 2.775 ;
      RECT 20.62 1.92 20.625 2.748 ;
      RECT 20.615 1.92 20.62 2.733 ;
      RECT 20.605 1.92 20.615 2.71 ;
      RECT 20.595 1.92 20.605 2.685 ;
      RECT 20.59 1.92 20.595 2.625 ;
      RECT 20.58 1.92 20.59 2.563 ;
      RECT 20.575 1.92 20.58 2.483 ;
      RECT 20.57 1.92 20.575 2.448 ;
      RECT 20.565 1.92 20.57 2.423 ;
      RECT 20.56 1.92 20.565 2.408 ;
      RECT 20.555 1.92 20.56 2.378 ;
      RECT 20.55 1.92 20.555 2.355 ;
      RECT 20.545 1.92 20.55 2.328 ;
      RECT 20.515 1.92 20.53 2.315 ;
      RECT 19.67 3.455 19.855 3.665 ;
      RECT 19.66 3.46 19.87 3.658 ;
      RECT 19.66 3.46 19.89 3.63 ;
      RECT 19.66 3.46 19.905 3.609 ;
      RECT 19.66 3.46 19.92 3.607 ;
      RECT 19.66 3.46 19.93 3.606 ;
      RECT 19.66 3.46 19.96 3.603 ;
      RECT 20.31 3.305 20.57 3.565 ;
      RECT 20.27 3.352 20.57 3.548 ;
      RECT 20.261 3.36 20.27 3.551 ;
      RECT 19.855 3.453 20.57 3.548 ;
      RECT 20.175 3.378 20.261 3.558 ;
      RECT 19.87 3.45 20.57 3.548 ;
      RECT 20.116 3.4 20.175 3.57 ;
      RECT 19.89 3.446 20.57 3.548 ;
      RECT 20.03 3.412 20.116 3.581 ;
      RECT 19.905 3.442 20.57 3.548 ;
      RECT 19.975 3.425 20.03 3.593 ;
      RECT 19.92 3.44 20.57 3.548 ;
      RECT 19.96 3.431 19.975 3.599 ;
      RECT 19.93 3.436 20.57 3.548 ;
      RECT 20.075 2.96 20.335 3.22 ;
      RECT 20.075 2.98 20.445 3.19 ;
      RECT 20.075 2.985 20.455 3.185 ;
      RECT 20.266 2.399 20.345 2.63 ;
      RECT 20.18 2.402 20.395 2.625 ;
      RECT 20.175 2.402 20.395 2.62 ;
      RECT 20.175 2.407 20.405 2.618 ;
      RECT 20.15 2.407 20.405 2.615 ;
      RECT 20.15 2.415 20.415 2.613 ;
      RECT 20.03 2.35 20.29 2.61 ;
      RECT 20.03 2.397 20.34 2.61 ;
      RECT 19.285 2.97 19.29 3.23 ;
      RECT 19.115 2.74 19.12 3.23 ;
      RECT 19 2.98 19.005 3.205 ;
      RECT 19.71 2.075 19.715 2.285 ;
      RECT 19.715 2.08 19.73 2.28 ;
      RECT 19.65 2.075 19.71 2.293 ;
      RECT 19.635 2.075 19.65 2.303 ;
      RECT 19.585 2.075 19.635 2.32 ;
      RECT 19.565 2.075 19.585 2.343 ;
      RECT 19.55 2.075 19.565 2.355 ;
      RECT 19.53 2.075 19.55 2.365 ;
      RECT 19.52 2.08 19.53 2.374 ;
      RECT 19.515 2.09 19.52 2.379 ;
      RECT 19.51 2.102 19.515 2.383 ;
      RECT 19.5 2.125 19.51 2.388 ;
      RECT 19.495 2.14 19.5 2.392 ;
      RECT 19.49 2.157 19.495 2.395 ;
      RECT 19.485 2.165 19.49 2.398 ;
      RECT 19.475 2.17 19.485 2.402 ;
      RECT 19.47 2.177 19.475 2.407 ;
      RECT 19.46 2.182 19.47 2.411 ;
      RECT 19.435 2.194 19.46 2.422 ;
      RECT 19.415 2.211 19.435 2.438 ;
      RECT 19.39 2.228 19.415 2.46 ;
      RECT 19.355 2.251 19.39 2.518 ;
      RECT 19.335 2.273 19.355 2.58 ;
      RECT 19.33 2.283 19.335 2.615 ;
      RECT 19.32 2.29 19.33 2.653 ;
      RECT 19.315 2.297 19.32 2.673 ;
      RECT 19.31 2.308 19.315 2.71 ;
      RECT 19.305 2.316 19.31 2.775 ;
      RECT 19.295 2.327 19.305 2.828 ;
      RECT 19.29 2.345 19.295 2.898 ;
      RECT 19.285 2.355 19.29 2.935 ;
      RECT 19.28 2.365 19.285 3.23 ;
      RECT 19.275 2.377 19.28 3.23 ;
      RECT 19.27 2.387 19.275 3.23 ;
      RECT 19.26 2.397 19.27 3.23 ;
      RECT 19.25 2.42 19.26 3.23 ;
      RECT 19.235 2.455 19.25 3.23 ;
      RECT 19.195 2.517 19.235 3.23 ;
      RECT 19.19 2.57 19.195 3.23 ;
      RECT 19.165 2.605 19.19 3.23 ;
      RECT 19.15 2.65 19.165 3.23 ;
      RECT 19.145 2.672 19.15 3.23 ;
      RECT 19.135 2.685 19.145 3.23 ;
      RECT 19.125 2.71 19.135 3.23 ;
      RECT 19.12 2.732 19.125 3.23 ;
      RECT 19.095 2.77 19.115 3.23 ;
      RECT 19.055 2.827 19.095 3.23 ;
      RECT 19.05 2.877 19.055 3.23 ;
      RECT 19.045 2.895 19.05 3.23 ;
      RECT 19.04 2.907 19.045 3.23 ;
      RECT 19.03 2.925 19.04 3.23 ;
      RECT 19.02 2.945 19.03 3.205 ;
      RECT 19.015 2.962 19.02 3.205 ;
      RECT 19.005 2.975 19.015 3.205 ;
      RECT 18.975 2.985 19 3.205 ;
      RECT 18.965 2.992 18.975 3.205 ;
      RECT 18.95 3.002 18.965 3.2 ;
      RECT 18.05 7.765 18.34 7.995 ;
      RECT 18.11 6.285 18.28 7.995 ;
      RECT 18.1 6.655 18.45 7.005 ;
      RECT 18.05 6.285 18.34 6.515 ;
      RECT 18.05 2.365 18.34 2.595 ;
      RECT 18.11 0.885 18.28 2.595 ;
      RECT 18.05 0.885 18.34 1.115 ;
      RECT 17.64 2.735 17.97 2.965 ;
      RECT 17.64 2.765 18.14 2.935 ;
      RECT 17.64 2.395 17.83 2.965 ;
      RECT 17.06 2.365 17.35 2.595 ;
      RECT 17.06 2.395 17.83 2.565 ;
      RECT 17.12 0.885 17.29 2.595 ;
      RECT 17.06 0.885 17.35 1.115 ;
      RECT 17.06 7.765 17.35 7.995 ;
      RECT 17.12 6.285 17.29 7.995 ;
      RECT 17.06 6.285 17.35 6.515 ;
      RECT 17.06 6.325 17.91 6.485 ;
      RECT 17.74 5.915 17.91 6.485 ;
      RECT 17.06 6.32 17.45 6.485 ;
      RECT 17.68 5.915 17.97 6.145 ;
      RECT 17.68 5.945 18.14 6.115 ;
      RECT 16.69 2.735 16.98 2.965 ;
      RECT 16.69 2.765 17.15 2.935 ;
      RECT 16.75 1.655 16.915 2.965 ;
      RECT 15.265 1.625 15.555 1.855 ;
      RECT 15.265 1.655 16.915 1.825 ;
      RECT 15.325 0.885 15.495 1.855 ;
      RECT 15.265 0.885 15.555 1.115 ;
      RECT 15.265 7.765 15.555 7.995 ;
      RECT 15.325 7.025 15.495 7.995 ;
      RECT 15.325 7.12 16.915 7.29 ;
      RECT 16.745 5.915 16.915 7.29 ;
      RECT 15.265 7.025 15.555 7.255 ;
      RECT 16.69 5.915 16.98 6.145 ;
      RECT 16.69 5.945 17.15 6.115 ;
      RECT 15.695 1.965 16.045 2.315 ;
      RECT 13.36 2.025 16.045 2.195 ;
      RECT 13.36 1.34 13.53 2.195 ;
      RECT 13.26 1.34 13.61 1.69 ;
      RECT 15.72 6.655 16.045 6.98 ;
      RECT 11.115 6.605 11.465 6.955 ;
      RECT 15.695 6.655 16.045 6.885 ;
      RECT 10.915 6.655 11.465 6.885 ;
      RECT 10.745 6.685 16.045 6.855 ;
      RECT 14.92 2.365 15.24 2.685 ;
      RECT 14.89 2.365 15.24 2.595 ;
      RECT 14.72 2.395 15.24 2.565 ;
      RECT 14.92 6.255 15.24 6.545 ;
      RECT 14.89 6.285 15.24 6.515 ;
      RECT 14.72 6.315 15.24 6.485 ;
      RECT 13.865 2.705 14.215 3.055 ;
      RECT 13.865 2.765 14.355 2.935 ;
      RECT 13.87 5.855 14.22 6.205 ;
      RECT 9.115 5.915 9.405 6.145 ;
      RECT 9.115 5.945 14.355 6.115 ;
      RECT 11.555 2.465 11.74 2.675 ;
      RECT 11.545 2.47 11.755 2.668 ;
      RECT 11.545 2.47 11.841 2.645 ;
      RECT 11.545 2.47 11.9 2.62 ;
      RECT 11.545 2.47 11.955 2.6 ;
      RECT 11.545 2.47 11.965 2.588 ;
      RECT 11.545 2.47 12.16 2.527 ;
      RECT 11.545 2.47 12.19 2.51 ;
      RECT 11.545 2.47 12.21 2.5 ;
      RECT 12.09 2.235 12.35 2.495 ;
      RECT 12.075 2.325 12.09 2.542 ;
      RECT 11.61 2.457 12.35 2.495 ;
      RECT 12.061 2.336 12.075 2.548 ;
      RECT 11.65 2.45 12.35 2.495 ;
      RECT 11.975 2.376 12.061 2.567 ;
      RECT 11.9 2.437 12.35 2.495 ;
      RECT 11.97 2.412 11.975 2.584 ;
      RECT 11.955 2.422 12.35 2.495 ;
      RECT 11.965 2.417 11.97 2.586 ;
      RECT 12.26 2.922 12.265 3.014 ;
      RECT 12.255 2.9 12.26 3.031 ;
      RECT 12.25 2.89 12.255 3.043 ;
      RECT 12.24 2.881 12.25 3.053 ;
      RECT 12.235 2.876 12.24 3.061 ;
      RECT 12.23 2.735 12.235 3.064 ;
      RECT 12.196 2.735 12.23 3.075 ;
      RECT 12.11 2.735 12.196 3.11 ;
      RECT 12.03 2.735 12.11 3.158 ;
      RECT 12.001 2.735 12.03 3.182 ;
      RECT 11.915 2.735 12.001 3.188 ;
      RECT 11.91 2.919 11.915 3.193 ;
      RECT 11.875 2.93 11.91 3.196 ;
      RECT 11.85 2.945 11.875 3.2 ;
      RECT 11.836 2.954 11.85 3.202 ;
      RECT 11.75 2.981 11.836 3.208 ;
      RECT 11.685 3.022 11.75 3.217 ;
      RECT 11.67 3.042 11.685 3.222 ;
      RECT 11.64 3.052 11.67 3.225 ;
      RECT 11.635 3.062 11.64 3.228 ;
      RECT 11.605 3.067 11.635 3.23 ;
      RECT 11.585 3.072 11.605 3.234 ;
      RECT 11.5 3.075 11.585 3.241 ;
      RECT 11.485 3.072 11.5 3.247 ;
      RECT 11.475 3.069 11.485 3.249 ;
      RECT 11.455 3.066 11.475 3.251 ;
      RECT 11.435 3.062 11.455 3.252 ;
      RECT 11.42 3.058 11.435 3.254 ;
      RECT 11.41 3.055 11.42 3.255 ;
      RECT 11.37 3.049 11.41 3.253 ;
      RECT 11.36 3.044 11.37 3.251 ;
      RECT 11.345 3.041 11.36 3.247 ;
      RECT 11.32 3.036 11.345 3.24 ;
      RECT 11.27 3.027 11.32 3.228 ;
      RECT 11.2 3.013 11.27 3.21 ;
      RECT 11.142 2.998 11.2 3.192 ;
      RECT 11.056 2.981 11.142 3.172 ;
      RECT 10.97 2.96 11.056 3.147 ;
      RECT 10.92 2.945 10.97 3.128 ;
      RECT 10.916 2.939 10.92 3.12 ;
      RECT 10.83 2.929 10.916 3.107 ;
      RECT 10.795 2.914 10.83 3.09 ;
      RECT 10.78 2.907 10.795 3.083 ;
      RECT 10.72 2.895 10.78 3.071 ;
      RECT 10.7 2.882 10.72 3.059 ;
      RECT 10.66 2.873 10.7 3.051 ;
      RECT 10.655 2.865 10.66 3.044 ;
      RECT 10.575 2.855 10.655 3.03 ;
      RECT 10.56 2.842 10.575 3.015 ;
      RECT 10.555 2.84 10.56 3.013 ;
      RECT 10.476 2.828 10.555 3 ;
      RECT 10.39 2.803 10.476 2.975 ;
      RECT 10.375 2.772 10.39 2.96 ;
      RECT 10.36 2.747 10.375 2.956 ;
      RECT 10.345 2.74 10.36 2.952 ;
      RECT 10.17 2.745 10.175 2.948 ;
      RECT 10.165 2.75 10.17 2.943 ;
      RECT 10.175 2.74 10.345 2.95 ;
      RECT 10.89 2.5 10.995 2.76 ;
      RECT 11.705 2.025 11.71 2.25 ;
      RECT 11.835 2.025 11.89 2.235 ;
      RECT 11.89 2.03 11.9 2.228 ;
      RECT 11.796 2.025 11.835 2.238 ;
      RECT 11.71 2.025 11.796 2.245 ;
      RECT 11.69 2.03 11.705 2.251 ;
      RECT 11.68 2.07 11.69 2.253 ;
      RECT 11.65 2.08 11.68 2.255 ;
      RECT 11.645 2.085 11.65 2.257 ;
      RECT 11.62 2.09 11.645 2.259 ;
      RECT 11.605 2.095 11.62 2.261 ;
      RECT 11.59 2.097 11.605 2.263 ;
      RECT 11.585 2.102 11.59 2.265 ;
      RECT 11.535 2.11 11.585 2.268 ;
      RECT 11.51 2.119 11.535 2.273 ;
      RECT 11.5 2.126 11.51 2.278 ;
      RECT 11.495 2.129 11.5 2.282 ;
      RECT 11.475 2.132 11.495 2.291 ;
      RECT 11.445 2.14 11.475 2.311 ;
      RECT 11.416 2.153 11.445 2.333 ;
      RECT 11.33 2.187 11.416 2.377 ;
      RECT 11.325 2.213 11.33 2.415 ;
      RECT 11.32 2.217 11.325 2.424 ;
      RECT 11.285 2.23 11.32 2.457 ;
      RECT 11.275 2.244 11.285 2.495 ;
      RECT 11.27 2.248 11.275 2.508 ;
      RECT 11.265 2.252 11.27 2.513 ;
      RECT 11.255 2.26 11.265 2.525 ;
      RECT 11.25 2.267 11.255 2.54 ;
      RECT 11.225 2.28 11.25 2.565 ;
      RECT 11.185 2.309 11.225 2.62 ;
      RECT 11.17 2.334 11.185 2.675 ;
      RECT 11.16 2.345 11.17 2.698 ;
      RECT 11.155 2.352 11.16 2.71 ;
      RECT 11.15 2.356 11.155 2.718 ;
      RECT 11.095 2.384 11.15 2.76 ;
      RECT 11.075 2.42 11.095 2.76 ;
      RECT 11.06 2.435 11.075 2.76 ;
      RECT 11.005 2.467 11.06 2.76 ;
      RECT 10.995 2.497 11.005 2.76 ;
      RECT 10.605 2.112 10.79 2.35 ;
      RECT 10.59 2.114 10.8 2.345 ;
      RECT 10.475 2.06 10.735 2.32 ;
      RECT 10.47 2.097 10.735 2.274 ;
      RECT 10.465 2.107 10.735 2.271 ;
      RECT 10.46 2.147 10.8 2.265 ;
      RECT 10.455 2.18 10.8 2.255 ;
      RECT 10.465 2.122 10.815 2.193 ;
      RECT 10.762 3.22 10.775 3.75 ;
      RECT 10.676 3.22 10.775 3.749 ;
      RECT 10.676 3.22 10.78 3.748 ;
      RECT 10.59 3.22 10.78 3.746 ;
      RECT 10.585 3.22 10.78 3.743 ;
      RECT 10.585 3.22 10.79 3.741 ;
      RECT 10.58 3.512 10.79 3.738 ;
      RECT 10.58 3.522 10.795 3.735 ;
      RECT 10.58 3.59 10.8 3.731 ;
      RECT 10.57 3.595 10.8 3.73 ;
      RECT 10.57 3.687 10.805 3.727 ;
      RECT 10.555 3.22 10.815 3.48 ;
      RECT 10.485 7.765 10.775 7.995 ;
      RECT 10.545 7.025 10.715 7.995 ;
      RECT 10.46 7.055 10.8 7.4 ;
      RECT 10.485 7.025 10.775 7.4 ;
      RECT 9.785 2.21 9.83 3.745 ;
      RECT 9.985 2.21 10.015 2.425 ;
      RECT 8.36 1.95 8.48 2.16 ;
      RECT 8.02 1.9 8.28 2.16 ;
      RECT 8.02 1.945 8.315 2.15 ;
      RECT 10.025 2.226 10.03 2.28 ;
      RECT 10.02 2.219 10.025 2.413 ;
      RECT 10.015 2.213 10.02 2.42 ;
      RECT 9.97 2.21 9.985 2.433 ;
      RECT 9.965 2.21 9.97 2.455 ;
      RECT 9.96 2.21 9.965 2.503 ;
      RECT 9.955 2.21 9.96 2.523 ;
      RECT 9.945 2.21 9.955 2.63 ;
      RECT 9.94 2.21 9.945 2.693 ;
      RECT 9.935 2.21 9.94 2.75 ;
      RECT 9.93 2.21 9.935 2.758 ;
      RECT 9.915 2.21 9.93 2.865 ;
      RECT 9.905 2.21 9.915 3 ;
      RECT 9.895 2.21 9.905 3.11 ;
      RECT 9.885 2.21 9.895 3.167 ;
      RECT 9.88 2.21 9.885 3.207 ;
      RECT 9.875 2.21 9.88 3.243 ;
      RECT 9.865 2.21 9.875 3.283 ;
      RECT 9.86 2.21 9.865 3.325 ;
      RECT 9.84 2.21 9.86 3.39 ;
      RECT 9.845 3.535 9.85 3.715 ;
      RECT 9.84 3.517 9.845 3.723 ;
      RECT 9.835 2.21 9.84 3.453 ;
      RECT 9.835 3.497 9.84 3.73 ;
      RECT 9.83 2.21 9.835 3.74 ;
      RECT 9.775 2.21 9.785 2.51 ;
      RECT 9.78 2.757 9.785 3.745 ;
      RECT 9.775 2.822 9.78 3.745 ;
      RECT 9.77 2.211 9.775 2.5 ;
      RECT 9.765 2.887 9.775 3.745 ;
      RECT 9.76 2.212 9.77 2.49 ;
      RECT 9.75 3 9.765 3.745 ;
      RECT 9.755 2.213 9.76 2.48 ;
      RECT 9.735 2.214 9.755 2.458 ;
      RECT 9.74 3.097 9.75 3.745 ;
      RECT 9.735 3.172 9.74 3.745 ;
      RECT 9.725 2.213 9.735 2.435 ;
      RECT 9.73 3.215 9.735 3.745 ;
      RECT 9.725 3.242 9.73 3.745 ;
      RECT 9.715 2.211 9.725 2.423 ;
      RECT 9.72 3.285 9.725 3.745 ;
      RECT 9.715 3.312 9.72 3.745 ;
      RECT 9.705 2.21 9.715 2.41 ;
      RECT 9.71 3.327 9.715 3.745 ;
      RECT 9.67 3.385 9.71 3.745 ;
      RECT 9.7 2.209 9.705 2.395 ;
      RECT 9.695 2.207 9.7 2.388 ;
      RECT 9.685 2.204 9.695 2.378 ;
      RECT 9.68 2.201 9.685 2.363 ;
      RECT 9.665 2.197 9.68 2.356 ;
      RECT 9.66 3.44 9.67 3.745 ;
      RECT 9.66 2.194 9.665 2.351 ;
      RECT 9.645 2.19 9.66 2.345 ;
      RECT 9.655 3.457 9.66 3.745 ;
      RECT 9.645 3.52 9.655 3.745 ;
      RECT 9.565 2.175 9.645 2.325 ;
      RECT 9.64 3.527 9.645 3.74 ;
      RECT 9.635 3.535 9.64 3.73 ;
      RECT 9.555 2.161 9.565 2.309 ;
      RECT 9.54 2.157 9.555 2.307 ;
      RECT 9.53 2.152 9.54 2.303 ;
      RECT 9.505 2.145 9.53 2.295 ;
      RECT 9.5 2.14 9.505 2.29 ;
      RECT 9.49 2.14 9.5 2.288 ;
      RECT 9.48 2.138 9.49 2.286 ;
      RECT 9.45 2.13 9.48 2.28 ;
      RECT 9.435 2.122 9.45 2.273 ;
      RECT 9.415 2.117 9.435 2.266 ;
      RECT 9.41 2.113 9.415 2.261 ;
      RECT 9.38 2.106 9.41 2.255 ;
      RECT 9.355 2.097 9.38 2.245 ;
      RECT 9.325 2.09 9.355 2.237 ;
      RECT 9.3 2.08 9.325 2.228 ;
      RECT 9.285 2.072 9.3 2.222 ;
      RECT 9.26 2.067 9.285 2.217 ;
      RECT 9.25 2.063 9.26 2.212 ;
      RECT 9.23 2.058 9.25 2.207 ;
      RECT 9.195 2.053 9.23 2.2 ;
      RECT 9.135 2.048 9.195 2.193 ;
      RECT 9.122 2.044 9.135 2.191 ;
      RECT 9.036 2.039 9.122 2.188 ;
      RECT 8.95 2.029 9.036 2.184 ;
      RECT 8.909 2.022 8.95 2.181 ;
      RECT 8.823 2.015 8.909 2.178 ;
      RECT 8.737 2.005 8.823 2.174 ;
      RECT 8.651 1.995 8.737 2.169 ;
      RECT 8.565 1.985 8.651 2.165 ;
      RECT 8.555 1.97 8.565 2.163 ;
      RECT 8.545 1.955 8.555 2.163 ;
      RECT 8.48 1.95 8.545 2.162 ;
      RECT 8.315 1.947 8.36 2.155 ;
      RECT 9.56 2.852 9.565 3.043 ;
      RECT 9.555 2.847 9.56 3.05 ;
      RECT 9.541 2.845 9.555 3.056 ;
      RECT 9.455 2.845 9.541 3.058 ;
      RECT 9.451 2.845 9.455 3.061 ;
      RECT 9.365 2.845 9.451 3.079 ;
      RECT 9.355 2.85 9.365 3.098 ;
      RECT 9.345 2.905 9.355 3.102 ;
      RECT 9.32 2.92 9.345 3.109 ;
      RECT 9.28 2.94 9.32 3.122 ;
      RECT 9.275 2.952 9.28 3.132 ;
      RECT 9.26 2.958 9.275 3.137 ;
      RECT 9.255 2.963 9.26 3.141 ;
      RECT 9.235 2.97 9.255 3.146 ;
      RECT 9.165 2.995 9.235 3.163 ;
      RECT 9.125 3.023 9.165 3.183 ;
      RECT 9.12 3.033 9.125 3.191 ;
      RECT 9.1 3.04 9.12 3.193 ;
      RECT 9.095 3.047 9.1 3.196 ;
      RECT 9.065 3.055 9.095 3.199 ;
      RECT 9.06 3.06 9.065 3.203 ;
      RECT 8.986 3.064 9.06 3.211 ;
      RECT 8.9 3.073 8.986 3.227 ;
      RECT 8.896 3.078 8.9 3.236 ;
      RECT 8.81 3.083 8.896 3.246 ;
      RECT 8.77 3.091 8.81 3.258 ;
      RECT 8.72 3.097 8.77 3.265 ;
      RECT 8.635 3.106 8.72 3.28 ;
      RECT 8.56 3.117 8.635 3.298 ;
      RECT 8.525 3.124 8.56 3.308 ;
      RECT 8.45 3.132 8.525 3.313 ;
      RECT 8.395 3.141 8.45 3.313 ;
      RECT 8.37 3.146 8.395 3.311 ;
      RECT 8.36 3.149 8.37 3.309 ;
      RECT 8.325 3.151 8.36 3.307 ;
      RECT 8.295 3.153 8.325 3.303 ;
      RECT 8.25 3.152 8.295 3.299 ;
      RECT 8.23 3.147 8.25 3.296 ;
      RECT 8.18 3.132 8.23 3.293 ;
      RECT 8.17 3.117 8.18 3.288 ;
      RECT 8.12 3.102 8.17 3.278 ;
      RECT 8.07 3.077 8.12 3.258 ;
      RECT 8.06 3.062 8.07 3.24 ;
      RECT 8.055 3.06 8.06 3.234 ;
      RECT 8.035 3.055 8.055 3.229 ;
      RECT 8.03 3.047 8.035 3.223 ;
      RECT 8.015 3.041 8.03 3.216 ;
      RECT 8.01 3.036 8.015 3.208 ;
      RECT 7.99 3.031 8.01 3.2 ;
      RECT 7.975 3.024 7.99 3.193 ;
      RECT 7.96 3.018 7.975 3.184 ;
      RECT 7.955 3.012 7.96 3.177 ;
      RECT 7.91 2.987 7.955 3.163 ;
      RECT 7.895 2.957 7.91 3.145 ;
      RECT 7.88 2.94 7.895 3.136 ;
      RECT 7.855 2.92 7.88 3.124 ;
      RECT 7.815 2.89 7.855 3.104 ;
      RECT 7.805 2.86 7.815 3.089 ;
      RECT 7.79 2.85 7.805 3.082 ;
      RECT 7.735 2.815 7.79 3.061 ;
      RECT 7.72 2.778 7.735 3.04 ;
      RECT 7.71 2.765 7.72 3.032 ;
      RECT 7.66 2.735 7.71 3.014 ;
      RECT 7.645 2.665 7.66 2.995 ;
      RECT 7.6 2.665 7.645 2.978 ;
      RECT 7.575 2.665 7.6 2.96 ;
      RECT 7.565 2.665 7.575 2.953 ;
      RECT 7.486 2.665 7.565 2.946 ;
      RECT 7.4 2.665 7.486 2.938 ;
      RECT 7.385 2.697 7.4 2.933 ;
      RECT 7.31 2.707 7.385 2.929 ;
      RECT 7.29 2.717 7.31 2.924 ;
      RECT 7.265 2.717 7.29 2.921 ;
      RECT 7.255 2.707 7.265 2.92 ;
      RECT 7.245 2.68 7.255 2.919 ;
      RECT 7.205 2.675 7.245 2.917 ;
      RECT 7.16 2.675 7.205 2.913 ;
      RECT 7.135 2.675 7.16 2.908 ;
      RECT 7.085 2.675 7.135 2.895 ;
      RECT 7.045 2.68 7.055 2.88 ;
      RECT 7.055 2.675 7.085 2.885 ;
      RECT 9.04 2.455 9.3 2.715 ;
      RECT 9.035 2.477 9.3 2.673 ;
      RECT 8.275 2.305 8.495 2.67 ;
      RECT 8.257 2.392 8.495 2.669 ;
      RECT 8.24 2.397 8.495 2.666 ;
      RECT 8.24 2.397 8.515 2.665 ;
      RECT 8.21 2.407 8.515 2.663 ;
      RECT 8.205 2.422 8.515 2.659 ;
      RECT 8.205 2.422 8.52 2.658 ;
      RECT 8.2 2.48 8.52 2.656 ;
      RECT 8.2 2.48 8.53 2.653 ;
      RECT 8.195 2.545 8.53 2.648 ;
      RECT 8.275 2.305 8.535 2.565 ;
      RECT 7.02 2.135 7.28 2.395 ;
      RECT 7.02 2.178 7.366 2.369 ;
      RECT 7.02 2.178 7.41 2.368 ;
      RECT 7.02 2.178 7.43 2.366 ;
      RECT 7.02 2.178 7.53 2.365 ;
      RECT 7.02 2.178 7.55 2.363 ;
      RECT 7.02 2.178 7.56 2.358 ;
      RECT 7.43 2.145 7.62 2.355 ;
      RECT 7.43 2.147 7.625 2.353 ;
      RECT 7.42 2.152 7.63 2.345 ;
      RECT 7.366 2.176 7.63 2.345 ;
      RECT 7.41 2.17 7.42 2.367 ;
      RECT 7.42 2.15 7.625 2.353 ;
      RECT 6.375 3.21 6.58 3.44 ;
      RECT 6.315 3.16 6.37 3.42 ;
      RECT 6.375 3.16 6.575 3.44 ;
      RECT 7.345 3.475 7.35 3.502 ;
      RECT 7.335 3.385 7.345 3.507 ;
      RECT 7.33 3.307 7.335 3.513 ;
      RECT 7.32 3.297 7.33 3.52 ;
      RECT 7.315 3.287 7.32 3.526 ;
      RECT 7.305 3.282 7.315 3.528 ;
      RECT 7.29 3.274 7.305 3.536 ;
      RECT 7.275 3.265 7.29 3.548 ;
      RECT 7.265 3.257 7.275 3.558 ;
      RECT 7.23 3.175 7.265 3.576 ;
      RECT 7.195 3.175 7.23 3.595 ;
      RECT 7.18 3.175 7.195 3.603 ;
      RECT 7.125 3.175 7.18 3.603 ;
      RECT 7.091 3.175 7.125 3.594 ;
      RECT 7.005 3.175 7.091 3.57 ;
      RECT 6.995 3.235 7.005 3.552 ;
      RECT 6.955 3.237 6.995 3.543 ;
      RECT 6.95 3.239 6.955 3.533 ;
      RECT 6.93 3.241 6.95 3.528 ;
      RECT 6.92 3.244 6.93 3.523 ;
      RECT 6.91 3.245 6.92 3.518 ;
      RECT 6.886 3.246 6.91 3.51 ;
      RECT 6.8 3.251 6.886 3.488 ;
      RECT 6.745 3.25 6.8 3.461 ;
      RECT 6.73 3.243 6.745 3.448 ;
      RECT 6.695 3.238 6.73 3.444 ;
      RECT 6.64 3.23 6.695 3.443 ;
      RECT 6.58 3.217 6.64 3.441 ;
      RECT 6.37 3.16 6.375 3.428 ;
      RECT 6.445 2.53 6.63 2.74 ;
      RECT 6.435 2.535 6.645 2.733 ;
      RECT 6.475 2.44 6.735 2.7 ;
      RECT 6.43 2.597 6.735 2.623 ;
      RECT 5.775 2.39 5.78 3.19 ;
      RECT 5.72 2.44 5.75 3.19 ;
      RECT 5.71 2.44 5.715 2.75 ;
      RECT 5.695 2.44 5.7 2.745 ;
      RECT 5.24 2.485 5.255 2.7 ;
      RECT 5.17 2.485 5.255 2.695 ;
      RECT 6.435 2.065 6.505 2.275 ;
      RECT 6.505 2.072 6.515 2.27 ;
      RECT 6.401 2.065 6.435 2.282 ;
      RECT 6.315 2.065 6.401 2.306 ;
      RECT 6.305 2.07 6.315 2.325 ;
      RECT 6.3 2.082 6.305 2.328 ;
      RECT 6.285 2.097 6.3 2.332 ;
      RECT 6.28 2.115 6.285 2.336 ;
      RECT 6.24 2.125 6.28 2.345 ;
      RECT 6.225 2.132 6.24 2.357 ;
      RECT 6.21 2.137 6.225 2.362 ;
      RECT 6.195 2.14 6.21 2.367 ;
      RECT 6.185 2.142 6.195 2.371 ;
      RECT 6.15 2.149 6.185 2.379 ;
      RECT 6.115 2.157 6.15 2.393 ;
      RECT 6.105 2.163 6.115 2.402 ;
      RECT 6.1 2.165 6.105 2.404 ;
      RECT 6.08 2.168 6.1 2.41 ;
      RECT 6.05 2.175 6.08 2.421 ;
      RECT 6.04 2.181 6.05 2.428 ;
      RECT 6.015 2.184 6.04 2.435 ;
      RECT 6.005 2.188 6.015 2.443 ;
      RECT 6 2.189 6.005 2.465 ;
      RECT 5.995 2.19 6 2.48 ;
      RECT 5.99 2.191 5.995 2.495 ;
      RECT 5.985 2.192 5.99 2.51 ;
      RECT 5.98 2.193 5.985 2.54 ;
      RECT 5.97 2.195 5.98 2.573 ;
      RECT 5.955 2.199 5.97 2.62 ;
      RECT 5.945 2.202 5.955 2.665 ;
      RECT 5.94 2.205 5.945 2.693 ;
      RECT 5.93 2.207 5.94 2.72 ;
      RECT 5.925 2.21 5.93 2.755 ;
      RECT 5.895 2.215 5.925 2.813 ;
      RECT 5.89 2.22 5.895 2.898 ;
      RECT 5.885 2.222 5.89 2.933 ;
      RECT 5.88 2.224 5.885 3.015 ;
      RECT 5.875 2.226 5.88 3.103 ;
      RECT 5.865 2.228 5.875 3.185 ;
      RECT 5.85 2.242 5.865 3.19 ;
      RECT 5.815 2.287 5.85 3.19 ;
      RECT 5.805 2.327 5.815 3.19 ;
      RECT 5.79 2.355 5.805 3.19 ;
      RECT 5.785 2.372 5.79 3.19 ;
      RECT 5.78 2.38 5.785 3.19 ;
      RECT 5.77 2.395 5.775 3.19 ;
      RECT 5.765 2.402 5.77 3.19 ;
      RECT 5.755 2.422 5.765 3.19 ;
      RECT 5.75 2.435 5.755 3.19 ;
      RECT 5.715 2.44 5.72 2.775 ;
      RECT 5.7 2.83 5.72 3.19 ;
      RECT 5.7 2.44 5.71 2.748 ;
      RECT 5.695 2.87 5.7 3.19 ;
      RECT 5.645 2.44 5.695 2.743 ;
      RECT 5.69 2.907 5.695 3.19 ;
      RECT 5.68 2.93 5.69 3.19 ;
      RECT 5.675 2.975 5.68 3.19 ;
      RECT 5.665 2.985 5.675 3.183 ;
      RECT 5.591 2.44 5.645 2.737 ;
      RECT 5.505 2.44 5.591 2.73 ;
      RECT 5.456 2.487 5.505 2.723 ;
      RECT 5.37 2.495 5.456 2.716 ;
      RECT 5.355 2.492 5.37 2.711 ;
      RECT 5.341 2.485 5.355 2.71 ;
      RECT 5.255 2.485 5.341 2.705 ;
      RECT 5.16 2.49 5.17 2.69 ;
      RECT 4.75 1.92 4.765 2.32 ;
      RECT 4.945 1.92 4.95 2.18 ;
      RECT 4.69 1.92 4.735 2.18 ;
      RECT 5.145 3.225 5.15 3.43 ;
      RECT 5.14 3.215 5.145 3.435 ;
      RECT 5.135 3.202 5.14 3.44 ;
      RECT 5.13 3.182 5.135 3.44 ;
      RECT 5.105 3.135 5.13 3.44 ;
      RECT 5.07 3.05 5.105 3.44 ;
      RECT 5.065 2.987 5.07 3.44 ;
      RECT 5.06 2.972 5.065 3.44 ;
      RECT 5.045 2.932 5.06 3.44 ;
      RECT 5.04 2.907 5.045 3.44 ;
      RECT 5.03 2.89 5.04 3.44 ;
      RECT 4.995 2.812 5.03 3.44 ;
      RECT 4.99 2.755 4.995 3.44 ;
      RECT 4.985 2.742 4.99 3.44 ;
      RECT 4.975 2.72 4.985 3.44 ;
      RECT 4.965 2.685 4.975 3.44 ;
      RECT 4.955 2.655 4.965 3.44 ;
      RECT 4.945 2.57 4.955 3.083 ;
      RECT 4.952 3.215 4.955 3.44 ;
      RECT 4.95 3.225 4.952 3.44 ;
      RECT 4.94 3.235 4.95 3.435 ;
      RECT 4.935 1.92 4.945 2.315 ;
      RECT 4.94 2.447 4.945 3.058 ;
      RECT 4.935 2.345 4.94 3.041 ;
      RECT 4.925 1.92 4.935 3.017 ;
      RECT 4.92 1.92 4.925 2.988 ;
      RECT 4.915 1.92 4.92 2.978 ;
      RECT 4.895 1.92 4.915 2.94 ;
      RECT 4.89 1.92 4.895 2.898 ;
      RECT 4.885 1.92 4.89 2.878 ;
      RECT 4.855 1.92 4.885 2.828 ;
      RECT 4.845 1.92 4.855 2.775 ;
      RECT 4.84 1.92 4.845 2.748 ;
      RECT 4.835 1.92 4.84 2.733 ;
      RECT 4.825 1.92 4.835 2.71 ;
      RECT 4.815 1.92 4.825 2.685 ;
      RECT 4.81 1.92 4.815 2.625 ;
      RECT 4.8 1.92 4.81 2.563 ;
      RECT 4.795 1.92 4.8 2.483 ;
      RECT 4.79 1.92 4.795 2.448 ;
      RECT 4.785 1.92 4.79 2.423 ;
      RECT 4.78 1.92 4.785 2.408 ;
      RECT 4.775 1.92 4.78 2.378 ;
      RECT 4.77 1.92 4.775 2.355 ;
      RECT 4.765 1.92 4.77 2.328 ;
      RECT 4.735 1.92 4.75 2.315 ;
      RECT 3.89 3.455 4.075 3.665 ;
      RECT 3.88 3.46 4.09 3.658 ;
      RECT 3.88 3.46 4.11 3.63 ;
      RECT 3.88 3.46 4.125 3.609 ;
      RECT 3.88 3.46 4.14 3.607 ;
      RECT 3.88 3.46 4.15 3.606 ;
      RECT 3.88 3.46 4.18 3.603 ;
      RECT 4.53 3.305 4.79 3.565 ;
      RECT 4.49 3.352 4.79 3.548 ;
      RECT 4.481 3.36 4.49 3.551 ;
      RECT 4.075 3.453 4.79 3.548 ;
      RECT 4.395 3.378 4.481 3.558 ;
      RECT 4.09 3.45 4.79 3.548 ;
      RECT 4.336 3.4 4.395 3.57 ;
      RECT 4.11 3.446 4.79 3.548 ;
      RECT 4.25 3.412 4.336 3.581 ;
      RECT 4.125 3.442 4.79 3.548 ;
      RECT 4.195 3.425 4.25 3.593 ;
      RECT 4.14 3.44 4.79 3.548 ;
      RECT 4.18 3.431 4.195 3.599 ;
      RECT 4.15 3.436 4.79 3.548 ;
      RECT 4.295 2.96 4.555 3.22 ;
      RECT 4.295 2.98 4.665 3.19 ;
      RECT 4.295 2.985 4.675 3.185 ;
      RECT 4.486 2.399 4.565 2.63 ;
      RECT 4.4 2.402 4.615 2.625 ;
      RECT 4.395 2.402 4.615 2.62 ;
      RECT 4.395 2.407 4.625 2.618 ;
      RECT 4.37 2.407 4.625 2.615 ;
      RECT 4.37 2.415 4.635 2.613 ;
      RECT 4.25 2.35 4.51 2.61 ;
      RECT 4.25 2.397 4.56 2.61 ;
      RECT 3.505 2.97 3.51 3.23 ;
      RECT 3.335 2.74 3.34 3.23 ;
      RECT 3.22 2.98 3.225 3.205 ;
      RECT 3.93 2.075 3.935 2.285 ;
      RECT 3.935 2.08 3.95 2.28 ;
      RECT 3.87 2.075 3.93 2.293 ;
      RECT 3.855 2.075 3.87 2.303 ;
      RECT 3.805 2.075 3.855 2.32 ;
      RECT 3.785 2.075 3.805 2.343 ;
      RECT 3.77 2.075 3.785 2.355 ;
      RECT 3.75 2.075 3.77 2.365 ;
      RECT 3.74 2.08 3.75 2.374 ;
      RECT 3.735 2.09 3.74 2.379 ;
      RECT 3.73 2.102 3.735 2.383 ;
      RECT 3.72 2.125 3.73 2.388 ;
      RECT 3.715 2.14 3.72 2.392 ;
      RECT 3.71 2.157 3.715 2.395 ;
      RECT 3.705 2.165 3.71 2.398 ;
      RECT 3.695 2.17 3.705 2.402 ;
      RECT 3.69 2.177 3.695 2.407 ;
      RECT 3.68 2.182 3.69 2.411 ;
      RECT 3.655 2.194 3.68 2.422 ;
      RECT 3.635 2.211 3.655 2.438 ;
      RECT 3.61 2.228 3.635 2.46 ;
      RECT 3.575 2.251 3.61 2.518 ;
      RECT 3.555 2.273 3.575 2.58 ;
      RECT 3.55 2.283 3.555 2.615 ;
      RECT 3.54 2.29 3.55 2.653 ;
      RECT 3.535 2.297 3.54 2.673 ;
      RECT 3.53 2.308 3.535 2.71 ;
      RECT 3.525 2.316 3.53 2.775 ;
      RECT 3.515 2.327 3.525 2.828 ;
      RECT 3.51 2.345 3.515 2.898 ;
      RECT 3.505 2.355 3.51 2.935 ;
      RECT 3.5 2.365 3.505 3.23 ;
      RECT 3.495 2.377 3.5 3.23 ;
      RECT 3.49 2.387 3.495 3.23 ;
      RECT 3.48 2.397 3.49 3.23 ;
      RECT 3.47 2.42 3.48 3.23 ;
      RECT 3.455 2.455 3.47 3.23 ;
      RECT 3.415 2.517 3.455 3.23 ;
      RECT 3.41 2.57 3.415 3.23 ;
      RECT 3.385 2.605 3.41 3.23 ;
      RECT 3.37 2.65 3.385 3.23 ;
      RECT 3.365 2.672 3.37 3.23 ;
      RECT 3.355 2.685 3.365 3.23 ;
      RECT 3.345 2.71 3.355 3.23 ;
      RECT 3.34 2.732 3.345 3.23 ;
      RECT 3.315 2.77 3.335 3.23 ;
      RECT 3.275 2.827 3.315 3.23 ;
      RECT 3.27 2.877 3.275 3.23 ;
      RECT 3.265 2.895 3.27 3.23 ;
      RECT 3.26 2.907 3.265 3.23 ;
      RECT 3.25 2.925 3.26 3.23 ;
      RECT 3.24 2.945 3.25 3.205 ;
      RECT 3.235 2.962 3.24 3.205 ;
      RECT 3.225 2.975 3.235 3.205 ;
      RECT 3.195 2.985 3.22 3.205 ;
      RECT 3.185 2.992 3.195 3.205 ;
      RECT 3.17 3.002 3.185 3.2 ;
      RECT 1.98 6.655 2.27 6.885 ;
      RECT 1.81 6.685 2.27 6.855 ;
      RECT 1.55 7.765 1.84 7.995 ;
      RECT 1.61 7.025 1.78 7.995 ;
      RECT 1.52 7.025 1.87 7.315 ;
      RECT 1.145 6.285 1.495 6.575 ;
      RECT 1.005 6.315 1.495 6.485 ;
      RECT 0.18 5.915 0.47 6.145 ;
      RECT 0.18 5.945 0.64 6.115 ;
      RECT 76.06 2.85 76.43 3.22 ;
      RECT 60.275 2.85 60.645 3.22 ;
      RECT 44.49 2.85 44.86 3.22 ;
      RECT 28.715 2.85 29.085 3.22 ;
      RECT 12.935 2.85 13.305 3.22 ;
    LAYER mcon ;
      RECT 0.355 8.64 0.525 8.81 ;
      RECT 0.31 8.605 0.48 8.775 ;
      RECT 81.235 0.915 81.405 1.085 ;
      RECT 81.235 2.395 81.405 2.565 ;
      RECT 81.235 6.315 81.405 6.485 ;
      RECT 81.235 7.795 81.405 7.965 ;
      RECT 80.885 0.105 81.055 0.275 ;
      RECT 80.885 4.165 81.055 4.335 ;
      RECT 80.885 4.545 81.055 4.715 ;
      RECT 80.885 8.605 81.055 8.775 ;
      RECT 80.865 2.765 81.035 2.935 ;
      RECT 80.865 5.945 81.035 6.115 ;
      RECT 80.245 0.915 80.415 1.085 ;
      RECT 80.245 2.395 80.415 2.565 ;
      RECT 80.245 6.315 80.415 6.485 ;
      RECT 80.245 7.795 80.415 7.965 ;
      RECT 79.895 0.105 80.065 0.275 ;
      RECT 79.895 4.165 80.065 4.335 ;
      RECT 79.895 4.545 80.065 4.715 ;
      RECT 79.895 8.605 80.065 8.775 ;
      RECT 79.875 2.765 80.045 2.935 ;
      RECT 79.875 5.945 80.045 6.115 ;
      RECT 79.19 0.105 79.36 0.275 ;
      RECT 79.19 4.165 79.36 4.335 ;
      RECT 79.19 4.545 79.36 4.715 ;
      RECT 79.19 8.605 79.36 8.775 ;
      RECT 78.88 2.025 79.05 2.195 ;
      RECT 78.88 6.685 79.05 6.855 ;
      RECT 78.51 0.105 78.68 0.275 ;
      RECT 78.51 8.605 78.68 8.775 ;
      RECT 78.45 0.915 78.62 1.085 ;
      RECT 78.45 1.655 78.62 1.825 ;
      RECT 78.45 7.055 78.62 7.225 ;
      RECT 78.45 7.795 78.62 7.965 ;
      RECT 78.075 2.395 78.245 2.565 ;
      RECT 78.075 6.315 78.245 6.485 ;
      RECT 77.83 0.105 78 0.275 ;
      RECT 77.83 8.605 78 8.775 ;
      RECT 77.15 0.105 77.32 0.275 ;
      RECT 77.15 8.605 77.32 8.775 ;
      RECT 77.08 2.765 77.25 2.935 ;
      RECT 77.08 5.945 77.25 6.115 ;
      RECT 75.525 1.415 75.695 1.585 ;
      RECT 75.525 4.135 75.695 4.305 ;
      RECT 75.155 2.875 75.325 3.045 ;
      RECT 75.065 1.415 75.235 1.585 ;
      RECT 75.065 4.135 75.235 4.305 ;
      RECT 74.835 2.045 75.005 2.215 ;
      RECT 74.69 2.485 74.86 2.655 ;
      RECT 74.605 1.415 74.775 1.585 ;
      RECT 74.605 4.135 74.775 4.305 ;
      RECT 74.41 4.545 74.58 4.715 ;
      RECT 74.41 8.605 74.58 8.775 ;
      RECT 74.145 1.415 74.315 1.585 ;
      RECT 74.145 4.135 74.315 4.305 ;
      RECT 74.1 6.685 74.27 6.855 ;
      RECT 74.08 2.525 74.25 2.695 ;
      RECT 73.735 2.16 73.905 2.33 ;
      RECT 73.73 8.605 73.9 8.775 ;
      RECT 73.725 3.52 73.895 3.69 ;
      RECT 73.685 1.415 73.855 1.585 ;
      RECT 73.685 4.135 73.855 4.305 ;
      RECT 73.67 7.055 73.84 7.225 ;
      RECT 73.67 7.795 73.84 7.965 ;
      RECT 73.31 2.76 73.48 2.93 ;
      RECT 73.295 6.315 73.465 6.485 ;
      RECT 73.225 1.415 73.395 1.585 ;
      RECT 73.225 4.135 73.395 4.305 ;
      RECT 73.05 8.605 73.22 8.775 ;
      RECT 72.96 2.235 73.13 2.405 ;
      RECT 72.78 3.55 72.95 3.72 ;
      RECT 72.765 1.415 72.935 1.585 ;
      RECT 72.765 4.135 72.935 4.305 ;
      RECT 72.5 2.865 72.67 3.035 ;
      RECT 72.37 8.605 72.54 8.775 ;
      RECT 72.305 1.415 72.475 1.585 ;
      RECT 72.305 4.135 72.475 4.305 ;
      RECT 72.3 5.945 72.47 6.115 ;
      RECT 72.18 2.49 72.35 2.66 ;
      RECT 71.845 1.415 72.015 1.585 ;
      RECT 71.845 4.135 72.015 4.305 ;
      RECT 71.49 1.97 71.66 2.14 ;
      RECT 71.415 2.44 71.585 2.61 ;
      RECT 71.385 1.415 71.555 1.585 ;
      RECT 71.385 4.135 71.555 4.305 ;
      RECT 70.925 1.415 71.095 1.585 ;
      RECT 70.925 4.135 71.095 4.305 ;
      RECT 70.565 2.165 70.735 2.335 ;
      RECT 70.465 1.415 70.635 1.585 ;
      RECT 70.465 4.135 70.635 4.305 ;
      RECT 70.225 3.36 70.395 3.53 ;
      RECT 70.19 2.695 70.36 2.865 ;
      RECT 70.005 1.415 70.175 1.585 ;
      RECT 70.005 4.135 70.175 4.305 ;
      RECT 69.58 2.55 69.75 2.72 ;
      RECT 69.545 1.415 69.715 1.585 ;
      RECT 69.545 4.135 69.715 4.305 ;
      RECT 69.51 3.25 69.68 3.42 ;
      RECT 69.45 2.085 69.62 2.255 ;
      RECT 69.085 1.415 69.255 1.585 ;
      RECT 69.085 4.135 69.255 4.305 ;
      RECT 68.81 3 68.98 3.17 ;
      RECT 68.625 1.415 68.795 1.585 ;
      RECT 68.625 4.135 68.795 4.305 ;
      RECT 68.305 2.505 68.475 2.675 ;
      RECT 68.165 1.415 68.335 1.585 ;
      RECT 68.165 4.135 68.335 4.305 ;
      RECT 68.085 3.25 68.255 3.42 ;
      RECT 67.88 2.13 68.05 2.3 ;
      RECT 67.705 1.415 67.875 1.585 ;
      RECT 67.705 4.135 67.875 4.305 ;
      RECT 67.61 3 67.78 3.17 ;
      RECT 67.57 2.43 67.74 2.6 ;
      RECT 67.245 1.415 67.415 1.585 ;
      RECT 67.245 4.135 67.415 4.305 ;
      RECT 67.025 3.475 67.195 3.645 ;
      RECT 66.885 2.095 67.055 2.265 ;
      RECT 66.785 1.415 66.955 1.585 ;
      RECT 66.785 4.135 66.955 4.305 ;
      RECT 66.325 1.415 66.495 1.585 ;
      RECT 66.325 4.135 66.495 4.305 ;
      RECT 66.315 3.015 66.485 3.185 ;
      RECT 65.45 0.915 65.62 1.085 ;
      RECT 65.45 2.395 65.62 2.565 ;
      RECT 65.45 6.315 65.62 6.485 ;
      RECT 65.45 7.795 65.62 7.965 ;
      RECT 65.1 0.105 65.27 0.275 ;
      RECT 65.1 4.165 65.27 4.335 ;
      RECT 65.1 4.545 65.27 4.715 ;
      RECT 65.1 8.605 65.27 8.775 ;
      RECT 65.08 2.765 65.25 2.935 ;
      RECT 65.08 5.945 65.25 6.115 ;
      RECT 64.46 0.915 64.63 1.085 ;
      RECT 64.46 2.395 64.63 2.565 ;
      RECT 64.46 6.315 64.63 6.485 ;
      RECT 64.46 7.795 64.63 7.965 ;
      RECT 64.11 0.105 64.28 0.275 ;
      RECT 64.11 4.165 64.28 4.335 ;
      RECT 64.11 4.545 64.28 4.715 ;
      RECT 64.11 8.605 64.28 8.775 ;
      RECT 64.09 2.765 64.26 2.935 ;
      RECT 64.09 5.945 64.26 6.115 ;
      RECT 63.405 0.105 63.575 0.275 ;
      RECT 63.405 4.165 63.575 4.335 ;
      RECT 63.405 4.545 63.575 4.715 ;
      RECT 63.405 8.605 63.575 8.775 ;
      RECT 63.095 2.025 63.265 2.195 ;
      RECT 63.095 6.685 63.265 6.855 ;
      RECT 62.725 0.105 62.895 0.275 ;
      RECT 62.725 8.605 62.895 8.775 ;
      RECT 62.665 0.915 62.835 1.085 ;
      RECT 62.665 1.655 62.835 1.825 ;
      RECT 62.665 7.055 62.835 7.225 ;
      RECT 62.665 7.795 62.835 7.965 ;
      RECT 62.29 2.395 62.46 2.565 ;
      RECT 62.29 6.315 62.46 6.485 ;
      RECT 62.045 0.105 62.215 0.275 ;
      RECT 62.045 8.605 62.215 8.775 ;
      RECT 61.365 0.105 61.535 0.275 ;
      RECT 61.365 8.605 61.535 8.775 ;
      RECT 61.295 2.765 61.465 2.935 ;
      RECT 61.295 5.945 61.465 6.115 ;
      RECT 59.74 1.415 59.91 1.585 ;
      RECT 59.74 4.135 59.91 4.305 ;
      RECT 59.37 2.875 59.54 3.045 ;
      RECT 59.28 1.415 59.45 1.585 ;
      RECT 59.28 4.135 59.45 4.305 ;
      RECT 59.05 2.045 59.22 2.215 ;
      RECT 58.905 2.485 59.075 2.655 ;
      RECT 58.82 1.415 58.99 1.585 ;
      RECT 58.82 4.135 58.99 4.305 ;
      RECT 58.625 4.545 58.795 4.715 ;
      RECT 58.625 8.605 58.795 8.775 ;
      RECT 58.36 1.415 58.53 1.585 ;
      RECT 58.36 4.135 58.53 4.305 ;
      RECT 58.315 6.685 58.485 6.855 ;
      RECT 58.295 2.525 58.465 2.695 ;
      RECT 57.95 2.16 58.12 2.33 ;
      RECT 57.945 8.605 58.115 8.775 ;
      RECT 57.94 3.52 58.11 3.69 ;
      RECT 57.9 1.415 58.07 1.585 ;
      RECT 57.9 4.135 58.07 4.305 ;
      RECT 57.885 7.055 58.055 7.225 ;
      RECT 57.885 7.795 58.055 7.965 ;
      RECT 57.525 2.76 57.695 2.93 ;
      RECT 57.51 6.315 57.68 6.485 ;
      RECT 57.44 1.415 57.61 1.585 ;
      RECT 57.44 4.135 57.61 4.305 ;
      RECT 57.265 8.605 57.435 8.775 ;
      RECT 57.175 2.235 57.345 2.405 ;
      RECT 56.995 3.55 57.165 3.72 ;
      RECT 56.98 1.415 57.15 1.585 ;
      RECT 56.98 4.135 57.15 4.305 ;
      RECT 56.715 2.865 56.885 3.035 ;
      RECT 56.585 8.605 56.755 8.775 ;
      RECT 56.52 1.415 56.69 1.585 ;
      RECT 56.52 4.135 56.69 4.305 ;
      RECT 56.515 5.945 56.685 6.115 ;
      RECT 56.395 2.49 56.565 2.66 ;
      RECT 56.06 1.415 56.23 1.585 ;
      RECT 56.06 4.135 56.23 4.305 ;
      RECT 55.705 1.97 55.875 2.14 ;
      RECT 55.63 2.44 55.8 2.61 ;
      RECT 55.6 1.415 55.77 1.585 ;
      RECT 55.6 4.135 55.77 4.305 ;
      RECT 55.14 1.415 55.31 1.585 ;
      RECT 55.14 4.135 55.31 4.305 ;
      RECT 54.78 2.165 54.95 2.335 ;
      RECT 54.68 1.415 54.85 1.585 ;
      RECT 54.68 4.135 54.85 4.305 ;
      RECT 54.44 3.36 54.61 3.53 ;
      RECT 54.405 2.695 54.575 2.865 ;
      RECT 54.22 1.415 54.39 1.585 ;
      RECT 54.22 4.135 54.39 4.305 ;
      RECT 53.795 2.55 53.965 2.72 ;
      RECT 53.76 1.415 53.93 1.585 ;
      RECT 53.76 4.135 53.93 4.305 ;
      RECT 53.725 3.25 53.895 3.42 ;
      RECT 53.665 2.085 53.835 2.255 ;
      RECT 53.3 1.415 53.47 1.585 ;
      RECT 53.3 4.135 53.47 4.305 ;
      RECT 53.025 3 53.195 3.17 ;
      RECT 52.84 1.415 53.01 1.585 ;
      RECT 52.84 4.135 53.01 4.305 ;
      RECT 52.52 2.505 52.69 2.675 ;
      RECT 52.38 1.415 52.55 1.585 ;
      RECT 52.38 4.135 52.55 4.305 ;
      RECT 52.3 3.25 52.47 3.42 ;
      RECT 52.095 2.13 52.265 2.3 ;
      RECT 51.92 1.415 52.09 1.585 ;
      RECT 51.92 4.135 52.09 4.305 ;
      RECT 51.825 3 51.995 3.17 ;
      RECT 51.785 2.43 51.955 2.6 ;
      RECT 51.46 1.415 51.63 1.585 ;
      RECT 51.46 4.135 51.63 4.305 ;
      RECT 51.24 3.475 51.41 3.645 ;
      RECT 51.1 2.095 51.27 2.265 ;
      RECT 51 1.415 51.17 1.585 ;
      RECT 51 4.135 51.17 4.305 ;
      RECT 50.54 1.415 50.71 1.585 ;
      RECT 50.54 4.135 50.71 4.305 ;
      RECT 50.53 3.015 50.7 3.185 ;
      RECT 49.665 0.915 49.835 1.085 ;
      RECT 49.665 2.395 49.835 2.565 ;
      RECT 49.665 6.315 49.835 6.485 ;
      RECT 49.665 7.795 49.835 7.965 ;
      RECT 49.315 0.105 49.485 0.275 ;
      RECT 49.315 4.165 49.485 4.335 ;
      RECT 49.315 4.545 49.485 4.715 ;
      RECT 49.315 8.605 49.485 8.775 ;
      RECT 49.295 2.765 49.465 2.935 ;
      RECT 49.295 5.945 49.465 6.115 ;
      RECT 48.675 0.915 48.845 1.085 ;
      RECT 48.675 2.395 48.845 2.565 ;
      RECT 48.675 6.315 48.845 6.485 ;
      RECT 48.675 7.795 48.845 7.965 ;
      RECT 48.325 0.105 48.495 0.275 ;
      RECT 48.325 4.165 48.495 4.335 ;
      RECT 48.325 4.545 48.495 4.715 ;
      RECT 48.325 8.605 48.495 8.775 ;
      RECT 48.305 2.765 48.475 2.935 ;
      RECT 48.305 5.945 48.475 6.115 ;
      RECT 47.62 0.105 47.79 0.275 ;
      RECT 47.62 4.165 47.79 4.335 ;
      RECT 47.62 4.545 47.79 4.715 ;
      RECT 47.62 8.605 47.79 8.775 ;
      RECT 47.31 2.025 47.48 2.195 ;
      RECT 47.31 6.685 47.48 6.855 ;
      RECT 46.94 0.105 47.11 0.275 ;
      RECT 46.94 8.605 47.11 8.775 ;
      RECT 46.88 0.915 47.05 1.085 ;
      RECT 46.88 1.655 47.05 1.825 ;
      RECT 46.88 7.055 47.05 7.225 ;
      RECT 46.88 7.795 47.05 7.965 ;
      RECT 46.505 2.395 46.675 2.565 ;
      RECT 46.505 6.315 46.675 6.485 ;
      RECT 46.26 0.105 46.43 0.275 ;
      RECT 46.26 8.605 46.43 8.775 ;
      RECT 45.58 0.105 45.75 0.275 ;
      RECT 45.58 8.605 45.75 8.775 ;
      RECT 45.51 2.765 45.68 2.935 ;
      RECT 45.51 5.945 45.68 6.115 ;
      RECT 43.955 1.415 44.125 1.585 ;
      RECT 43.955 4.135 44.125 4.305 ;
      RECT 43.585 2.875 43.755 3.045 ;
      RECT 43.495 1.415 43.665 1.585 ;
      RECT 43.495 4.135 43.665 4.305 ;
      RECT 43.265 2.045 43.435 2.215 ;
      RECT 43.12 2.485 43.29 2.655 ;
      RECT 43.035 1.415 43.205 1.585 ;
      RECT 43.035 4.135 43.205 4.305 ;
      RECT 42.84 4.545 43.01 4.715 ;
      RECT 42.84 8.605 43.01 8.775 ;
      RECT 42.575 1.415 42.745 1.585 ;
      RECT 42.575 4.135 42.745 4.305 ;
      RECT 42.53 6.685 42.7 6.855 ;
      RECT 42.51 2.525 42.68 2.695 ;
      RECT 42.165 2.16 42.335 2.33 ;
      RECT 42.16 8.605 42.33 8.775 ;
      RECT 42.155 3.52 42.325 3.69 ;
      RECT 42.115 1.415 42.285 1.585 ;
      RECT 42.115 4.135 42.285 4.305 ;
      RECT 42.1 7.055 42.27 7.225 ;
      RECT 42.1 7.795 42.27 7.965 ;
      RECT 41.74 2.76 41.91 2.93 ;
      RECT 41.725 6.315 41.895 6.485 ;
      RECT 41.655 1.415 41.825 1.585 ;
      RECT 41.655 4.135 41.825 4.305 ;
      RECT 41.48 8.605 41.65 8.775 ;
      RECT 41.39 2.235 41.56 2.405 ;
      RECT 41.21 3.55 41.38 3.72 ;
      RECT 41.195 1.415 41.365 1.585 ;
      RECT 41.195 4.135 41.365 4.305 ;
      RECT 40.93 2.865 41.1 3.035 ;
      RECT 40.8 8.605 40.97 8.775 ;
      RECT 40.735 1.415 40.905 1.585 ;
      RECT 40.735 4.135 40.905 4.305 ;
      RECT 40.73 5.945 40.9 6.115 ;
      RECT 40.61 2.49 40.78 2.66 ;
      RECT 40.275 1.415 40.445 1.585 ;
      RECT 40.275 4.135 40.445 4.305 ;
      RECT 39.92 1.97 40.09 2.14 ;
      RECT 39.845 2.44 40.015 2.61 ;
      RECT 39.815 1.415 39.985 1.585 ;
      RECT 39.815 4.135 39.985 4.305 ;
      RECT 39.355 1.415 39.525 1.585 ;
      RECT 39.355 4.135 39.525 4.305 ;
      RECT 38.995 2.165 39.165 2.335 ;
      RECT 38.895 1.415 39.065 1.585 ;
      RECT 38.895 4.135 39.065 4.305 ;
      RECT 38.655 3.36 38.825 3.53 ;
      RECT 38.62 2.695 38.79 2.865 ;
      RECT 38.435 1.415 38.605 1.585 ;
      RECT 38.435 4.135 38.605 4.305 ;
      RECT 38.01 2.55 38.18 2.72 ;
      RECT 37.975 1.415 38.145 1.585 ;
      RECT 37.975 4.135 38.145 4.305 ;
      RECT 37.94 3.25 38.11 3.42 ;
      RECT 37.88 2.085 38.05 2.255 ;
      RECT 37.515 1.415 37.685 1.585 ;
      RECT 37.515 4.135 37.685 4.305 ;
      RECT 37.24 3 37.41 3.17 ;
      RECT 37.055 1.415 37.225 1.585 ;
      RECT 37.055 4.135 37.225 4.305 ;
      RECT 36.735 2.505 36.905 2.675 ;
      RECT 36.595 1.415 36.765 1.585 ;
      RECT 36.595 4.135 36.765 4.305 ;
      RECT 36.515 3.25 36.685 3.42 ;
      RECT 36.31 2.13 36.48 2.3 ;
      RECT 36.135 1.415 36.305 1.585 ;
      RECT 36.135 4.135 36.305 4.305 ;
      RECT 36.04 3 36.21 3.17 ;
      RECT 36 2.43 36.17 2.6 ;
      RECT 35.675 1.415 35.845 1.585 ;
      RECT 35.675 4.135 35.845 4.305 ;
      RECT 35.455 3.475 35.625 3.645 ;
      RECT 35.315 2.095 35.485 2.265 ;
      RECT 35.215 1.415 35.385 1.585 ;
      RECT 35.215 4.135 35.385 4.305 ;
      RECT 34.755 1.415 34.925 1.585 ;
      RECT 34.755 4.135 34.925 4.305 ;
      RECT 34.745 3.015 34.915 3.185 ;
      RECT 33.89 0.915 34.06 1.085 ;
      RECT 33.89 2.395 34.06 2.565 ;
      RECT 33.89 6.315 34.06 6.485 ;
      RECT 33.89 7.795 34.06 7.965 ;
      RECT 33.54 0.105 33.71 0.275 ;
      RECT 33.54 4.165 33.71 4.335 ;
      RECT 33.54 4.545 33.71 4.715 ;
      RECT 33.54 8.605 33.71 8.775 ;
      RECT 33.52 2.765 33.69 2.935 ;
      RECT 33.52 5.945 33.69 6.115 ;
      RECT 32.9 0.915 33.07 1.085 ;
      RECT 32.9 2.395 33.07 2.565 ;
      RECT 32.9 6.315 33.07 6.485 ;
      RECT 32.9 7.795 33.07 7.965 ;
      RECT 32.55 0.105 32.72 0.275 ;
      RECT 32.55 4.165 32.72 4.335 ;
      RECT 32.55 4.545 32.72 4.715 ;
      RECT 32.55 8.605 32.72 8.775 ;
      RECT 32.53 2.765 32.7 2.935 ;
      RECT 32.53 5.945 32.7 6.115 ;
      RECT 31.845 0.105 32.015 0.275 ;
      RECT 31.845 4.165 32.015 4.335 ;
      RECT 31.845 4.545 32.015 4.715 ;
      RECT 31.845 8.605 32.015 8.775 ;
      RECT 31.535 2.025 31.705 2.195 ;
      RECT 31.535 6.685 31.705 6.855 ;
      RECT 31.165 0.105 31.335 0.275 ;
      RECT 31.165 8.605 31.335 8.775 ;
      RECT 31.105 0.915 31.275 1.085 ;
      RECT 31.105 1.655 31.275 1.825 ;
      RECT 31.105 7.055 31.275 7.225 ;
      RECT 31.105 7.795 31.275 7.965 ;
      RECT 30.73 2.395 30.9 2.565 ;
      RECT 30.73 6.315 30.9 6.485 ;
      RECT 30.485 0.105 30.655 0.275 ;
      RECT 30.485 8.605 30.655 8.775 ;
      RECT 29.805 0.105 29.975 0.275 ;
      RECT 29.805 8.605 29.975 8.775 ;
      RECT 29.735 2.765 29.905 2.935 ;
      RECT 29.735 5.945 29.905 6.115 ;
      RECT 28.18 1.415 28.35 1.585 ;
      RECT 28.18 4.135 28.35 4.305 ;
      RECT 27.81 2.875 27.98 3.045 ;
      RECT 27.72 1.415 27.89 1.585 ;
      RECT 27.72 4.135 27.89 4.305 ;
      RECT 27.49 2.045 27.66 2.215 ;
      RECT 27.345 2.485 27.515 2.655 ;
      RECT 27.26 1.415 27.43 1.585 ;
      RECT 27.26 4.135 27.43 4.305 ;
      RECT 27.065 4.545 27.235 4.715 ;
      RECT 27.065 8.605 27.235 8.775 ;
      RECT 26.8 1.415 26.97 1.585 ;
      RECT 26.8 4.135 26.97 4.305 ;
      RECT 26.755 6.685 26.925 6.855 ;
      RECT 26.735 2.525 26.905 2.695 ;
      RECT 26.39 2.16 26.56 2.33 ;
      RECT 26.385 8.605 26.555 8.775 ;
      RECT 26.38 3.52 26.55 3.69 ;
      RECT 26.34 1.415 26.51 1.585 ;
      RECT 26.34 4.135 26.51 4.305 ;
      RECT 26.325 7.055 26.495 7.225 ;
      RECT 26.325 7.795 26.495 7.965 ;
      RECT 25.965 2.76 26.135 2.93 ;
      RECT 25.95 6.315 26.12 6.485 ;
      RECT 25.88 1.415 26.05 1.585 ;
      RECT 25.88 4.135 26.05 4.305 ;
      RECT 25.705 8.605 25.875 8.775 ;
      RECT 25.615 2.235 25.785 2.405 ;
      RECT 25.435 3.55 25.605 3.72 ;
      RECT 25.42 1.415 25.59 1.585 ;
      RECT 25.42 4.135 25.59 4.305 ;
      RECT 25.155 2.865 25.325 3.035 ;
      RECT 25.025 8.605 25.195 8.775 ;
      RECT 24.96 1.415 25.13 1.585 ;
      RECT 24.96 4.135 25.13 4.305 ;
      RECT 24.955 5.945 25.125 6.115 ;
      RECT 24.835 2.49 25.005 2.66 ;
      RECT 24.5 1.415 24.67 1.585 ;
      RECT 24.5 4.135 24.67 4.305 ;
      RECT 24.145 1.97 24.315 2.14 ;
      RECT 24.07 2.44 24.24 2.61 ;
      RECT 24.04 1.415 24.21 1.585 ;
      RECT 24.04 4.135 24.21 4.305 ;
      RECT 23.58 1.415 23.75 1.585 ;
      RECT 23.58 4.135 23.75 4.305 ;
      RECT 23.22 2.165 23.39 2.335 ;
      RECT 23.12 1.415 23.29 1.585 ;
      RECT 23.12 4.135 23.29 4.305 ;
      RECT 22.88 3.36 23.05 3.53 ;
      RECT 22.845 2.695 23.015 2.865 ;
      RECT 22.66 1.415 22.83 1.585 ;
      RECT 22.66 4.135 22.83 4.305 ;
      RECT 22.235 2.55 22.405 2.72 ;
      RECT 22.2 1.415 22.37 1.585 ;
      RECT 22.2 4.135 22.37 4.305 ;
      RECT 22.165 3.25 22.335 3.42 ;
      RECT 22.105 2.085 22.275 2.255 ;
      RECT 21.74 1.415 21.91 1.585 ;
      RECT 21.74 4.135 21.91 4.305 ;
      RECT 21.465 3 21.635 3.17 ;
      RECT 21.28 1.415 21.45 1.585 ;
      RECT 21.28 4.135 21.45 4.305 ;
      RECT 20.96 2.505 21.13 2.675 ;
      RECT 20.82 1.415 20.99 1.585 ;
      RECT 20.82 4.135 20.99 4.305 ;
      RECT 20.74 3.25 20.91 3.42 ;
      RECT 20.535 2.13 20.705 2.3 ;
      RECT 20.36 1.415 20.53 1.585 ;
      RECT 20.36 4.135 20.53 4.305 ;
      RECT 20.265 3 20.435 3.17 ;
      RECT 20.225 2.43 20.395 2.6 ;
      RECT 19.9 1.415 20.07 1.585 ;
      RECT 19.9 4.135 20.07 4.305 ;
      RECT 19.68 3.475 19.85 3.645 ;
      RECT 19.54 2.095 19.71 2.265 ;
      RECT 19.44 1.415 19.61 1.585 ;
      RECT 19.44 4.135 19.61 4.305 ;
      RECT 18.98 1.415 19.15 1.585 ;
      RECT 18.98 4.135 19.15 4.305 ;
      RECT 18.97 3.015 19.14 3.185 ;
      RECT 18.11 0.915 18.28 1.085 ;
      RECT 18.11 2.395 18.28 2.565 ;
      RECT 18.11 6.315 18.28 6.485 ;
      RECT 18.11 7.795 18.28 7.965 ;
      RECT 17.76 0.105 17.93 0.275 ;
      RECT 17.76 4.165 17.93 4.335 ;
      RECT 17.76 4.545 17.93 4.715 ;
      RECT 17.76 8.605 17.93 8.775 ;
      RECT 17.74 2.765 17.91 2.935 ;
      RECT 17.74 5.945 17.91 6.115 ;
      RECT 17.12 0.915 17.29 1.085 ;
      RECT 17.12 2.395 17.29 2.565 ;
      RECT 17.12 6.315 17.29 6.485 ;
      RECT 17.12 7.795 17.29 7.965 ;
      RECT 16.77 0.105 16.94 0.275 ;
      RECT 16.77 4.165 16.94 4.335 ;
      RECT 16.77 4.545 16.94 4.715 ;
      RECT 16.77 8.605 16.94 8.775 ;
      RECT 16.75 2.765 16.92 2.935 ;
      RECT 16.75 5.945 16.92 6.115 ;
      RECT 16.065 0.105 16.235 0.275 ;
      RECT 16.065 4.165 16.235 4.335 ;
      RECT 16.065 4.545 16.235 4.715 ;
      RECT 16.065 8.605 16.235 8.775 ;
      RECT 15.755 2.025 15.925 2.195 ;
      RECT 15.755 6.685 15.925 6.855 ;
      RECT 15.385 0.105 15.555 0.275 ;
      RECT 15.385 8.605 15.555 8.775 ;
      RECT 15.325 0.915 15.495 1.085 ;
      RECT 15.325 1.655 15.495 1.825 ;
      RECT 15.325 7.055 15.495 7.225 ;
      RECT 15.325 7.795 15.495 7.965 ;
      RECT 14.95 2.395 15.12 2.565 ;
      RECT 14.95 6.315 15.12 6.485 ;
      RECT 14.705 0.105 14.875 0.275 ;
      RECT 14.705 8.605 14.875 8.775 ;
      RECT 14.025 0.105 14.195 0.275 ;
      RECT 14.025 8.605 14.195 8.775 ;
      RECT 13.955 2.765 14.125 2.935 ;
      RECT 13.955 5.945 14.125 6.115 ;
      RECT 12.4 1.415 12.57 1.585 ;
      RECT 12.4 4.135 12.57 4.305 ;
      RECT 12.03 2.875 12.2 3.045 ;
      RECT 11.94 1.415 12.11 1.585 ;
      RECT 11.94 4.135 12.11 4.305 ;
      RECT 11.71 2.045 11.88 2.215 ;
      RECT 11.565 2.485 11.735 2.655 ;
      RECT 11.48 1.415 11.65 1.585 ;
      RECT 11.48 4.135 11.65 4.305 ;
      RECT 11.285 4.545 11.455 4.715 ;
      RECT 11.285 8.605 11.455 8.775 ;
      RECT 11.02 1.415 11.19 1.585 ;
      RECT 11.02 4.135 11.19 4.305 ;
      RECT 10.975 6.685 11.145 6.855 ;
      RECT 10.955 2.525 11.125 2.695 ;
      RECT 10.61 2.16 10.78 2.33 ;
      RECT 10.605 8.605 10.775 8.775 ;
      RECT 10.6 3.52 10.77 3.69 ;
      RECT 10.56 1.415 10.73 1.585 ;
      RECT 10.56 4.135 10.73 4.305 ;
      RECT 10.545 7.055 10.715 7.225 ;
      RECT 10.545 7.795 10.715 7.965 ;
      RECT 10.185 2.76 10.355 2.93 ;
      RECT 10.17 6.315 10.34 6.485 ;
      RECT 10.1 1.415 10.27 1.585 ;
      RECT 10.1 4.135 10.27 4.305 ;
      RECT 9.925 8.605 10.095 8.775 ;
      RECT 9.835 2.235 10.005 2.405 ;
      RECT 9.655 3.55 9.825 3.72 ;
      RECT 9.64 1.415 9.81 1.585 ;
      RECT 9.64 4.135 9.81 4.305 ;
      RECT 9.375 2.865 9.545 3.035 ;
      RECT 9.245 8.605 9.415 8.775 ;
      RECT 9.18 1.415 9.35 1.585 ;
      RECT 9.18 4.135 9.35 4.305 ;
      RECT 9.175 5.945 9.345 6.115 ;
      RECT 9.055 2.49 9.225 2.66 ;
      RECT 8.72 1.415 8.89 1.585 ;
      RECT 8.72 4.135 8.89 4.305 ;
      RECT 8.365 1.97 8.535 2.14 ;
      RECT 8.29 2.44 8.46 2.61 ;
      RECT 8.26 1.415 8.43 1.585 ;
      RECT 8.26 4.135 8.43 4.305 ;
      RECT 7.8 1.415 7.97 1.585 ;
      RECT 7.8 4.135 7.97 4.305 ;
      RECT 7.44 2.165 7.61 2.335 ;
      RECT 7.34 1.415 7.51 1.585 ;
      RECT 7.34 4.135 7.51 4.305 ;
      RECT 7.1 3.36 7.27 3.53 ;
      RECT 7.065 2.695 7.235 2.865 ;
      RECT 6.88 1.415 7.05 1.585 ;
      RECT 6.88 4.135 7.05 4.305 ;
      RECT 6.455 2.55 6.625 2.72 ;
      RECT 6.42 1.415 6.59 1.585 ;
      RECT 6.42 4.135 6.59 4.305 ;
      RECT 6.385 3.25 6.555 3.42 ;
      RECT 6.325 2.085 6.495 2.255 ;
      RECT 5.96 1.415 6.13 1.585 ;
      RECT 5.96 4.135 6.13 4.305 ;
      RECT 5.685 3 5.855 3.17 ;
      RECT 5.5 1.415 5.67 1.585 ;
      RECT 5.5 4.135 5.67 4.305 ;
      RECT 5.18 2.505 5.35 2.675 ;
      RECT 5.04 1.415 5.21 1.585 ;
      RECT 5.04 4.135 5.21 4.305 ;
      RECT 4.96 3.25 5.13 3.42 ;
      RECT 4.755 2.13 4.925 2.3 ;
      RECT 4.58 1.415 4.75 1.585 ;
      RECT 4.58 4.135 4.75 4.305 ;
      RECT 4.485 3 4.655 3.17 ;
      RECT 4.445 2.43 4.615 2.6 ;
      RECT 4.12 1.415 4.29 1.585 ;
      RECT 4.12 4.135 4.29 4.305 ;
      RECT 3.9 3.475 4.07 3.645 ;
      RECT 3.76 2.095 3.93 2.265 ;
      RECT 3.66 1.415 3.83 1.585 ;
      RECT 3.66 4.135 3.83 4.305 ;
      RECT 3.2 1.415 3.37 1.585 ;
      RECT 3.2 4.135 3.37 4.305 ;
      RECT 3.19 3.015 3.36 3.185 ;
      RECT 2.35 4.545 2.52 4.715 ;
      RECT 2.35 8.605 2.52 8.775 ;
      RECT 2.04 6.685 2.21 6.855 ;
      RECT 1.67 8.605 1.84 8.775 ;
      RECT 1.61 7.055 1.78 7.225 ;
      RECT 1.61 7.795 1.78 7.965 ;
      RECT 1.235 6.315 1.405 6.485 ;
      RECT 0.99 8.605 1.16 8.775 ;
      RECT 0.94 4.335 1.11 4.505 ;
      RECT 0.885 0.065 1.055 0.235 ;
      RECT 0.24 5.945 0.41 6.115 ;
    LAYER li ;
      RECT 74.31 0 74.48 2.085 ;
      RECT 72.35 0 72.52 2.085 ;
      RECT 69.91 0 70.08 2.085 ;
      RECT 68.95 0 69.12 2.085 ;
      RECT 68.43 0 68.6 2.085 ;
      RECT 67.47 0 67.64 2.085 ;
      RECT 66.51 0 66.68 2.085 ;
      RECT 58.525 0 58.695 2.085 ;
      RECT 56.565 0 56.735 2.085 ;
      RECT 54.125 0 54.295 2.085 ;
      RECT 53.165 0 53.335 2.085 ;
      RECT 52.645 0 52.815 2.085 ;
      RECT 51.685 0 51.855 2.085 ;
      RECT 50.725 0 50.895 2.085 ;
      RECT 42.74 0 42.91 2.085 ;
      RECT 40.78 0 40.95 2.085 ;
      RECT 38.34 0 38.51 2.085 ;
      RECT 37.38 0 37.55 2.085 ;
      RECT 36.86 0 37.03 2.085 ;
      RECT 35.9 0 36.07 2.085 ;
      RECT 34.94 0 35.11 2.085 ;
      RECT 26.965 0 27.135 2.085 ;
      RECT 25.005 0 25.175 2.085 ;
      RECT 22.565 0 22.735 2.085 ;
      RECT 21.605 0 21.775 2.085 ;
      RECT 21.085 0 21.255 2.085 ;
      RECT 20.125 0 20.295 2.085 ;
      RECT 19.165 0 19.335 2.085 ;
      RECT 11.185 0 11.355 2.085 ;
      RECT 9.225 0 9.395 2.085 ;
      RECT 6.785 0 6.955 2.085 ;
      RECT 5.825 0 5.995 2.085 ;
      RECT 5.305 0 5.475 2.085 ;
      RECT 4.345 0 4.515 2.085 ;
      RECT 3.385 0 3.555 2.085 ;
      RECT 66.295 0 75.895 1.59 ;
      RECT 50.51 0 60.11 1.59 ;
      RECT 34.725 0 44.325 1.59 ;
      RECT 18.95 0 28.55 1.59 ;
      RECT 3.17 0 12.77 1.59 ;
      RECT 66.18 1.415 76.01 1.585 ;
      RECT 66.295 0 76.01 1.585 ;
      RECT 50.395 1.415 60.225 1.585 ;
      RECT 50.51 0 60.225 1.585 ;
      RECT 34.61 1.415 44.44 1.585 ;
      RECT 34.725 0 44.44 1.585 ;
      RECT 18.835 1.415 28.665 1.585 ;
      RECT 18.95 0 28.665 1.585 ;
      RECT 3.055 1.415 12.885 1.585 ;
      RECT 3.17 0 12.885 1.585 ;
      RECT 80.805 0 80.975 0.935 ;
      RECT 79.815 0 79.985 0.935 ;
      RECT 77.07 0 77.24 0.935 ;
      RECT 65.02 0 65.19 0.935 ;
      RECT 64.03 0 64.2 0.935 ;
      RECT 61.285 0 61.455 0.935 ;
      RECT 49.235 0 49.405 0.935 ;
      RECT 48.245 0 48.415 0.935 ;
      RECT 45.5 0 45.67 0.935 ;
      RECT 33.46 0 33.63 0.935 ;
      RECT 32.47 0 32.64 0.935 ;
      RECT 29.725 0 29.895 0.935 ;
      RECT 17.68 0 17.85 0.935 ;
      RECT 16.69 0 16.86 0.935 ;
      RECT 13.945 0 14.115 0.935 ;
      RECT 0.885 0 1.055 0.355 ;
      RECT 0 0 81.775 0.305 ;
      RECT 2.04 4.135 2.21 8.305 ;
      RECT 80.805 3.405 80.975 5.475 ;
      RECT 79.815 3.405 79.985 5.475 ;
      RECT 77.07 3.405 77.24 5.475 ;
      RECT 72.29 4.135 72.46 5.475 ;
      RECT 65.02 3.405 65.19 5.475 ;
      RECT 64.03 3.405 64.2 5.475 ;
      RECT 61.285 3.405 61.455 5.475 ;
      RECT 56.505 4.135 56.675 5.475 ;
      RECT 49.235 3.405 49.405 5.475 ;
      RECT 48.245 3.405 48.415 5.475 ;
      RECT 45.5 3.405 45.67 5.475 ;
      RECT 40.72 4.135 40.89 5.475 ;
      RECT 33.46 3.405 33.63 5.475 ;
      RECT 32.47 3.405 32.64 5.475 ;
      RECT 29.725 3.405 29.895 5.475 ;
      RECT 24.945 4.135 25.115 5.475 ;
      RECT 17.68 3.405 17.85 5.475 ;
      RECT 16.69 3.405 16.86 5.475 ;
      RECT 13.945 3.405 14.115 5.475 ;
      RECT 9.165 4.135 9.335 5.475 ;
      RECT 0.23 4.135 0.4 5.475 ;
      RECT 0 4.135 81.775 4.745 ;
      RECT 75.27 3.635 75.44 4.745 ;
      RECT 74.31 3.635 74.48 4.745 ;
      RECT 71.87 3.635 72.04 4.745 ;
      RECT 70.87 3.635 71.04 4.745 ;
      RECT 69.91 3.635 70.08 4.745 ;
      RECT 67.47 3.635 67.64 4.745 ;
      RECT 59.485 3.635 59.655 4.745 ;
      RECT 58.525 3.635 58.695 4.745 ;
      RECT 56.085 3.635 56.255 4.745 ;
      RECT 55.085 3.635 55.255 4.745 ;
      RECT 54.125 3.635 54.295 4.745 ;
      RECT 51.685 3.635 51.855 4.745 ;
      RECT 43.7 3.635 43.87 4.745 ;
      RECT 42.74 3.635 42.91 4.745 ;
      RECT 40.3 3.635 40.47 4.745 ;
      RECT 39.3 3.635 39.47 4.745 ;
      RECT 38.34 3.635 38.51 4.745 ;
      RECT 35.9 3.635 36.07 4.745 ;
      RECT 27.925 3.635 28.095 4.745 ;
      RECT 26.965 3.635 27.135 4.745 ;
      RECT 24.525 3.635 24.695 4.745 ;
      RECT 23.525 3.635 23.695 4.745 ;
      RECT 22.565 3.635 22.735 4.745 ;
      RECT 20.125 3.635 20.295 4.745 ;
      RECT 12.145 3.635 12.315 4.745 ;
      RECT 11.185 3.635 11.355 4.745 ;
      RECT 8.745 3.635 8.915 4.745 ;
      RECT 7.745 3.635 7.915 4.745 ;
      RECT 6.785 3.635 6.955 4.745 ;
      RECT 4.345 3.635 4.515 4.745 ;
      RECT -0.005 8.575 81.775 8.88 ;
      RECT 80.805 7.945 80.975 8.88 ;
      RECT 79.815 7.945 79.985 8.88 ;
      RECT 77.07 7.945 77.24 8.88 ;
      RECT 72.29 7.945 72.46 8.88 ;
      RECT 65.02 7.945 65.19 8.88 ;
      RECT 64.03 7.945 64.2 8.88 ;
      RECT 61.285 7.945 61.455 8.88 ;
      RECT 56.505 7.945 56.675 8.88 ;
      RECT 49.235 7.945 49.405 8.88 ;
      RECT 48.245 7.945 48.415 8.88 ;
      RECT 45.5 7.945 45.67 8.88 ;
      RECT 40.72 7.945 40.89 8.88 ;
      RECT 33.46 7.945 33.63 8.88 ;
      RECT 32.47 7.945 32.64 8.88 ;
      RECT 29.725 7.945 29.895 8.88 ;
      RECT 24.945 7.945 25.115 8.88 ;
      RECT 17.68 7.945 17.85 8.88 ;
      RECT 16.69 7.945 16.86 8.88 ;
      RECT 13.945 7.945 14.115 8.88 ;
      RECT 9.165 7.945 9.335 8.88 ;
      RECT 0.23 7.945 0.4 8.88 ;
      RECT 80.865 1.74 81.035 2.935 ;
      RECT 80.865 1.74 81.33 1.91 ;
      RECT 80.865 6.97 81.33 7.14 ;
      RECT 80.865 5.945 81.035 7.14 ;
      RECT 79.875 1.74 80.045 2.935 ;
      RECT 79.875 1.74 80.34 1.91 ;
      RECT 79.875 6.97 80.34 7.14 ;
      RECT 79.875 5.945 80.045 7.14 ;
      RECT 78.02 2.635 78.19 3.865 ;
      RECT 78.075 0.855 78.245 2.805 ;
      RECT 78.02 0.575 78.19 1.025 ;
      RECT 78.02 7.855 78.19 8.305 ;
      RECT 78.075 6.075 78.245 8.025 ;
      RECT 78.02 5.015 78.19 6.245 ;
      RECT 77.5 0.575 77.67 3.865 ;
      RECT 77.5 2.075 77.905 2.405 ;
      RECT 77.5 1.235 77.905 1.565 ;
      RECT 77.5 5.015 77.67 8.305 ;
      RECT 77.5 7.315 77.905 7.645 ;
      RECT 77.5 6.475 77.905 6.805 ;
      RECT 74.835 1.975 75.565 2.215 ;
      RECT 75.377 1.77 75.565 2.215 ;
      RECT 75.205 1.782 75.58 2.209 ;
      RECT 75.12 1.797 75.6 2.194 ;
      RECT 75.12 1.812 75.605 2.184 ;
      RECT 75.075 1.832 75.62 2.176 ;
      RECT 75.052 1.867 75.635 2.13 ;
      RECT 74.966 1.89 75.64 2.09 ;
      RECT 74.966 1.908 75.65 2.06 ;
      RECT 74.835 1.977 75.655 2.023 ;
      RECT 74.88 1.92 75.65 2.06 ;
      RECT 74.966 1.872 75.635 2.13 ;
      RECT 75.052 1.841 75.62 2.176 ;
      RECT 75.075 1.822 75.605 2.184 ;
      RECT 75.12 1.795 75.58 2.209 ;
      RECT 75.205 1.777 75.565 2.215 ;
      RECT 75.291 1.771 75.565 2.215 ;
      RECT 75.377 1.766 75.51 2.215 ;
      RECT 75.463 1.761 75.51 2.215 ;
      RECT 75.155 2.659 75.325 3.045 ;
      RECT 75.15 2.659 75.325 3.04 ;
      RECT 75.125 2.659 75.325 3.005 ;
      RECT 75.125 2.687 75.335 2.995 ;
      RECT 75.105 2.687 75.335 2.955 ;
      RECT 75.1 2.687 75.335 2.928 ;
      RECT 75.1 2.705 75.34 2.92 ;
      RECT 75.045 2.705 75.34 2.855 ;
      RECT 75.045 2.722 75.35 2.838 ;
      RECT 75.035 2.722 75.35 2.778 ;
      RECT 75.035 2.739 75.355 2.775 ;
      RECT 75.03 2.575 75.2 2.753 ;
      RECT 75.03 2.609 75.286 2.753 ;
      RECT 75.025 3.375 75.03 3.388 ;
      RECT 75.02 3.27 75.025 3.393 ;
      RECT 74.995 3.13 75.02 3.408 ;
      RECT 74.96 3.081 74.995 3.44 ;
      RECT 74.955 3.049 74.96 3.46 ;
      RECT 74.95 3.04 74.955 3.46 ;
      RECT 74.87 3.005 74.95 3.46 ;
      RECT 74.807 2.975 74.87 3.46 ;
      RECT 74.721 2.963 74.807 3.46 ;
      RECT 74.635 2.949 74.721 3.46 ;
      RECT 74.555 2.936 74.635 3.446 ;
      RECT 74.52 2.928 74.555 3.426 ;
      RECT 74.51 2.925 74.52 3.417 ;
      RECT 74.48 2.92 74.51 3.404 ;
      RECT 74.43 2.895 74.48 3.38 ;
      RECT 74.416 2.869 74.43 3.362 ;
      RECT 74.33 2.829 74.416 3.338 ;
      RECT 74.285 2.777 74.33 3.307 ;
      RECT 74.275 2.752 74.285 3.294 ;
      RECT 74.27 2.533 74.275 2.555 ;
      RECT 74.265 2.735 74.275 3.29 ;
      RECT 74.265 2.531 74.27 2.645 ;
      RECT 74.255 2.527 74.265 3.286 ;
      RECT 74.211 2.525 74.255 3.274 ;
      RECT 74.125 2.525 74.211 3.245 ;
      RECT 74.095 2.525 74.125 3.218 ;
      RECT 74.08 2.525 74.095 3.206 ;
      RECT 74.04 2.537 74.08 3.191 ;
      RECT 74.02 2.556 74.04 3.17 ;
      RECT 74.01 2.566 74.02 3.154 ;
      RECT 74 2.572 74.01 3.143 ;
      RECT 73.98 2.582 74 3.126 ;
      RECT 73.975 2.591 73.98 3.113 ;
      RECT 73.97 2.595 73.975 3.063 ;
      RECT 73.96 2.601 73.97 2.98 ;
      RECT 73.955 2.605 73.96 2.894 ;
      RECT 73.95 2.625 73.955 2.831 ;
      RECT 73.945 2.648 73.95 2.778 ;
      RECT 73.94 2.666 73.945 2.723 ;
      RECT 74.55 2.485 74.72 2.745 ;
      RECT 74.72 2.45 74.765 2.731 ;
      RECT 74.681 2.452 74.77 2.714 ;
      RECT 74.57 2.469 74.856 2.685 ;
      RECT 74.57 2.484 74.86 2.657 ;
      RECT 74.57 2.465 74.77 2.714 ;
      RECT 74.595 2.453 74.72 2.745 ;
      RECT 74.681 2.451 74.765 2.731 ;
      RECT 73.735 1.84 73.905 2.33 ;
      RECT 73.735 1.84 73.94 2.31 ;
      RECT 73.87 1.76 73.98 2.27 ;
      RECT 73.851 1.764 74 2.24 ;
      RECT 73.765 1.772 74.02 2.223 ;
      RECT 73.765 1.778 74.025 2.213 ;
      RECT 73.765 1.787 74.045 2.201 ;
      RECT 73.74 1.812 74.075 2.179 ;
      RECT 73.74 1.832 74.08 2.159 ;
      RECT 73.735 1.845 74.09 2.139 ;
      RECT 73.735 1.912 74.095 2.12 ;
      RECT 73.735 2.045 74.1 2.107 ;
      RECT 73.73 1.85 74.09 1.94 ;
      RECT 73.74 1.807 74.045 2.201 ;
      RECT 73.851 1.762 73.98 2.27 ;
      RECT 73.725 3.515 74.025 3.77 ;
      RECT 73.81 3.481 74.025 3.77 ;
      RECT 73.81 3.484 74.03 3.63 ;
      RECT 73.745 3.505 74.03 3.63 ;
      RECT 73.78 3.495 74.025 3.77 ;
      RECT 73.775 3.5 74.03 3.63 ;
      RECT 73.81 3.479 74.011 3.77 ;
      RECT 73.896 3.47 74.011 3.77 ;
      RECT 73.896 3.464 73.925 3.77 ;
      RECT 73.385 3.105 73.395 3.595 ;
      RECT 73.045 3.04 73.055 3.34 ;
      RECT 73.56 3.212 73.565 3.431 ;
      RECT 73.55 3.192 73.56 3.448 ;
      RECT 73.54 3.172 73.55 3.478 ;
      RECT 73.535 3.162 73.54 3.493 ;
      RECT 73.53 3.158 73.535 3.498 ;
      RECT 73.515 3.15 73.53 3.505 ;
      RECT 73.475 3.13 73.515 3.53 ;
      RECT 73.45 3.112 73.475 3.563 ;
      RECT 73.445 3.11 73.45 3.576 ;
      RECT 73.425 3.107 73.445 3.58 ;
      RECT 73.395 3.105 73.425 3.59 ;
      RECT 73.325 3.107 73.385 3.591 ;
      RECT 73.305 3.107 73.325 3.585 ;
      RECT 73.28 3.105 73.305 3.582 ;
      RECT 73.245 3.1 73.28 3.578 ;
      RECT 73.225 3.094 73.245 3.565 ;
      RECT 73.215 3.091 73.225 3.553 ;
      RECT 73.195 3.088 73.215 3.538 ;
      RECT 73.175 3.084 73.195 3.52 ;
      RECT 73.17 3.081 73.175 3.51 ;
      RECT 73.165 3.08 73.17 3.508 ;
      RECT 73.155 3.077 73.165 3.5 ;
      RECT 73.145 3.071 73.155 3.483 ;
      RECT 73.135 3.065 73.145 3.465 ;
      RECT 73.125 3.059 73.135 3.453 ;
      RECT 73.115 3.053 73.125 3.433 ;
      RECT 73.11 3.049 73.115 3.418 ;
      RECT 73.105 3.047 73.11 3.41 ;
      RECT 73.1 3.045 73.105 3.403 ;
      RECT 73.095 3.043 73.1 3.393 ;
      RECT 73.09 3.041 73.095 3.387 ;
      RECT 73.08 3.04 73.09 3.377 ;
      RECT 73.07 3.04 73.08 3.368 ;
      RECT 73.055 3.04 73.07 3.353 ;
      RECT 73.015 3.04 73.045 3.337 ;
      RECT 72.995 3.042 73.015 3.332 ;
      RECT 72.99 3.047 72.995 3.33 ;
      RECT 72.96 3.055 72.99 3.328 ;
      RECT 72.93 3.07 72.96 3.327 ;
      RECT 72.885 3.092 72.93 3.332 ;
      RECT 72.88 3.107 72.885 3.336 ;
      RECT 72.865 3.112 72.88 3.338 ;
      RECT 72.86 3.116 72.865 3.34 ;
      RECT 72.8 3.139 72.86 3.349 ;
      RECT 72.78 3.165 72.8 3.362 ;
      RECT 72.77 3.172 72.78 3.366 ;
      RECT 72.755 3.179 72.77 3.369 ;
      RECT 72.735 3.189 72.755 3.372 ;
      RECT 72.73 3.197 72.735 3.375 ;
      RECT 72.685 3.202 72.73 3.382 ;
      RECT 72.675 3.205 72.685 3.389 ;
      RECT 72.665 3.205 72.675 3.393 ;
      RECT 72.63 3.207 72.665 3.405 ;
      RECT 72.61 3.21 72.63 3.418 ;
      RECT 72.57 3.213 72.61 3.429 ;
      RECT 72.555 3.215 72.57 3.442 ;
      RECT 72.545 3.215 72.555 3.447 ;
      RECT 72.52 3.216 72.545 3.455 ;
      RECT 72.51 3.218 72.52 3.46 ;
      RECT 72.505 3.219 72.51 3.463 ;
      RECT 72.48 3.217 72.505 3.466 ;
      RECT 72.465 3.215 72.48 3.467 ;
      RECT 72.445 3.212 72.465 3.469 ;
      RECT 72.425 3.207 72.445 3.469 ;
      RECT 72.365 3.202 72.425 3.466 ;
      RECT 72.33 3.177 72.365 3.462 ;
      RECT 72.32 3.154 72.33 3.46 ;
      RECT 72.29 3.131 72.32 3.46 ;
      RECT 72.28 3.11 72.29 3.46 ;
      RECT 72.255 3.092 72.28 3.458 ;
      RECT 72.24 3.07 72.255 3.455 ;
      RECT 72.225 3.052 72.24 3.453 ;
      RECT 72.205 3.042 72.225 3.451 ;
      RECT 72.19 3.037 72.205 3.45 ;
      RECT 72.175 3.035 72.19 3.449 ;
      RECT 72.145 3.036 72.175 3.447 ;
      RECT 72.125 3.039 72.145 3.445 ;
      RECT 72.068 3.043 72.125 3.445 ;
      RECT 71.982 3.052 72.068 3.445 ;
      RECT 71.896 3.063 71.982 3.445 ;
      RECT 71.81 3.074 71.896 3.445 ;
      RECT 71.79 3.081 71.81 3.453 ;
      RECT 71.78 3.084 71.79 3.46 ;
      RECT 71.715 3.089 71.78 3.478 ;
      RECT 71.685 3.096 71.715 3.503 ;
      RECT 71.675 3.099 71.685 3.51 ;
      RECT 71.63 3.103 71.675 3.515 ;
      RECT 71.6 3.108 71.63 3.52 ;
      RECT 71.599 3.11 71.6 3.52 ;
      RECT 71.513 3.116 71.599 3.52 ;
      RECT 71.427 3.127 71.513 3.52 ;
      RECT 71.341 3.139 71.427 3.52 ;
      RECT 71.255 3.15 71.341 3.52 ;
      RECT 71.24 3.157 71.255 3.515 ;
      RECT 71.235 3.159 71.24 3.509 ;
      RECT 71.215 3.17 71.235 3.504 ;
      RECT 71.205 3.188 71.215 3.498 ;
      RECT 71.2 3.2 71.205 3.298 ;
      RECT 73.495 1.953 73.515 2.04 ;
      RECT 73.49 1.888 73.495 2.072 ;
      RECT 73.48 1.855 73.49 2.077 ;
      RECT 73.475 1.835 73.48 2.083 ;
      RECT 73.445 1.835 73.475 2.1 ;
      RECT 73.396 1.835 73.445 2.136 ;
      RECT 73.31 1.835 73.396 2.194 ;
      RECT 73.281 1.845 73.31 2.243 ;
      RECT 73.195 1.887 73.281 2.296 ;
      RECT 73.175 1.925 73.195 2.343 ;
      RECT 73.15 1.942 73.175 2.363 ;
      RECT 73.14 1.956 73.15 2.383 ;
      RECT 73.135 1.962 73.14 2.393 ;
      RECT 73.13 1.966 73.135 2.4 ;
      RECT 73.08 1.986 73.13 2.405 ;
      RECT 73.015 2.03 73.08 2.405 ;
      RECT 72.99 2.08 73.015 2.405 ;
      RECT 72.98 2.11 72.99 2.405 ;
      RECT 72.975 2.137 72.98 2.405 ;
      RECT 72.97 2.155 72.975 2.405 ;
      RECT 72.96 2.197 72.97 2.405 ;
      RECT 73.31 2.755 73.48 2.93 ;
      RECT 73.25 2.583 73.31 2.918 ;
      RECT 73.24 2.576 73.25 2.901 ;
      RECT 73.195 2.755 73.48 2.881 ;
      RECT 73.176 2.755 73.48 2.859 ;
      RECT 73.09 2.755 73.48 2.824 ;
      RECT 73.07 2.575 73.24 2.78 ;
      RECT 73.07 2.722 73.475 2.78 ;
      RECT 73.07 2.67 73.45 2.78 ;
      RECT 73.07 2.625 73.415 2.78 ;
      RECT 73.07 2.607 73.38 2.78 ;
      RECT 73.07 2.597 73.375 2.78 ;
      RECT 73.24 7.855 73.41 8.305 ;
      RECT 73.295 6.075 73.465 8.025 ;
      RECT 73.24 5.015 73.41 6.245 ;
      RECT 72.72 5.015 72.89 8.305 ;
      RECT 72.72 7.315 73.125 7.645 ;
      RECT 72.72 6.475 73.125 6.805 ;
      RECT 72.79 3.555 72.98 3.78 ;
      RECT 72.78 3.556 72.985 3.775 ;
      RECT 72.78 3.558 72.995 3.755 ;
      RECT 72.78 3.562 73 3.74 ;
      RECT 72.78 3.549 72.95 3.775 ;
      RECT 72.78 3.552 72.975 3.775 ;
      RECT 72.79 3.548 72.95 3.78 ;
      RECT 72.876 3.546 72.95 3.78 ;
      RECT 72.5 2.797 72.67 3.035 ;
      RECT 72.5 2.797 72.756 2.949 ;
      RECT 72.5 2.797 72.76 2.859 ;
      RECT 72.55 2.57 72.77 2.838 ;
      RECT 72.545 2.587 72.775 2.811 ;
      RECT 72.51 2.745 72.775 2.811 ;
      RECT 72.53 2.595 72.67 3.035 ;
      RECT 72.52 2.677 72.78 2.794 ;
      RECT 72.515 2.725 72.78 2.794 ;
      RECT 72.52 2.635 72.775 2.811 ;
      RECT 72.545 2.572 72.77 2.838 ;
      RECT 72.11 2.547 72.28 2.745 ;
      RECT 72.11 2.547 72.325 2.72 ;
      RECT 72.18 2.49 72.35 2.678 ;
      RECT 72.155 2.505 72.35 2.678 ;
      RECT 71.77 2.551 71.8 2.745 ;
      RECT 71.765 2.523 71.77 2.745 ;
      RECT 71.735 2.497 71.765 2.747 ;
      RECT 71.71 2.455 71.735 2.75 ;
      RECT 71.7 2.427 71.71 2.752 ;
      RECT 71.665 2.407 71.7 2.754 ;
      RECT 71.6 2.392 71.665 2.76 ;
      RECT 71.55 2.39 71.6 2.766 ;
      RECT 71.527 2.392 71.55 2.771 ;
      RECT 71.441 2.403 71.527 2.777 ;
      RECT 71.355 2.421 71.441 2.787 ;
      RECT 71.34 2.432 71.355 2.793 ;
      RECT 71.27 2.455 71.34 2.799 ;
      RECT 71.215 2.487 71.27 2.807 ;
      RECT 71.175 2.51 71.215 2.813 ;
      RECT 71.161 2.523 71.175 2.816 ;
      RECT 71.075 2.545 71.161 2.822 ;
      RECT 71.06 2.57 71.075 2.828 ;
      RECT 71.02 2.585 71.06 2.832 ;
      RECT 70.97 2.6 71.02 2.837 ;
      RECT 70.945 2.607 70.97 2.841 ;
      RECT 70.885 2.602 70.945 2.845 ;
      RECT 70.87 2.593 70.885 2.849 ;
      RECT 70.8 2.583 70.87 2.845 ;
      RECT 70.775 2.575 70.795 2.835 ;
      RECT 70.716 2.575 70.775 2.813 ;
      RECT 70.63 2.575 70.716 2.77 ;
      RECT 70.795 2.575 70.8 2.84 ;
      RECT 71.49 1.806 71.66 2.14 ;
      RECT 71.46 1.806 71.66 2.135 ;
      RECT 71.4 1.773 71.46 2.123 ;
      RECT 71.4 1.829 71.67 2.118 ;
      RECT 71.375 1.829 71.67 2.112 ;
      RECT 71.37 1.77 71.4 2.109 ;
      RECT 71.355 1.776 71.49 2.107 ;
      RECT 71.35 1.784 71.575 2.095 ;
      RECT 71.35 1.836 71.685 2.048 ;
      RECT 71.335 1.792 71.575 2.043 ;
      RECT 71.335 1.862 71.695 1.984 ;
      RECT 71.305 1.812 71.66 1.945 ;
      RECT 71.305 1.902 71.705 1.941 ;
      RECT 71.355 1.781 71.575 2.107 ;
      RECT 70.695 2.111 70.75 2.375 ;
      RECT 70.695 2.111 70.815 2.374 ;
      RECT 70.695 2.111 70.84 2.373 ;
      RECT 70.695 2.111 70.905 2.372 ;
      RECT 70.84 2.077 70.92 2.371 ;
      RECT 70.655 2.121 71.065 2.37 ;
      RECT 70.695 2.118 71.065 2.37 ;
      RECT 70.655 2.126 71.07 2.363 ;
      RECT 70.64 2.128 71.07 2.362 ;
      RECT 70.64 2.135 71.075 2.358 ;
      RECT 70.62 2.134 71.07 2.354 ;
      RECT 70.62 2.142 71.08 2.353 ;
      RECT 70.615 2.139 71.075 2.349 ;
      RECT 70.615 2.152 71.09 2.348 ;
      RECT 70.6 2.142 71.08 2.347 ;
      RECT 70.565 2.155 71.09 2.34 ;
      RECT 70.75 2.11 71.06 2.37 ;
      RECT 70.75 2.095 71.01 2.37 ;
      RECT 70.815 2.082 70.945 2.37 ;
      RECT 70.36 3.171 70.375 3.564 ;
      RECT 70.325 3.176 70.375 3.563 ;
      RECT 70.36 3.175 70.42 3.562 ;
      RECT 70.305 3.186 70.42 3.561 ;
      RECT 70.32 3.182 70.42 3.561 ;
      RECT 70.285 3.192 70.495 3.558 ;
      RECT 70.285 3.211 70.54 3.556 ;
      RECT 70.285 3.218 70.545 3.553 ;
      RECT 70.27 3.195 70.495 3.55 ;
      RECT 70.25 3.2 70.495 3.543 ;
      RECT 70.245 3.204 70.495 3.539 ;
      RECT 70.245 3.221 70.555 3.538 ;
      RECT 70.225 3.215 70.54 3.534 ;
      RECT 70.225 3.224 70.56 3.528 ;
      RECT 70.22 3.23 70.56 3.3 ;
      RECT 70.285 3.19 70.42 3.558 ;
      RECT 70.16 2.553 70.36 2.865 ;
      RECT 70.235 2.531 70.36 2.865 ;
      RECT 70.175 2.55 70.365 2.85 ;
      RECT 70.145 2.561 70.365 2.848 ;
      RECT 70.16 2.556 70.37 2.814 ;
      RECT 70.145 2.66 70.375 2.781 ;
      RECT 70.175 2.532 70.36 2.865 ;
      RECT 70.235 2.51 70.335 2.865 ;
      RECT 70.26 2.507 70.335 2.865 ;
      RECT 70.26 2.502 70.28 2.865 ;
      RECT 69.665 2.57 69.84 2.745 ;
      RECT 69.66 2.57 69.84 2.743 ;
      RECT 69.635 2.57 69.84 2.738 ;
      RECT 69.58 2.55 69.75 2.728 ;
      RECT 69.58 2.557 69.815 2.728 ;
      RECT 69.665 3.237 69.68 3.42 ;
      RECT 69.655 3.215 69.665 3.42 ;
      RECT 69.64 3.195 69.655 3.42 ;
      RECT 69.63 3.17 69.64 3.42 ;
      RECT 69.6 3.135 69.63 3.42 ;
      RECT 69.565 3.075 69.6 3.42 ;
      RECT 69.56 3.037 69.565 3.42 ;
      RECT 69.51 2.988 69.56 3.42 ;
      RECT 69.5 2.938 69.51 3.408 ;
      RECT 69.485 2.917 69.5 3.368 ;
      RECT 69.465 2.885 69.485 3.318 ;
      RECT 69.44 2.841 69.465 3.258 ;
      RECT 69.435 2.813 69.44 3.213 ;
      RECT 69.43 2.804 69.435 3.199 ;
      RECT 69.425 2.797 69.43 3.186 ;
      RECT 69.42 2.792 69.425 3.175 ;
      RECT 69.415 2.777 69.42 3.165 ;
      RECT 69.41 2.755 69.415 3.152 ;
      RECT 69.4 2.715 69.41 3.127 ;
      RECT 69.375 2.645 69.4 3.083 ;
      RECT 69.37 2.585 69.375 3.048 ;
      RECT 69.355 2.565 69.37 3.015 ;
      RECT 69.35 2.565 69.355 2.99 ;
      RECT 69.32 2.565 69.35 2.945 ;
      RECT 69.275 2.565 69.32 2.885 ;
      RECT 69.2 2.565 69.275 2.833 ;
      RECT 69.195 2.565 69.2 2.798 ;
      RECT 69.19 2.565 69.195 2.788 ;
      RECT 69.185 2.565 69.19 2.768 ;
      RECT 69.45 1.785 69.62 2.255 ;
      RECT 69.395 1.778 69.59 2.239 ;
      RECT 69.395 1.792 69.625 2.238 ;
      RECT 69.38 1.793 69.625 2.219 ;
      RECT 69.375 1.811 69.625 2.205 ;
      RECT 69.38 1.794 69.63 2.203 ;
      RECT 69.365 1.825 69.63 2.188 ;
      RECT 69.38 1.8 69.635 2.173 ;
      RECT 69.36 1.84 69.635 2.17 ;
      RECT 69.375 1.812 69.64 2.155 ;
      RECT 69.375 1.824 69.645 2.135 ;
      RECT 69.36 1.84 69.65 2.118 ;
      RECT 69.36 1.85 69.655 1.973 ;
      RECT 69.355 1.85 69.655 1.93 ;
      RECT 69.355 1.865 69.66 1.908 ;
      RECT 69.45 1.775 69.59 2.255 ;
      RECT 69.45 1.773 69.56 2.255 ;
      RECT 69.536 1.77 69.56 2.255 ;
      RECT 69.195 3.437 69.2 3.483 ;
      RECT 69.185 3.285 69.195 3.507 ;
      RECT 69.18 3.13 69.185 3.532 ;
      RECT 69.165 3.092 69.18 3.543 ;
      RECT 69.16 3.075 69.165 3.55 ;
      RECT 69.15 3.063 69.16 3.557 ;
      RECT 69.145 3.054 69.15 3.559 ;
      RECT 69.14 3.052 69.145 3.563 ;
      RECT 69.095 3.043 69.14 3.578 ;
      RECT 69.09 3.035 69.095 3.592 ;
      RECT 69.085 3.032 69.09 3.596 ;
      RECT 69.07 3.027 69.085 3.604 ;
      RECT 69.015 3.017 69.07 3.615 ;
      RECT 68.98 3.005 69.015 3.616 ;
      RECT 68.971 3 68.98 3.61 ;
      RECT 68.885 3 68.971 3.6 ;
      RECT 68.855 3 68.885 3.578 ;
      RECT 68.845 3 68.85 3.558 ;
      RECT 68.84 3 68.845 3.52 ;
      RECT 68.835 3 68.84 3.478 ;
      RECT 68.83 3 68.835 3.438 ;
      RECT 68.825 3 68.83 3.368 ;
      RECT 68.815 3 68.825 3.29 ;
      RECT 68.81 3 68.815 3.19 ;
      RECT 68.85 3 68.855 3.56 ;
      RECT 68.345 3.082 68.435 3.56 ;
      RECT 68.33 3.085 68.45 3.558 ;
      RECT 68.345 3.084 68.45 3.558 ;
      RECT 68.31 3.091 68.475 3.548 ;
      RECT 68.33 3.085 68.475 3.548 ;
      RECT 68.295 3.097 68.475 3.536 ;
      RECT 68.33 3.088 68.525 3.529 ;
      RECT 68.281 3.105 68.525 3.527 ;
      RECT 68.31 3.095 68.535 3.515 ;
      RECT 68.281 3.116 68.565 3.506 ;
      RECT 68.195 3.14 68.565 3.5 ;
      RECT 68.195 3.153 68.605 3.483 ;
      RECT 68.19 3.175 68.605 3.476 ;
      RECT 68.16 3.19 68.605 3.466 ;
      RECT 68.155 3.201 68.605 3.456 ;
      RECT 68.125 3.214 68.605 3.447 ;
      RECT 68.11 3.232 68.605 3.436 ;
      RECT 68.085 3.245 68.605 3.426 ;
      RECT 68.345 3.081 68.355 3.56 ;
      RECT 68.391 2.505 68.43 2.75 ;
      RECT 68.305 2.505 68.44 2.748 ;
      RECT 68.19 2.53 68.44 2.745 ;
      RECT 68.19 2.53 68.445 2.743 ;
      RECT 68.19 2.53 68.46 2.738 ;
      RECT 68.296 2.505 68.475 2.718 ;
      RECT 68.21 2.513 68.475 2.718 ;
      RECT 67.88 1.865 68.05 2.3 ;
      RECT 67.87 1.899 68.05 2.283 ;
      RECT 67.95 1.835 68.12 2.27 ;
      RECT 67.855 1.91 68.12 2.248 ;
      RECT 67.95 1.845 68.125 2.238 ;
      RECT 67.88 1.897 68.155 2.223 ;
      RECT 67.84 1.923 68.155 2.208 ;
      RECT 67.84 1.965 68.165 2.188 ;
      RECT 67.835 1.99 68.17 2.17 ;
      RECT 67.835 2 68.175 2.155 ;
      RECT 67.83 1.937 68.155 2.153 ;
      RECT 67.83 2.01 68.18 2.138 ;
      RECT 67.825 1.947 68.155 2.135 ;
      RECT 67.82 2.031 68.185 2.118 ;
      RECT 67.82 2.063 68.19 2.098 ;
      RECT 67.815 1.977 68.165 2.09 ;
      RECT 67.82 1.962 68.155 2.118 ;
      RECT 67.835 1.932 68.155 2.17 ;
      RECT 67.68 2.519 67.905 2.775 ;
      RECT 67.68 2.552 67.925 2.765 ;
      RECT 67.645 2.552 67.925 2.763 ;
      RECT 67.645 2.565 67.93 2.753 ;
      RECT 67.645 2.585 67.94 2.745 ;
      RECT 67.645 2.682 67.945 2.738 ;
      RECT 67.625 2.43 67.755 2.728 ;
      RECT 67.58 2.585 67.94 2.67 ;
      RECT 67.57 2.43 67.755 2.615 ;
      RECT 67.57 2.462 67.841 2.615 ;
      RECT 67.535 2.992 67.555 3.17 ;
      RECT 67.5 2.945 67.535 3.17 ;
      RECT 67.485 2.885 67.5 3.17 ;
      RECT 67.46 2.832 67.485 3.17 ;
      RECT 67.445 2.785 67.46 3.17 ;
      RECT 67.425 2.762 67.445 3.17 ;
      RECT 67.4 2.727 67.425 3.17 ;
      RECT 67.39 2.573 67.4 3.17 ;
      RECT 67.36 2.568 67.39 3.161 ;
      RECT 67.355 2.565 67.36 3.151 ;
      RECT 67.34 2.565 67.355 3.125 ;
      RECT 67.335 2.565 67.34 3.088 ;
      RECT 67.31 2.565 67.335 3.04 ;
      RECT 67.29 2.565 67.31 2.965 ;
      RECT 67.28 2.565 67.29 2.925 ;
      RECT 67.275 2.565 67.28 2.9 ;
      RECT 67.27 2.565 67.275 2.883 ;
      RECT 67.265 2.565 67.27 2.865 ;
      RECT 67.26 2.566 67.265 2.855 ;
      RECT 67.25 2.568 67.26 2.823 ;
      RECT 67.24 2.57 67.25 2.79 ;
      RECT 67.23 2.573 67.24 2.763 ;
      RECT 67.555 3 67.78 3.17 ;
      RECT 66.885 1.812 67.055 2.265 ;
      RECT 66.885 1.812 67.145 2.231 ;
      RECT 66.885 1.812 67.175 2.215 ;
      RECT 66.885 1.812 67.205 2.188 ;
      RECT 67.141 1.79 67.22 2.17 ;
      RECT 66.92 1.797 67.225 2.155 ;
      RECT 66.92 1.805 67.235 2.118 ;
      RECT 66.88 1.832 67.235 2.09 ;
      RECT 66.865 1.845 67.235 2.055 ;
      RECT 66.885 1.82 67.255 2.045 ;
      RECT 66.86 1.885 67.255 2.015 ;
      RECT 66.86 1.915 67.26 1.998 ;
      RECT 66.855 1.945 67.26 1.985 ;
      RECT 66.92 1.794 67.22 2.17 ;
      RECT 67.055 1.791 67.141 2.249 ;
      RECT 67.006 1.792 67.22 2.17 ;
      RECT 67.15 3.452 67.195 3.645 ;
      RECT 67.14 3.422 67.15 3.645 ;
      RECT 67.135 3.407 67.14 3.645 ;
      RECT 67.095 3.317 67.135 3.645 ;
      RECT 67.09 3.23 67.095 3.645 ;
      RECT 67.08 3.2 67.09 3.645 ;
      RECT 67.075 3.16 67.08 3.645 ;
      RECT 67.065 3.122 67.075 3.645 ;
      RECT 67.06 3.087 67.065 3.645 ;
      RECT 67.04 3.04 67.06 3.645 ;
      RECT 67.025 2.965 67.04 3.645 ;
      RECT 67.02 2.92 67.025 3.64 ;
      RECT 67.015 2.9 67.02 3.613 ;
      RECT 67.01 2.88 67.015 3.598 ;
      RECT 67.005 2.855 67.01 3.578 ;
      RECT 67 2.833 67.005 3.563 ;
      RECT 66.995 2.811 67 3.545 ;
      RECT 66.99 2.79 66.995 3.535 ;
      RECT 66.98 2.762 66.99 3.505 ;
      RECT 66.97 2.725 66.98 3.473 ;
      RECT 66.96 2.685 66.97 3.44 ;
      RECT 66.95 2.663 66.96 3.41 ;
      RECT 66.92 2.615 66.95 3.342 ;
      RECT 66.905 2.575 66.92 3.269 ;
      RECT 66.895 2.575 66.905 3.235 ;
      RECT 66.89 2.575 66.895 3.21 ;
      RECT 66.885 2.575 66.89 3.195 ;
      RECT 66.88 2.575 66.885 3.173 ;
      RECT 66.875 2.575 66.88 3.16 ;
      RECT 66.86 2.575 66.875 3.125 ;
      RECT 66.84 2.575 66.86 3.065 ;
      RECT 66.83 2.575 66.84 3.015 ;
      RECT 66.81 2.575 66.83 2.963 ;
      RECT 66.79 2.575 66.81 2.92 ;
      RECT 66.78 2.575 66.79 2.908 ;
      RECT 66.75 2.575 66.78 2.895 ;
      RECT 66.72 2.596 66.75 2.875 ;
      RECT 66.71 2.624 66.72 2.855 ;
      RECT 66.695 2.641 66.71 2.823 ;
      RECT 66.69 2.655 66.695 2.79 ;
      RECT 66.685 2.663 66.69 2.763 ;
      RECT 66.68 2.671 66.685 2.725 ;
      RECT 66.685 3.195 66.69 3.53 ;
      RECT 66.65 3.182 66.685 3.529 ;
      RECT 66.58 3.122 66.65 3.528 ;
      RECT 66.5 3.065 66.58 3.527 ;
      RECT 66.365 3.025 66.5 3.526 ;
      RECT 66.365 3.212 66.7 3.515 ;
      RECT 66.325 3.212 66.7 3.505 ;
      RECT 66.325 3.23 66.705 3.5 ;
      RECT 66.325 3.32 66.71 3.49 ;
      RECT 66.32 3.015 66.485 3.47 ;
      RECT 66.315 3.015 66.485 3.213 ;
      RECT 66.315 3.172 66.68 3.213 ;
      RECT 66.315 3.16 66.675 3.213 ;
      RECT 65.08 1.74 65.25 2.935 ;
      RECT 65.08 1.74 65.545 1.91 ;
      RECT 65.08 6.97 65.545 7.14 ;
      RECT 65.08 5.945 65.25 7.14 ;
      RECT 64.09 1.74 64.26 2.935 ;
      RECT 64.09 1.74 64.555 1.91 ;
      RECT 64.09 6.97 64.555 7.14 ;
      RECT 64.09 5.945 64.26 7.14 ;
      RECT 62.235 2.635 62.405 3.865 ;
      RECT 62.29 0.855 62.46 2.805 ;
      RECT 62.235 0.575 62.405 1.025 ;
      RECT 62.235 7.855 62.405 8.305 ;
      RECT 62.29 6.075 62.46 8.025 ;
      RECT 62.235 5.015 62.405 6.245 ;
      RECT 61.715 0.575 61.885 3.865 ;
      RECT 61.715 2.075 62.12 2.405 ;
      RECT 61.715 1.235 62.12 1.565 ;
      RECT 61.715 5.015 61.885 8.305 ;
      RECT 61.715 7.315 62.12 7.645 ;
      RECT 61.715 6.475 62.12 6.805 ;
      RECT 59.05 1.975 59.78 2.215 ;
      RECT 59.592 1.77 59.78 2.215 ;
      RECT 59.42 1.782 59.795 2.209 ;
      RECT 59.335 1.797 59.815 2.194 ;
      RECT 59.335 1.812 59.82 2.184 ;
      RECT 59.29 1.832 59.835 2.176 ;
      RECT 59.267 1.867 59.85 2.13 ;
      RECT 59.181 1.89 59.855 2.09 ;
      RECT 59.181 1.908 59.865 2.06 ;
      RECT 59.05 1.977 59.87 2.023 ;
      RECT 59.095 1.92 59.865 2.06 ;
      RECT 59.181 1.872 59.85 2.13 ;
      RECT 59.267 1.841 59.835 2.176 ;
      RECT 59.29 1.822 59.82 2.184 ;
      RECT 59.335 1.795 59.795 2.209 ;
      RECT 59.42 1.777 59.78 2.215 ;
      RECT 59.506 1.771 59.78 2.215 ;
      RECT 59.592 1.766 59.725 2.215 ;
      RECT 59.678 1.761 59.725 2.215 ;
      RECT 59.37 2.659 59.54 3.045 ;
      RECT 59.365 2.659 59.54 3.04 ;
      RECT 59.34 2.659 59.54 3.005 ;
      RECT 59.34 2.687 59.55 2.995 ;
      RECT 59.32 2.687 59.55 2.955 ;
      RECT 59.315 2.687 59.55 2.928 ;
      RECT 59.315 2.705 59.555 2.92 ;
      RECT 59.26 2.705 59.555 2.855 ;
      RECT 59.26 2.722 59.565 2.838 ;
      RECT 59.25 2.722 59.565 2.778 ;
      RECT 59.25 2.739 59.57 2.775 ;
      RECT 59.245 2.575 59.415 2.753 ;
      RECT 59.245 2.609 59.501 2.753 ;
      RECT 59.24 3.375 59.245 3.388 ;
      RECT 59.235 3.27 59.24 3.393 ;
      RECT 59.21 3.13 59.235 3.408 ;
      RECT 59.175 3.081 59.21 3.44 ;
      RECT 59.17 3.049 59.175 3.46 ;
      RECT 59.165 3.04 59.17 3.46 ;
      RECT 59.085 3.005 59.165 3.46 ;
      RECT 59.022 2.975 59.085 3.46 ;
      RECT 58.936 2.963 59.022 3.46 ;
      RECT 58.85 2.949 58.936 3.46 ;
      RECT 58.77 2.936 58.85 3.446 ;
      RECT 58.735 2.928 58.77 3.426 ;
      RECT 58.725 2.925 58.735 3.417 ;
      RECT 58.695 2.92 58.725 3.404 ;
      RECT 58.645 2.895 58.695 3.38 ;
      RECT 58.631 2.869 58.645 3.362 ;
      RECT 58.545 2.829 58.631 3.338 ;
      RECT 58.5 2.777 58.545 3.307 ;
      RECT 58.49 2.752 58.5 3.294 ;
      RECT 58.485 2.533 58.49 2.555 ;
      RECT 58.48 2.735 58.49 3.29 ;
      RECT 58.48 2.531 58.485 2.645 ;
      RECT 58.47 2.527 58.48 3.286 ;
      RECT 58.426 2.525 58.47 3.274 ;
      RECT 58.34 2.525 58.426 3.245 ;
      RECT 58.31 2.525 58.34 3.218 ;
      RECT 58.295 2.525 58.31 3.206 ;
      RECT 58.255 2.537 58.295 3.191 ;
      RECT 58.235 2.556 58.255 3.17 ;
      RECT 58.225 2.566 58.235 3.154 ;
      RECT 58.215 2.572 58.225 3.143 ;
      RECT 58.195 2.582 58.215 3.126 ;
      RECT 58.19 2.591 58.195 3.113 ;
      RECT 58.185 2.595 58.19 3.063 ;
      RECT 58.175 2.601 58.185 2.98 ;
      RECT 58.17 2.605 58.175 2.894 ;
      RECT 58.165 2.625 58.17 2.831 ;
      RECT 58.16 2.648 58.165 2.778 ;
      RECT 58.155 2.666 58.16 2.723 ;
      RECT 58.765 2.485 58.935 2.745 ;
      RECT 58.935 2.45 58.98 2.731 ;
      RECT 58.896 2.452 58.985 2.714 ;
      RECT 58.785 2.469 59.071 2.685 ;
      RECT 58.785 2.484 59.075 2.657 ;
      RECT 58.785 2.465 58.985 2.714 ;
      RECT 58.81 2.453 58.935 2.745 ;
      RECT 58.896 2.451 58.98 2.731 ;
      RECT 57.95 1.84 58.12 2.33 ;
      RECT 57.95 1.84 58.155 2.31 ;
      RECT 58.085 1.76 58.195 2.27 ;
      RECT 58.066 1.764 58.215 2.24 ;
      RECT 57.98 1.772 58.235 2.223 ;
      RECT 57.98 1.778 58.24 2.213 ;
      RECT 57.98 1.787 58.26 2.201 ;
      RECT 57.955 1.812 58.29 2.179 ;
      RECT 57.955 1.832 58.295 2.159 ;
      RECT 57.95 1.845 58.305 2.139 ;
      RECT 57.95 1.912 58.31 2.12 ;
      RECT 57.95 2.045 58.315 2.107 ;
      RECT 57.945 1.85 58.305 1.94 ;
      RECT 57.955 1.807 58.26 2.201 ;
      RECT 58.066 1.762 58.195 2.27 ;
      RECT 57.94 3.515 58.24 3.77 ;
      RECT 58.025 3.481 58.24 3.77 ;
      RECT 58.025 3.484 58.245 3.63 ;
      RECT 57.96 3.505 58.245 3.63 ;
      RECT 57.995 3.495 58.24 3.77 ;
      RECT 57.99 3.5 58.245 3.63 ;
      RECT 58.025 3.479 58.226 3.77 ;
      RECT 58.111 3.47 58.226 3.77 ;
      RECT 58.111 3.464 58.14 3.77 ;
      RECT 57.6 3.105 57.61 3.595 ;
      RECT 57.26 3.04 57.27 3.34 ;
      RECT 57.775 3.212 57.78 3.431 ;
      RECT 57.765 3.192 57.775 3.448 ;
      RECT 57.755 3.172 57.765 3.478 ;
      RECT 57.75 3.162 57.755 3.493 ;
      RECT 57.745 3.158 57.75 3.498 ;
      RECT 57.73 3.15 57.745 3.505 ;
      RECT 57.69 3.13 57.73 3.53 ;
      RECT 57.665 3.112 57.69 3.563 ;
      RECT 57.66 3.11 57.665 3.576 ;
      RECT 57.64 3.107 57.66 3.58 ;
      RECT 57.61 3.105 57.64 3.59 ;
      RECT 57.54 3.107 57.6 3.591 ;
      RECT 57.52 3.107 57.54 3.585 ;
      RECT 57.495 3.105 57.52 3.582 ;
      RECT 57.46 3.1 57.495 3.578 ;
      RECT 57.44 3.094 57.46 3.565 ;
      RECT 57.43 3.091 57.44 3.553 ;
      RECT 57.41 3.088 57.43 3.538 ;
      RECT 57.39 3.084 57.41 3.52 ;
      RECT 57.385 3.081 57.39 3.51 ;
      RECT 57.38 3.08 57.385 3.508 ;
      RECT 57.37 3.077 57.38 3.5 ;
      RECT 57.36 3.071 57.37 3.483 ;
      RECT 57.35 3.065 57.36 3.465 ;
      RECT 57.34 3.059 57.35 3.453 ;
      RECT 57.33 3.053 57.34 3.433 ;
      RECT 57.325 3.049 57.33 3.418 ;
      RECT 57.32 3.047 57.325 3.41 ;
      RECT 57.315 3.045 57.32 3.403 ;
      RECT 57.31 3.043 57.315 3.393 ;
      RECT 57.305 3.041 57.31 3.387 ;
      RECT 57.295 3.04 57.305 3.377 ;
      RECT 57.285 3.04 57.295 3.368 ;
      RECT 57.27 3.04 57.285 3.353 ;
      RECT 57.23 3.04 57.26 3.337 ;
      RECT 57.21 3.042 57.23 3.332 ;
      RECT 57.205 3.047 57.21 3.33 ;
      RECT 57.175 3.055 57.205 3.328 ;
      RECT 57.145 3.07 57.175 3.327 ;
      RECT 57.1 3.092 57.145 3.332 ;
      RECT 57.095 3.107 57.1 3.336 ;
      RECT 57.08 3.112 57.095 3.338 ;
      RECT 57.075 3.116 57.08 3.34 ;
      RECT 57.015 3.139 57.075 3.349 ;
      RECT 56.995 3.165 57.015 3.362 ;
      RECT 56.985 3.172 56.995 3.366 ;
      RECT 56.97 3.179 56.985 3.369 ;
      RECT 56.95 3.189 56.97 3.372 ;
      RECT 56.945 3.197 56.95 3.375 ;
      RECT 56.9 3.202 56.945 3.382 ;
      RECT 56.89 3.205 56.9 3.389 ;
      RECT 56.88 3.205 56.89 3.393 ;
      RECT 56.845 3.207 56.88 3.405 ;
      RECT 56.825 3.21 56.845 3.418 ;
      RECT 56.785 3.213 56.825 3.429 ;
      RECT 56.77 3.215 56.785 3.442 ;
      RECT 56.76 3.215 56.77 3.447 ;
      RECT 56.735 3.216 56.76 3.455 ;
      RECT 56.725 3.218 56.735 3.46 ;
      RECT 56.72 3.219 56.725 3.463 ;
      RECT 56.695 3.217 56.72 3.466 ;
      RECT 56.68 3.215 56.695 3.467 ;
      RECT 56.66 3.212 56.68 3.469 ;
      RECT 56.64 3.207 56.66 3.469 ;
      RECT 56.58 3.202 56.64 3.466 ;
      RECT 56.545 3.177 56.58 3.462 ;
      RECT 56.535 3.154 56.545 3.46 ;
      RECT 56.505 3.131 56.535 3.46 ;
      RECT 56.495 3.11 56.505 3.46 ;
      RECT 56.47 3.092 56.495 3.458 ;
      RECT 56.455 3.07 56.47 3.455 ;
      RECT 56.44 3.052 56.455 3.453 ;
      RECT 56.42 3.042 56.44 3.451 ;
      RECT 56.405 3.037 56.42 3.45 ;
      RECT 56.39 3.035 56.405 3.449 ;
      RECT 56.36 3.036 56.39 3.447 ;
      RECT 56.34 3.039 56.36 3.445 ;
      RECT 56.283 3.043 56.34 3.445 ;
      RECT 56.197 3.052 56.283 3.445 ;
      RECT 56.111 3.063 56.197 3.445 ;
      RECT 56.025 3.074 56.111 3.445 ;
      RECT 56.005 3.081 56.025 3.453 ;
      RECT 55.995 3.084 56.005 3.46 ;
      RECT 55.93 3.089 55.995 3.478 ;
      RECT 55.9 3.096 55.93 3.503 ;
      RECT 55.89 3.099 55.9 3.51 ;
      RECT 55.845 3.103 55.89 3.515 ;
      RECT 55.815 3.108 55.845 3.52 ;
      RECT 55.814 3.11 55.815 3.52 ;
      RECT 55.728 3.116 55.814 3.52 ;
      RECT 55.642 3.127 55.728 3.52 ;
      RECT 55.556 3.139 55.642 3.52 ;
      RECT 55.47 3.15 55.556 3.52 ;
      RECT 55.455 3.157 55.47 3.515 ;
      RECT 55.45 3.159 55.455 3.509 ;
      RECT 55.43 3.17 55.45 3.504 ;
      RECT 55.42 3.188 55.43 3.498 ;
      RECT 55.415 3.2 55.42 3.298 ;
      RECT 57.71 1.953 57.73 2.04 ;
      RECT 57.705 1.888 57.71 2.072 ;
      RECT 57.695 1.855 57.705 2.077 ;
      RECT 57.69 1.835 57.695 2.083 ;
      RECT 57.66 1.835 57.69 2.1 ;
      RECT 57.611 1.835 57.66 2.136 ;
      RECT 57.525 1.835 57.611 2.194 ;
      RECT 57.496 1.845 57.525 2.243 ;
      RECT 57.41 1.887 57.496 2.296 ;
      RECT 57.39 1.925 57.41 2.343 ;
      RECT 57.365 1.942 57.39 2.363 ;
      RECT 57.355 1.956 57.365 2.383 ;
      RECT 57.35 1.962 57.355 2.393 ;
      RECT 57.345 1.966 57.35 2.4 ;
      RECT 57.295 1.986 57.345 2.405 ;
      RECT 57.23 2.03 57.295 2.405 ;
      RECT 57.205 2.08 57.23 2.405 ;
      RECT 57.195 2.11 57.205 2.405 ;
      RECT 57.19 2.137 57.195 2.405 ;
      RECT 57.185 2.155 57.19 2.405 ;
      RECT 57.175 2.197 57.185 2.405 ;
      RECT 57.525 2.755 57.695 2.93 ;
      RECT 57.465 2.583 57.525 2.918 ;
      RECT 57.455 2.576 57.465 2.901 ;
      RECT 57.41 2.755 57.695 2.881 ;
      RECT 57.391 2.755 57.695 2.859 ;
      RECT 57.305 2.755 57.695 2.824 ;
      RECT 57.285 2.575 57.455 2.78 ;
      RECT 57.285 2.722 57.69 2.78 ;
      RECT 57.285 2.67 57.665 2.78 ;
      RECT 57.285 2.625 57.63 2.78 ;
      RECT 57.285 2.607 57.595 2.78 ;
      RECT 57.285 2.597 57.59 2.78 ;
      RECT 57.455 7.855 57.625 8.305 ;
      RECT 57.51 6.075 57.68 8.025 ;
      RECT 57.455 5.015 57.625 6.245 ;
      RECT 56.935 5.015 57.105 8.305 ;
      RECT 56.935 7.315 57.34 7.645 ;
      RECT 56.935 6.475 57.34 6.805 ;
      RECT 57.005 3.555 57.195 3.78 ;
      RECT 56.995 3.556 57.2 3.775 ;
      RECT 56.995 3.558 57.21 3.755 ;
      RECT 56.995 3.562 57.215 3.74 ;
      RECT 56.995 3.549 57.165 3.775 ;
      RECT 56.995 3.552 57.19 3.775 ;
      RECT 57.005 3.548 57.165 3.78 ;
      RECT 57.091 3.546 57.165 3.78 ;
      RECT 56.715 2.797 56.885 3.035 ;
      RECT 56.715 2.797 56.971 2.949 ;
      RECT 56.715 2.797 56.975 2.859 ;
      RECT 56.765 2.57 56.985 2.838 ;
      RECT 56.76 2.587 56.99 2.811 ;
      RECT 56.725 2.745 56.99 2.811 ;
      RECT 56.745 2.595 56.885 3.035 ;
      RECT 56.735 2.677 56.995 2.794 ;
      RECT 56.73 2.725 56.995 2.794 ;
      RECT 56.735 2.635 56.99 2.811 ;
      RECT 56.76 2.572 56.985 2.838 ;
      RECT 56.325 2.547 56.495 2.745 ;
      RECT 56.325 2.547 56.54 2.72 ;
      RECT 56.395 2.49 56.565 2.678 ;
      RECT 56.37 2.505 56.565 2.678 ;
      RECT 55.985 2.551 56.015 2.745 ;
      RECT 55.98 2.523 55.985 2.745 ;
      RECT 55.95 2.497 55.98 2.747 ;
      RECT 55.925 2.455 55.95 2.75 ;
      RECT 55.915 2.427 55.925 2.752 ;
      RECT 55.88 2.407 55.915 2.754 ;
      RECT 55.815 2.392 55.88 2.76 ;
      RECT 55.765 2.39 55.815 2.766 ;
      RECT 55.742 2.392 55.765 2.771 ;
      RECT 55.656 2.403 55.742 2.777 ;
      RECT 55.57 2.421 55.656 2.787 ;
      RECT 55.555 2.432 55.57 2.793 ;
      RECT 55.485 2.455 55.555 2.799 ;
      RECT 55.43 2.487 55.485 2.807 ;
      RECT 55.39 2.51 55.43 2.813 ;
      RECT 55.376 2.523 55.39 2.816 ;
      RECT 55.29 2.545 55.376 2.822 ;
      RECT 55.275 2.57 55.29 2.828 ;
      RECT 55.235 2.585 55.275 2.832 ;
      RECT 55.185 2.6 55.235 2.837 ;
      RECT 55.16 2.607 55.185 2.841 ;
      RECT 55.1 2.602 55.16 2.845 ;
      RECT 55.085 2.593 55.1 2.849 ;
      RECT 55.015 2.583 55.085 2.845 ;
      RECT 54.99 2.575 55.01 2.835 ;
      RECT 54.931 2.575 54.99 2.813 ;
      RECT 54.845 2.575 54.931 2.77 ;
      RECT 55.01 2.575 55.015 2.84 ;
      RECT 55.705 1.806 55.875 2.14 ;
      RECT 55.675 1.806 55.875 2.135 ;
      RECT 55.615 1.773 55.675 2.123 ;
      RECT 55.615 1.829 55.885 2.118 ;
      RECT 55.59 1.829 55.885 2.112 ;
      RECT 55.585 1.77 55.615 2.109 ;
      RECT 55.57 1.776 55.705 2.107 ;
      RECT 55.565 1.784 55.79 2.095 ;
      RECT 55.565 1.836 55.9 2.048 ;
      RECT 55.55 1.792 55.79 2.043 ;
      RECT 55.55 1.862 55.91 1.984 ;
      RECT 55.52 1.812 55.875 1.945 ;
      RECT 55.52 1.902 55.92 1.941 ;
      RECT 55.57 1.781 55.79 2.107 ;
      RECT 54.91 2.111 54.965 2.375 ;
      RECT 54.91 2.111 55.03 2.374 ;
      RECT 54.91 2.111 55.055 2.373 ;
      RECT 54.91 2.111 55.12 2.372 ;
      RECT 55.055 2.077 55.135 2.371 ;
      RECT 54.87 2.121 55.28 2.37 ;
      RECT 54.91 2.118 55.28 2.37 ;
      RECT 54.87 2.126 55.285 2.363 ;
      RECT 54.855 2.128 55.285 2.362 ;
      RECT 54.855 2.135 55.29 2.358 ;
      RECT 54.835 2.134 55.285 2.354 ;
      RECT 54.835 2.142 55.295 2.353 ;
      RECT 54.83 2.139 55.29 2.349 ;
      RECT 54.83 2.152 55.305 2.348 ;
      RECT 54.815 2.142 55.295 2.347 ;
      RECT 54.78 2.155 55.305 2.34 ;
      RECT 54.965 2.11 55.275 2.37 ;
      RECT 54.965 2.095 55.225 2.37 ;
      RECT 55.03 2.082 55.16 2.37 ;
      RECT 54.575 3.171 54.59 3.564 ;
      RECT 54.54 3.176 54.59 3.563 ;
      RECT 54.575 3.175 54.635 3.562 ;
      RECT 54.52 3.186 54.635 3.561 ;
      RECT 54.535 3.182 54.635 3.561 ;
      RECT 54.5 3.192 54.71 3.558 ;
      RECT 54.5 3.211 54.755 3.556 ;
      RECT 54.5 3.218 54.76 3.553 ;
      RECT 54.485 3.195 54.71 3.55 ;
      RECT 54.465 3.2 54.71 3.543 ;
      RECT 54.46 3.204 54.71 3.539 ;
      RECT 54.46 3.221 54.77 3.538 ;
      RECT 54.44 3.215 54.755 3.534 ;
      RECT 54.44 3.224 54.775 3.528 ;
      RECT 54.435 3.23 54.775 3.3 ;
      RECT 54.5 3.19 54.635 3.558 ;
      RECT 54.375 2.553 54.575 2.865 ;
      RECT 54.45 2.531 54.575 2.865 ;
      RECT 54.39 2.55 54.58 2.85 ;
      RECT 54.36 2.561 54.58 2.848 ;
      RECT 54.375 2.556 54.585 2.814 ;
      RECT 54.36 2.66 54.59 2.781 ;
      RECT 54.39 2.532 54.575 2.865 ;
      RECT 54.45 2.51 54.55 2.865 ;
      RECT 54.475 2.507 54.55 2.865 ;
      RECT 54.475 2.502 54.495 2.865 ;
      RECT 53.88 2.57 54.055 2.745 ;
      RECT 53.875 2.57 54.055 2.743 ;
      RECT 53.85 2.57 54.055 2.738 ;
      RECT 53.795 2.55 53.965 2.728 ;
      RECT 53.795 2.557 54.03 2.728 ;
      RECT 53.88 3.237 53.895 3.42 ;
      RECT 53.87 3.215 53.88 3.42 ;
      RECT 53.855 3.195 53.87 3.42 ;
      RECT 53.845 3.17 53.855 3.42 ;
      RECT 53.815 3.135 53.845 3.42 ;
      RECT 53.78 3.075 53.815 3.42 ;
      RECT 53.775 3.037 53.78 3.42 ;
      RECT 53.725 2.988 53.775 3.42 ;
      RECT 53.715 2.938 53.725 3.408 ;
      RECT 53.7 2.917 53.715 3.368 ;
      RECT 53.68 2.885 53.7 3.318 ;
      RECT 53.655 2.841 53.68 3.258 ;
      RECT 53.65 2.813 53.655 3.213 ;
      RECT 53.645 2.804 53.65 3.199 ;
      RECT 53.64 2.797 53.645 3.186 ;
      RECT 53.635 2.792 53.64 3.175 ;
      RECT 53.63 2.777 53.635 3.165 ;
      RECT 53.625 2.755 53.63 3.152 ;
      RECT 53.615 2.715 53.625 3.127 ;
      RECT 53.59 2.645 53.615 3.083 ;
      RECT 53.585 2.585 53.59 3.048 ;
      RECT 53.57 2.565 53.585 3.015 ;
      RECT 53.565 2.565 53.57 2.99 ;
      RECT 53.535 2.565 53.565 2.945 ;
      RECT 53.49 2.565 53.535 2.885 ;
      RECT 53.415 2.565 53.49 2.833 ;
      RECT 53.41 2.565 53.415 2.798 ;
      RECT 53.405 2.565 53.41 2.788 ;
      RECT 53.4 2.565 53.405 2.768 ;
      RECT 53.665 1.785 53.835 2.255 ;
      RECT 53.61 1.778 53.805 2.239 ;
      RECT 53.61 1.792 53.84 2.238 ;
      RECT 53.595 1.793 53.84 2.219 ;
      RECT 53.59 1.811 53.84 2.205 ;
      RECT 53.595 1.794 53.845 2.203 ;
      RECT 53.58 1.825 53.845 2.188 ;
      RECT 53.595 1.8 53.85 2.173 ;
      RECT 53.575 1.84 53.85 2.17 ;
      RECT 53.59 1.812 53.855 2.155 ;
      RECT 53.59 1.824 53.86 2.135 ;
      RECT 53.575 1.84 53.865 2.118 ;
      RECT 53.575 1.85 53.87 1.973 ;
      RECT 53.57 1.85 53.87 1.93 ;
      RECT 53.57 1.865 53.875 1.908 ;
      RECT 53.665 1.775 53.805 2.255 ;
      RECT 53.665 1.773 53.775 2.255 ;
      RECT 53.751 1.77 53.775 2.255 ;
      RECT 53.41 3.437 53.415 3.483 ;
      RECT 53.4 3.285 53.41 3.507 ;
      RECT 53.395 3.13 53.4 3.532 ;
      RECT 53.38 3.092 53.395 3.543 ;
      RECT 53.375 3.075 53.38 3.55 ;
      RECT 53.365 3.063 53.375 3.557 ;
      RECT 53.36 3.054 53.365 3.559 ;
      RECT 53.355 3.052 53.36 3.563 ;
      RECT 53.31 3.043 53.355 3.578 ;
      RECT 53.305 3.035 53.31 3.592 ;
      RECT 53.3 3.032 53.305 3.596 ;
      RECT 53.285 3.027 53.3 3.604 ;
      RECT 53.23 3.017 53.285 3.615 ;
      RECT 53.195 3.005 53.23 3.616 ;
      RECT 53.186 3 53.195 3.61 ;
      RECT 53.1 3 53.186 3.6 ;
      RECT 53.07 3 53.1 3.578 ;
      RECT 53.06 3 53.065 3.558 ;
      RECT 53.055 3 53.06 3.52 ;
      RECT 53.05 3 53.055 3.478 ;
      RECT 53.045 3 53.05 3.438 ;
      RECT 53.04 3 53.045 3.368 ;
      RECT 53.03 3 53.04 3.29 ;
      RECT 53.025 3 53.03 3.19 ;
      RECT 53.065 3 53.07 3.56 ;
      RECT 52.56 3.082 52.65 3.56 ;
      RECT 52.545 3.085 52.665 3.558 ;
      RECT 52.56 3.084 52.665 3.558 ;
      RECT 52.525 3.091 52.69 3.548 ;
      RECT 52.545 3.085 52.69 3.548 ;
      RECT 52.51 3.097 52.69 3.536 ;
      RECT 52.545 3.088 52.74 3.529 ;
      RECT 52.496 3.105 52.74 3.527 ;
      RECT 52.525 3.095 52.75 3.515 ;
      RECT 52.496 3.116 52.78 3.506 ;
      RECT 52.41 3.14 52.78 3.5 ;
      RECT 52.41 3.153 52.82 3.483 ;
      RECT 52.405 3.175 52.82 3.476 ;
      RECT 52.375 3.19 52.82 3.466 ;
      RECT 52.37 3.201 52.82 3.456 ;
      RECT 52.34 3.214 52.82 3.447 ;
      RECT 52.325 3.232 52.82 3.436 ;
      RECT 52.3 3.245 52.82 3.426 ;
      RECT 52.56 3.081 52.57 3.56 ;
      RECT 52.606 2.505 52.645 2.75 ;
      RECT 52.52 2.505 52.655 2.748 ;
      RECT 52.405 2.53 52.655 2.745 ;
      RECT 52.405 2.53 52.66 2.743 ;
      RECT 52.405 2.53 52.675 2.738 ;
      RECT 52.511 2.505 52.69 2.718 ;
      RECT 52.425 2.513 52.69 2.718 ;
      RECT 52.095 1.865 52.265 2.3 ;
      RECT 52.085 1.899 52.265 2.283 ;
      RECT 52.165 1.835 52.335 2.27 ;
      RECT 52.07 1.91 52.335 2.248 ;
      RECT 52.165 1.845 52.34 2.238 ;
      RECT 52.095 1.897 52.37 2.223 ;
      RECT 52.055 1.923 52.37 2.208 ;
      RECT 52.055 1.965 52.38 2.188 ;
      RECT 52.05 1.99 52.385 2.17 ;
      RECT 52.05 2 52.39 2.155 ;
      RECT 52.045 1.937 52.37 2.153 ;
      RECT 52.045 2.01 52.395 2.138 ;
      RECT 52.04 1.947 52.37 2.135 ;
      RECT 52.035 2.031 52.4 2.118 ;
      RECT 52.035 2.063 52.405 2.098 ;
      RECT 52.03 1.977 52.38 2.09 ;
      RECT 52.035 1.962 52.37 2.118 ;
      RECT 52.05 1.932 52.37 2.17 ;
      RECT 51.895 2.519 52.12 2.775 ;
      RECT 51.895 2.552 52.14 2.765 ;
      RECT 51.86 2.552 52.14 2.763 ;
      RECT 51.86 2.565 52.145 2.753 ;
      RECT 51.86 2.585 52.155 2.745 ;
      RECT 51.86 2.682 52.16 2.738 ;
      RECT 51.84 2.43 51.97 2.728 ;
      RECT 51.795 2.585 52.155 2.67 ;
      RECT 51.785 2.43 51.97 2.615 ;
      RECT 51.785 2.462 52.056 2.615 ;
      RECT 51.75 2.992 51.77 3.17 ;
      RECT 51.715 2.945 51.75 3.17 ;
      RECT 51.7 2.885 51.715 3.17 ;
      RECT 51.675 2.832 51.7 3.17 ;
      RECT 51.66 2.785 51.675 3.17 ;
      RECT 51.64 2.762 51.66 3.17 ;
      RECT 51.615 2.727 51.64 3.17 ;
      RECT 51.605 2.573 51.615 3.17 ;
      RECT 51.575 2.568 51.605 3.161 ;
      RECT 51.57 2.565 51.575 3.151 ;
      RECT 51.555 2.565 51.57 3.125 ;
      RECT 51.55 2.565 51.555 3.088 ;
      RECT 51.525 2.565 51.55 3.04 ;
      RECT 51.505 2.565 51.525 2.965 ;
      RECT 51.495 2.565 51.505 2.925 ;
      RECT 51.49 2.565 51.495 2.9 ;
      RECT 51.485 2.565 51.49 2.883 ;
      RECT 51.48 2.565 51.485 2.865 ;
      RECT 51.475 2.566 51.48 2.855 ;
      RECT 51.465 2.568 51.475 2.823 ;
      RECT 51.455 2.57 51.465 2.79 ;
      RECT 51.445 2.573 51.455 2.763 ;
      RECT 51.77 3 51.995 3.17 ;
      RECT 51.1 1.812 51.27 2.265 ;
      RECT 51.1 1.812 51.36 2.231 ;
      RECT 51.1 1.812 51.39 2.215 ;
      RECT 51.1 1.812 51.42 2.188 ;
      RECT 51.356 1.79 51.435 2.17 ;
      RECT 51.135 1.797 51.44 2.155 ;
      RECT 51.135 1.805 51.45 2.118 ;
      RECT 51.095 1.832 51.45 2.09 ;
      RECT 51.08 1.845 51.45 2.055 ;
      RECT 51.1 1.82 51.47 2.045 ;
      RECT 51.075 1.885 51.47 2.015 ;
      RECT 51.075 1.915 51.475 1.998 ;
      RECT 51.07 1.945 51.475 1.985 ;
      RECT 51.135 1.794 51.435 2.17 ;
      RECT 51.27 1.791 51.356 2.249 ;
      RECT 51.221 1.792 51.435 2.17 ;
      RECT 51.365 3.452 51.41 3.645 ;
      RECT 51.355 3.422 51.365 3.645 ;
      RECT 51.35 3.407 51.355 3.645 ;
      RECT 51.31 3.317 51.35 3.645 ;
      RECT 51.305 3.23 51.31 3.645 ;
      RECT 51.295 3.2 51.305 3.645 ;
      RECT 51.29 3.16 51.295 3.645 ;
      RECT 51.28 3.122 51.29 3.645 ;
      RECT 51.275 3.087 51.28 3.645 ;
      RECT 51.255 3.04 51.275 3.645 ;
      RECT 51.24 2.965 51.255 3.645 ;
      RECT 51.235 2.92 51.24 3.64 ;
      RECT 51.23 2.9 51.235 3.613 ;
      RECT 51.225 2.88 51.23 3.598 ;
      RECT 51.22 2.855 51.225 3.578 ;
      RECT 51.215 2.833 51.22 3.563 ;
      RECT 51.21 2.811 51.215 3.545 ;
      RECT 51.205 2.79 51.21 3.535 ;
      RECT 51.195 2.762 51.205 3.505 ;
      RECT 51.185 2.725 51.195 3.473 ;
      RECT 51.175 2.685 51.185 3.44 ;
      RECT 51.165 2.663 51.175 3.41 ;
      RECT 51.135 2.615 51.165 3.342 ;
      RECT 51.12 2.575 51.135 3.269 ;
      RECT 51.11 2.575 51.12 3.235 ;
      RECT 51.105 2.575 51.11 3.21 ;
      RECT 51.1 2.575 51.105 3.195 ;
      RECT 51.095 2.575 51.1 3.173 ;
      RECT 51.09 2.575 51.095 3.16 ;
      RECT 51.075 2.575 51.09 3.125 ;
      RECT 51.055 2.575 51.075 3.065 ;
      RECT 51.045 2.575 51.055 3.015 ;
      RECT 51.025 2.575 51.045 2.963 ;
      RECT 51.005 2.575 51.025 2.92 ;
      RECT 50.995 2.575 51.005 2.908 ;
      RECT 50.965 2.575 50.995 2.895 ;
      RECT 50.935 2.596 50.965 2.875 ;
      RECT 50.925 2.624 50.935 2.855 ;
      RECT 50.91 2.641 50.925 2.823 ;
      RECT 50.905 2.655 50.91 2.79 ;
      RECT 50.9 2.663 50.905 2.763 ;
      RECT 50.895 2.671 50.9 2.725 ;
      RECT 50.9 3.195 50.905 3.53 ;
      RECT 50.865 3.182 50.9 3.529 ;
      RECT 50.795 3.122 50.865 3.528 ;
      RECT 50.715 3.065 50.795 3.527 ;
      RECT 50.58 3.025 50.715 3.526 ;
      RECT 50.58 3.212 50.915 3.515 ;
      RECT 50.54 3.212 50.915 3.505 ;
      RECT 50.54 3.23 50.92 3.5 ;
      RECT 50.54 3.32 50.925 3.49 ;
      RECT 50.535 3.015 50.7 3.47 ;
      RECT 50.53 3.015 50.7 3.213 ;
      RECT 50.53 3.172 50.895 3.213 ;
      RECT 50.53 3.16 50.89 3.213 ;
      RECT 49.295 1.74 49.465 2.935 ;
      RECT 49.295 1.74 49.76 1.91 ;
      RECT 49.295 6.97 49.76 7.14 ;
      RECT 49.295 5.945 49.465 7.14 ;
      RECT 48.305 1.74 48.475 2.935 ;
      RECT 48.305 1.74 48.77 1.91 ;
      RECT 48.305 6.97 48.77 7.14 ;
      RECT 48.305 5.945 48.475 7.14 ;
      RECT 46.45 2.635 46.62 3.865 ;
      RECT 46.505 0.855 46.675 2.805 ;
      RECT 46.45 0.575 46.62 1.025 ;
      RECT 46.45 7.855 46.62 8.305 ;
      RECT 46.505 6.075 46.675 8.025 ;
      RECT 46.45 5.015 46.62 6.245 ;
      RECT 45.93 0.575 46.1 3.865 ;
      RECT 45.93 2.075 46.335 2.405 ;
      RECT 45.93 1.235 46.335 1.565 ;
      RECT 45.93 5.015 46.1 8.305 ;
      RECT 45.93 7.315 46.335 7.645 ;
      RECT 45.93 6.475 46.335 6.805 ;
      RECT 43.265 1.975 43.995 2.215 ;
      RECT 43.807 1.77 43.995 2.215 ;
      RECT 43.635 1.782 44.01 2.209 ;
      RECT 43.55 1.797 44.03 2.194 ;
      RECT 43.55 1.812 44.035 2.184 ;
      RECT 43.505 1.832 44.05 2.176 ;
      RECT 43.482 1.867 44.065 2.13 ;
      RECT 43.396 1.89 44.07 2.09 ;
      RECT 43.396 1.908 44.08 2.06 ;
      RECT 43.265 1.977 44.085 2.023 ;
      RECT 43.31 1.92 44.08 2.06 ;
      RECT 43.396 1.872 44.065 2.13 ;
      RECT 43.482 1.841 44.05 2.176 ;
      RECT 43.505 1.822 44.035 2.184 ;
      RECT 43.55 1.795 44.01 2.209 ;
      RECT 43.635 1.777 43.995 2.215 ;
      RECT 43.721 1.771 43.995 2.215 ;
      RECT 43.807 1.766 43.94 2.215 ;
      RECT 43.893 1.761 43.94 2.215 ;
      RECT 43.585 2.659 43.755 3.045 ;
      RECT 43.58 2.659 43.755 3.04 ;
      RECT 43.555 2.659 43.755 3.005 ;
      RECT 43.555 2.687 43.765 2.995 ;
      RECT 43.535 2.687 43.765 2.955 ;
      RECT 43.53 2.687 43.765 2.928 ;
      RECT 43.53 2.705 43.77 2.92 ;
      RECT 43.475 2.705 43.77 2.855 ;
      RECT 43.475 2.722 43.78 2.838 ;
      RECT 43.465 2.722 43.78 2.778 ;
      RECT 43.465 2.739 43.785 2.775 ;
      RECT 43.46 2.575 43.63 2.753 ;
      RECT 43.46 2.609 43.716 2.753 ;
      RECT 43.455 3.375 43.46 3.388 ;
      RECT 43.45 3.27 43.455 3.393 ;
      RECT 43.425 3.13 43.45 3.408 ;
      RECT 43.39 3.081 43.425 3.44 ;
      RECT 43.385 3.049 43.39 3.46 ;
      RECT 43.38 3.04 43.385 3.46 ;
      RECT 43.3 3.005 43.38 3.46 ;
      RECT 43.237 2.975 43.3 3.46 ;
      RECT 43.151 2.963 43.237 3.46 ;
      RECT 43.065 2.949 43.151 3.46 ;
      RECT 42.985 2.936 43.065 3.446 ;
      RECT 42.95 2.928 42.985 3.426 ;
      RECT 42.94 2.925 42.95 3.417 ;
      RECT 42.91 2.92 42.94 3.404 ;
      RECT 42.86 2.895 42.91 3.38 ;
      RECT 42.846 2.869 42.86 3.362 ;
      RECT 42.76 2.829 42.846 3.338 ;
      RECT 42.715 2.777 42.76 3.307 ;
      RECT 42.705 2.752 42.715 3.294 ;
      RECT 42.7 2.533 42.705 2.555 ;
      RECT 42.695 2.735 42.705 3.29 ;
      RECT 42.695 2.531 42.7 2.645 ;
      RECT 42.685 2.527 42.695 3.286 ;
      RECT 42.641 2.525 42.685 3.274 ;
      RECT 42.555 2.525 42.641 3.245 ;
      RECT 42.525 2.525 42.555 3.218 ;
      RECT 42.51 2.525 42.525 3.206 ;
      RECT 42.47 2.537 42.51 3.191 ;
      RECT 42.45 2.556 42.47 3.17 ;
      RECT 42.44 2.566 42.45 3.154 ;
      RECT 42.43 2.572 42.44 3.143 ;
      RECT 42.41 2.582 42.43 3.126 ;
      RECT 42.405 2.591 42.41 3.113 ;
      RECT 42.4 2.595 42.405 3.063 ;
      RECT 42.39 2.601 42.4 2.98 ;
      RECT 42.385 2.605 42.39 2.894 ;
      RECT 42.38 2.625 42.385 2.831 ;
      RECT 42.375 2.648 42.38 2.778 ;
      RECT 42.37 2.666 42.375 2.723 ;
      RECT 42.98 2.485 43.15 2.745 ;
      RECT 43.15 2.45 43.195 2.731 ;
      RECT 43.111 2.452 43.2 2.714 ;
      RECT 43 2.469 43.286 2.685 ;
      RECT 43 2.484 43.29 2.657 ;
      RECT 43 2.465 43.2 2.714 ;
      RECT 43.025 2.453 43.15 2.745 ;
      RECT 43.111 2.451 43.195 2.731 ;
      RECT 42.165 1.84 42.335 2.33 ;
      RECT 42.165 1.84 42.37 2.31 ;
      RECT 42.3 1.76 42.41 2.27 ;
      RECT 42.281 1.764 42.43 2.24 ;
      RECT 42.195 1.772 42.45 2.223 ;
      RECT 42.195 1.778 42.455 2.213 ;
      RECT 42.195 1.787 42.475 2.201 ;
      RECT 42.17 1.812 42.505 2.179 ;
      RECT 42.17 1.832 42.51 2.159 ;
      RECT 42.165 1.845 42.52 2.139 ;
      RECT 42.165 1.912 42.525 2.12 ;
      RECT 42.165 2.045 42.53 2.107 ;
      RECT 42.16 1.85 42.52 1.94 ;
      RECT 42.17 1.807 42.475 2.201 ;
      RECT 42.281 1.762 42.41 2.27 ;
      RECT 42.155 3.515 42.455 3.77 ;
      RECT 42.24 3.481 42.455 3.77 ;
      RECT 42.24 3.484 42.46 3.63 ;
      RECT 42.175 3.505 42.46 3.63 ;
      RECT 42.21 3.495 42.455 3.77 ;
      RECT 42.205 3.5 42.46 3.63 ;
      RECT 42.24 3.479 42.441 3.77 ;
      RECT 42.326 3.47 42.441 3.77 ;
      RECT 42.326 3.464 42.355 3.77 ;
      RECT 41.815 3.105 41.825 3.595 ;
      RECT 41.475 3.04 41.485 3.34 ;
      RECT 41.99 3.212 41.995 3.431 ;
      RECT 41.98 3.192 41.99 3.448 ;
      RECT 41.97 3.172 41.98 3.478 ;
      RECT 41.965 3.162 41.97 3.493 ;
      RECT 41.96 3.158 41.965 3.498 ;
      RECT 41.945 3.15 41.96 3.505 ;
      RECT 41.905 3.13 41.945 3.53 ;
      RECT 41.88 3.112 41.905 3.563 ;
      RECT 41.875 3.11 41.88 3.576 ;
      RECT 41.855 3.107 41.875 3.58 ;
      RECT 41.825 3.105 41.855 3.59 ;
      RECT 41.755 3.107 41.815 3.591 ;
      RECT 41.735 3.107 41.755 3.585 ;
      RECT 41.71 3.105 41.735 3.582 ;
      RECT 41.675 3.1 41.71 3.578 ;
      RECT 41.655 3.094 41.675 3.565 ;
      RECT 41.645 3.091 41.655 3.553 ;
      RECT 41.625 3.088 41.645 3.538 ;
      RECT 41.605 3.084 41.625 3.52 ;
      RECT 41.6 3.081 41.605 3.51 ;
      RECT 41.595 3.08 41.6 3.508 ;
      RECT 41.585 3.077 41.595 3.5 ;
      RECT 41.575 3.071 41.585 3.483 ;
      RECT 41.565 3.065 41.575 3.465 ;
      RECT 41.555 3.059 41.565 3.453 ;
      RECT 41.545 3.053 41.555 3.433 ;
      RECT 41.54 3.049 41.545 3.418 ;
      RECT 41.535 3.047 41.54 3.41 ;
      RECT 41.53 3.045 41.535 3.403 ;
      RECT 41.525 3.043 41.53 3.393 ;
      RECT 41.52 3.041 41.525 3.387 ;
      RECT 41.51 3.04 41.52 3.377 ;
      RECT 41.5 3.04 41.51 3.368 ;
      RECT 41.485 3.04 41.5 3.353 ;
      RECT 41.445 3.04 41.475 3.337 ;
      RECT 41.425 3.042 41.445 3.332 ;
      RECT 41.42 3.047 41.425 3.33 ;
      RECT 41.39 3.055 41.42 3.328 ;
      RECT 41.36 3.07 41.39 3.327 ;
      RECT 41.315 3.092 41.36 3.332 ;
      RECT 41.31 3.107 41.315 3.336 ;
      RECT 41.295 3.112 41.31 3.338 ;
      RECT 41.29 3.116 41.295 3.34 ;
      RECT 41.23 3.139 41.29 3.349 ;
      RECT 41.21 3.165 41.23 3.362 ;
      RECT 41.2 3.172 41.21 3.366 ;
      RECT 41.185 3.179 41.2 3.369 ;
      RECT 41.165 3.189 41.185 3.372 ;
      RECT 41.16 3.197 41.165 3.375 ;
      RECT 41.115 3.202 41.16 3.382 ;
      RECT 41.105 3.205 41.115 3.389 ;
      RECT 41.095 3.205 41.105 3.393 ;
      RECT 41.06 3.207 41.095 3.405 ;
      RECT 41.04 3.21 41.06 3.418 ;
      RECT 41 3.213 41.04 3.429 ;
      RECT 40.985 3.215 41 3.442 ;
      RECT 40.975 3.215 40.985 3.447 ;
      RECT 40.95 3.216 40.975 3.455 ;
      RECT 40.94 3.218 40.95 3.46 ;
      RECT 40.935 3.219 40.94 3.463 ;
      RECT 40.91 3.217 40.935 3.466 ;
      RECT 40.895 3.215 40.91 3.467 ;
      RECT 40.875 3.212 40.895 3.469 ;
      RECT 40.855 3.207 40.875 3.469 ;
      RECT 40.795 3.202 40.855 3.466 ;
      RECT 40.76 3.177 40.795 3.462 ;
      RECT 40.75 3.154 40.76 3.46 ;
      RECT 40.72 3.131 40.75 3.46 ;
      RECT 40.71 3.11 40.72 3.46 ;
      RECT 40.685 3.092 40.71 3.458 ;
      RECT 40.67 3.07 40.685 3.455 ;
      RECT 40.655 3.052 40.67 3.453 ;
      RECT 40.635 3.042 40.655 3.451 ;
      RECT 40.62 3.037 40.635 3.45 ;
      RECT 40.605 3.035 40.62 3.449 ;
      RECT 40.575 3.036 40.605 3.447 ;
      RECT 40.555 3.039 40.575 3.445 ;
      RECT 40.498 3.043 40.555 3.445 ;
      RECT 40.412 3.052 40.498 3.445 ;
      RECT 40.326 3.063 40.412 3.445 ;
      RECT 40.24 3.074 40.326 3.445 ;
      RECT 40.22 3.081 40.24 3.453 ;
      RECT 40.21 3.084 40.22 3.46 ;
      RECT 40.145 3.089 40.21 3.478 ;
      RECT 40.115 3.096 40.145 3.503 ;
      RECT 40.105 3.099 40.115 3.51 ;
      RECT 40.06 3.103 40.105 3.515 ;
      RECT 40.03 3.108 40.06 3.52 ;
      RECT 40.029 3.11 40.03 3.52 ;
      RECT 39.943 3.116 40.029 3.52 ;
      RECT 39.857 3.127 39.943 3.52 ;
      RECT 39.771 3.139 39.857 3.52 ;
      RECT 39.685 3.15 39.771 3.52 ;
      RECT 39.67 3.157 39.685 3.515 ;
      RECT 39.665 3.159 39.67 3.509 ;
      RECT 39.645 3.17 39.665 3.504 ;
      RECT 39.635 3.188 39.645 3.498 ;
      RECT 39.63 3.2 39.635 3.298 ;
      RECT 41.925 1.953 41.945 2.04 ;
      RECT 41.92 1.888 41.925 2.072 ;
      RECT 41.91 1.855 41.92 2.077 ;
      RECT 41.905 1.835 41.91 2.083 ;
      RECT 41.875 1.835 41.905 2.1 ;
      RECT 41.826 1.835 41.875 2.136 ;
      RECT 41.74 1.835 41.826 2.194 ;
      RECT 41.711 1.845 41.74 2.243 ;
      RECT 41.625 1.887 41.711 2.296 ;
      RECT 41.605 1.925 41.625 2.343 ;
      RECT 41.58 1.942 41.605 2.363 ;
      RECT 41.57 1.956 41.58 2.383 ;
      RECT 41.565 1.962 41.57 2.393 ;
      RECT 41.56 1.966 41.565 2.4 ;
      RECT 41.51 1.986 41.56 2.405 ;
      RECT 41.445 2.03 41.51 2.405 ;
      RECT 41.42 2.08 41.445 2.405 ;
      RECT 41.41 2.11 41.42 2.405 ;
      RECT 41.405 2.137 41.41 2.405 ;
      RECT 41.4 2.155 41.405 2.405 ;
      RECT 41.39 2.197 41.4 2.405 ;
      RECT 41.74 2.755 41.91 2.93 ;
      RECT 41.68 2.583 41.74 2.918 ;
      RECT 41.67 2.576 41.68 2.901 ;
      RECT 41.625 2.755 41.91 2.881 ;
      RECT 41.606 2.755 41.91 2.859 ;
      RECT 41.52 2.755 41.91 2.824 ;
      RECT 41.5 2.575 41.67 2.78 ;
      RECT 41.5 2.722 41.905 2.78 ;
      RECT 41.5 2.67 41.88 2.78 ;
      RECT 41.5 2.625 41.845 2.78 ;
      RECT 41.5 2.607 41.81 2.78 ;
      RECT 41.5 2.597 41.805 2.78 ;
      RECT 41.67 7.855 41.84 8.305 ;
      RECT 41.725 6.075 41.895 8.025 ;
      RECT 41.67 5.015 41.84 6.245 ;
      RECT 41.15 5.015 41.32 8.305 ;
      RECT 41.15 7.315 41.555 7.645 ;
      RECT 41.15 6.475 41.555 6.805 ;
      RECT 41.22 3.555 41.41 3.78 ;
      RECT 41.21 3.556 41.415 3.775 ;
      RECT 41.21 3.558 41.425 3.755 ;
      RECT 41.21 3.562 41.43 3.74 ;
      RECT 41.21 3.549 41.38 3.775 ;
      RECT 41.21 3.552 41.405 3.775 ;
      RECT 41.22 3.548 41.38 3.78 ;
      RECT 41.306 3.546 41.38 3.78 ;
      RECT 40.93 2.797 41.1 3.035 ;
      RECT 40.93 2.797 41.186 2.949 ;
      RECT 40.93 2.797 41.19 2.859 ;
      RECT 40.98 2.57 41.2 2.838 ;
      RECT 40.975 2.587 41.205 2.811 ;
      RECT 40.94 2.745 41.205 2.811 ;
      RECT 40.96 2.595 41.1 3.035 ;
      RECT 40.95 2.677 41.21 2.794 ;
      RECT 40.945 2.725 41.21 2.794 ;
      RECT 40.95 2.635 41.205 2.811 ;
      RECT 40.975 2.572 41.2 2.838 ;
      RECT 40.54 2.547 40.71 2.745 ;
      RECT 40.54 2.547 40.755 2.72 ;
      RECT 40.61 2.49 40.78 2.678 ;
      RECT 40.585 2.505 40.78 2.678 ;
      RECT 40.2 2.551 40.23 2.745 ;
      RECT 40.195 2.523 40.2 2.745 ;
      RECT 40.165 2.497 40.195 2.747 ;
      RECT 40.14 2.455 40.165 2.75 ;
      RECT 40.13 2.427 40.14 2.752 ;
      RECT 40.095 2.407 40.13 2.754 ;
      RECT 40.03 2.392 40.095 2.76 ;
      RECT 39.98 2.39 40.03 2.766 ;
      RECT 39.957 2.392 39.98 2.771 ;
      RECT 39.871 2.403 39.957 2.777 ;
      RECT 39.785 2.421 39.871 2.787 ;
      RECT 39.77 2.432 39.785 2.793 ;
      RECT 39.7 2.455 39.77 2.799 ;
      RECT 39.645 2.487 39.7 2.807 ;
      RECT 39.605 2.51 39.645 2.813 ;
      RECT 39.591 2.523 39.605 2.816 ;
      RECT 39.505 2.545 39.591 2.822 ;
      RECT 39.49 2.57 39.505 2.828 ;
      RECT 39.45 2.585 39.49 2.832 ;
      RECT 39.4 2.6 39.45 2.837 ;
      RECT 39.375 2.607 39.4 2.841 ;
      RECT 39.315 2.602 39.375 2.845 ;
      RECT 39.3 2.593 39.315 2.849 ;
      RECT 39.23 2.583 39.3 2.845 ;
      RECT 39.205 2.575 39.225 2.835 ;
      RECT 39.146 2.575 39.205 2.813 ;
      RECT 39.06 2.575 39.146 2.77 ;
      RECT 39.225 2.575 39.23 2.84 ;
      RECT 39.92 1.806 40.09 2.14 ;
      RECT 39.89 1.806 40.09 2.135 ;
      RECT 39.83 1.773 39.89 2.123 ;
      RECT 39.83 1.829 40.1 2.118 ;
      RECT 39.805 1.829 40.1 2.112 ;
      RECT 39.8 1.77 39.83 2.109 ;
      RECT 39.785 1.776 39.92 2.107 ;
      RECT 39.78 1.784 40.005 2.095 ;
      RECT 39.78 1.836 40.115 2.048 ;
      RECT 39.765 1.792 40.005 2.043 ;
      RECT 39.765 1.862 40.125 1.984 ;
      RECT 39.735 1.812 40.09 1.945 ;
      RECT 39.735 1.902 40.135 1.941 ;
      RECT 39.785 1.781 40.005 2.107 ;
      RECT 39.125 2.111 39.18 2.375 ;
      RECT 39.125 2.111 39.245 2.374 ;
      RECT 39.125 2.111 39.27 2.373 ;
      RECT 39.125 2.111 39.335 2.372 ;
      RECT 39.27 2.077 39.35 2.371 ;
      RECT 39.085 2.121 39.495 2.37 ;
      RECT 39.125 2.118 39.495 2.37 ;
      RECT 39.085 2.126 39.5 2.363 ;
      RECT 39.07 2.128 39.5 2.362 ;
      RECT 39.07 2.135 39.505 2.358 ;
      RECT 39.05 2.134 39.5 2.354 ;
      RECT 39.05 2.142 39.51 2.353 ;
      RECT 39.045 2.139 39.505 2.349 ;
      RECT 39.045 2.152 39.52 2.348 ;
      RECT 39.03 2.142 39.51 2.347 ;
      RECT 38.995 2.155 39.52 2.34 ;
      RECT 39.18 2.11 39.49 2.37 ;
      RECT 39.18 2.095 39.44 2.37 ;
      RECT 39.245 2.082 39.375 2.37 ;
      RECT 38.79 3.171 38.805 3.564 ;
      RECT 38.755 3.176 38.805 3.563 ;
      RECT 38.79 3.175 38.85 3.562 ;
      RECT 38.735 3.186 38.85 3.561 ;
      RECT 38.75 3.182 38.85 3.561 ;
      RECT 38.715 3.192 38.925 3.558 ;
      RECT 38.715 3.211 38.97 3.556 ;
      RECT 38.715 3.218 38.975 3.553 ;
      RECT 38.7 3.195 38.925 3.55 ;
      RECT 38.68 3.2 38.925 3.543 ;
      RECT 38.675 3.204 38.925 3.539 ;
      RECT 38.675 3.221 38.985 3.538 ;
      RECT 38.655 3.215 38.97 3.534 ;
      RECT 38.655 3.224 38.99 3.528 ;
      RECT 38.65 3.23 38.99 3.3 ;
      RECT 38.715 3.19 38.85 3.558 ;
      RECT 38.59 2.553 38.79 2.865 ;
      RECT 38.665 2.531 38.79 2.865 ;
      RECT 38.605 2.55 38.795 2.85 ;
      RECT 38.575 2.561 38.795 2.848 ;
      RECT 38.59 2.556 38.8 2.814 ;
      RECT 38.575 2.66 38.805 2.781 ;
      RECT 38.605 2.532 38.79 2.865 ;
      RECT 38.665 2.51 38.765 2.865 ;
      RECT 38.69 2.507 38.765 2.865 ;
      RECT 38.69 2.502 38.71 2.865 ;
      RECT 38.095 2.57 38.27 2.745 ;
      RECT 38.09 2.57 38.27 2.743 ;
      RECT 38.065 2.57 38.27 2.738 ;
      RECT 38.01 2.55 38.18 2.728 ;
      RECT 38.01 2.557 38.245 2.728 ;
      RECT 38.095 3.237 38.11 3.42 ;
      RECT 38.085 3.215 38.095 3.42 ;
      RECT 38.07 3.195 38.085 3.42 ;
      RECT 38.06 3.17 38.07 3.42 ;
      RECT 38.03 3.135 38.06 3.42 ;
      RECT 37.995 3.075 38.03 3.42 ;
      RECT 37.99 3.037 37.995 3.42 ;
      RECT 37.94 2.988 37.99 3.42 ;
      RECT 37.93 2.938 37.94 3.408 ;
      RECT 37.915 2.917 37.93 3.368 ;
      RECT 37.895 2.885 37.915 3.318 ;
      RECT 37.87 2.841 37.895 3.258 ;
      RECT 37.865 2.813 37.87 3.213 ;
      RECT 37.86 2.804 37.865 3.199 ;
      RECT 37.855 2.797 37.86 3.186 ;
      RECT 37.85 2.792 37.855 3.175 ;
      RECT 37.845 2.777 37.85 3.165 ;
      RECT 37.84 2.755 37.845 3.152 ;
      RECT 37.83 2.715 37.84 3.127 ;
      RECT 37.805 2.645 37.83 3.083 ;
      RECT 37.8 2.585 37.805 3.048 ;
      RECT 37.785 2.565 37.8 3.015 ;
      RECT 37.78 2.565 37.785 2.99 ;
      RECT 37.75 2.565 37.78 2.945 ;
      RECT 37.705 2.565 37.75 2.885 ;
      RECT 37.63 2.565 37.705 2.833 ;
      RECT 37.625 2.565 37.63 2.798 ;
      RECT 37.62 2.565 37.625 2.788 ;
      RECT 37.615 2.565 37.62 2.768 ;
      RECT 37.88 1.785 38.05 2.255 ;
      RECT 37.825 1.778 38.02 2.239 ;
      RECT 37.825 1.792 38.055 2.238 ;
      RECT 37.81 1.793 38.055 2.219 ;
      RECT 37.805 1.811 38.055 2.205 ;
      RECT 37.81 1.794 38.06 2.203 ;
      RECT 37.795 1.825 38.06 2.188 ;
      RECT 37.81 1.8 38.065 2.173 ;
      RECT 37.79 1.84 38.065 2.17 ;
      RECT 37.805 1.812 38.07 2.155 ;
      RECT 37.805 1.824 38.075 2.135 ;
      RECT 37.79 1.84 38.08 2.118 ;
      RECT 37.79 1.85 38.085 1.973 ;
      RECT 37.785 1.85 38.085 1.93 ;
      RECT 37.785 1.865 38.09 1.908 ;
      RECT 37.88 1.775 38.02 2.255 ;
      RECT 37.88 1.773 37.99 2.255 ;
      RECT 37.966 1.77 37.99 2.255 ;
      RECT 37.625 3.437 37.63 3.483 ;
      RECT 37.615 3.285 37.625 3.507 ;
      RECT 37.61 3.13 37.615 3.532 ;
      RECT 37.595 3.092 37.61 3.543 ;
      RECT 37.59 3.075 37.595 3.55 ;
      RECT 37.58 3.063 37.59 3.557 ;
      RECT 37.575 3.054 37.58 3.559 ;
      RECT 37.57 3.052 37.575 3.563 ;
      RECT 37.525 3.043 37.57 3.578 ;
      RECT 37.52 3.035 37.525 3.592 ;
      RECT 37.515 3.032 37.52 3.596 ;
      RECT 37.5 3.027 37.515 3.604 ;
      RECT 37.445 3.017 37.5 3.615 ;
      RECT 37.41 3.005 37.445 3.616 ;
      RECT 37.401 3 37.41 3.61 ;
      RECT 37.315 3 37.401 3.6 ;
      RECT 37.285 3 37.315 3.578 ;
      RECT 37.275 3 37.28 3.558 ;
      RECT 37.27 3 37.275 3.52 ;
      RECT 37.265 3 37.27 3.478 ;
      RECT 37.26 3 37.265 3.438 ;
      RECT 37.255 3 37.26 3.368 ;
      RECT 37.245 3 37.255 3.29 ;
      RECT 37.24 3 37.245 3.19 ;
      RECT 37.28 3 37.285 3.56 ;
      RECT 36.775 3.082 36.865 3.56 ;
      RECT 36.76 3.085 36.88 3.558 ;
      RECT 36.775 3.084 36.88 3.558 ;
      RECT 36.74 3.091 36.905 3.548 ;
      RECT 36.76 3.085 36.905 3.548 ;
      RECT 36.725 3.097 36.905 3.536 ;
      RECT 36.76 3.088 36.955 3.529 ;
      RECT 36.711 3.105 36.955 3.527 ;
      RECT 36.74 3.095 36.965 3.515 ;
      RECT 36.711 3.116 36.995 3.506 ;
      RECT 36.625 3.14 36.995 3.5 ;
      RECT 36.625 3.153 37.035 3.483 ;
      RECT 36.62 3.175 37.035 3.476 ;
      RECT 36.59 3.19 37.035 3.466 ;
      RECT 36.585 3.201 37.035 3.456 ;
      RECT 36.555 3.214 37.035 3.447 ;
      RECT 36.54 3.232 37.035 3.436 ;
      RECT 36.515 3.245 37.035 3.426 ;
      RECT 36.775 3.081 36.785 3.56 ;
      RECT 36.821 2.505 36.86 2.75 ;
      RECT 36.735 2.505 36.87 2.748 ;
      RECT 36.62 2.53 36.87 2.745 ;
      RECT 36.62 2.53 36.875 2.743 ;
      RECT 36.62 2.53 36.89 2.738 ;
      RECT 36.726 2.505 36.905 2.718 ;
      RECT 36.64 2.513 36.905 2.718 ;
      RECT 36.31 1.865 36.48 2.3 ;
      RECT 36.3 1.899 36.48 2.283 ;
      RECT 36.38 1.835 36.55 2.27 ;
      RECT 36.285 1.91 36.55 2.248 ;
      RECT 36.38 1.845 36.555 2.238 ;
      RECT 36.31 1.897 36.585 2.223 ;
      RECT 36.27 1.923 36.585 2.208 ;
      RECT 36.27 1.965 36.595 2.188 ;
      RECT 36.265 1.99 36.6 2.17 ;
      RECT 36.265 2 36.605 2.155 ;
      RECT 36.26 1.937 36.585 2.153 ;
      RECT 36.26 2.01 36.61 2.138 ;
      RECT 36.255 1.947 36.585 2.135 ;
      RECT 36.25 2.031 36.615 2.118 ;
      RECT 36.25 2.063 36.62 2.098 ;
      RECT 36.245 1.977 36.595 2.09 ;
      RECT 36.25 1.962 36.585 2.118 ;
      RECT 36.265 1.932 36.585 2.17 ;
      RECT 36.11 2.519 36.335 2.775 ;
      RECT 36.11 2.552 36.355 2.765 ;
      RECT 36.075 2.552 36.355 2.763 ;
      RECT 36.075 2.565 36.36 2.753 ;
      RECT 36.075 2.585 36.37 2.745 ;
      RECT 36.075 2.682 36.375 2.738 ;
      RECT 36.055 2.43 36.185 2.728 ;
      RECT 36.01 2.585 36.37 2.67 ;
      RECT 36 2.43 36.185 2.615 ;
      RECT 36 2.462 36.271 2.615 ;
      RECT 35.965 2.992 35.985 3.17 ;
      RECT 35.93 2.945 35.965 3.17 ;
      RECT 35.915 2.885 35.93 3.17 ;
      RECT 35.89 2.832 35.915 3.17 ;
      RECT 35.875 2.785 35.89 3.17 ;
      RECT 35.855 2.762 35.875 3.17 ;
      RECT 35.83 2.727 35.855 3.17 ;
      RECT 35.82 2.573 35.83 3.17 ;
      RECT 35.79 2.568 35.82 3.161 ;
      RECT 35.785 2.565 35.79 3.151 ;
      RECT 35.77 2.565 35.785 3.125 ;
      RECT 35.765 2.565 35.77 3.088 ;
      RECT 35.74 2.565 35.765 3.04 ;
      RECT 35.72 2.565 35.74 2.965 ;
      RECT 35.71 2.565 35.72 2.925 ;
      RECT 35.705 2.565 35.71 2.9 ;
      RECT 35.7 2.565 35.705 2.883 ;
      RECT 35.695 2.565 35.7 2.865 ;
      RECT 35.69 2.566 35.695 2.855 ;
      RECT 35.68 2.568 35.69 2.823 ;
      RECT 35.67 2.57 35.68 2.79 ;
      RECT 35.66 2.573 35.67 2.763 ;
      RECT 35.985 3 36.21 3.17 ;
      RECT 35.315 1.812 35.485 2.265 ;
      RECT 35.315 1.812 35.575 2.231 ;
      RECT 35.315 1.812 35.605 2.215 ;
      RECT 35.315 1.812 35.635 2.188 ;
      RECT 35.571 1.79 35.65 2.17 ;
      RECT 35.35 1.797 35.655 2.155 ;
      RECT 35.35 1.805 35.665 2.118 ;
      RECT 35.31 1.832 35.665 2.09 ;
      RECT 35.295 1.845 35.665 2.055 ;
      RECT 35.315 1.82 35.685 2.045 ;
      RECT 35.29 1.885 35.685 2.015 ;
      RECT 35.29 1.915 35.69 1.998 ;
      RECT 35.285 1.945 35.69 1.985 ;
      RECT 35.35 1.794 35.65 2.17 ;
      RECT 35.485 1.791 35.571 2.249 ;
      RECT 35.436 1.792 35.65 2.17 ;
      RECT 35.58 3.452 35.625 3.645 ;
      RECT 35.57 3.422 35.58 3.645 ;
      RECT 35.565 3.407 35.57 3.645 ;
      RECT 35.525 3.317 35.565 3.645 ;
      RECT 35.52 3.23 35.525 3.645 ;
      RECT 35.51 3.2 35.52 3.645 ;
      RECT 35.505 3.16 35.51 3.645 ;
      RECT 35.495 3.122 35.505 3.645 ;
      RECT 35.49 3.087 35.495 3.645 ;
      RECT 35.47 3.04 35.49 3.645 ;
      RECT 35.455 2.965 35.47 3.645 ;
      RECT 35.45 2.92 35.455 3.64 ;
      RECT 35.445 2.9 35.45 3.613 ;
      RECT 35.44 2.88 35.445 3.598 ;
      RECT 35.435 2.855 35.44 3.578 ;
      RECT 35.43 2.833 35.435 3.563 ;
      RECT 35.425 2.811 35.43 3.545 ;
      RECT 35.42 2.79 35.425 3.535 ;
      RECT 35.41 2.762 35.42 3.505 ;
      RECT 35.4 2.725 35.41 3.473 ;
      RECT 35.39 2.685 35.4 3.44 ;
      RECT 35.38 2.663 35.39 3.41 ;
      RECT 35.35 2.615 35.38 3.342 ;
      RECT 35.335 2.575 35.35 3.269 ;
      RECT 35.325 2.575 35.335 3.235 ;
      RECT 35.32 2.575 35.325 3.21 ;
      RECT 35.315 2.575 35.32 3.195 ;
      RECT 35.31 2.575 35.315 3.173 ;
      RECT 35.305 2.575 35.31 3.16 ;
      RECT 35.29 2.575 35.305 3.125 ;
      RECT 35.27 2.575 35.29 3.065 ;
      RECT 35.26 2.575 35.27 3.015 ;
      RECT 35.24 2.575 35.26 2.963 ;
      RECT 35.22 2.575 35.24 2.92 ;
      RECT 35.21 2.575 35.22 2.908 ;
      RECT 35.18 2.575 35.21 2.895 ;
      RECT 35.15 2.596 35.18 2.875 ;
      RECT 35.14 2.624 35.15 2.855 ;
      RECT 35.125 2.641 35.14 2.823 ;
      RECT 35.12 2.655 35.125 2.79 ;
      RECT 35.115 2.663 35.12 2.763 ;
      RECT 35.11 2.671 35.115 2.725 ;
      RECT 35.115 3.195 35.12 3.53 ;
      RECT 35.08 3.182 35.115 3.529 ;
      RECT 35.01 3.122 35.08 3.528 ;
      RECT 34.93 3.065 35.01 3.527 ;
      RECT 34.795 3.025 34.93 3.526 ;
      RECT 34.795 3.212 35.13 3.515 ;
      RECT 34.755 3.212 35.13 3.505 ;
      RECT 34.755 3.23 35.135 3.5 ;
      RECT 34.755 3.32 35.14 3.49 ;
      RECT 34.75 3.015 34.915 3.47 ;
      RECT 34.745 3.015 34.915 3.213 ;
      RECT 34.745 3.172 35.11 3.213 ;
      RECT 34.745 3.16 35.105 3.213 ;
      RECT 33.52 1.74 33.69 2.935 ;
      RECT 33.52 1.74 33.985 1.91 ;
      RECT 33.52 6.97 33.985 7.14 ;
      RECT 33.52 5.945 33.69 7.14 ;
      RECT 32.53 1.74 32.7 2.935 ;
      RECT 32.53 1.74 32.995 1.91 ;
      RECT 32.53 6.97 32.995 7.14 ;
      RECT 32.53 5.945 32.7 7.14 ;
      RECT 30.675 2.635 30.845 3.865 ;
      RECT 30.73 0.855 30.9 2.805 ;
      RECT 30.675 0.575 30.845 1.025 ;
      RECT 30.675 7.855 30.845 8.305 ;
      RECT 30.73 6.075 30.9 8.025 ;
      RECT 30.675 5.015 30.845 6.245 ;
      RECT 30.155 0.575 30.325 3.865 ;
      RECT 30.155 2.075 30.56 2.405 ;
      RECT 30.155 1.235 30.56 1.565 ;
      RECT 30.155 5.015 30.325 8.305 ;
      RECT 30.155 7.315 30.56 7.645 ;
      RECT 30.155 6.475 30.56 6.805 ;
      RECT 27.49 1.975 28.22 2.215 ;
      RECT 28.032 1.77 28.22 2.215 ;
      RECT 27.86 1.782 28.235 2.209 ;
      RECT 27.775 1.797 28.255 2.194 ;
      RECT 27.775 1.812 28.26 2.184 ;
      RECT 27.73 1.832 28.275 2.176 ;
      RECT 27.707 1.867 28.29 2.13 ;
      RECT 27.621 1.89 28.295 2.09 ;
      RECT 27.621 1.908 28.305 2.06 ;
      RECT 27.49 1.977 28.31 2.023 ;
      RECT 27.535 1.92 28.305 2.06 ;
      RECT 27.621 1.872 28.29 2.13 ;
      RECT 27.707 1.841 28.275 2.176 ;
      RECT 27.73 1.822 28.26 2.184 ;
      RECT 27.775 1.795 28.235 2.209 ;
      RECT 27.86 1.777 28.22 2.215 ;
      RECT 27.946 1.771 28.22 2.215 ;
      RECT 28.032 1.766 28.165 2.215 ;
      RECT 28.118 1.761 28.165 2.215 ;
      RECT 27.81 2.659 27.98 3.045 ;
      RECT 27.805 2.659 27.98 3.04 ;
      RECT 27.78 2.659 27.98 3.005 ;
      RECT 27.78 2.687 27.99 2.995 ;
      RECT 27.76 2.687 27.99 2.955 ;
      RECT 27.755 2.687 27.99 2.928 ;
      RECT 27.755 2.705 27.995 2.92 ;
      RECT 27.7 2.705 27.995 2.855 ;
      RECT 27.7 2.722 28.005 2.838 ;
      RECT 27.69 2.722 28.005 2.778 ;
      RECT 27.69 2.739 28.01 2.775 ;
      RECT 27.685 2.575 27.855 2.753 ;
      RECT 27.685 2.609 27.941 2.753 ;
      RECT 27.68 3.375 27.685 3.388 ;
      RECT 27.675 3.27 27.68 3.393 ;
      RECT 27.65 3.13 27.675 3.408 ;
      RECT 27.615 3.081 27.65 3.44 ;
      RECT 27.61 3.049 27.615 3.46 ;
      RECT 27.605 3.04 27.61 3.46 ;
      RECT 27.525 3.005 27.605 3.46 ;
      RECT 27.462 2.975 27.525 3.46 ;
      RECT 27.376 2.963 27.462 3.46 ;
      RECT 27.29 2.949 27.376 3.46 ;
      RECT 27.21 2.936 27.29 3.446 ;
      RECT 27.175 2.928 27.21 3.426 ;
      RECT 27.165 2.925 27.175 3.417 ;
      RECT 27.135 2.92 27.165 3.404 ;
      RECT 27.085 2.895 27.135 3.38 ;
      RECT 27.071 2.869 27.085 3.362 ;
      RECT 26.985 2.829 27.071 3.338 ;
      RECT 26.94 2.777 26.985 3.307 ;
      RECT 26.93 2.752 26.94 3.294 ;
      RECT 26.925 2.533 26.93 2.555 ;
      RECT 26.92 2.735 26.93 3.29 ;
      RECT 26.92 2.531 26.925 2.645 ;
      RECT 26.91 2.527 26.92 3.286 ;
      RECT 26.866 2.525 26.91 3.274 ;
      RECT 26.78 2.525 26.866 3.245 ;
      RECT 26.75 2.525 26.78 3.218 ;
      RECT 26.735 2.525 26.75 3.206 ;
      RECT 26.695 2.537 26.735 3.191 ;
      RECT 26.675 2.556 26.695 3.17 ;
      RECT 26.665 2.566 26.675 3.154 ;
      RECT 26.655 2.572 26.665 3.143 ;
      RECT 26.635 2.582 26.655 3.126 ;
      RECT 26.63 2.591 26.635 3.113 ;
      RECT 26.625 2.595 26.63 3.063 ;
      RECT 26.615 2.601 26.625 2.98 ;
      RECT 26.61 2.605 26.615 2.894 ;
      RECT 26.605 2.625 26.61 2.831 ;
      RECT 26.6 2.648 26.605 2.778 ;
      RECT 26.595 2.666 26.6 2.723 ;
      RECT 27.205 2.485 27.375 2.745 ;
      RECT 27.375 2.45 27.42 2.731 ;
      RECT 27.336 2.452 27.425 2.714 ;
      RECT 27.225 2.469 27.511 2.685 ;
      RECT 27.225 2.484 27.515 2.657 ;
      RECT 27.225 2.465 27.425 2.714 ;
      RECT 27.25 2.453 27.375 2.745 ;
      RECT 27.336 2.451 27.42 2.731 ;
      RECT 26.39 1.84 26.56 2.33 ;
      RECT 26.39 1.84 26.595 2.31 ;
      RECT 26.525 1.76 26.635 2.27 ;
      RECT 26.506 1.764 26.655 2.24 ;
      RECT 26.42 1.772 26.675 2.223 ;
      RECT 26.42 1.778 26.68 2.213 ;
      RECT 26.42 1.787 26.7 2.201 ;
      RECT 26.395 1.812 26.73 2.179 ;
      RECT 26.395 1.832 26.735 2.159 ;
      RECT 26.39 1.845 26.745 2.139 ;
      RECT 26.39 1.912 26.75 2.12 ;
      RECT 26.39 2.045 26.755 2.107 ;
      RECT 26.385 1.85 26.745 1.94 ;
      RECT 26.395 1.807 26.7 2.201 ;
      RECT 26.506 1.762 26.635 2.27 ;
      RECT 26.38 3.515 26.68 3.77 ;
      RECT 26.465 3.481 26.68 3.77 ;
      RECT 26.465 3.484 26.685 3.63 ;
      RECT 26.4 3.505 26.685 3.63 ;
      RECT 26.435 3.495 26.68 3.77 ;
      RECT 26.43 3.5 26.685 3.63 ;
      RECT 26.465 3.479 26.666 3.77 ;
      RECT 26.551 3.47 26.666 3.77 ;
      RECT 26.551 3.464 26.58 3.77 ;
      RECT 26.04 3.105 26.05 3.595 ;
      RECT 25.7 3.04 25.71 3.34 ;
      RECT 26.215 3.212 26.22 3.431 ;
      RECT 26.205 3.192 26.215 3.448 ;
      RECT 26.195 3.172 26.205 3.478 ;
      RECT 26.19 3.162 26.195 3.493 ;
      RECT 26.185 3.158 26.19 3.498 ;
      RECT 26.17 3.15 26.185 3.505 ;
      RECT 26.13 3.13 26.17 3.53 ;
      RECT 26.105 3.112 26.13 3.563 ;
      RECT 26.1 3.11 26.105 3.576 ;
      RECT 26.08 3.107 26.1 3.58 ;
      RECT 26.05 3.105 26.08 3.59 ;
      RECT 25.98 3.107 26.04 3.591 ;
      RECT 25.96 3.107 25.98 3.585 ;
      RECT 25.935 3.105 25.96 3.582 ;
      RECT 25.9 3.1 25.935 3.578 ;
      RECT 25.88 3.094 25.9 3.565 ;
      RECT 25.87 3.091 25.88 3.553 ;
      RECT 25.85 3.088 25.87 3.538 ;
      RECT 25.83 3.084 25.85 3.52 ;
      RECT 25.825 3.081 25.83 3.51 ;
      RECT 25.82 3.08 25.825 3.508 ;
      RECT 25.81 3.077 25.82 3.5 ;
      RECT 25.8 3.071 25.81 3.483 ;
      RECT 25.79 3.065 25.8 3.465 ;
      RECT 25.78 3.059 25.79 3.453 ;
      RECT 25.77 3.053 25.78 3.433 ;
      RECT 25.765 3.049 25.77 3.418 ;
      RECT 25.76 3.047 25.765 3.41 ;
      RECT 25.755 3.045 25.76 3.403 ;
      RECT 25.75 3.043 25.755 3.393 ;
      RECT 25.745 3.041 25.75 3.387 ;
      RECT 25.735 3.04 25.745 3.377 ;
      RECT 25.725 3.04 25.735 3.368 ;
      RECT 25.71 3.04 25.725 3.353 ;
      RECT 25.67 3.04 25.7 3.337 ;
      RECT 25.65 3.042 25.67 3.332 ;
      RECT 25.645 3.047 25.65 3.33 ;
      RECT 25.615 3.055 25.645 3.328 ;
      RECT 25.585 3.07 25.615 3.327 ;
      RECT 25.54 3.092 25.585 3.332 ;
      RECT 25.535 3.107 25.54 3.336 ;
      RECT 25.52 3.112 25.535 3.338 ;
      RECT 25.515 3.116 25.52 3.34 ;
      RECT 25.455 3.139 25.515 3.349 ;
      RECT 25.435 3.165 25.455 3.362 ;
      RECT 25.425 3.172 25.435 3.366 ;
      RECT 25.41 3.179 25.425 3.369 ;
      RECT 25.39 3.189 25.41 3.372 ;
      RECT 25.385 3.197 25.39 3.375 ;
      RECT 25.34 3.202 25.385 3.382 ;
      RECT 25.33 3.205 25.34 3.389 ;
      RECT 25.32 3.205 25.33 3.393 ;
      RECT 25.285 3.207 25.32 3.405 ;
      RECT 25.265 3.21 25.285 3.418 ;
      RECT 25.225 3.213 25.265 3.429 ;
      RECT 25.21 3.215 25.225 3.442 ;
      RECT 25.2 3.215 25.21 3.447 ;
      RECT 25.175 3.216 25.2 3.455 ;
      RECT 25.165 3.218 25.175 3.46 ;
      RECT 25.16 3.219 25.165 3.463 ;
      RECT 25.135 3.217 25.16 3.466 ;
      RECT 25.12 3.215 25.135 3.467 ;
      RECT 25.1 3.212 25.12 3.469 ;
      RECT 25.08 3.207 25.1 3.469 ;
      RECT 25.02 3.202 25.08 3.466 ;
      RECT 24.985 3.177 25.02 3.462 ;
      RECT 24.975 3.154 24.985 3.46 ;
      RECT 24.945 3.131 24.975 3.46 ;
      RECT 24.935 3.11 24.945 3.46 ;
      RECT 24.91 3.092 24.935 3.458 ;
      RECT 24.895 3.07 24.91 3.455 ;
      RECT 24.88 3.052 24.895 3.453 ;
      RECT 24.86 3.042 24.88 3.451 ;
      RECT 24.845 3.037 24.86 3.45 ;
      RECT 24.83 3.035 24.845 3.449 ;
      RECT 24.8 3.036 24.83 3.447 ;
      RECT 24.78 3.039 24.8 3.445 ;
      RECT 24.723 3.043 24.78 3.445 ;
      RECT 24.637 3.052 24.723 3.445 ;
      RECT 24.551 3.063 24.637 3.445 ;
      RECT 24.465 3.074 24.551 3.445 ;
      RECT 24.445 3.081 24.465 3.453 ;
      RECT 24.435 3.084 24.445 3.46 ;
      RECT 24.37 3.089 24.435 3.478 ;
      RECT 24.34 3.096 24.37 3.503 ;
      RECT 24.33 3.099 24.34 3.51 ;
      RECT 24.285 3.103 24.33 3.515 ;
      RECT 24.255 3.108 24.285 3.52 ;
      RECT 24.254 3.11 24.255 3.52 ;
      RECT 24.168 3.116 24.254 3.52 ;
      RECT 24.082 3.127 24.168 3.52 ;
      RECT 23.996 3.139 24.082 3.52 ;
      RECT 23.91 3.15 23.996 3.52 ;
      RECT 23.895 3.157 23.91 3.515 ;
      RECT 23.89 3.159 23.895 3.509 ;
      RECT 23.87 3.17 23.89 3.504 ;
      RECT 23.86 3.188 23.87 3.498 ;
      RECT 23.855 3.2 23.86 3.298 ;
      RECT 26.15 1.953 26.17 2.04 ;
      RECT 26.145 1.888 26.15 2.072 ;
      RECT 26.135 1.855 26.145 2.077 ;
      RECT 26.13 1.835 26.135 2.083 ;
      RECT 26.1 1.835 26.13 2.1 ;
      RECT 26.051 1.835 26.1 2.136 ;
      RECT 25.965 1.835 26.051 2.194 ;
      RECT 25.936 1.845 25.965 2.243 ;
      RECT 25.85 1.887 25.936 2.296 ;
      RECT 25.83 1.925 25.85 2.343 ;
      RECT 25.805 1.942 25.83 2.363 ;
      RECT 25.795 1.956 25.805 2.383 ;
      RECT 25.79 1.962 25.795 2.393 ;
      RECT 25.785 1.966 25.79 2.4 ;
      RECT 25.735 1.986 25.785 2.405 ;
      RECT 25.67 2.03 25.735 2.405 ;
      RECT 25.645 2.08 25.67 2.405 ;
      RECT 25.635 2.11 25.645 2.405 ;
      RECT 25.63 2.137 25.635 2.405 ;
      RECT 25.625 2.155 25.63 2.405 ;
      RECT 25.615 2.197 25.625 2.405 ;
      RECT 25.965 2.755 26.135 2.93 ;
      RECT 25.905 2.583 25.965 2.918 ;
      RECT 25.895 2.576 25.905 2.901 ;
      RECT 25.85 2.755 26.135 2.881 ;
      RECT 25.831 2.755 26.135 2.859 ;
      RECT 25.745 2.755 26.135 2.824 ;
      RECT 25.725 2.575 25.895 2.78 ;
      RECT 25.725 2.722 26.13 2.78 ;
      RECT 25.725 2.67 26.105 2.78 ;
      RECT 25.725 2.625 26.07 2.78 ;
      RECT 25.725 2.607 26.035 2.78 ;
      RECT 25.725 2.597 26.03 2.78 ;
      RECT 25.895 7.855 26.065 8.305 ;
      RECT 25.95 6.075 26.12 8.025 ;
      RECT 25.895 5.015 26.065 6.245 ;
      RECT 25.375 5.015 25.545 8.305 ;
      RECT 25.375 7.315 25.78 7.645 ;
      RECT 25.375 6.475 25.78 6.805 ;
      RECT 25.445 3.555 25.635 3.78 ;
      RECT 25.435 3.556 25.64 3.775 ;
      RECT 25.435 3.558 25.65 3.755 ;
      RECT 25.435 3.562 25.655 3.74 ;
      RECT 25.435 3.549 25.605 3.775 ;
      RECT 25.435 3.552 25.63 3.775 ;
      RECT 25.445 3.548 25.605 3.78 ;
      RECT 25.531 3.546 25.605 3.78 ;
      RECT 25.155 2.797 25.325 3.035 ;
      RECT 25.155 2.797 25.411 2.949 ;
      RECT 25.155 2.797 25.415 2.859 ;
      RECT 25.205 2.57 25.425 2.838 ;
      RECT 25.2 2.587 25.43 2.811 ;
      RECT 25.165 2.745 25.43 2.811 ;
      RECT 25.185 2.595 25.325 3.035 ;
      RECT 25.175 2.677 25.435 2.794 ;
      RECT 25.17 2.725 25.435 2.794 ;
      RECT 25.175 2.635 25.43 2.811 ;
      RECT 25.2 2.572 25.425 2.838 ;
      RECT 24.765 2.547 24.935 2.745 ;
      RECT 24.765 2.547 24.98 2.72 ;
      RECT 24.835 2.49 25.005 2.678 ;
      RECT 24.81 2.505 25.005 2.678 ;
      RECT 24.425 2.551 24.455 2.745 ;
      RECT 24.42 2.523 24.425 2.745 ;
      RECT 24.39 2.497 24.42 2.747 ;
      RECT 24.365 2.455 24.39 2.75 ;
      RECT 24.355 2.427 24.365 2.752 ;
      RECT 24.32 2.407 24.355 2.754 ;
      RECT 24.255 2.392 24.32 2.76 ;
      RECT 24.205 2.39 24.255 2.766 ;
      RECT 24.182 2.392 24.205 2.771 ;
      RECT 24.096 2.403 24.182 2.777 ;
      RECT 24.01 2.421 24.096 2.787 ;
      RECT 23.995 2.432 24.01 2.793 ;
      RECT 23.925 2.455 23.995 2.799 ;
      RECT 23.87 2.487 23.925 2.807 ;
      RECT 23.83 2.51 23.87 2.813 ;
      RECT 23.816 2.523 23.83 2.816 ;
      RECT 23.73 2.545 23.816 2.822 ;
      RECT 23.715 2.57 23.73 2.828 ;
      RECT 23.675 2.585 23.715 2.832 ;
      RECT 23.625 2.6 23.675 2.837 ;
      RECT 23.6 2.607 23.625 2.841 ;
      RECT 23.54 2.602 23.6 2.845 ;
      RECT 23.525 2.593 23.54 2.849 ;
      RECT 23.455 2.583 23.525 2.845 ;
      RECT 23.43 2.575 23.45 2.835 ;
      RECT 23.371 2.575 23.43 2.813 ;
      RECT 23.285 2.575 23.371 2.77 ;
      RECT 23.45 2.575 23.455 2.84 ;
      RECT 24.145 1.806 24.315 2.14 ;
      RECT 24.115 1.806 24.315 2.135 ;
      RECT 24.055 1.773 24.115 2.123 ;
      RECT 24.055 1.829 24.325 2.118 ;
      RECT 24.03 1.829 24.325 2.112 ;
      RECT 24.025 1.77 24.055 2.109 ;
      RECT 24.01 1.776 24.145 2.107 ;
      RECT 24.005 1.784 24.23 2.095 ;
      RECT 24.005 1.836 24.34 2.048 ;
      RECT 23.99 1.792 24.23 2.043 ;
      RECT 23.99 1.862 24.35 1.984 ;
      RECT 23.96 1.812 24.315 1.945 ;
      RECT 23.96 1.902 24.36 1.941 ;
      RECT 24.01 1.781 24.23 2.107 ;
      RECT 23.35 2.111 23.405 2.375 ;
      RECT 23.35 2.111 23.47 2.374 ;
      RECT 23.35 2.111 23.495 2.373 ;
      RECT 23.35 2.111 23.56 2.372 ;
      RECT 23.495 2.077 23.575 2.371 ;
      RECT 23.31 2.121 23.72 2.37 ;
      RECT 23.35 2.118 23.72 2.37 ;
      RECT 23.31 2.126 23.725 2.363 ;
      RECT 23.295 2.128 23.725 2.362 ;
      RECT 23.295 2.135 23.73 2.358 ;
      RECT 23.275 2.134 23.725 2.354 ;
      RECT 23.275 2.142 23.735 2.353 ;
      RECT 23.27 2.139 23.73 2.349 ;
      RECT 23.27 2.152 23.745 2.348 ;
      RECT 23.255 2.142 23.735 2.347 ;
      RECT 23.22 2.155 23.745 2.34 ;
      RECT 23.405 2.11 23.715 2.37 ;
      RECT 23.405 2.095 23.665 2.37 ;
      RECT 23.47 2.082 23.6 2.37 ;
      RECT 23.015 3.171 23.03 3.564 ;
      RECT 22.98 3.176 23.03 3.563 ;
      RECT 23.015 3.175 23.075 3.562 ;
      RECT 22.96 3.186 23.075 3.561 ;
      RECT 22.975 3.182 23.075 3.561 ;
      RECT 22.94 3.192 23.15 3.558 ;
      RECT 22.94 3.211 23.195 3.556 ;
      RECT 22.94 3.218 23.2 3.553 ;
      RECT 22.925 3.195 23.15 3.55 ;
      RECT 22.905 3.2 23.15 3.543 ;
      RECT 22.9 3.204 23.15 3.539 ;
      RECT 22.9 3.221 23.21 3.538 ;
      RECT 22.88 3.215 23.195 3.534 ;
      RECT 22.88 3.224 23.215 3.528 ;
      RECT 22.875 3.23 23.215 3.3 ;
      RECT 22.94 3.19 23.075 3.558 ;
      RECT 22.815 2.553 23.015 2.865 ;
      RECT 22.89 2.531 23.015 2.865 ;
      RECT 22.83 2.55 23.02 2.85 ;
      RECT 22.8 2.561 23.02 2.848 ;
      RECT 22.815 2.556 23.025 2.814 ;
      RECT 22.8 2.66 23.03 2.781 ;
      RECT 22.83 2.532 23.015 2.865 ;
      RECT 22.89 2.51 22.99 2.865 ;
      RECT 22.915 2.507 22.99 2.865 ;
      RECT 22.915 2.502 22.935 2.865 ;
      RECT 22.32 2.57 22.495 2.745 ;
      RECT 22.315 2.57 22.495 2.743 ;
      RECT 22.29 2.57 22.495 2.738 ;
      RECT 22.235 2.55 22.405 2.728 ;
      RECT 22.235 2.557 22.47 2.728 ;
      RECT 22.32 3.237 22.335 3.42 ;
      RECT 22.31 3.215 22.32 3.42 ;
      RECT 22.295 3.195 22.31 3.42 ;
      RECT 22.285 3.17 22.295 3.42 ;
      RECT 22.255 3.135 22.285 3.42 ;
      RECT 22.22 3.075 22.255 3.42 ;
      RECT 22.215 3.037 22.22 3.42 ;
      RECT 22.165 2.988 22.215 3.42 ;
      RECT 22.155 2.938 22.165 3.408 ;
      RECT 22.14 2.917 22.155 3.368 ;
      RECT 22.12 2.885 22.14 3.318 ;
      RECT 22.095 2.841 22.12 3.258 ;
      RECT 22.09 2.813 22.095 3.213 ;
      RECT 22.085 2.804 22.09 3.199 ;
      RECT 22.08 2.797 22.085 3.186 ;
      RECT 22.075 2.792 22.08 3.175 ;
      RECT 22.07 2.777 22.075 3.165 ;
      RECT 22.065 2.755 22.07 3.152 ;
      RECT 22.055 2.715 22.065 3.127 ;
      RECT 22.03 2.645 22.055 3.083 ;
      RECT 22.025 2.585 22.03 3.048 ;
      RECT 22.01 2.565 22.025 3.015 ;
      RECT 22.005 2.565 22.01 2.99 ;
      RECT 21.975 2.565 22.005 2.945 ;
      RECT 21.93 2.565 21.975 2.885 ;
      RECT 21.855 2.565 21.93 2.833 ;
      RECT 21.85 2.565 21.855 2.798 ;
      RECT 21.845 2.565 21.85 2.788 ;
      RECT 21.84 2.565 21.845 2.768 ;
      RECT 22.105 1.785 22.275 2.255 ;
      RECT 22.05 1.778 22.245 2.239 ;
      RECT 22.05 1.792 22.28 2.238 ;
      RECT 22.035 1.793 22.28 2.219 ;
      RECT 22.03 1.811 22.28 2.205 ;
      RECT 22.035 1.794 22.285 2.203 ;
      RECT 22.02 1.825 22.285 2.188 ;
      RECT 22.035 1.8 22.29 2.173 ;
      RECT 22.015 1.84 22.29 2.17 ;
      RECT 22.03 1.812 22.295 2.155 ;
      RECT 22.03 1.824 22.3 2.135 ;
      RECT 22.015 1.84 22.305 2.118 ;
      RECT 22.015 1.85 22.31 1.973 ;
      RECT 22.01 1.85 22.31 1.93 ;
      RECT 22.01 1.865 22.315 1.908 ;
      RECT 22.105 1.775 22.245 2.255 ;
      RECT 22.105 1.773 22.215 2.255 ;
      RECT 22.191 1.77 22.215 2.255 ;
      RECT 21.85 3.437 21.855 3.483 ;
      RECT 21.84 3.285 21.85 3.507 ;
      RECT 21.835 3.13 21.84 3.532 ;
      RECT 21.82 3.092 21.835 3.543 ;
      RECT 21.815 3.075 21.82 3.55 ;
      RECT 21.805 3.063 21.815 3.557 ;
      RECT 21.8 3.054 21.805 3.559 ;
      RECT 21.795 3.052 21.8 3.563 ;
      RECT 21.75 3.043 21.795 3.578 ;
      RECT 21.745 3.035 21.75 3.592 ;
      RECT 21.74 3.032 21.745 3.596 ;
      RECT 21.725 3.027 21.74 3.604 ;
      RECT 21.67 3.017 21.725 3.615 ;
      RECT 21.635 3.005 21.67 3.616 ;
      RECT 21.626 3 21.635 3.61 ;
      RECT 21.54 3 21.626 3.6 ;
      RECT 21.51 3 21.54 3.578 ;
      RECT 21.5 3 21.505 3.558 ;
      RECT 21.495 3 21.5 3.52 ;
      RECT 21.49 3 21.495 3.478 ;
      RECT 21.485 3 21.49 3.438 ;
      RECT 21.48 3 21.485 3.368 ;
      RECT 21.47 3 21.48 3.29 ;
      RECT 21.465 3 21.47 3.19 ;
      RECT 21.505 3 21.51 3.56 ;
      RECT 21 3.082 21.09 3.56 ;
      RECT 20.985 3.085 21.105 3.558 ;
      RECT 21 3.084 21.105 3.558 ;
      RECT 20.965 3.091 21.13 3.548 ;
      RECT 20.985 3.085 21.13 3.548 ;
      RECT 20.95 3.097 21.13 3.536 ;
      RECT 20.985 3.088 21.18 3.529 ;
      RECT 20.936 3.105 21.18 3.527 ;
      RECT 20.965 3.095 21.19 3.515 ;
      RECT 20.936 3.116 21.22 3.506 ;
      RECT 20.85 3.14 21.22 3.5 ;
      RECT 20.85 3.153 21.26 3.483 ;
      RECT 20.845 3.175 21.26 3.476 ;
      RECT 20.815 3.19 21.26 3.466 ;
      RECT 20.81 3.201 21.26 3.456 ;
      RECT 20.78 3.214 21.26 3.447 ;
      RECT 20.765 3.232 21.26 3.436 ;
      RECT 20.74 3.245 21.26 3.426 ;
      RECT 21 3.081 21.01 3.56 ;
      RECT 21.046 2.505 21.085 2.75 ;
      RECT 20.96 2.505 21.095 2.748 ;
      RECT 20.845 2.53 21.095 2.745 ;
      RECT 20.845 2.53 21.1 2.743 ;
      RECT 20.845 2.53 21.115 2.738 ;
      RECT 20.951 2.505 21.13 2.718 ;
      RECT 20.865 2.513 21.13 2.718 ;
      RECT 20.535 1.865 20.705 2.3 ;
      RECT 20.525 1.899 20.705 2.283 ;
      RECT 20.605 1.835 20.775 2.27 ;
      RECT 20.51 1.91 20.775 2.248 ;
      RECT 20.605 1.845 20.78 2.238 ;
      RECT 20.535 1.897 20.81 2.223 ;
      RECT 20.495 1.923 20.81 2.208 ;
      RECT 20.495 1.965 20.82 2.188 ;
      RECT 20.49 1.99 20.825 2.17 ;
      RECT 20.49 2 20.83 2.155 ;
      RECT 20.485 1.937 20.81 2.153 ;
      RECT 20.485 2.01 20.835 2.138 ;
      RECT 20.48 1.947 20.81 2.135 ;
      RECT 20.475 2.031 20.84 2.118 ;
      RECT 20.475 2.063 20.845 2.098 ;
      RECT 20.47 1.977 20.82 2.09 ;
      RECT 20.475 1.962 20.81 2.118 ;
      RECT 20.49 1.932 20.81 2.17 ;
      RECT 20.335 2.519 20.56 2.775 ;
      RECT 20.335 2.552 20.58 2.765 ;
      RECT 20.3 2.552 20.58 2.763 ;
      RECT 20.3 2.565 20.585 2.753 ;
      RECT 20.3 2.585 20.595 2.745 ;
      RECT 20.3 2.682 20.6 2.738 ;
      RECT 20.28 2.43 20.41 2.728 ;
      RECT 20.235 2.585 20.595 2.67 ;
      RECT 20.225 2.43 20.41 2.615 ;
      RECT 20.225 2.462 20.496 2.615 ;
      RECT 20.19 2.992 20.21 3.17 ;
      RECT 20.155 2.945 20.19 3.17 ;
      RECT 20.14 2.885 20.155 3.17 ;
      RECT 20.115 2.832 20.14 3.17 ;
      RECT 20.1 2.785 20.115 3.17 ;
      RECT 20.08 2.762 20.1 3.17 ;
      RECT 20.055 2.727 20.08 3.17 ;
      RECT 20.045 2.573 20.055 3.17 ;
      RECT 20.015 2.568 20.045 3.161 ;
      RECT 20.01 2.565 20.015 3.151 ;
      RECT 19.995 2.565 20.01 3.125 ;
      RECT 19.99 2.565 19.995 3.088 ;
      RECT 19.965 2.565 19.99 3.04 ;
      RECT 19.945 2.565 19.965 2.965 ;
      RECT 19.935 2.565 19.945 2.925 ;
      RECT 19.93 2.565 19.935 2.9 ;
      RECT 19.925 2.565 19.93 2.883 ;
      RECT 19.92 2.565 19.925 2.865 ;
      RECT 19.915 2.566 19.92 2.855 ;
      RECT 19.905 2.568 19.915 2.823 ;
      RECT 19.895 2.57 19.905 2.79 ;
      RECT 19.885 2.573 19.895 2.763 ;
      RECT 20.21 3 20.435 3.17 ;
      RECT 19.54 1.812 19.71 2.265 ;
      RECT 19.54 1.812 19.8 2.231 ;
      RECT 19.54 1.812 19.83 2.215 ;
      RECT 19.54 1.812 19.86 2.188 ;
      RECT 19.796 1.79 19.875 2.17 ;
      RECT 19.575 1.797 19.88 2.155 ;
      RECT 19.575 1.805 19.89 2.118 ;
      RECT 19.535 1.832 19.89 2.09 ;
      RECT 19.52 1.845 19.89 2.055 ;
      RECT 19.54 1.82 19.91 2.045 ;
      RECT 19.515 1.885 19.91 2.015 ;
      RECT 19.515 1.915 19.915 1.998 ;
      RECT 19.51 1.945 19.915 1.985 ;
      RECT 19.575 1.794 19.875 2.17 ;
      RECT 19.71 1.791 19.796 2.249 ;
      RECT 19.661 1.792 19.875 2.17 ;
      RECT 19.805 3.452 19.85 3.645 ;
      RECT 19.795 3.422 19.805 3.645 ;
      RECT 19.79 3.407 19.795 3.645 ;
      RECT 19.75 3.317 19.79 3.645 ;
      RECT 19.745 3.23 19.75 3.645 ;
      RECT 19.735 3.2 19.745 3.645 ;
      RECT 19.73 3.16 19.735 3.645 ;
      RECT 19.72 3.122 19.73 3.645 ;
      RECT 19.715 3.087 19.72 3.645 ;
      RECT 19.695 3.04 19.715 3.645 ;
      RECT 19.68 2.965 19.695 3.645 ;
      RECT 19.675 2.92 19.68 3.64 ;
      RECT 19.67 2.9 19.675 3.613 ;
      RECT 19.665 2.88 19.67 3.598 ;
      RECT 19.66 2.855 19.665 3.578 ;
      RECT 19.655 2.833 19.66 3.563 ;
      RECT 19.65 2.811 19.655 3.545 ;
      RECT 19.645 2.79 19.65 3.535 ;
      RECT 19.635 2.762 19.645 3.505 ;
      RECT 19.625 2.725 19.635 3.473 ;
      RECT 19.615 2.685 19.625 3.44 ;
      RECT 19.605 2.663 19.615 3.41 ;
      RECT 19.575 2.615 19.605 3.342 ;
      RECT 19.56 2.575 19.575 3.269 ;
      RECT 19.55 2.575 19.56 3.235 ;
      RECT 19.545 2.575 19.55 3.21 ;
      RECT 19.54 2.575 19.545 3.195 ;
      RECT 19.535 2.575 19.54 3.173 ;
      RECT 19.53 2.575 19.535 3.16 ;
      RECT 19.515 2.575 19.53 3.125 ;
      RECT 19.495 2.575 19.515 3.065 ;
      RECT 19.485 2.575 19.495 3.015 ;
      RECT 19.465 2.575 19.485 2.963 ;
      RECT 19.445 2.575 19.465 2.92 ;
      RECT 19.435 2.575 19.445 2.908 ;
      RECT 19.405 2.575 19.435 2.895 ;
      RECT 19.375 2.596 19.405 2.875 ;
      RECT 19.365 2.624 19.375 2.855 ;
      RECT 19.35 2.641 19.365 2.823 ;
      RECT 19.345 2.655 19.35 2.79 ;
      RECT 19.34 2.663 19.345 2.763 ;
      RECT 19.335 2.671 19.34 2.725 ;
      RECT 19.34 3.195 19.345 3.53 ;
      RECT 19.305 3.182 19.34 3.529 ;
      RECT 19.235 3.122 19.305 3.528 ;
      RECT 19.155 3.065 19.235 3.527 ;
      RECT 19.02 3.025 19.155 3.526 ;
      RECT 19.02 3.212 19.355 3.515 ;
      RECT 18.98 3.212 19.355 3.505 ;
      RECT 18.98 3.23 19.36 3.5 ;
      RECT 18.98 3.32 19.365 3.49 ;
      RECT 18.975 3.015 19.14 3.47 ;
      RECT 18.97 3.015 19.14 3.213 ;
      RECT 18.97 3.172 19.335 3.213 ;
      RECT 18.97 3.16 19.33 3.213 ;
      RECT 17.74 1.74 17.91 2.935 ;
      RECT 17.74 1.74 18.205 1.91 ;
      RECT 17.74 6.97 18.205 7.14 ;
      RECT 17.74 5.945 17.91 7.14 ;
      RECT 16.75 1.74 16.92 2.935 ;
      RECT 16.75 1.74 17.215 1.91 ;
      RECT 16.75 6.97 17.215 7.14 ;
      RECT 16.75 5.945 16.92 7.14 ;
      RECT 14.895 2.635 15.065 3.865 ;
      RECT 14.95 0.855 15.12 2.805 ;
      RECT 14.895 0.575 15.065 1.025 ;
      RECT 14.895 7.855 15.065 8.305 ;
      RECT 14.95 6.075 15.12 8.025 ;
      RECT 14.895 5.015 15.065 6.245 ;
      RECT 14.375 0.575 14.545 3.865 ;
      RECT 14.375 2.075 14.78 2.405 ;
      RECT 14.375 1.235 14.78 1.565 ;
      RECT 14.375 5.015 14.545 8.305 ;
      RECT 14.375 7.315 14.78 7.645 ;
      RECT 14.375 6.475 14.78 6.805 ;
      RECT 11.71 1.975 12.44 2.215 ;
      RECT 12.252 1.77 12.44 2.215 ;
      RECT 12.08 1.782 12.455 2.209 ;
      RECT 11.995 1.797 12.475 2.194 ;
      RECT 11.995 1.812 12.48 2.184 ;
      RECT 11.95 1.832 12.495 2.176 ;
      RECT 11.927 1.867 12.51 2.13 ;
      RECT 11.841 1.89 12.515 2.09 ;
      RECT 11.841 1.908 12.525 2.06 ;
      RECT 11.71 1.977 12.53 2.023 ;
      RECT 11.755 1.92 12.525 2.06 ;
      RECT 11.841 1.872 12.51 2.13 ;
      RECT 11.927 1.841 12.495 2.176 ;
      RECT 11.95 1.822 12.48 2.184 ;
      RECT 11.995 1.795 12.455 2.209 ;
      RECT 12.08 1.777 12.44 2.215 ;
      RECT 12.166 1.771 12.44 2.215 ;
      RECT 12.252 1.766 12.385 2.215 ;
      RECT 12.338 1.761 12.385 2.215 ;
      RECT 12.03 2.659 12.2 3.045 ;
      RECT 12.025 2.659 12.2 3.04 ;
      RECT 12 2.659 12.2 3.005 ;
      RECT 12 2.687 12.21 2.995 ;
      RECT 11.98 2.687 12.21 2.955 ;
      RECT 11.975 2.687 12.21 2.928 ;
      RECT 11.975 2.705 12.215 2.92 ;
      RECT 11.92 2.705 12.215 2.855 ;
      RECT 11.92 2.722 12.225 2.838 ;
      RECT 11.91 2.722 12.225 2.778 ;
      RECT 11.91 2.739 12.23 2.775 ;
      RECT 11.905 2.575 12.075 2.753 ;
      RECT 11.905 2.609 12.161 2.753 ;
      RECT 11.9 3.375 11.905 3.388 ;
      RECT 11.895 3.27 11.9 3.393 ;
      RECT 11.87 3.13 11.895 3.408 ;
      RECT 11.835 3.081 11.87 3.44 ;
      RECT 11.83 3.049 11.835 3.46 ;
      RECT 11.825 3.04 11.83 3.46 ;
      RECT 11.745 3.005 11.825 3.46 ;
      RECT 11.682 2.975 11.745 3.46 ;
      RECT 11.596 2.963 11.682 3.46 ;
      RECT 11.51 2.949 11.596 3.46 ;
      RECT 11.43 2.936 11.51 3.446 ;
      RECT 11.395 2.928 11.43 3.426 ;
      RECT 11.385 2.925 11.395 3.417 ;
      RECT 11.355 2.92 11.385 3.404 ;
      RECT 11.305 2.895 11.355 3.38 ;
      RECT 11.291 2.869 11.305 3.362 ;
      RECT 11.205 2.829 11.291 3.338 ;
      RECT 11.16 2.777 11.205 3.307 ;
      RECT 11.15 2.752 11.16 3.294 ;
      RECT 11.145 2.533 11.15 2.555 ;
      RECT 11.14 2.735 11.15 3.29 ;
      RECT 11.14 2.531 11.145 2.645 ;
      RECT 11.13 2.527 11.14 3.286 ;
      RECT 11.086 2.525 11.13 3.274 ;
      RECT 11 2.525 11.086 3.245 ;
      RECT 10.97 2.525 11 3.218 ;
      RECT 10.955 2.525 10.97 3.206 ;
      RECT 10.915 2.537 10.955 3.191 ;
      RECT 10.895 2.556 10.915 3.17 ;
      RECT 10.885 2.566 10.895 3.154 ;
      RECT 10.875 2.572 10.885 3.143 ;
      RECT 10.855 2.582 10.875 3.126 ;
      RECT 10.85 2.591 10.855 3.113 ;
      RECT 10.845 2.595 10.85 3.063 ;
      RECT 10.835 2.601 10.845 2.98 ;
      RECT 10.83 2.605 10.835 2.894 ;
      RECT 10.825 2.625 10.83 2.831 ;
      RECT 10.82 2.648 10.825 2.778 ;
      RECT 10.815 2.666 10.82 2.723 ;
      RECT 11.425 2.485 11.595 2.745 ;
      RECT 11.595 2.45 11.64 2.731 ;
      RECT 11.556 2.452 11.645 2.714 ;
      RECT 11.445 2.469 11.731 2.685 ;
      RECT 11.445 2.484 11.735 2.657 ;
      RECT 11.445 2.465 11.645 2.714 ;
      RECT 11.47 2.453 11.595 2.745 ;
      RECT 11.556 2.451 11.64 2.731 ;
      RECT 10.61 1.84 10.78 2.33 ;
      RECT 10.61 1.84 10.815 2.31 ;
      RECT 10.745 1.76 10.855 2.27 ;
      RECT 10.726 1.764 10.875 2.24 ;
      RECT 10.64 1.772 10.895 2.223 ;
      RECT 10.64 1.778 10.9 2.213 ;
      RECT 10.64 1.787 10.92 2.201 ;
      RECT 10.615 1.812 10.95 2.179 ;
      RECT 10.615 1.832 10.955 2.159 ;
      RECT 10.61 1.845 10.965 2.139 ;
      RECT 10.61 1.912 10.97 2.12 ;
      RECT 10.61 2.045 10.975 2.107 ;
      RECT 10.605 1.85 10.965 1.94 ;
      RECT 10.615 1.807 10.92 2.201 ;
      RECT 10.726 1.762 10.855 2.27 ;
      RECT 10.6 3.515 10.9 3.77 ;
      RECT 10.685 3.481 10.9 3.77 ;
      RECT 10.685 3.484 10.905 3.63 ;
      RECT 10.62 3.505 10.905 3.63 ;
      RECT 10.655 3.495 10.9 3.77 ;
      RECT 10.65 3.5 10.905 3.63 ;
      RECT 10.685 3.479 10.886 3.77 ;
      RECT 10.771 3.47 10.886 3.77 ;
      RECT 10.771 3.464 10.8 3.77 ;
      RECT 10.26 3.105 10.27 3.595 ;
      RECT 9.92 3.04 9.93 3.34 ;
      RECT 10.435 3.212 10.44 3.431 ;
      RECT 10.425 3.192 10.435 3.448 ;
      RECT 10.415 3.172 10.425 3.478 ;
      RECT 10.41 3.162 10.415 3.493 ;
      RECT 10.405 3.158 10.41 3.498 ;
      RECT 10.39 3.15 10.405 3.505 ;
      RECT 10.35 3.13 10.39 3.53 ;
      RECT 10.325 3.112 10.35 3.563 ;
      RECT 10.32 3.11 10.325 3.576 ;
      RECT 10.3 3.107 10.32 3.58 ;
      RECT 10.27 3.105 10.3 3.59 ;
      RECT 10.2 3.107 10.26 3.591 ;
      RECT 10.18 3.107 10.2 3.585 ;
      RECT 10.155 3.105 10.18 3.582 ;
      RECT 10.12 3.1 10.155 3.578 ;
      RECT 10.1 3.094 10.12 3.565 ;
      RECT 10.09 3.091 10.1 3.553 ;
      RECT 10.07 3.088 10.09 3.538 ;
      RECT 10.05 3.084 10.07 3.52 ;
      RECT 10.045 3.081 10.05 3.51 ;
      RECT 10.04 3.08 10.045 3.508 ;
      RECT 10.03 3.077 10.04 3.5 ;
      RECT 10.02 3.071 10.03 3.483 ;
      RECT 10.01 3.065 10.02 3.465 ;
      RECT 10 3.059 10.01 3.453 ;
      RECT 9.99 3.053 10 3.433 ;
      RECT 9.985 3.049 9.99 3.418 ;
      RECT 9.98 3.047 9.985 3.41 ;
      RECT 9.975 3.045 9.98 3.403 ;
      RECT 9.97 3.043 9.975 3.393 ;
      RECT 9.965 3.041 9.97 3.387 ;
      RECT 9.955 3.04 9.965 3.377 ;
      RECT 9.945 3.04 9.955 3.368 ;
      RECT 9.93 3.04 9.945 3.353 ;
      RECT 9.89 3.04 9.92 3.337 ;
      RECT 9.87 3.042 9.89 3.332 ;
      RECT 9.865 3.047 9.87 3.33 ;
      RECT 9.835 3.055 9.865 3.328 ;
      RECT 9.805 3.07 9.835 3.327 ;
      RECT 9.76 3.092 9.805 3.332 ;
      RECT 9.755 3.107 9.76 3.336 ;
      RECT 9.74 3.112 9.755 3.338 ;
      RECT 9.735 3.116 9.74 3.34 ;
      RECT 9.675 3.139 9.735 3.349 ;
      RECT 9.655 3.165 9.675 3.362 ;
      RECT 9.645 3.172 9.655 3.366 ;
      RECT 9.63 3.179 9.645 3.369 ;
      RECT 9.61 3.189 9.63 3.372 ;
      RECT 9.605 3.197 9.61 3.375 ;
      RECT 9.56 3.202 9.605 3.382 ;
      RECT 9.55 3.205 9.56 3.389 ;
      RECT 9.54 3.205 9.55 3.393 ;
      RECT 9.505 3.207 9.54 3.405 ;
      RECT 9.485 3.21 9.505 3.418 ;
      RECT 9.445 3.213 9.485 3.429 ;
      RECT 9.43 3.215 9.445 3.442 ;
      RECT 9.42 3.215 9.43 3.447 ;
      RECT 9.395 3.216 9.42 3.455 ;
      RECT 9.385 3.218 9.395 3.46 ;
      RECT 9.38 3.219 9.385 3.463 ;
      RECT 9.355 3.217 9.38 3.466 ;
      RECT 9.34 3.215 9.355 3.467 ;
      RECT 9.32 3.212 9.34 3.469 ;
      RECT 9.3 3.207 9.32 3.469 ;
      RECT 9.24 3.202 9.3 3.466 ;
      RECT 9.205 3.177 9.24 3.462 ;
      RECT 9.195 3.154 9.205 3.46 ;
      RECT 9.165 3.131 9.195 3.46 ;
      RECT 9.155 3.11 9.165 3.46 ;
      RECT 9.13 3.092 9.155 3.458 ;
      RECT 9.115 3.07 9.13 3.455 ;
      RECT 9.1 3.052 9.115 3.453 ;
      RECT 9.08 3.042 9.1 3.451 ;
      RECT 9.065 3.037 9.08 3.45 ;
      RECT 9.05 3.035 9.065 3.449 ;
      RECT 9.02 3.036 9.05 3.447 ;
      RECT 9 3.039 9.02 3.445 ;
      RECT 8.943 3.043 9 3.445 ;
      RECT 8.857 3.052 8.943 3.445 ;
      RECT 8.771 3.063 8.857 3.445 ;
      RECT 8.685 3.074 8.771 3.445 ;
      RECT 8.665 3.081 8.685 3.453 ;
      RECT 8.655 3.084 8.665 3.46 ;
      RECT 8.59 3.089 8.655 3.478 ;
      RECT 8.56 3.096 8.59 3.503 ;
      RECT 8.55 3.099 8.56 3.51 ;
      RECT 8.505 3.103 8.55 3.515 ;
      RECT 8.475 3.108 8.505 3.52 ;
      RECT 8.474 3.11 8.475 3.52 ;
      RECT 8.388 3.116 8.474 3.52 ;
      RECT 8.302 3.127 8.388 3.52 ;
      RECT 8.216 3.139 8.302 3.52 ;
      RECT 8.13 3.15 8.216 3.52 ;
      RECT 8.115 3.157 8.13 3.515 ;
      RECT 8.11 3.159 8.115 3.509 ;
      RECT 8.09 3.17 8.11 3.504 ;
      RECT 8.08 3.188 8.09 3.498 ;
      RECT 8.075 3.2 8.08 3.298 ;
      RECT 10.37 1.953 10.39 2.04 ;
      RECT 10.365 1.888 10.37 2.072 ;
      RECT 10.355 1.855 10.365 2.077 ;
      RECT 10.35 1.835 10.355 2.083 ;
      RECT 10.32 1.835 10.35 2.1 ;
      RECT 10.271 1.835 10.32 2.136 ;
      RECT 10.185 1.835 10.271 2.194 ;
      RECT 10.156 1.845 10.185 2.243 ;
      RECT 10.07 1.887 10.156 2.296 ;
      RECT 10.05 1.925 10.07 2.343 ;
      RECT 10.025 1.942 10.05 2.363 ;
      RECT 10.015 1.956 10.025 2.383 ;
      RECT 10.01 1.962 10.015 2.393 ;
      RECT 10.005 1.966 10.01 2.4 ;
      RECT 9.955 1.986 10.005 2.405 ;
      RECT 9.89 2.03 9.955 2.405 ;
      RECT 9.865 2.08 9.89 2.405 ;
      RECT 9.855 2.11 9.865 2.405 ;
      RECT 9.85 2.137 9.855 2.405 ;
      RECT 9.845 2.155 9.85 2.405 ;
      RECT 9.835 2.197 9.845 2.405 ;
      RECT 10.185 2.755 10.355 2.93 ;
      RECT 10.125 2.583 10.185 2.918 ;
      RECT 10.115 2.576 10.125 2.901 ;
      RECT 10.07 2.755 10.355 2.881 ;
      RECT 10.051 2.755 10.355 2.859 ;
      RECT 9.965 2.755 10.355 2.824 ;
      RECT 9.945 2.575 10.115 2.78 ;
      RECT 9.945 2.722 10.35 2.78 ;
      RECT 9.945 2.67 10.325 2.78 ;
      RECT 9.945 2.625 10.29 2.78 ;
      RECT 9.945 2.607 10.255 2.78 ;
      RECT 9.945 2.597 10.25 2.78 ;
      RECT 10.115 7.855 10.285 8.305 ;
      RECT 10.17 6.075 10.34 8.025 ;
      RECT 10.115 5.015 10.285 6.245 ;
      RECT 9.595 5.015 9.765 8.305 ;
      RECT 9.595 7.315 10 7.645 ;
      RECT 9.595 6.475 10 6.805 ;
      RECT 9.665 3.555 9.855 3.78 ;
      RECT 9.655 3.556 9.86 3.775 ;
      RECT 9.655 3.558 9.87 3.755 ;
      RECT 9.655 3.562 9.875 3.74 ;
      RECT 9.655 3.549 9.825 3.775 ;
      RECT 9.655 3.552 9.85 3.775 ;
      RECT 9.665 3.548 9.825 3.78 ;
      RECT 9.751 3.546 9.825 3.78 ;
      RECT 9.375 2.797 9.545 3.035 ;
      RECT 9.375 2.797 9.631 2.949 ;
      RECT 9.375 2.797 9.635 2.859 ;
      RECT 9.425 2.57 9.645 2.838 ;
      RECT 9.42 2.587 9.65 2.811 ;
      RECT 9.385 2.745 9.65 2.811 ;
      RECT 9.405 2.595 9.545 3.035 ;
      RECT 9.395 2.677 9.655 2.794 ;
      RECT 9.39 2.725 9.655 2.794 ;
      RECT 9.395 2.635 9.65 2.811 ;
      RECT 9.42 2.572 9.645 2.838 ;
      RECT 8.985 2.547 9.155 2.745 ;
      RECT 8.985 2.547 9.2 2.72 ;
      RECT 9.055 2.49 9.225 2.678 ;
      RECT 9.03 2.505 9.225 2.678 ;
      RECT 8.645 2.551 8.675 2.745 ;
      RECT 8.64 2.523 8.645 2.745 ;
      RECT 8.61 2.497 8.64 2.747 ;
      RECT 8.585 2.455 8.61 2.75 ;
      RECT 8.575 2.427 8.585 2.752 ;
      RECT 8.54 2.407 8.575 2.754 ;
      RECT 8.475 2.392 8.54 2.76 ;
      RECT 8.425 2.39 8.475 2.766 ;
      RECT 8.402 2.392 8.425 2.771 ;
      RECT 8.316 2.403 8.402 2.777 ;
      RECT 8.23 2.421 8.316 2.787 ;
      RECT 8.215 2.432 8.23 2.793 ;
      RECT 8.145 2.455 8.215 2.799 ;
      RECT 8.09 2.487 8.145 2.807 ;
      RECT 8.05 2.51 8.09 2.813 ;
      RECT 8.036 2.523 8.05 2.816 ;
      RECT 7.95 2.545 8.036 2.822 ;
      RECT 7.935 2.57 7.95 2.828 ;
      RECT 7.895 2.585 7.935 2.832 ;
      RECT 7.845 2.6 7.895 2.837 ;
      RECT 7.82 2.607 7.845 2.841 ;
      RECT 7.76 2.602 7.82 2.845 ;
      RECT 7.745 2.593 7.76 2.849 ;
      RECT 7.675 2.583 7.745 2.845 ;
      RECT 7.65 2.575 7.67 2.835 ;
      RECT 7.591 2.575 7.65 2.813 ;
      RECT 7.505 2.575 7.591 2.77 ;
      RECT 7.67 2.575 7.675 2.84 ;
      RECT 8.365 1.806 8.535 2.14 ;
      RECT 8.335 1.806 8.535 2.135 ;
      RECT 8.275 1.773 8.335 2.123 ;
      RECT 8.275 1.829 8.545 2.118 ;
      RECT 8.25 1.829 8.545 2.112 ;
      RECT 8.245 1.77 8.275 2.109 ;
      RECT 8.23 1.776 8.365 2.107 ;
      RECT 8.225 1.784 8.45 2.095 ;
      RECT 8.225 1.836 8.56 2.048 ;
      RECT 8.21 1.792 8.45 2.043 ;
      RECT 8.21 1.862 8.57 1.984 ;
      RECT 8.18 1.812 8.535 1.945 ;
      RECT 8.18 1.902 8.58 1.941 ;
      RECT 8.23 1.781 8.45 2.107 ;
      RECT 7.57 2.111 7.625 2.375 ;
      RECT 7.57 2.111 7.69 2.374 ;
      RECT 7.57 2.111 7.715 2.373 ;
      RECT 7.57 2.111 7.78 2.372 ;
      RECT 7.715 2.077 7.795 2.371 ;
      RECT 7.53 2.121 7.94 2.37 ;
      RECT 7.57 2.118 7.94 2.37 ;
      RECT 7.53 2.126 7.945 2.363 ;
      RECT 7.515 2.128 7.945 2.362 ;
      RECT 7.515 2.135 7.95 2.358 ;
      RECT 7.495 2.134 7.945 2.354 ;
      RECT 7.495 2.142 7.955 2.353 ;
      RECT 7.49 2.139 7.95 2.349 ;
      RECT 7.49 2.152 7.965 2.348 ;
      RECT 7.475 2.142 7.955 2.347 ;
      RECT 7.44 2.155 7.965 2.34 ;
      RECT 7.625 2.11 7.935 2.37 ;
      RECT 7.625 2.095 7.885 2.37 ;
      RECT 7.69 2.082 7.82 2.37 ;
      RECT 7.235 3.171 7.25 3.564 ;
      RECT 7.2 3.176 7.25 3.563 ;
      RECT 7.235 3.175 7.295 3.562 ;
      RECT 7.18 3.186 7.295 3.561 ;
      RECT 7.195 3.182 7.295 3.561 ;
      RECT 7.16 3.192 7.37 3.558 ;
      RECT 7.16 3.211 7.415 3.556 ;
      RECT 7.16 3.218 7.42 3.553 ;
      RECT 7.145 3.195 7.37 3.55 ;
      RECT 7.125 3.2 7.37 3.543 ;
      RECT 7.12 3.204 7.37 3.539 ;
      RECT 7.12 3.221 7.43 3.538 ;
      RECT 7.1 3.215 7.415 3.534 ;
      RECT 7.1 3.224 7.435 3.528 ;
      RECT 7.095 3.23 7.435 3.3 ;
      RECT 7.16 3.19 7.295 3.558 ;
      RECT 7.035 2.553 7.235 2.865 ;
      RECT 7.11 2.531 7.235 2.865 ;
      RECT 7.05 2.55 7.24 2.85 ;
      RECT 7.02 2.561 7.24 2.848 ;
      RECT 7.035 2.556 7.245 2.814 ;
      RECT 7.02 2.66 7.25 2.781 ;
      RECT 7.05 2.532 7.235 2.865 ;
      RECT 7.11 2.51 7.21 2.865 ;
      RECT 7.135 2.507 7.21 2.865 ;
      RECT 7.135 2.502 7.155 2.865 ;
      RECT 6.54 2.57 6.715 2.745 ;
      RECT 6.535 2.57 6.715 2.743 ;
      RECT 6.51 2.57 6.715 2.738 ;
      RECT 6.455 2.55 6.625 2.728 ;
      RECT 6.455 2.557 6.69 2.728 ;
      RECT 6.54 3.237 6.555 3.42 ;
      RECT 6.53 3.215 6.54 3.42 ;
      RECT 6.515 3.195 6.53 3.42 ;
      RECT 6.505 3.17 6.515 3.42 ;
      RECT 6.475 3.135 6.505 3.42 ;
      RECT 6.44 3.075 6.475 3.42 ;
      RECT 6.435 3.037 6.44 3.42 ;
      RECT 6.385 2.988 6.435 3.42 ;
      RECT 6.375 2.938 6.385 3.408 ;
      RECT 6.36 2.917 6.375 3.368 ;
      RECT 6.34 2.885 6.36 3.318 ;
      RECT 6.315 2.841 6.34 3.258 ;
      RECT 6.31 2.813 6.315 3.213 ;
      RECT 6.305 2.804 6.31 3.199 ;
      RECT 6.3 2.797 6.305 3.186 ;
      RECT 6.295 2.792 6.3 3.175 ;
      RECT 6.29 2.777 6.295 3.165 ;
      RECT 6.285 2.755 6.29 3.152 ;
      RECT 6.275 2.715 6.285 3.127 ;
      RECT 6.25 2.645 6.275 3.083 ;
      RECT 6.245 2.585 6.25 3.048 ;
      RECT 6.23 2.565 6.245 3.015 ;
      RECT 6.225 2.565 6.23 2.99 ;
      RECT 6.195 2.565 6.225 2.945 ;
      RECT 6.15 2.565 6.195 2.885 ;
      RECT 6.075 2.565 6.15 2.833 ;
      RECT 6.07 2.565 6.075 2.798 ;
      RECT 6.065 2.565 6.07 2.788 ;
      RECT 6.06 2.565 6.065 2.768 ;
      RECT 6.325 1.785 6.495 2.255 ;
      RECT 6.27 1.778 6.465 2.239 ;
      RECT 6.27 1.792 6.5 2.238 ;
      RECT 6.255 1.793 6.5 2.219 ;
      RECT 6.25 1.811 6.5 2.205 ;
      RECT 6.255 1.794 6.505 2.203 ;
      RECT 6.24 1.825 6.505 2.188 ;
      RECT 6.255 1.8 6.51 2.173 ;
      RECT 6.235 1.84 6.51 2.17 ;
      RECT 6.25 1.812 6.515 2.155 ;
      RECT 6.25 1.824 6.52 2.135 ;
      RECT 6.235 1.84 6.525 2.118 ;
      RECT 6.235 1.85 6.53 1.973 ;
      RECT 6.23 1.85 6.53 1.93 ;
      RECT 6.23 1.865 6.535 1.908 ;
      RECT 6.325 1.775 6.465 2.255 ;
      RECT 6.325 1.773 6.435 2.255 ;
      RECT 6.411 1.77 6.435 2.255 ;
      RECT 6.07 3.437 6.075 3.483 ;
      RECT 6.06 3.285 6.07 3.507 ;
      RECT 6.055 3.13 6.06 3.532 ;
      RECT 6.04 3.092 6.055 3.543 ;
      RECT 6.035 3.075 6.04 3.55 ;
      RECT 6.025 3.063 6.035 3.557 ;
      RECT 6.02 3.054 6.025 3.559 ;
      RECT 6.015 3.052 6.02 3.563 ;
      RECT 5.97 3.043 6.015 3.578 ;
      RECT 5.965 3.035 5.97 3.592 ;
      RECT 5.96 3.032 5.965 3.596 ;
      RECT 5.945 3.027 5.96 3.604 ;
      RECT 5.89 3.017 5.945 3.615 ;
      RECT 5.855 3.005 5.89 3.616 ;
      RECT 5.846 3 5.855 3.61 ;
      RECT 5.76 3 5.846 3.6 ;
      RECT 5.73 3 5.76 3.578 ;
      RECT 5.72 3 5.725 3.558 ;
      RECT 5.715 3 5.72 3.52 ;
      RECT 5.71 3 5.715 3.478 ;
      RECT 5.705 3 5.71 3.438 ;
      RECT 5.7 3 5.705 3.368 ;
      RECT 5.69 3 5.7 3.29 ;
      RECT 5.685 3 5.69 3.19 ;
      RECT 5.725 3 5.73 3.56 ;
      RECT 5.22 3.082 5.31 3.56 ;
      RECT 5.205 3.085 5.325 3.558 ;
      RECT 5.22 3.084 5.325 3.558 ;
      RECT 5.185 3.091 5.35 3.548 ;
      RECT 5.205 3.085 5.35 3.548 ;
      RECT 5.17 3.097 5.35 3.536 ;
      RECT 5.205 3.088 5.4 3.529 ;
      RECT 5.156 3.105 5.4 3.527 ;
      RECT 5.185 3.095 5.41 3.515 ;
      RECT 5.156 3.116 5.44 3.506 ;
      RECT 5.07 3.14 5.44 3.5 ;
      RECT 5.07 3.153 5.48 3.483 ;
      RECT 5.065 3.175 5.48 3.476 ;
      RECT 5.035 3.19 5.48 3.466 ;
      RECT 5.03 3.201 5.48 3.456 ;
      RECT 5 3.214 5.48 3.447 ;
      RECT 4.985 3.232 5.48 3.436 ;
      RECT 4.96 3.245 5.48 3.426 ;
      RECT 5.22 3.081 5.23 3.56 ;
      RECT 5.266 2.505 5.305 2.75 ;
      RECT 5.18 2.505 5.315 2.748 ;
      RECT 5.065 2.53 5.315 2.745 ;
      RECT 5.065 2.53 5.32 2.743 ;
      RECT 5.065 2.53 5.335 2.738 ;
      RECT 5.171 2.505 5.35 2.718 ;
      RECT 5.085 2.513 5.35 2.718 ;
      RECT 4.755 1.865 4.925 2.3 ;
      RECT 4.745 1.899 4.925 2.283 ;
      RECT 4.825 1.835 4.995 2.27 ;
      RECT 4.73 1.91 4.995 2.248 ;
      RECT 4.825 1.845 5 2.238 ;
      RECT 4.755 1.897 5.03 2.223 ;
      RECT 4.715 1.923 5.03 2.208 ;
      RECT 4.715 1.965 5.04 2.188 ;
      RECT 4.71 1.99 5.045 2.17 ;
      RECT 4.71 2 5.05 2.155 ;
      RECT 4.705 1.937 5.03 2.153 ;
      RECT 4.705 2.01 5.055 2.138 ;
      RECT 4.7 1.947 5.03 2.135 ;
      RECT 4.695 2.031 5.06 2.118 ;
      RECT 4.695 2.063 5.065 2.098 ;
      RECT 4.69 1.977 5.04 2.09 ;
      RECT 4.695 1.962 5.03 2.118 ;
      RECT 4.71 1.932 5.03 2.17 ;
      RECT 4.555 2.519 4.78 2.775 ;
      RECT 4.555 2.552 4.8 2.765 ;
      RECT 4.52 2.552 4.8 2.763 ;
      RECT 4.52 2.565 4.805 2.753 ;
      RECT 4.52 2.585 4.815 2.745 ;
      RECT 4.52 2.682 4.82 2.738 ;
      RECT 4.5 2.43 4.63 2.728 ;
      RECT 4.455 2.585 4.815 2.67 ;
      RECT 4.445 2.43 4.63 2.615 ;
      RECT 4.445 2.462 4.716 2.615 ;
      RECT 4.41 2.992 4.43 3.17 ;
      RECT 4.375 2.945 4.41 3.17 ;
      RECT 4.36 2.885 4.375 3.17 ;
      RECT 4.335 2.832 4.36 3.17 ;
      RECT 4.32 2.785 4.335 3.17 ;
      RECT 4.3 2.762 4.32 3.17 ;
      RECT 4.275 2.727 4.3 3.17 ;
      RECT 4.265 2.573 4.275 3.17 ;
      RECT 4.235 2.568 4.265 3.161 ;
      RECT 4.23 2.565 4.235 3.151 ;
      RECT 4.215 2.565 4.23 3.125 ;
      RECT 4.21 2.565 4.215 3.088 ;
      RECT 4.185 2.565 4.21 3.04 ;
      RECT 4.165 2.565 4.185 2.965 ;
      RECT 4.155 2.565 4.165 2.925 ;
      RECT 4.15 2.565 4.155 2.9 ;
      RECT 4.145 2.565 4.15 2.883 ;
      RECT 4.14 2.565 4.145 2.865 ;
      RECT 4.135 2.566 4.14 2.855 ;
      RECT 4.125 2.568 4.135 2.823 ;
      RECT 4.115 2.57 4.125 2.79 ;
      RECT 4.105 2.573 4.115 2.763 ;
      RECT 4.43 3 4.655 3.17 ;
      RECT 3.76 1.812 3.93 2.265 ;
      RECT 3.76 1.812 4.02 2.231 ;
      RECT 3.76 1.812 4.05 2.215 ;
      RECT 3.76 1.812 4.08 2.188 ;
      RECT 4.016 1.79 4.095 2.17 ;
      RECT 3.795 1.797 4.1 2.155 ;
      RECT 3.795 1.805 4.11 2.118 ;
      RECT 3.755 1.832 4.11 2.09 ;
      RECT 3.74 1.845 4.11 2.055 ;
      RECT 3.76 1.82 4.13 2.045 ;
      RECT 3.735 1.885 4.13 2.015 ;
      RECT 3.735 1.915 4.135 1.998 ;
      RECT 3.73 1.945 4.135 1.985 ;
      RECT 3.795 1.794 4.095 2.17 ;
      RECT 3.93 1.791 4.016 2.249 ;
      RECT 3.881 1.792 4.095 2.17 ;
      RECT 4.025 3.452 4.07 3.645 ;
      RECT 4.015 3.422 4.025 3.645 ;
      RECT 4.01 3.407 4.015 3.645 ;
      RECT 3.97 3.317 4.01 3.645 ;
      RECT 3.965 3.23 3.97 3.645 ;
      RECT 3.955 3.2 3.965 3.645 ;
      RECT 3.95 3.16 3.955 3.645 ;
      RECT 3.94 3.122 3.95 3.645 ;
      RECT 3.935 3.087 3.94 3.645 ;
      RECT 3.915 3.04 3.935 3.645 ;
      RECT 3.9 2.965 3.915 3.645 ;
      RECT 3.895 2.92 3.9 3.64 ;
      RECT 3.89 2.9 3.895 3.613 ;
      RECT 3.885 2.88 3.89 3.598 ;
      RECT 3.88 2.855 3.885 3.578 ;
      RECT 3.875 2.833 3.88 3.563 ;
      RECT 3.87 2.811 3.875 3.545 ;
      RECT 3.865 2.79 3.87 3.535 ;
      RECT 3.855 2.762 3.865 3.505 ;
      RECT 3.845 2.725 3.855 3.473 ;
      RECT 3.835 2.685 3.845 3.44 ;
      RECT 3.825 2.663 3.835 3.41 ;
      RECT 3.795 2.615 3.825 3.342 ;
      RECT 3.78 2.575 3.795 3.269 ;
      RECT 3.77 2.575 3.78 3.235 ;
      RECT 3.765 2.575 3.77 3.21 ;
      RECT 3.76 2.575 3.765 3.195 ;
      RECT 3.755 2.575 3.76 3.173 ;
      RECT 3.75 2.575 3.755 3.16 ;
      RECT 3.735 2.575 3.75 3.125 ;
      RECT 3.715 2.575 3.735 3.065 ;
      RECT 3.705 2.575 3.715 3.015 ;
      RECT 3.685 2.575 3.705 2.963 ;
      RECT 3.665 2.575 3.685 2.92 ;
      RECT 3.655 2.575 3.665 2.908 ;
      RECT 3.625 2.575 3.655 2.895 ;
      RECT 3.595 2.596 3.625 2.875 ;
      RECT 3.585 2.624 3.595 2.855 ;
      RECT 3.57 2.641 3.585 2.823 ;
      RECT 3.565 2.655 3.57 2.79 ;
      RECT 3.56 2.663 3.565 2.763 ;
      RECT 3.555 2.671 3.56 2.725 ;
      RECT 3.56 3.195 3.565 3.53 ;
      RECT 3.525 3.182 3.56 3.529 ;
      RECT 3.455 3.122 3.525 3.528 ;
      RECT 3.375 3.065 3.455 3.527 ;
      RECT 3.24 3.025 3.375 3.526 ;
      RECT 3.24 3.212 3.575 3.515 ;
      RECT 3.2 3.212 3.575 3.505 ;
      RECT 3.2 3.23 3.58 3.5 ;
      RECT 3.2 3.32 3.585 3.49 ;
      RECT 3.195 3.015 3.36 3.47 ;
      RECT 3.19 3.015 3.36 3.213 ;
      RECT 3.19 3.172 3.555 3.213 ;
      RECT 3.19 3.16 3.55 3.213 ;
      RECT 1.18 7.855 1.35 8.305 ;
      RECT 1.235 6.075 1.405 8.025 ;
      RECT 1.18 5.015 1.35 6.245 ;
      RECT 0.66 5.015 0.83 8.305 ;
      RECT 0.66 7.315 1.065 7.645 ;
      RECT 0.66 6.475 1.065 6.805 ;
      RECT 81.235 0.575 81.405 1.085 ;
      RECT 81.235 2.395 81.405 3.865 ;
      RECT 81.235 5.015 81.405 6.485 ;
      RECT 81.235 7.795 81.405 8.305 ;
      RECT 80.245 0.575 80.415 1.085 ;
      RECT 80.245 2.395 80.415 3.865 ;
      RECT 80.245 5.015 80.415 6.485 ;
      RECT 80.245 7.795 80.415 8.305 ;
      RECT 78.88 0.575 79.05 3.865 ;
      RECT 78.88 5.015 79.05 8.305 ;
      RECT 78.45 0.575 78.62 1.085 ;
      RECT 78.45 1.655 78.62 3.865 ;
      RECT 78.45 5.015 78.62 7.225 ;
      RECT 78.45 7.795 78.62 8.305 ;
      RECT 77.08 1.66 77.25 2.935 ;
      RECT 77.08 5.945 77.25 7.22 ;
      RECT 76.06 2.85 76.43 3.22 ;
      RECT 74.1 5.015 74.27 8.305 ;
      RECT 73.67 5.015 73.84 7.225 ;
      RECT 73.67 7.795 73.84 8.305 ;
      RECT 72.3 5.945 72.47 7.22 ;
      RECT 65.45 0.575 65.62 1.085 ;
      RECT 65.45 2.395 65.62 3.865 ;
      RECT 65.45 5.015 65.62 6.485 ;
      RECT 65.45 7.795 65.62 8.305 ;
      RECT 64.46 0.575 64.63 1.085 ;
      RECT 64.46 2.395 64.63 3.865 ;
      RECT 64.46 5.015 64.63 6.485 ;
      RECT 64.46 7.795 64.63 8.305 ;
      RECT 63.095 0.575 63.265 3.865 ;
      RECT 63.095 5.015 63.265 8.305 ;
      RECT 62.665 0.575 62.835 1.085 ;
      RECT 62.665 1.655 62.835 3.865 ;
      RECT 62.665 5.015 62.835 7.225 ;
      RECT 62.665 7.795 62.835 8.305 ;
      RECT 61.295 1.66 61.465 2.935 ;
      RECT 61.295 5.945 61.465 7.22 ;
      RECT 60.275 2.85 60.645 3.22 ;
      RECT 58.315 5.015 58.485 8.305 ;
      RECT 57.885 5.015 58.055 7.225 ;
      RECT 57.885 7.795 58.055 8.305 ;
      RECT 56.515 5.945 56.685 7.22 ;
      RECT 49.665 0.575 49.835 1.085 ;
      RECT 49.665 2.395 49.835 3.865 ;
      RECT 49.665 5.015 49.835 6.485 ;
      RECT 49.665 7.795 49.835 8.305 ;
      RECT 48.675 0.575 48.845 1.085 ;
      RECT 48.675 2.395 48.845 3.865 ;
      RECT 48.675 5.015 48.845 6.485 ;
      RECT 48.675 7.795 48.845 8.305 ;
      RECT 47.31 0.575 47.48 3.865 ;
      RECT 47.31 5.015 47.48 8.305 ;
      RECT 46.88 0.575 47.05 1.085 ;
      RECT 46.88 1.655 47.05 3.865 ;
      RECT 46.88 5.015 47.05 7.225 ;
      RECT 46.88 7.795 47.05 8.305 ;
      RECT 45.51 1.66 45.68 2.935 ;
      RECT 45.51 5.945 45.68 7.22 ;
      RECT 44.49 2.85 44.86 3.22 ;
      RECT 42.53 5.015 42.7 8.305 ;
      RECT 42.1 5.015 42.27 7.225 ;
      RECT 42.1 7.795 42.27 8.305 ;
      RECT 40.73 5.945 40.9 7.22 ;
      RECT 33.89 0.575 34.06 1.085 ;
      RECT 33.89 2.395 34.06 3.865 ;
      RECT 33.89 5.015 34.06 6.485 ;
      RECT 33.89 7.795 34.06 8.305 ;
      RECT 32.9 0.575 33.07 1.085 ;
      RECT 32.9 2.395 33.07 3.865 ;
      RECT 32.9 5.015 33.07 6.485 ;
      RECT 32.9 7.795 33.07 8.305 ;
      RECT 31.535 0.575 31.705 3.865 ;
      RECT 31.535 5.015 31.705 8.305 ;
      RECT 31.105 0.575 31.275 1.085 ;
      RECT 31.105 1.655 31.275 3.865 ;
      RECT 31.105 5.015 31.275 7.225 ;
      RECT 31.105 7.795 31.275 8.305 ;
      RECT 29.735 1.66 29.905 2.935 ;
      RECT 29.735 5.945 29.905 7.22 ;
      RECT 28.715 2.85 29.085 3.22 ;
      RECT 26.755 5.015 26.925 8.305 ;
      RECT 26.325 5.015 26.495 7.225 ;
      RECT 26.325 7.795 26.495 8.305 ;
      RECT 24.955 5.945 25.125 7.22 ;
      RECT 18.11 0.575 18.28 1.085 ;
      RECT 18.11 2.395 18.28 3.865 ;
      RECT 18.11 5.015 18.28 6.485 ;
      RECT 18.11 7.795 18.28 8.305 ;
      RECT 17.12 0.575 17.29 1.085 ;
      RECT 17.12 2.395 17.29 3.865 ;
      RECT 17.12 5.015 17.29 6.485 ;
      RECT 17.12 7.795 17.29 8.305 ;
      RECT 15.755 0.575 15.925 3.865 ;
      RECT 15.755 5.015 15.925 8.305 ;
      RECT 15.325 0.575 15.495 1.085 ;
      RECT 15.325 1.655 15.495 3.865 ;
      RECT 15.325 5.015 15.495 7.225 ;
      RECT 15.325 7.795 15.495 8.305 ;
      RECT 13.955 1.66 14.125 2.935 ;
      RECT 13.955 5.945 14.125 7.22 ;
      RECT 12.935 2.85 13.305 3.22 ;
      RECT 10.975 5.015 11.145 8.305 ;
      RECT 10.545 5.015 10.715 7.225 ;
      RECT 10.545 7.795 10.715 8.305 ;
      RECT 9.175 5.945 9.345 7.22 ;
      RECT 1.61 5.015 1.78 7.225 ;
      RECT 1.61 7.795 1.78 8.305 ;
      RECT 0.24 5.945 0.41 7.22 ;
  END
END sky130_osu_ring_oscillator_mpr2aa_8_b0r1

MACRO sky130_osu_ring_oscillator_mpr2aa_8_b0r2
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 2.79 0 ;
  SIZE 81.765 BY 8.88 ;
  SYMMETRY X Y R90 ;
  SITE CoreSite ;
  OBS
    LAYER met3 ;
      RECT 70.77 7.04 71.14 7.41 ;
      RECT 70.81 6.72 71.14 7.41 ;
      RECT 70.81 6.72 73.6 7.025 ;
      RECT 73.295 2.85 73.6 7.025 ;
      RECT 73.26 2.85 73.63 3.22 ;
      RECT 72.52 0.815 72.825 4.02 ;
      RECT 72.27 2.975 72.825 3.705 ;
      RECT 72.48 0.815 72.85 1.185 ;
      RECT 68.63 1.85 68.96 2.745 ;
      RECT 67.75 2.015 68.08 2.745 ;
      RECT 68.625 1.85 68.995 2.65 ;
      RECT 71.79 1.85 72.12 2.58 ;
      RECT 71.75 1.735 71.93 2.385 ;
      RECT 67.76 1.85 72.12 2.22 ;
      RECT 68.25 3.535 68.58 3.865 ;
      RECT 67.045 3.55 68.58 3.85 ;
      RECT 67.045 2.43 67.345 3.85 ;
      RECT 66.79 2.415 67.12 2.745 ;
      RECT 54.985 7.04 55.355 7.41 ;
      RECT 55.025 6.72 55.355 7.41 ;
      RECT 55.025 6.72 57.815 7.025 ;
      RECT 57.51 2.85 57.815 7.025 ;
      RECT 57.475 2.85 57.845 3.22 ;
      RECT 56.735 0.815 57.04 4.02 ;
      RECT 56.485 2.975 57.04 3.705 ;
      RECT 56.695 0.815 57.065 1.185 ;
      RECT 52.845 1.85 53.175 2.745 ;
      RECT 51.965 2.015 52.295 2.745 ;
      RECT 52.84 1.85 53.21 2.65 ;
      RECT 56.005 1.85 56.335 2.58 ;
      RECT 55.965 1.735 56.145 2.385 ;
      RECT 51.975 1.85 56.335 2.22 ;
      RECT 52.465 3.535 52.795 3.865 ;
      RECT 51.26 3.55 52.795 3.85 ;
      RECT 51.26 2.43 51.56 3.85 ;
      RECT 51.005 2.415 51.335 2.745 ;
      RECT 39.2 7.04 39.57 7.41 ;
      RECT 39.24 6.72 39.57 7.41 ;
      RECT 39.24 6.72 42.03 7.025 ;
      RECT 41.725 2.85 42.03 7.025 ;
      RECT 41.69 2.85 42.06 3.22 ;
      RECT 40.95 0.815 41.255 4.02 ;
      RECT 40.7 2.975 41.255 3.705 ;
      RECT 40.91 0.815 41.28 1.185 ;
      RECT 37.06 1.85 37.39 2.745 ;
      RECT 36.18 2.015 36.51 2.745 ;
      RECT 37.055 1.85 37.425 2.65 ;
      RECT 40.22 1.85 40.55 2.58 ;
      RECT 40.18 1.735 40.36 2.385 ;
      RECT 36.19 1.85 40.55 2.22 ;
      RECT 36.68 3.535 37.01 3.865 ;
      RECT 35.475 3.55 37.01 3.85 ;
      RECT 35.475 2.43 35.775 3.85 ;
      RECT 35.22 2.415 35.55 2.745 ;
      RECT 23.425 7.04 23.795 7.41 ;
      RECT 23.465 6.72 23.795 7.41 ;
      RECT 23.465 6.72 26.255 7.025 ;
      RECT 25.95 2.85 26.255 7.025 ;
      RECT 25.915 2.85 26.285 3.22 ;
      RECT 25.175 0.815 25.48 4.02 ;
      RECT 24.925 2.975 25.48 3.705 ;
      RECT 25.135 0.815 25.505 1.185 ;
      RECT 21.285 1.85 21.615 2.745 ;
      RECT 20.405 2.015 20.735 2.745 ;
      RECT 21.28 1.85 21.65 2.65 ;
      RECT 24.445 1.85 24.775 2.58 ;
      RECT 24.405 1.735 24.585 2.385 ;
      RECT 20.415 1.85 24.775 2.22 ;
      RECT 20.905 3.535 21.235 3.865 ;
      RECT 19.7 3.55 21.235 3.85 ;
      RECT 19.7 2.43 20 3.85 ;
      RECT 19.445 2.415 19.775 2.745 ;
      RECT 7.645 7.04 8.015 7.41 ;
      RECT 7.685 6.72 8.015 7.41 ;
      RECT 7.685 6.72 10.475 7.025 ;
      RECT 10.17 2.85 10.475 7.025 ;
      RECT 10.135 2.85 10.505 3.22 ;
      RECT 9.395 0.815 9.7 4.02 ;
      RECT 9.145 2.975 9.7 3.705 ;
      RECT 9.355 0.815 9.725 1.185 ;
      RECT 5.505 1.85 5.835 2.745 ;
      RECT 4.625 2.015 4.955 2.745 ;
      RECT 5.5 1.85 5.87 2.65 ;
      RECT 8.665 1.85 8.995 2.58 ;
      RECT 8.625 1.735 8.805 2.385 ;
      RECT 4.635 1.85 8.995 2.22 ;
      RECT 5.125 3.535 5.455 3.865 ;
      RECT 3.92 3.55 5.455 3.85 ;
      RECT 3.92 2.43 4.22 3.85 ;
      RECT 3.665 2.415 3.995 2.745 ;
      RECT 70.19 2.575 70.52 3.305 ;
      RECT 66.07 2.415 66.4 3.145 ;
      RECT 65.07 1.855 65.4 2.585 ;
      RECT 63.63 2.575 63.96 3.305 ;
      RECT 54.405 2.575 54.735 3.305 ;
      RECT 50.285 2.415 50.615 3.145 ;
      RECT 49.285 1.855 49.615 2.585 ;
      RECT 47.845 2.575 48.175 3.305 ;
      RECT 38.62 2.575 38.95 3.305 ;
      RECT 34.5 2.415 34.83 3.145 ;
      RECT 33.5 1.855 33.83 2.585 ;
      RECT 32.06 2.575 32.39 3.305 ;
      RECT 22.845 2.575 23.175 3.305 ;
      RECT 18.725 2.415 19.055 3.145 ;
      RECT 17.725 1.855 18.055 2.585 ;
      RECT 16.285 2.575 16.615 3.305 ;
      RECT 7.065 2.575 7.395 3.305 ;
      RECT 2.945 2.415 3.275 3.145 ;
      RECT 1.945 1.855 2.275 2.585 ;
      RECT 0.505 2.575 0.835 3.305 ;
    LAYER via2 ;
      RECT 73.345 2.935 73.545 3.135 ;
      RECT 72.565 0.9 72.765 1.1 ;
      RECT 72.335 3.04 72.535 3.24 ;
      RECT 71.855 2.315 72.055 2.515 ;
      RECT 70.855 7.125 71.055 7.325 ;
      RECT 70.255 3.04 70.455 3.24 ;
      RECT 68.695 2.48 68.895 2.68 ;
      RECT 68.315 3.6 68.515 3.8 ;
      RECT 67.815 2.48 68.015 2.68 ;
      RECT 66.855 2.48 67.055 2.68 ;
      RECT 66.135 2.48 66.335 2.68 ;
      RECT 65.135 1.92 65.335 2.12 ;
      RECT 63.695 3.04 63.895 3.24 ;
      RECT 57.56 2.935 57.76 3.135 ;
      RECT 56.78 0.9 56.98 1.1 ;
      RECT 56.55 3.04 56.75 3.24 ;
      RECT 56.07 2.315 56.27 2.515 ;
      RECT 55.07 7.125 55.27 7.325 ;
      RECT 54.47 3.04 54.67 3.24 ;
      RECT 52.91 2.48 53.11 2.68 ;
      RECT 52.53 3.6 52.73 3.8 ;
      RECT 52.03 2.48 52.23 2.68 ;
      RECT 51.07 2.48 51.27 2.68 ;
      RECT 50.35 2.48 50.55 2.68 ;
      RECT 49.35 1.92 49.55 2.12 ;
      RECT 47.91 3.04 48.11 3.24 ;
      RECT 41.775 2.935 41.975 3.135 ;
      RECT 40.995 0.9 41.195 1.1 ;
      RECT 40.765 3.04 40.965 3.24 ;
      RECT 40.285 2.315 40.485 2.515 ;
      RECT 39.285 7.125 39.485 7.325 ;
      RECT 38.685 3.04 38.885 3.24 ;
      RECT 37.125 2.48 37.325 2.68 ;
      RECT 36.745 3.6 36.945 3.8 ;
      RECT 36.245 2.48 36.445 2.68 ;
      RECT 35.285 2.48 35.485 2.68 ;
      RECT 34.565 2.48 34.765 2.68 ;
      RECT 33.565 1.92 33.765 2.12 ;
      RECT 32.125 3.04 32.325 3.24 ;
      RECT 26 2.935 26.2 3.135 ;
      RECT 25.22 0.9 25.42 1.1 ;
      RECT 24.99 3.04 25.19 3.24 ;
      RECT 24.51 2.315 24.71 2.515 ;
      RECT 23.51 7.125 23.71 7.325 ;
      RECT 22.91 3.04 23.11 3.24 ;
      RECT 21.35 2.48 21.55 2.68 ;
      RECT 20.97 3.6 21.17 3.8 ;
      RECT 20.47 2.48 20.67 2.68 ;
      RECT 19.51 2.48 19.71 2.68 ;
      RECT 18.79 2.48 18.99 2.68 ;
      RECT 17.79 1.92 17.99 2.12 ;
      RECT 16.35 3.04 16.55 3.24 ;
      RECT 10.22 2.935 10.42 3.135 ;
      RECT 9.44 0.9 9.64 1.1 ;
      RECT 9.21 3.04 9.41 3.24 ;
      RECT 8.73 2.315 8.93 2.515 ;
      RECT 7.73 7.125 7.93 7.325 ;
      RECT 7.13 3.04 7.33 3.24 ;
      RECT 5.57 2.48 5.77 2.68 ;
      RECT 5.19 3.6 5.39 3.8 ;
      RECT 4.69 2.48 4.89 2.68 ;
      RECT 3.73 2.48 3.93 2.68 ;
      RECT 3.01 2.48 3.21 2.68 ;
      RECT 2.01 1.92 2.21 2.12 ;
      RECT 0.57 3.04 0.77 3.24 ;
    LAYER met2 ;
      RECT -1.565 8.4 78.605 8.57 ;
      RECT 78.435 7.275 78.605 8.57 ;
      RECT -1.565 6.255 -1.395 8.57 ;
      RECT 78.405 7.275 78.755 7.625 ;
      RECT -1.625 6.255 -1.335 6.605 ;
      RECT 75.245 6.22 75.565 6.545 ;
      RECT 75.275 5.695 75.445 6.545 ;
      RECT 75.275 5.695 75.45 6.045 ;
      RECT 75.275 5.695 76.25 5.87 ;
      RECT 76.075 1.965 76.25 5.87 ;
      RECT 76.02 1.965 76.37 2.315 ;
      RECT 76.045 6.655 76.37 6.98 ;
      RECT 74.93 6.745 76.37 6.915 ;
      RECT 74.93 2.395 75.09 6.915 ;
      RECT 75.245 2.365 75.565 2.685 ;
      RECT 74.93 2.395 75.565 2.565 ;
      RECT 74.195 5.855 74.545 6.205 ;
      RECT 74.265 2.705 74.44 6.205 ;
      RECT 74.19 2.705 74.54 3.055 ;
      RECT 63.655 3 63.935 3.28 ;
      RECT 63.625 3 63.935 3.265 ;
      RECT 63.62 3 63.935 3.263 ;
      RECT 63.615 1.33 63.785 3.257 ;
      RECT 63.61 2.967 63.88 3.25 ;
      RECT 63.605 3 63.935 3.243 ;
      RECT 63.575 2.97 63.88 3.23 ;
      RECT 63.575 2.997 63.9 3.23 ;
      RECT 63.575 2.987 63.895 3.23 ;
      RECT 63.575 2.972 63.89 3.23 ;
      RECT 63.615 2.962 63.88 3.257 ;
      RECT 63.615 2.957 63.87 3.257 ;
      RECT 63.615 2.956 63.855 3.257 ;
      RECT 73.585 1.34 73.935 1.69 ;
      RECT 73.58 1.34 73.935 1.595 ;
      RECT 63.615 1.33 73.825 1.5 ;
      RECT 73.26 2.85 73.63 3.22 ;
      RECT 73.345 2.235 73.515 3.22 ;
      RECT 69.365 2.455 69.6 2.715 ;
      RECT 72.51 2.235 72.675 2.495 ;
      RECT 72.415 2.225 72.43 2.495 ;
      RECT 72.51 2.235 73.515 2.415 ;
      RECT 71.015 1.795 71.055 1.935 ;
      RECT 72.43 2.23 72.51 2.495 ;
      RECT 72.375 2.225 72.415 2.461 ;
      RECT 72.361 2.225 72.375 2.461 ;
      RECT 72.275 2.23 72.361 2.463 ;
      RECT 72.23 2.237 72.275 2.465 ;
      RECT 72.2 2.237 72.23 2.467 ;
      RECT 72.175 2.232 72.2 2.469 ;
      RECT 72.145 2.228 72.175 2.478 ;
      RECT 72.135 2.225 72.145 2.49 ;
      RECT 72.13 2.225 72.135 2.498 ;
      RECT 72.125 2.225 72.13 2.503 ;
      RECT 72.115 2.224 72.125 2.513 ;
      RECT 72.11 2.223 72.115 2.523 ;
      RECT 72.095 2.222 72.11 2.528 ;
      RECT 72.067 2.219 72.095 2.555 ;
      RECT 71.981 2.211 72.067 2.555 ;
      RECT 71.895 2.2 71.981 2.555 ;
      RECT 71.855 2.185 71.895 2.555 ;
      RECT 71.815 2.159 71.855 2.555 ;
      RECT 71.81 2.141 71.815 2.367 ;
      RECT 71.8 2.137 71.81 2.357 ;
      RECT 71.785 2.127 71.8 2.344 ;
      RECT 71.765 2.111 71.785 2.329 ;
      RECT 71.75 2.096 71.765 2.314 ;
      RECT 71.74 2.085 71.75 2.304 ;
      RECT 71.715 2.069 71.74 2.293 ;
      RECT 71.71 2.056 71.715 2.283 ;
      RECT 71.705 2.052 71.71 2.278 ;
      RECT 71.65 2.038 71.705 2.256 ;
      RECT 71.611 2.019 71.65 2.22 ;
      RECT 71.525 1.993 71.611 2.173 ;
      RECT 71.521 1.975 71.525 2.139 ;
      RECT 71.435 1.956 71.521 2.117 ;
      RECT 71.43 1.938 71.435 2.095 ;
      RECT 71.425 1.936 71.43 2.093 ;
      RECT 71.415 1.935 71.425 2.088 ;
      RECT 71.355 1.922 71.415 2.074 ;
      RECT 71.31 1.9 71.355 2.053 ;
      RECT 71.25 1.877 71.31 2.032 ;
      RECT 71.186 1.852 71.25 2.007 ;
      RECT 71.1 1.822 71.186 1.976 ;
      RECT 71.085 1.802 71.1 1.955 ;
      RECT 71.055 1.797 71.085 1.946 ;
      RECT 71.002 1.795 71.015 1.935 ;
      RECT 70.916 1.795 71.002 1.937 ;
      RECT 70.83 1.795 70.916 1.939 ;
      RECT 70.81 1.795 70.83 1.943 ;
      RECT 70.765 1.797 70.81 1.954 ;
      RECT 70.725 1.807 70.765 1.97 ;
      RECT 70.721 1.816 70.725 1.978 ;
      RECT 70.635 1.836 70.721 1.994 ;
      RECT 70.625 1.855 70.635 2.012 ;
      RECT 70.62 1.857 70.625 2.015 ;
      RECT 70.61 1.861 70.62 2.018 ;
      RECT 70.59 1.866 70.61 2.028 ;
      RECT 70.56 1.876 70.59 2.048 ;
      RECT 70.555 1.883 70.56 2.062 ;
      RECT 70.545 1.887 70.555 2.069 ;
      RECT 70.53 1.895 70.545 2.08 ;
      RECT 70.52 1.905 70.53 2.091 ;
      RECT 70.51 1.912 70.52 2.099 ;
      RECT 70.485 1.925 70.51 2.114 ;
      RECT 70.421 1.961 70.485 2.153 ;
      RECT 70.335 2.024 70.421 2.217 ;
      RECT 70.3 2.075 70.335 2.27 ;
      RECT 70.295 2.092 70.3 2.287 ;
      RECT 70.28 2.101 70.295 2.294 ;
      RECT 70.26 2.116 70.28 2.308 ;
      RECT 70.255 2.127 70.26 2.318 ;
      RECT 70.235 2.14 70.255 2.328 ;
      RECT 70.23 2.15 70.235 2.338 ;
      RECT 70.215 2.155 70.23 2.347 ;
      RECT 70.205 2.165 70.215 2.358 ;
      RECT 70.175 2.182 70.205 2.375 ;
      RECT 70.165 2.2 70.175 2.393 ;
      RECT 70.15 2.211 70.165 2.404 ;
      RECT 70.11 2.235 70.15 2.42 ;
      RECT 70.075 2.269 70.11 2.437 ;
      RECT 70.045 2.292 70.075 2.449 ;
      RECT 70.03 2.302 70.045 2.458 ;
      RECT 69.99 2.312 70.03 2.469 ;
      RECT 69.97 2.323 69.99 2.481 ;
      RECT 69.965 2.327 69.97 2.488 ;
      RECT 69.95 2.331 69.965 2.493 ;
      RECT 69.94 2.336 69.95 2.498 ;
      RECT 69.935 2.339 69.94 2.501 ;
      RECT 69.905 2.345 69.935 2.508 ;
      RECT 69.87 2.355 69.905 2.522 ;
      RECT 69.81 2.37 69.87 2.542 ;
      RECT 69.755 2.39 69.81 2.566 ;
      RECT 69.726 2.405 69.755 2.584 ;
      RECT 69.64 2.425 69.726 2.609 ;
      RECT 69.635 2.44 69.64 2.629 ;
      RECT 69.625 2.443 69.635 2.63 ;
      RECT 69.6 2.45 69.625 2.715 ;
      RECT 72.295 2.943 72.575 3.28 ;
      RECT 72.295 2.953 72.58 3.238 ;
      RECT 72.295 2.962 72.585 3.135 ;
      RECT 72.295 2.977 72.59 3.003 ;
      RECT 72.295 2.805 72.555 3.28 ;
      RECT 62.595 6.655 62.945 7.005 ;
      RECT 71.42 6.61 71.77 6.96 ;
      RECT 62.595 6.685 71.77 6.885 ;
      RECT 70.015 3.685 70.025 3.875 ;
      RECT 68.275 3.56 68.555 3.84 ;
      RECT 71.32 2.5 71.325 2.985 ;
      RECT 71.215 2.5 71.275 2.76 ;
      RECT 71.54 3.47 71.545 3.545 ;
      RECT 71.53 3.337 71.54 3.58 ;
      RECT 71.52 3.172 71.53 3.601 ;
      RECT 71.515 3.042 71.52 3.617 ;
      RECT 71.505 2.932 71.515 3.633 ;
      RECT 71.5 2.831 71.505 3.65 ;
      RECT 71.495 2.813 71.5 3.66 ;
      RECT 71.49 2.795 71.495 3.67 ;
      RECT 71.48 2.77 71.49 3.685 ;
      RECT 71.475 2.75 71.48 3.7 ;
      RECT 71.455 2.5 71.475 3.725 ;
      RECT 71.44 2.5 71.455 3.758 ;
      RECT 71.41 2.5 71.44 3.78 ;
      RECT 71.39 2.5 71.41 3.794 ;
      RECT 71.37 2.5 71.39 3.31 ;
      RECT 71.385 3.377 71.39 3.799 ;
      RECT 71.38 3.407 71.385 3.801 ;
      RECT 71.375 3.42 71.38 3.804 ;
      RECT 71.37 3.43 71.375 3.808 ;
      RECT 71.365 2.5 71.37 3.228 ;
      RECT 71.365 3.44 71.37 3.81 ;
      RECT 71.36 2.5 71.365 3.205 ;
      RECT 71.35 3.462 71.365 3.81 ;
      RECT 71.345 2.5 71.36 3.15 ;
      RECT 71.34 3.487 71.35 3.81 ;
      RECT 71.34 2.5 71.345 3.095 ;
      RECT 71.33 2.5 71.34 3.043 ;
      RECT 71.335 3.5 71.34 3.811 ;
      RECT 71.33 3.512 71.335 3.812 ;
      RECT 71.325 2.5 71.33 3.003 ;
      RECT 71.325 3.525 71.33 3.813 ;
      RECT 71.31 3.54 71.325 3.814 ;
      RECT 71.315 2.5 71.32 2.965 ;
      RECT 71.31 2.5 71.315 2.93 ;
      RECT 71.305 2.5 71.31 2.905 ;
      RECT 71.3 3.567 71.31 3.816 ;
      RECT 71.295 2.5 71.305 2.863 ;
      RECT 71.295 3.585 71.3 3.817 ;
      RECT 71.29 2.5 71.295 2.823 ;
      RECT 71.29 3.592 71.295 3.818 ;
      RECT 71.285 2.5 71.29 2.795 ;
      RECT 71.28 3.61 71.29 3.819 ;
      RECT 71.275 2.5 71.285 2.775 ;
      RECT 71.27 3.63 71.28 3.821 ;
      RECT 71.26 3.647 71.27 3.822 ;
      RECT 71.225 3.67 71.26 3.825 ;
      RECT 71.17 3.688 71.225 3.831 ;
      RECT 71.084 3.696 71.17 3.84 ;
      RECT 70.998 3.707 71.084 3.851 ;
      RECT 70.912 3.717 70.998 3.862 ;
      RECT 70.826 3.727 70.912 3.874 ;
      RECT 70.74 3.737 70.826 3.885 ;
      RECT 70.72 3.743 70.74 3.891 ;
      RECT 70.64 3.745 70.72 3.895 ;
      RECT 70.635 3.744 70.64 3.9 ;
      RECT 70.627 3.743 70.635 3.9 ;
      RECT 70.541 3.739 70.627 3.898 ;
      RECT 70.455 3.731 70.541 3.895 ;
      RECT 70.369 3.722 70.455 3.891 ;
      RECT 70.283 3.714 70.369 3.888 ;
      RECT 70.197 3.706 70.283 3.884 ;
      RECT 70.111 3.697 70.197 3.881 ;
      RECT 70.025 3.689 70.111 3.877 ;
      RECT 69.97 3.682 70.015 3.875 ;
      RECT 69.885 3.675 69.97 3.873 ;
      RECT 69.811 3.667 69.885 3.869 ;
      RECT 69.725 3.659 69.811 3.866 ;
      RECT 69.722 3.655 69.725 3.864 ;
      RECT 69.636 3.651 69.722 3.863 ;
      RECT 69.55 3.643 69.636 3.86 ;
      RECT 69.465 3.638 69.55 3.857 ;
      RECT 69.379 3.635 69.465 3.854 ;
      RECT 69.293 3.633 69.379 3.851 ;
      RECT 69.207 3.63 69.293 3.848 ;
      RECT 69.121 3.627 69.207 3.845 ;
      RECT 69.035 3.624 69.121 3.842 ;
      RECT 68.959 3.622 69.035 3.839 ;
      RECT 68.873 3.619 68.959 3.836 ;
      RECT 68.787 3.616 68.873 3.834 ;
      RECT 68.701 3.614 68.787 3.831 ;
      RECT 68.615 3.611 68.701 3.828 ;
      RECT 68.555 3.602 68.615 3.826 ;
      RECT 71.065 3.22 71.14 3.48 ;
      RECT 71.045 3.2 71.05 3.48 ;
      RECT 70.365 2.985 70.47 3.28 ;
      RECT 64.81 2.96 64.88 3.22 ;
      RECT 70.705 2.835 70.71 3.206 ;
      RECT 70.695 2.89 70.7 3.206 ;
      RECT 71 2.06 71.06 2.32 ;
      RECT 71.055 3.215 71.065 3.48 ;
      RECT 71.05 3.205 71.055 3.48 ;
      RECT 70.97 3.152 71.045 3.48 ;
      RECT 70.995 2.06 71 2.34 ;
      RECT 70.985 2.06 70.995 2.36 ;
      RECT 70.97 2.06 70.985 2.39 ;
      RECT 70.955 2.06 70.97 2.433 ;
      RECT 70.95 3.095 70.97 3.48 ;
      RECT 70.94 2.06 70.955 2.47 ;
      RECT 70.935 3.075 70.95 3.48 ;
      RECT 70.935 2.06 70.94 2.493 ;
      RECT 70.925 2.06 70.935 2.518 ;
      RECT 70.895 3.042 70.935 3.48 ;
      RECT 70.9 2.06 70.925 2.568 ;
      RECT 70.895 2.06 70.9 2.623 ;
      RECT 70.89 2.06 70.895 2.665 ;
      RECT 70.88 3.005 70.895 3.48 ;
      RECT 70.885 2.06 70.89 2.708 ;
      RECT 70.88 2.06 70.885 2.773 ;
      RECT 70.875 2.06 70.88 2.795 ;
      RECT 70.875 2.993 70.88 3.345 ;
      RECT 70.87 2.06 70.875 2.863 ;
      RECT 70.87 2.985 70.875 3.328 ;
      RECT 70.865 2.06 70.87 2.908 ;
      RECT 70.86 2.967 70.87 3.305 ;
      RECT 70.86 2.06 70.865 2.945 ;
      RECT 70.85 2.06 70.86 3.285 ;
      RECT 70.845 2.06 70.85 3.268 ;
      RECT 70.84 2.06 70.845 3.253 ;
      RECT 70.835 2.06 70.84 3.238 ;
      RECT 70.815 2.06 70.835 3.228 ;
      RECT 70.81 2.06 70.815 3.218 ;
      RECT 70.8 2.06 70.81 3.214 ;
      RECT 70.795 2.337 70.8 3.213 ;
      RECT 70.79 2.36 70.795 3.212 ;
      RECT 70.785 2.39 70.79 3.211 ;
      RECT 70.78 2.417 70.785 3.21 ;
      RECT 70.775 2.445 70.78 3.21 ;
      RECT 70.77 2.472 70.775 3.21 ;
      RECT 70.765 2.492 70.77 3.21 ;
      RECT 70.76 2.52 70.765 3.21 ;
      RECT 70.75 2.562 70.76 3.21 ;
      RECT 70.74 2.607 70.75 3.209 ;
      RECT 70.735 2.66 70.74 3.208 ;
      RECT 70.73 2.692 70.735 3.207 ;
      RECT 70.725 2.712 70.73 3.206 ;
      RECT 70.72 2.75 70.725 3.206 ;
      RECT 70.715 2.772 70.72 3.206 ;
      RECT 70.71 2.797 70.715 3.206 ;
      RECT 70.7 2.862 70.705 3.206 ;
      RECT 70.685 2.922 70.695 3.206 ;
      RECT 70.67 2.932 70.685 3.206 ;
      RECT 70.65 2.942 70.67 3.206 ;
      RECT 70.62 2.947 70.65 3.203 ;
      RECT 70.56 2.957 70.62 3.2 ;
      RECT 70.54 2.966 70.56 3.205 ;
      RECT 70.515 2.972 70.54 3.218 ;
      RECT 70.495 2.977 70.515 3.233 ;
      RECT 70.47 2.982 70.495 3.28 ;
      RECT 70.341 2.984 70.365 3.28 ;
      RECT 70.255 2.979 70.341 3.28 ;
      RECT 70.215 2.976 70.255 3.28 ;
      RECT 70.165 2.978 70.215 3.26 ;
      RECT 70.135 2.982 70.165 3.26 ;
      RECT 70.056 2.992 70.135 3.26 ;
      RECT 69.97 3.007 70.056 3.261 ;
      RECT 69.92 3.017 69.97 3.262 ;
      RECT 69.912 3.02 69.92 3.262 ;
      RECT 69.826 3.022 69.912 3.263 ;
      RECT 69.74 3.026 69.826 3.263 ;
      RECT 69.654 3.03 69.74 3.264 ;
      RECT 69.568 3.033 69.654 3.265 ;
      RECT 69.482 3.037 69.568 3.265 ;
      RECT 69.396 3.041 69.482 3.266 ;
      RECT 69.31 3.044 69.396 3.267 ;
      RECT 69.224 3.048 69.31 3.267 ;
      RECT 69.138 3.052 69.224 3.268 ;
      RECT 69.052 3.056 69.138 3.269 ;
      RECT 68.966 3.059 69.052 3.269 ;
      RECT 68.88 3.063 68.966 3.27 ;
      RECT 68.85 3.065 68.88 3.27 ;
      RECT 68.764 3.068 68.85 3.271 ;
      RECT 68.678 3.072 68.764 3.272 ;
      RECT 68.592 3.076 68.678 3.273 ;
      RECT 68.506 3.079 68.592 3.273 ;
      RECT 68.42 3.083 68.506 3.274 ;
      RECT 68.385 3.088 68.42 3.275 ;
      RECT 68.33 3.098 68.385 3.282 ;
      RECT 68.305 3.11 68.33 3.292 ;
      RECT 68.27 3.123 68.305 3.3 ;
      RECT 68.23 3.14 68.27 3.323 ;
      RECT 68.21 3.153 68.23 3.35 ;
      RECT 68.18 3.165 68.21 3.378 ;
      RECT 68.175 3.173 68.18 3.398 ;
      RECT 68.17 3.176 68.175 3.408 ;
      RECT 68.12 3.188 68.17 3.442 ;
      RECT 68.11 3.203 68.12 3.475 ;
      RECT 68.1 3.209 68.11 3.488 ;
      RECT 68.09 3.216 68.1 3.5 ;
      RECT 68.065 3.229 68.09 3.518 ;
      RECT 68.05 3.244 68.065 3.54 ;
      RECT 68.04 3.252 68.05 3.556 ;
      RECT 68.025 3.261 68.04 3.571 ;
      RECT 68.015 3.271 68.025 3.585 ;
      RECT 67.996 3.284 68.015 3.602 ;
      RECT 67.91 3.329 67.996 3.667 ;
      RECT 67.895 3.374 67.91 3.725 ;
      RECT 67.89 3.383 67.895 3.738 ;
      RECT 67.88 3.39 67.89 3.743 ;
      RECT 67.875 3.395 67.88 3.747 ;
      RECT 67.855 3.405 67.875 3.754 ;
      RECT 67.83 3.425 67.855 3.768 ;
      RECT 67.795 3.45 67.83 3.788 ;
      RECT 67.78 3.473 67.795 3.803 ;
      RECT 67.77 3.483 67.78 3.808 ;
      RECT 67.76 3.491 67.77 3.815 ;
      RECT 67.75 3.5 67.76 3.821 ;
      RECT 67.73 3.512 67.75 3.823 ;
      RECT 67.72 3.525 67.73 3.825 ;
      RECT 67.695 3.54 67.72 3.828 ;
      RECT 67.675 3.557 67.695 3.832 ;
      RECT 67.635 3.585 67.675 3.838 ;
      RECT 67.57 3.632 67.635 3.847 ;
      RECT 67.555 3.665 67.57 3.855 ;
      RECT 67.55 3.672 67.555 3.857 ;
      RECT 67.5 3.697 67.55 3.862 ;
      RECT 67.485 3.721 67.5 3.869 ;
      RECT 67.435 3.726 67.485 3.87 ;
      RECT 67.349 3.73 67.435 3.87 ;
      RECT 67.263 3.73 67.349 3.87 ;
      RECT 67.177 3.73 67.263 3.871 ;
      RECT 67.091 3.73 67.177 3.871 ;
      RECT 67.005 3.73 67.091 3.871 ;
      RECT 66.939 3.73 67.005 3.871 ;
      RECT 66.853 3.73 66.939 3.872 ;
      RECT 66.767 3.73 66.853 3.872 ;
      RECT 66.681 3.731 66.767 3.873 ;
      RECT 66.595 3.731 66.681 3.873 ;
      RECT 66.509 3.731 66.595 3.873 ;
      RECT 66.423 3.731 66.509 3.874 ;
      RECT 66.337 3.731 66.423 3.874 ;
      RECT 66.251 3.732 66.337 3.875 ;
      RECT 66.165 3.732 66.251 3.875 ;
      RECT 66.145 3.732 66.165 3.875 ;
      RECT 66.059 3.732 66.145 3.875 ;
      RECT 65.973 3.732 66.059 3.875 ;
      RECT 65.887 3.733 65.973 3.875 ;
      RECT 65.801 3.733 65.887 3.875 ;
      RECT 65.715 3.733 65.801 3.875 ;
      RECT 65.629 3.734 65.715 3.875 ;
      RECT 65.543 3.734 65.629 3.875 ;
      RECT 65.457 3.734 65.543 3.875 ;
      RECT 65.371 3.734 65.457 3.875 ;
      RECT 65.285 3.735 65.371 3.875 ;
      RECT 65.235 3.732 65.285 3.875 ;
      RECT 65.225 3.73 65.235 3.874 ;
      RECT 65.221 3.73 65.225 3.873 ;
      RECT 65.135 3.725 65.221 3.868 ;
      RECT 65.113 3.718 65.135 3.862 ;
      RECT 65.027 3.709 65.113 3.856 ;
      RECT 64.941 3.696 65.027 3.847 ;
      RECT 64.855 3.682 64.941 3.837 ;
      RECT 64.81 3.672 64.855 3.83 ;
      RECT 64.79 2.96 64.81 3.238 ;
      RECT 64.79 3.665 64.81 3.826 ;
      RECT 64.76 2.96 64.79 3.26 ;
      RECT 64.75 3.632 64.79 3.823 ;
      RECT 64.745 2.96 64.76 3.28 ;
      RECT 64.745 3.597 64.75 3.821 ;
      RECT 64.74 2.96 64.745 3.405 ;
      RECT 64.74 3.557 64.745 3.821 ;
      RECT 64.73 2.96 64.74 3.821 ;
      RECT 64.655 2.96 64.73 3.815 ;
      RECT 64.625 2.96 64.655 3.805 ;
      RECT 64.62 2.96 64.625 3.797 ;
      RECT 64.615 3.002 64.62 3.79 ;
      RECT 64.605 3.071 64.615 3.781 ;
      RECT 64.6 3.141 64.605 3.733 ;
      RECT 64.595 3.205 64.6 3.63 ;
      RECT 64.59 3.24 64.595 3.585 ;
      RECT 64.588 3.277 64.59 3.477 ;
      RECT 64.585 3.285 64.588 3.47 ;
      RECT 64.58 3.35 64.585 3.413 ;
      RECT 68.655 2.44 68.935 2.72 ;
      RECT 68.645 2.44 68.935 2.583 ;
      RECT 68.6 2.305 68.86 2.565 ;
      RECT 68.6 2.42 68.915 2.565 ;
      RECT 68.6 2.39 68.91 2.565 ;
      RECT 68.6 2.377 68.9 2.565 ;
      RECT 68.6 2.367 68.895 2.565 ;
      RECT 64.575 2.35 64.835 2.61 ;
      RECT 68.345 1.9 68.605 2.16 ;
      RECT 68.335 1.925 68.605 2.12 ;
      RECT 68.33 1.925 68.335 2.119 ;
      RECT 68.26 1.92 68.33 2.111 ;
      RECT 68.175 1.907 68.26 2.094 ;
      RECT 68.171 1.899 68.175 2.084 ;
      RECT 68.085 1.892 68.171 2.074 ;
      RECT 68.076 1.884 68.085 2.064 ;
      RECT 67.99 1.877 68.076 2.052 ;
      RECT 67.97 1.868 67.99 2.038 ;
      RECT 67.915 1.863 67.97 2.03 ;
      RECT 67.905 1.857 67.915 2.024 ;
      RECT 67.885 1.855 67.905 2.02 ;
      RECT 67.877 1.854 67.885 2.016 ;
      RECT 67.791 1.846 67.877 2.005 ;
      RECT 67.705 1.832 67.791 1.985 ;
      RECT 67.645 1.82 67.705 1.97 ;
      RECT 67.635 1.815 67.645 1.965 ;
      RECT 67.585 1.815 67.635 1.967 ;
      RECT 67.538 1.817 67.585 1.971 ;
      RECT 67.452 1.824 67.538 1.976 ;
      RECT 67.366 1.832 67.452 1.982 ;
      RECT 67.28 1.841 67.366 1.988 ;
      RECT 67.221 1.847 67.28 1.993 ;
      RECT 67.135 1.852 67.221 1.999 ;
      RECT 67.06 1.857 67.135 2.005 ;
      RECT 67.021 1.859 67.06 2.01 ;
      RECT 66.935 1.856 67.021 2.015 ;
      RECT 66.85 1.854 66.935 2.022 ;
      RECT 66.818 1.853 66.85 2.025 ;
      RECT 66.732 1.852 66.818 2.026 ;
      RECT 66.646 1.851 66.732 2.027 ;
      RECT 66.56 1.85 66.646 2.027 ;
      RECT 66.474 1.849 66.56 2.028 ;
      RECT 66.388 1.848 66.474 2.029 ;
      RECT 66.302 1.847 66.388 2.03 ;
      RECT 66.216 1.846 66.302 2.03 ;
      RECT 66.13 1.845 66.216 2.031 ;
      RECT 66.08 1.845 66.13 2.032 ;
      RECT 66.066 1.846 66.08 2.032 ;
      RECT 65.98 1.853 66.066 2.033 ;
      RECT 65.906 1.864 65.98 2.034 ;
      RECT 65.82 1.873 65.906 2.035 ;
      RECT 65.785 1.88 65.82 2.05 ;
      RECT 65.76 1.883 65.785 2.08 ;
      RECT 65.735 1.892 65.76 2.109 ;
      RECT 65.725 1.903 65.735 2.129 ;
      RECT 65.715 1.911 65.725 2.143 ;
      RECT 65.71 1.917 65.715 2.153 ;
      RECT 65.685 1.934 65.71 2.17 ;
      RECT 65.67 1.956 65.685 2.198 ;
      RECT 65.64 1.982 65.67 2.228 ;
      RECT 65.62 2.011 65.64 2.258 ;
      RECT 65.615 2.026 65.62 2.275 ;
      RECT 65.595 2.041 65.615 2.29 ;
      RECT 65.585 2.059 65.595 2.308 ;
      RECT 65.575 2.07 65.585 2.323 ;
      RECT 65.525 2.102 65.575 2.349 ;
      RECT 65.52 2.132 65.525 2.369 ;
      RECT 65.51 2.145 65.52 2.375 ;
      RECT 65.501 2.155 65.51 2.383 ;
      RECT 65.49 2.166 65.501 2.391 ;
      RECT 65.485 2.176 65.49 2.397 ;
      RECT 65.47 2.197 65.485 2.404 ;
      RECT 65.455 2.227 65.47 2.412 ;
      RECT 65.42 2.257 65.455 2.418 ;
      RECT 65.395 2.275 65.42 2.425 ;
      RECT 65.345 2.283 65.395 2.434 ;
      RECT 65.32 2.288 65.345 2.443 ;
      RECT 65.265 2.294 65.32 2.453 ;
      RECT 65.26 2.299 65.265 2.461 ;
      RECT 65.246 2.302 65.26 2.463 ;
      RECT 65.16 2.314 65.246 2.475 ;
      RECT 65.15 2.326 65.16 2.488 ;
      RECT 65.065 2.339 65.15 2.5 ;
      RECT 65.021 2.356 65.065 2.514 ;
      RECT 64.935 2.373 65.021 2.53 ;
      RECT 64.905 2.387 64.935 2.544 ;
      RECT 64.895 2.392 64.905 2.549 ;
      RECT 64.835 2.395 64.895 2.558 ;
      RECT 67.725 2.665 67.985 2.925 ;
      RECT 67.725 2.665 68.005 2.778 ;
      RECT 67.725 2.665 68.03 2.745 ;
      RECT 67.725 2.665 68.035 2.725 ;
      RECT 67.775 2.44 68.055 2.72 ;
      RECT 67.33 3.175 67.59 3.435 ;
      RECT 67.32 3.032 67.515 3.373 ;
      RECT 67.315 3.14 67.53 3.365 ;
      RECT 67.31 3.19 67.59 3.355 ;
      RECT 67.3 3.267 67.59 3.34 ;
      RECT 67.32 3.115 67.53 3.373 ;
      RECT 67.33 2.99 67.515 3.435 ;
      RECT 67.33 2.885 67.495 3.435 ;
      RECT 67.34 2.872 67.495 3.435 ;
      RECT 67.34 2.83 67.485 3.435 ;
      RECT 67.345 2.755 67.485 3.435 ;
      RECT 67.375 2.405 67.485 3.435 ;
      RECT 67.38 2.135 67.505 2.758 ;
      RECT 67.35 2.71 67.505 2.758 ;
      RECT 67.365 2.512 67.485 3.435 ;
      RECT 67.355 2.622 67.505 2.758 ;
      RECT 67.38 2.135 67.52 2.615 ;
      RECT 67.38 2.135 67.54 2.49 ;
      RECT 67.345 2.135 67.605 2.395 ;
      RECT 66.815 2.44 67.095 2.72 ;
      RECT 66.8 2.44 67.095 2.7 ;
      RECT 64.855 3.305 65.115 3.565 ;
      RECT 66.64 3.16 66.9 3.42 ;
      RECT 66.62 3.18 66.9 3.395 ;
      RECT 66.577 3.18 66.62 3.394 ;
      RECT 66.491 3.181 66.577 3.391 ;
      RECT 66.405 3.182 66.491 3.387 ;
      RECT 66.33 3.184 66.405 3.384 ;
      RECT 66.307 3.185 66.33 3.382 ;
      RECT 66.221 3.186 66.307 3.38 ;
      RECT 66.135 3.187 66.221 3.377 ;
      RECT 66.111 3.188 66.135 3.375 ;
      RECT 66.025 3.19 66.111 3.372 ;
      RECT 65.94 3.192 66.025 3.373 ;
      RECT 65.883 3.193 65.94 3.379 ;
      RECT 65.797 3.195 65.883 3.389 ;
      RECT 65.711 3.198 65.797 3.402 ;
      RECT 65.625 3.2 65.711 3.414 ;
      RECT 65.611 3.201 65.625 3.421 ;
      RECT 65.525 3.202 65.611 3.429 ;
      RECT 65.485 3.204 65.525 3.438 ;
      RECT 65.476 3.205 65.485 3.441 ;
      RECT 65.39 3.213 65.476 3.447 ;
      RECT 65.37 3.222 65.39 3.455 ;
      RECT 65.285 3.237 65.37 3.463 ;
      RECT 65.225 3.26 65.285 3.474 ;
      RECT 65.215 3.272 65.225 3.479 ;
      RECT 65.175 3.282 65.215 3.483 ;
      RECT 65.12 3.299 65.175 3.491 ;
      RECT 65.115 3.309 65.12 3.495 ;
      RECT 66.181 2.44 66.24 2.837 ;
      RECT 66.095 2.44 66.3 2.828 ;
      RECT 66.09 2.47 66.3 2.823 ;
      RECT 66.056 2.47 66.3 2.821 ;
      RECT 65.97 2.47 66.3 2.815 ;
      RECT 65.925 2.47 66.32 2.793 ;
      RECT 65.925 2.47 66.34 2.748 ;
      RECT 65.885 2.47 66.34 2.738 ;
      RECT 66.095 2.44 66.375 2.72 ;
      RECT 65.83 2.44 66.09 2.7 ;
      RECT 65.015 1.92 65.275 2.18 ;
      RECT 65.095 1.88 65.375 2.16 ;
      RECT 59.46 6.22 59.78 6.545 ;
      RECT 59.49 5.695 59.66 6.545 ;
      RECT 59.49 5.695 59.665 6.045 ;
      RECT 59.49 5.695 60.465 5.87 ;
      RECT 60.29 1.965 60.465 5.87 ;
      RECT 60.235 1.965 60.585 2.315 ;
      RECT 60.26 6.655 60.585 6.98 ;
      RECT 59.145 6.745 60.585 6.915 ;
      RECT 59.145 2.395 59.305 6.915 ;
      RECT 59.46 2.365 59.78 2.685 ;
      RECT 59.145 2.395 59.78 2.565 ;
      RECT 58.41 5.855 58.76 6.205 ;
      RECT 58.48 2.705 58.655 6.205 ;
      RECT 58.405 2.705 58.755 3.055 ;
      RECT 47.87 3 48.15 3.28 ;
      RECT 47.84 3 48.15 3.265 ;
      RECT 47.835 3 48.15 3.263 ;
      RECT 47.83 1.33 48 3.257 ;
      RECT 47.825 2.967 48.095 3.25 ;
      RECT 47.82 3 48.15 3.243 ;
      RECT 47.79 2.97 48.095 3.23 ;
      RECT 47.79 2.997 48.115 3.23 ;
      RECT 47.79 2.987 48.11 3.23 ;
      RECT 47.79 2.972 48.105 3.23 ;
      RECT 47.83 2.962 48.095 3.257 ;
      RECT 47.83 2.957 48.085 3.257 ;
      RECT 47.83 2.956 48.07 3.257 ;
      RECT 57.8 1.34 58.15 1.69 ;
      RECT 57.795 1.34 58.15 1.595 ;
      RECT 47.83 1.33 58.04 1.5 ;
      RECT 57.475 2.85 57.845 3.22 ;
      RECT 57.56 2.235 57.73 3.22 ;
      RECT 53.58 2.455 53.815 2.715 ;
      RECT 56.725 2.235 56.89 2.495 ;
      RECT 56.63 2.225 56.645 2.495 ;
      RECT 56.725 2.235 57.73 2.415 ;
      RECT 55.23 1.795 55.27 1.935 ;
      RECT 56.645 2.23 56.725 2.495 ;
      RECT 56.59 2.225 56.63 2.461 ;
      RECT 56.576 2.225 56.59 2.461 ;
      RECT 56.49 2.23 56.576 2.463 ;
      RECT 56.445 2.237 56.49 2.465 ;
      RECT 56.415 2.237 56.445 2.467 ;
      RECT 56.39 2.232 56.415 2.469 ;
      RECT 56.36 2.228 56.39 2.478 ;
      RECT 56.35 2.225 56.36 2.49 ;
      RECT 56.345 2.225 56.35 2.498 ;
      RECT 56.34 2.225 56.345 2.503 ;
      RECT 56.33 2.224 56.34 2.513 ;
      RECT 56.325 2.223 56.33 2.523 ;
      RECT 56.31 2.222 56.325 2.528 ;
      RECT 56.282 2.219 56.31 2.555 ;
      RECT 56.196 2.211 56.282 2.555 ;
      RECT 56.11 2.2 56.196 2.555 ;
      RECT 56.07 2.185 56.11 2.555 ;
      RECT 56.03 2.159 56.07 2.555 ;
      RECT 56.025 2.141 56.03 2.367 ;
      RECT 56.015 2.137 56.025 2.357 ;
      RECT 56 2.127 56.015 2.344 ;
      RECT 55.98 2.111 56 2.329 ;
      RECT 55.965 2.096 55.98 2.314 ;
      RECT 55.955 2.085 55.965 2.304 ;
      RECT 55.93 2.069 55.955 2.293 ;
      RECT 55.925 2.056 55.93 2.283 ;
      RECT 55.92 2.052 55.925 2.278 ;
      RECT 55.865 2.038 55.92 2.256 ;
      RECT 55.826 2.019 55.865 2.22 ;
      RECT 55.74 1.993 55.826 2.173 ;
      RECT 55.736 1.975 55.74 2.139 ;
      RECT 55.65 1.956 55.736 2.117 ;
      RECT 55.645 1.938 55.65 2.095 ;
      RECT 55.64 1.936 55.645 2.093 ;
      RECT 55.63 1.935 55.64 2.088 ;
      RECT 55.57 1.922 55.63 2.074 ;
      RECT 55.525 1.9 55.57 2.053 ;
      RECT 55.465 1.877 55.525 2.032 ;
      RECT 55.401 1.852 55.465 2.007 ;
      RECT 55.315 1.822 55.401 1.976 ;
      RECT 55.3 1.802 55.315 1.955 ;
      RECT 55.27 1.797 55.3 1.946 ;
      RECT 55.217 1.795 55.23 1.935 ;
      RECT 55.131 1.795 55.217 1.937 ;
      RECT 55.045 1.795 55.131 1.939 ;
      RECT 55.025 1.795 55.045 1.943 ;
      RECT 54.98 1.797 55.025 1.954 ;
      RECT 54.94 1.807 54.98 1.97 ;
      RECT 54.936 1.816 54.94 1.978 ;
      RECT 54.85 1.836 54.936 1.994 ;
      RECT 54.84 1.855 54.85 2.012 ;
      RECT 54.835 1.857 54.84 2.015 ;
      RECT 54.825 1.861 54.835 2.018 ;
      RECT 54.805 1.866 54.825 2.028 ;
      RECT 54.775 1.876 54.805 2.048 ;
      RECT 54.77 1.883 54.775 2.062 ;
      RECT 54.76 1.887 54.77 2.069 ;
      RECT 54.745 1.895 54.76 2.08 ;
      RECT 54.735 1.905 54.745 2.091 ;
      RECT 54.725 1.912 54.735 2.099 ;
      RECT 54.7 1.925 54.725 2.114 ;
      RECT 54.636 1.961 54.7 2.153 ;
      RECT 54.55 2.024 54.636 2.217 ;
      RECT 54.515 2.075 54.55 2.27 ;
      RECT 54.51 2.092 54.515 2.287 ;
      RECT 54.495 2.101 54.51 2.294 ;
      RECT 54.475 2.116 54.495 2.308 ;
      RECT 54.47 2.127 54.475 2.318 ;
      RECT 54.45 2.14 54.47 2.328 ;
      RECT 54.445 2.15 54.45 2.338 ;
      RECT 54.43 2.155 54.445 2.347 ;
      RECT 54.42 2.165 54.43 2.358 ;
      RECT 54.39 2.182 54.42 2.375 ;
      RECT 54.38 2.2 54.39 2.393 ;
      RECT 54.365 2.211 54.38 2.404 ;
      RECT 54.325 2.235 54.365 2.42 ;
      RECT 54.29 2.269 54.325 2.437 ;
      RECT 54.26 2.292 54.29 2.449 ;
      RECT 54.245 2.302 54.26 2.458 ;
      RECT 54.205 2.312 54.245 2.469 ;
      RECT 54.185 2.323 54.205 2.481 ;
      RECT 54.18 2.327 54.185 2.488 ;
      RECT 54.165 2.331 54.18 2.493 ;
      RECT 54.155 2.336 54.165 2.498 ;
      RECT 54.15 2.339 54.155 2.501 ;
      RECT 54.12 2.345 54.15 2.508 ;
      RECT 54.085 2.355 54.12 2.522 ;
      RECT 54.025 2.37 54.085 2.542 ;
      RECT 53.97 2.39 54.025 2.566 ;
      RECT 53.941 2.405 53.97 2.584 ;
      RECT 53.855 2.425 53.941 2.609 ;
      RECT 53.85 2.44 53.855 2.629 ;
      RECT 53.84 2.443 53.85 2.63 ;
      RECT 53.815 2.45 53.84 2.715 ;
      RECT 56.51 2.943 56.79 3.28 ;
      RECT 56.51 2.953 56.795 3.238 ;
      RECT 56.51 2.962 56.8 3.135 ;
      RECT 56.51 2.977 56.805 3.003 ;
      RECT 56.51 2.805 56.77 3.28 ;
      RECT 46.81 6.655 47.16 7.005 ;
      RECT 55.635 6.61 55.985 6.96 ;
      RECT 46.81 6.685 55.985 6.885 ;
      RECT 54.23 3.685 54.24 3.875 ;
      RECT 52.49 3.56 52.77 3.84 ;
      RECT 55.535 2.5 55.54 2.985 ;
      RECT 55.43 2.5 55.49 2.76 ;
      RECT 55.755 3.47 55.76 3.545 ;
      RECT 55.745 3.337 55.755 3.58 ;
      RECT 55.735 3.172 55.745 3.601 ;
      RECT 55.73 3.042 55.735 3.617 ;
      RECT 55.72 2.932 55.73 3.633 ;
      RECT 55.715 2.831 55.72 3.65 ;
      RECT 55.71 2.813 55.715 3.66 ;
      RECT 55.705 2.795 55.71 3.67 ;
      RECT 55.695 2.77 55.705 3.685 ;
      RECT 55.69 2.75 55.695 3.7 ;
      RECT 55.67 2.5 55.69 3.725 ;
      RECT 55.655 2.5 55.67 3.758 ;
      RECT 55.625 2.5 55.655 3.78 ;
      RECT 55.605 2.5 55.625 3.794 ;
      RECT 55.585 2.5 55.605 3.31 ;
      RECT 55.6 3.377 55.605 3.799 ;
      RECT 55.595 3.407 55.6 3.801 ;
      RECT 55.59 3.42 55.595 3.804 ;
      RECT 55.585 3.43 55.59 3.808 ;
      RECT 55.58 2.5 55.585 3.228 ;
      RECT 55.58 3.44 55.585 3.81 ;
      RECT 55.575 2.5 55.58 3.205 ;
      RECT 55.565 3.462 55.58 3.81 ;
      RECT 55.56 2.5 55.575 3.15 ;
      RECT 55.555 3.487 55.565 3.81 ;
      RECT 55.555 2.5 55.56 3.095 ;
      RECT 55.545 2.5 55.555 3.043 ;
      RECT 55.55 3.5 55.555 3.811 ;
      RECT 55.545 3.512 55.55 3.812 ;
      RECT 55.54 2.5 55.545 3.003 ;
      RECT 55.54 3.525 55.545 3.813 ;
      RECT 55.525 3.54 55.54 3.814 ;
      RECT 55.53 2.5 55.535 2.965 ;
      RECT 55.525 2.5 55.53 2.93 ;
      RECT 55.52 2.5 55.525 2.905 ;
      RECT 55.515 3.567 55.525 3.816 ;
      RECT 55.51 2.5 55.52 2.863 ;
      RECT 55.51 3.585 55.515 3.817 ;
      RECT 55.505 2.5 55.51 2.823 ;
      RECT 55.505 3.592 55.51 3.818 ;
      RECT 55.5 2.5 55.505 2.795 ;
      RECT 55.495 3.61 55.505 3.819 ;
      RECT 55.49 2.5 55.5 2.775 ;
      RECT 55.485 3.63 55.495 3.821 ;
      RECT 55.475 3.647 55.485 3.822 ;
      RECT 55.44 3.67 55.475 3.825 ;
      RECT 55.385 3.688 55.44 3.831 ;
      RECT 55.299 3.696 55.385 3.84 ;
      RECT 55.213 3.707 55.299 3.851 ;
      RECT 55.127 3.717 55.213 3.862 ;
      RECT 55.041 3.727 55.127 3.874 ;
      RECT 54.955 3.737 55.041 3.885 ;
      RECT 54.935 3.743 54.955 3.891 ;
      RECT 54.855 3.745 54.935 3.895 ;
      RECT 54.85 3.744 54.855 3.9 ;
      RECT 54.842 3.743 54.85 3.9 ;
      RECT 54.756 3.739 54.842 3.898 ;
      RECT 54.67 3.731 54.756 3.895 ;
      RECT 54.584 3.722 54.67 3.891 ;
      RECT 54.498 3.714 54.584 3.888 ;
      RECT 54.412 3.706 54.498 3.884 ;
      RECT 54.326 3.697 54.412 3.881 ;
      RECT 54.24 3.689 54.326 3.877 ;
      RECT 54.185 3.682 54.23 3.875 ;
      RECT 54.1 3.675 54.185 3.873 ;
      RECT 54.026 3.667 54.1 3.869 ;
      RECT 53.94 3.659 54.026 3.866 ;
      RECT 53.937 3.655 53.94 3.864 ;
      RECT 53.851 3.651 53.937 3.863 ;
      RECT 53.765 3.643 53.851 3.86 ;
      RECT 53.68 3.638 53.765 3.857 ;
      RECT 53.594 3.635 53.68 3.854 ;
      RECT 53.508 3.633 53.594 3.851 ;
      RECT 53.422 3.63 53.508 3.848 ;
      RECT 53.336 3.627 53.422 3.845 ;
      RECT 53.25 3.624 53.336 3.842 ;
      RECT 53.174 3.622 53.25 3.839 ;
      RECT 53.088 3.619 53.174 3.836 ;
      RECT 53.002 3.616 53.088 3.834 ;
      RECT 52.916 3.614 53.002 3.831 ;
      RECT 52.83 3.611 52.916 3.828 ;
      RECT 52.77 3.602 52.83 3.826 ;
      RECT 55.28 3.22 55.355 3.48 ;
      RECT 55.26 3.2 55.265 3.48 ;
      RECT 54.58 2.985 54.685 3.28 ;
      RECT 49.025 2.96 49.095 3.22 ;
      RECT 54.92 2.835 54.925 3.206 ;
      RECT 54.91 2.89 54.915 3.206 ;
      RECT 55.215 2.06 55.275 2.32 ;
      RECT 55.27 3.215 55.28 3.48 ;
      RECT 55.265 3.205 55.27 3.48 ;
      RECT 55.185 3.152 55.26 3.48 ;
      RECT 55.21 2.06 55.215 2.34 ;
      RECT 55.2 2.06 55.21 2.36 ;
      RECT 55.185 2.06 55.2 2.39 ;
      RECT 55.17 2.06 55.185 2.433 ;
      RECT 55.165 3.095 55.185 3.48 ;
      RECT 55.155 2.06 55.17 2.47 ;
      RECT 55.15 3.075 55.165 3.48 ;
      RECT 55.15 2.06 55.155 2.493 ;
      RECT 55.14 2.06 55.15 2.518 ;
      RECT 55.11 3.042 55.15 3.48 ;
      RECT 55.115 2.06 55.14 2.568 ;
      RECT 55.11 2.06 55.115 2.623 ;
      RECT 55.105 2.06 55.11 2.665 ;
      RECT 55.095 3.005 55.11 3.48 ;
      RECT 55.1 2.06 55.105 2.708 ;
      RECT 55.095 2.06 55.1 2.773 ;
      RECT 55.09 2.06 55.095 2.795 ;
      RECT 55.09 2.993 55.095 3.345 ;
      RECT 55.085 2.06 55.09 2.863 ;
      RECT 55.085 2.985 55.09 3.328 ;
      RECT 55.08 2.06 55.085 2.908 ;
      RECT 55.075 2.967 55.085 3.305 ;
      RECT 55.075 2.06 55.08 2.945 ;
      RECT 55.065 2.06 55.075 3.285 ;
      RECT 55.06 2.06 55.065 3.268 ;
      RECT 55.055 2.06 55.06 3.253 ;
      RECT 55.05 2.06 55.055 3.238 ;
      RECT 55.03 2.06 55.05 3.228 ;
      RECT 55.025 2.06 55.03 3.218 ;
      RECT 55.015 2.06 55.025 3.214 ;
      RECT 55.01 2.337 55.015 3.213 ;
      RECT 55.005 2.36 55.01 3.212 ;
      RECT 55 2.39 55.005 3.211 ;
      RECT 54.995 2.417 55 3.21 ;
      RECT 54.99 2.445 54.995 3.21 ;
      RECT 54.985 2.472 54.99 3.21 ;
      RECT 54.98 2.492 54.985 3.21 ;
      RECT 54.975 2.52 54.98 3.21 ;
      RECT 54.965 2.562 54.975 3.21 ;
      RECT 54.955 2.607 54.965 3.209 ;
      RECT 54.95 2.66 54.955 3.208 ;
      RECT 54.945 2.692 54.95 3.207 ;
      RECT 54.94 2.712 54.945 3.206 ;
      RECT 54.935 2.75 54.94 3.206 ;
      RECT 54.93 2.772 54.935 3.206 ;
      RECT 54.925 2.797 54.93 3.206 ;
      RECT 54.915 2.862 54.92 3.206 ;
      RECT 54.9 2.922 54.91 3.206 ;
      RECT 54.885 2.932 54.9 3.206 ;
      RECT 54.865 2.942 54.885 3.206 ;
      RECT 54.835 2.947 54.865 3.203 ;
      RECT 54.775 2.957 54.835 3.2 ;
      RECT 54.755 2.966 54.775 3.205 ;
      RECT 54.73 2.972 54.755 3.218 ;
      RECT 54.71 2.977 54.73 3.233 ;
      RECT 54.685 2.982 54.71 3.28 ;
      RECT 54.556 2.984 54.58 3.28 ;
      RECT 54.47 2.979 54.556 3.28 ;
      RECT 54.43 2.976 54.47 3.28 ;
      RECT 54.38 2.978 54.43 3.26 ;
      RECT 54.35 2.982 54.38 3.26 ;
      RECT 54.271 2.992 54.35 3.26 ;
      RECT 54.185 3.007 54.271 3.261 ;
      RECT 54.135 3.017 54.185 3.262 ;
      RECT 54.127 3.02 54.135 3.262 ;
      RECT 54.041 3.022 54.127 3.263 ;
      RECT 53.955 3.026 54.041 3.263 ;
      RECT 53.869 3.03 53.955 3.264 ;
      RECT 53.783 3.033 53.869 3.265 ;
      RECT 53.697 3.037 53.783 3.265 ;
      RECT 53.611 3.041 53.697 3.266 ;
      RECT 53.525 3.044 53.611 3.267 ;
      RECT 53.439 3.048 53.525 3.267 ;
      RECT 53.353 3.052 53.439 3.268 ;
      RECT 53.267 3.056 53.353 3.269 ;
      RECT 53.181 3.059 53.267 3.269 ;
      RECT 53.095 3.063 53.181 3.27 ;
      RECT 53.065 3.065 53.095 3.27 ;
      RECT 52.979 3.068 53.065 3.271 ;
      RECT 52.893 3.072 52.979 3.272 ;
      RECT 52.807 3.076 52.893 3.273 ;
      RECT 52.721 3.079 52.807 3.273 ;
      RECT 52.635 3.083 52.721 3.274 ;
      RECT 52.6 3.088 52.635 3.275 ;
      RECT 52.545 3.098 52.6 3.282 ;
      RECT 52.52 3.11 52.545 3.292 ;
      RECT 52.485 3.123 52.52 3.3 ;
      RECT 52.445 3.14 52.485 3.323 ;
      RECT 52.425 3.153 52.445 3.35 ;
      RECT 52.395 3.165 52.425 3.378 ;
      RECT 52.39 3.173 52.395 3.398 ;
      RECT 52.385 3.176 52.39 3.408 ;
      RECT 52.335 3.188 52.385 3.442 ;
      RECT 52.325 3.203 52.335 3.475 ;
      RECT 52.315 3.209 52.325 3.488 ;
      RECT 52.305 3.216 52.315 3.5 ;
      RECT 52.28 3.229 52.305 3.518 ;
      RECT 52.265 3.244 52.28 3.54 ;
      RECT 52.255 3.252 52.265 3.556 ;
      RECT 52.24 3.261 52.255 3.571 ;
      RECT 52.23 3.271 52.24 3.585 ;
      RECT 52.211 3.284 52.23 3.602 ;
      RECT 52.125 3.329 52.211 3.667 ;
      RECT 52.11 3.374 52.125 3.725 ;
      RECT 52.105 3.383 52.11 3.738 ;
      RECT 52.095 3.39 52.105 3.743 ;
      RECT 52.09 3.395 52.095 3.747 ;
      RECT 52.07 3.405 52.09 3.754 ;
      RECT 52.045 3.425 52.07 3.768 ;
      RECT 52.01 3.45 52.045 3.788 ;
      RECT 51.995 3.473 52.01 3.803 ;
      RECT 51.985 3.483 51.995 3.808 ;
      RECT 51.975 3.491 51.985 3.815 ;
      RECT 51.965 3.5 51.975 3.821 ;
      RECT 51.945 3.512 51.965 3.823 ;
      RECT 51.935 3.525 51.945 3.825 ;
      RECT 51.91 3.54 51.935 3.828 ;
      RECT 51.89 3.557 51.91 3.832 ;
      RECT 51.85 3.585 51.89 3.838 ;
      RECT 51.785 3.632 51.85 3.847 ;
      RECT 51.77 3.665 51.785 3.855 ;
      RECT 51.765 3.672 51.77 3.857 ;
      RECT 51.715 3.697 51.765 3.862 ;
      RECT 51.7 3.721 51.715 3.869 ;
      RECT 51.65 3.726 51.7 3.87 ;
      RECT 51.564 3.73 51.65 3.87 ;
      RECT 51.478 3.73 51.564 3.87 ;
      RECT 51.392 3.73 51.478 3.871 ;
      RECT 51.306 3.73 51.392 3.871 ;
      RECT 51.22 3.73 51.306 3.871 ;
      RECT 51.154 3.73 51.22 3.871 ;
      RECT 51.068 3.73 51.154 3.872 ;
      RECT 50.982 3.73 51.068 3.872 ;
      RECT 50.896 3.731 50.982 3.873 ;
      RECT 50.81 3.731 50.896 3.873 ;
      RECT 50.724 3.731 50.81 3.873 ;
      RECT 50.638 3.731 50.724 3.874 ;
      RECT 50.552 3.731 50.638 3.874 ;
      RECT 50.466 3.732 50.552 3.875 ;
      RECT 50.38 3.732 50.466 3.875 ;
      RECT 50.36 3.732 50.38 3.875 ;
      RECT 50.274 3.732 50.36 3.875 ;
      RECT 50.188 3.732 50.274 3.875 ;
      RECT 50.102 3.733 50.188 3.875 ;
      RECT 50.016 3.733 50.102 3.875 ;
      RECT 49.93 3.733 50.016 3.875 ;
      RECT 49.844 3.734 49.93 3.875 ;
      RECT 49.758 3.734 49.844 3.875 ;
      RECT 49.672 3.734 49.758 3.875 ;
      RECT 49.586 3.734 49.672 3.875 ;
      RECT 49.5 3.735 49.586 3.875 ;
      RECT 49.45 3.732 49.5 3.875 ;
      RECT 49.44 3.73 49.45 3.874 ;
      RECT 49.436 3.73 49.44 3.873 ;
      RECT 49.35 3.725 49.436 3.868 ;
      RECT 49.328 3.718 49.35 3.862 ;
      RECT 49.242 3.709 49.328 3.856 ;
      RECT 49.156 3.696 49.242 3.847 ;
      RECT 49.07 3.682 49.156 3.837 ;
      RECT 49.025 3.672 49.07 3.83 ;
      RECT 49.005 2.96 49.025 3.238 ;
      RECT 49.005 3.665 49.025 3.826 ;
      RECT 48.975 2.96 49.005 3.26 ;
      RECT 48.965 3.632 49.005 3.823 ;
      RECT 48.96 2.96 48.975 3.28 ;
      RECT 48.96 3.597 48.965 3.821 ;
      RECT 48.955 2.96 48.96 3.405 ;
      RECT 48.955 3.557 48.96 3.821 ;
      RECT 48.945 2.96 48.955 3.821 ;
      RECT 48.87 2.96 48.945 3.815 ;
      RECT 48.84 2.96 48.87 3.805 ;
      RECT 48.835 2.96 48.84 3.797 ;
      RECT 48.83 3.002 48.835 3.79 ;
      RECT 48.82 3.071 48.83 3.781 ;
      RECT 48.815 3.141 48.82 3.733 ;
      RECT 48.81 3.205 48.815 3.63 ;
      RECT 48.805 3.24 48.81 3.585 ;
      RECT 48.803 3.277 48.805 3.477 ;
      RECT 48.8 3.285 48.803 3.47 ;
      RECT 48.795 3.35 48.8 3.413 ;
      RECT 52.87 2.44 53.15 2.72 ;
      RECT 52.86 2.44 53.15 2.583 ;
      RECT 52.815 2.305 53.075 2.565 ;
      RECT 52.815 2.42 53.13 2.565 ;
      RECT 52.815 2.39 53.125 2.565 ;
      RECT 52.815 2.377 53.115 2.565 ;
      RECT 52.815 2.367 53.11 2.565 ;
      RECT 48.79 2.35 49.05 2.61 ;
      RECT 52.56 1.9 52.82 2.16 ;
      RECT 52.55 1.925 52.82 2.12 ;
      RECT 52.545 1.925 52.55 2.119 ;
      RECT 52.475 1.92 52.545 2.111 ;
      RECT 52.39 1.907 52.475 2.094 ;
      RECT 52.386 1.899 52.39 2.084 ;
      RECT 52.3 1.892 52.386 2.074 ;
      RECT 52.291 1.884 52.3 2.064 ;
      RECT 52.205 1.877 52.291 2.052 ;
      RECT 52.185 1.868 52.205 2.038 ;
      RECT 52.13 1.863 52.185 2.03 ;
      RECT 52.12 1.857 52.13 2.024 ;
      RECT 52.1 1.855 52.12 2.02 ;
      RECT 52.092 1.854 52.1 2.016 ;
      RECT 52.006 1.846 52.092 2.005 ;
      RECT 51.92 1.832 52.006 1.985 ;
      RECT 51.86 1.82 51.92 1.97 ;
      RECT 51.85 1.815 51.86 1.965 ;
      RECT 51.8 1.815 51.85 1.967 ;
      RECT 51.753 1.817 51.8 1.971 ;
      RECT 51.667 1.824 51.753 1.976 ;
      RECT 51.581 1.832 51.667 1.982 ;
      RECT 51.495 1.841 51.581 1.988 ;
      RECT 51.436 1.847 51.495 1.993 ;
      RECT 51.35 1.852 51.436 1.999 ;
      RECT 51.275 1.857 51.35 2.005 ;
      RECT 51.236 1.859 51.275 2.01 ;
      RECT 51.15 1.856 51.236 2.015 ;
      RECT 51.065 1.854 51.15 2.022 ;
      RECT 51.033 1.853 51.065 2.025 ;
      RECT 50.947 1.852 51.033 2.026 ;
      RECT 50.861 1.851 50.947 2.027 ;
      RECT 50.775 1.85 50.861 2.027 ;
      RECT 50.689 1.849 50.775 2.028 ;
      RECT 50.603 1.848 50.689 2.029 ;
      RECT 50.517 1.847 50.603 2.03 ;
      RECT 50.431 1.846 50.517 2.03 ;
      RECT 50.345 1.845 50.431 2.031 ;
      RECT 50.295 1.845 50.345 2.032 ;
      RECT 50.281 1.846 50.295 2.032 ;
      RECT 50.195 1.853 50.281 2.033 ;
      RECT 50.121 1.864 50.195 2.034 ;
      RECT 50.035 1.873 50.121 2.035 ;
      RECT 50 1.88 50.035 2.05 ;
      RECT 49.975 1.883 50 2.08 ;
      RECT 49.95 1.892 49.975 2.109 ;
      RECT 49.94 1.903 49.95 2.129 ;
      RECT 49.93 1.911 49.94 2.143 ;
      RECT 49.925 1.917 49.93 2.153 ;
      RECT 49.9 1.934 49.925 2.17 ;
      RECT 49.885 1.956 49.9 2.198 ;
      RECT 49.855 1.982 49.885 2.228 ;
      RECT 49.835 2.011 49.855 2.258 ;
      RECT 49.83 2.026 49.835 2.275 ;
      RECT 49.81 2.041 49.83 2.29 ;
      RECT 49.8 2.059 49.81 2.308 ;
      RECT 49.79 2.07 49.8 2.323 ;
      RECT 49.74 2.102 49.79 2.349 ;
      RECT 49.735 2.132 49.74 2.369 ;
      RECT 49.725 2.145 49.735 2.375 ;
      RECT 49.716 2.155 49.725 2.383 ;
      RECT 49.705 2.166 49.716 2.391 ;
      RECT 49.7 2.176 49.705 2.397 ;
      RECT 49.685 2.197 49.7 2.404 ;
      RECT 49.67 2.227 49.685 2.412 ;
      RECT 49.635 2.257 49.67 2.418 ;
      RECT 49.61 2.275 49.635 2.425 ;
      RECT 49.56 2.283 49.61 2.434 ;
      RECT 49.535 2.288 49.56 2.443 ;
      RECT 49.48 2.294 49.535 2.453 ;
      RECT 49.475 2.299 49.48 2.461 ;
      RECT 49.461 2.302 49.475 2.463 ;
      RECT 49.375 2.314 49.461 2.475 ;
      RECT 49.365 2.326 49.375 2.488 ;
      RECT 49.28 2.339 49.365 2.5 ;
      RECT 49.236 2.356 49.28 2.514 ;
      RECT 49.15 2.373 49.236 2.53 ;
      RECT 49.12 2.387 49.15 2.544 ;
      RECT 49.11 2.392 49.12 2.549 ;
      RECT 49.05 2.395 49.11 2.558 ;
      RECT 51.94 2.665 52.2 2.925 ;
      RECT 51.94 2.665 52.22 2.778 ;
      RECT 51.94 2.665 52.245 2.745 ;
      RECT 51.94 2.665 52.25 2.725 ;
      RECT 51.99 2.44 52.27 2.72 ;
      RECT 51.545 3.175 51.805 3.435 ;
      RECT 51.535 3.032 51.73 3.373 ;
      RECT 51.53 3.14 51.745 3.365 ;
      RECT 51.525 3.19 51.805 3.355 ;
      RECT 51.515 3.267 51.805 3.34 ;
      RECT 51.535 3.115 51.745 3.373 ;
      RECT 51.545 2.99 51.73 3.435 ;
      RECT 51.545 2.885 51.71 3.435 ;
      RECT 51.555 2.872 51.71 3.435 ;
      RECT 51.555 2.83 51.7 3.435 ;
      RECT 51.56 2.755 51.7 3.435 ;
      RECT 51.59 2.405 51.7 3.435 ;
      RECT 51.595 2.135 51.72 2.758 ;
      RECT 51.565 2.71 51.72 2.758 ;
      RECT 51.58 2.512 51.7 3.435 ;
      RECT 51.57 2.622 51.72 2.758 ;
      RECT 51.595 2.135 51.735 2.615 ;
      RECT 51.595 2.135 51.755 2.49 ;
      RECT 51.56 2.135 51.82 2.395 ;
      RECT 51.03 2.44 51.31 2.72 ;
      RECT 51.015 2.44 51.31 2.7 ;
      RECT 49.07 3.305 49.33 3.565 ;
      RECT 50.855 3.16 51.115 3.42 ;
      RECT 50.835 3.18 51.115 3.395 ;
      RECT 50.792 3.18 50.835 3.394 ;
      RECT 50.706 3.181 50.792 3.391 ;
      RECT 50.62 3.182 50.706 3.387 ;
      RECT 50.545 3.184 50.62 3.384 ;
      RECT 50.522 3.185 50.545 3.382 ;
      RECT 50.436 3.186 50.522 3.38 ;
      RECT 50.35 3.187 50.436 3.377 ;
      RECT 50.326 3.188 50.35 3.375 ;
      RECT 50.24 3.19 50.326 3.372 ;
      RECT 50.155 3.192 50.24 3.373 ;
      RECT 50.098 3.193 50.155 3.379 ;
      RECT 50.012 3.195 50.098 3.389 ;
      RECT 49.926 3.198 50.012 3.402 ;
      RECT 49.84 3.2 49.926 3.414 ;
      RECT 49.826 3.201 49.84 3.421 ;
      RECT 49.74 3.202 49.826 3.429 ;
      RECT 49.7 3.204 49.74 3.438 ;
      RECT 49.691 3.205 49.7 3.441 ;
      RECT 49.605 3.213 49.691 3.447 ;
      RECT 49.585 3.222 49.605 3.455 ;
      RECT 49.5 3.237 49.585 3.463 ;
      RECT 49.44 3.26 49.5 3.474 ;
      RECT 49.43 3.272 49.44 3.479 ;
      RECT 49.39 3.282 49.43 3.483 ;
      RECT 49.335 3.299 49.39 3.491 ;
      RECT 49.33 3.309 49.335 3.495 ;
      RECT 50.396 2.44 50.455 2.837 ;
      RECT 50.31 2.44 50.515 2.828 ;
      RECT 50.305 2.47 50.515 2.823 ;
      RECT 50.271 2.47 50.515 2.821 ;
      RECT 50.185 2.47 50.515 2.815 ;
      RECT 50.14 2.47 50.535 2.793 ;
      RECT 50.14 2.47 50.555 2.748 ;
      RECT 50.1 2.47 50.555 2.738 ;
      RECT 50.31 2.44 50.59 2.72 ;
      RECT 50.045 2.44 50.305 2.7 ;
      RECT 49.23 1.92 49.49 2.18 ;
      RECT 49.31 1.88 49.59 2.16 ;
      RECT 43.675 6.22 43.995 6.545 ;
      RECT 43.705 5.695 43.875 6.545 ;
      RECT 43.705 5.695 43.88 6.045 ;
      RECT 43.705 5.695 44.68 5.87 ;
      RECT 44.505 1.965 44.68 5.87 ;
      RECT 44.45 1.965 44.8 2.315 ;
      RECT 44.475 6.655 44.8 6.98 ;
      RECT 43.36 6.745 44.8 6.915 ;
      RECT 43.36 2.395 43.52 6.915 ;
      RECT 43.675 2.365 43.995 2.685 ;
      RECT 43.36 2.395 43.995 2.565 ;
      RECT 42.625 5.855 42.975 6.205 ;
      RECT 42.695 2.705 42.87 6.205 ;
      RECT 42.62 2.705 42.97 3.055 ;
      RECT 32.085 3 32.365 3.28 ;
      RECT 32.055 3 32.365 3.265 ;
      RECT 32.05 3 32.365 3.263 ;
      RECT 32.045 1.33 32.215 3.257 ;
      RECT 32.04 2.967 32.31 3.25 ;
      RECT 32.035 3 32.365 3.243 ;
      RECT 32.005 2.97 32.31 3.23 ;
      RECT 32.005 2.997 32.33 3.23 ;
      RECT 32.005 2.987 32.325 3.23 ;
      RECT 32.005 2.972 32.32 3.23 ;
      RECT 32.045 2.962 32.31 3.257 ;
      RECT 32.045 2.957 32.3 3.257 ;
      RECT 32.045 2.956 32.285 3.257 ;
      RECT 42.015 1.34 42.365 1.69 ;
      RECT 42.01 1.34 42.365 1.595 ;
      RECT 32.045 1.33 42.255 1.5 ;
      RECT 41.69 2.85 42.06 3.22 ;
      RECT 41.775 2.235 41.945 3.22 ;
      RECT 37.795 2.455 38.03 2.715 ;
      RECT 40.94 2.235 41.105 2.495 ;
      RECT 40.845 2.225 40.86 2.495 ;
      RECT 40.94 2.235 41.945 2.415 ;
      RECT 39.445 1.795 39.485 1.935 ;
      RECT 40.86 2.23 40.94 2.495 ;
      RECT 40.805 2.225 40.845 2.461 ;
      RECT 40.791 2.225 40.805 2.461 ;
      RECT 40.705 2.23 40.791 2.463 ;
      RECT 40.66 2.237 40.705 2.465 ;
      RECT 40.63 2.237 40.66 2.467 ;
      RECT 40.605 2.232 40.63 2.469 ;
      RECT 40.575 2.228 40.605 2.478 ;
      RECT 40.565 2.225 40.575 2.49 ;
      RECT 40.56 2.225 40.565 2.498 ;
      RECT 40.555 2.225 40.56 2.503 ;
      RECT 40.545 2.224 40.555 2.513 ;
      RECT 40.54 2.223 40.545 2.523 ;
      RECT 40.525 2.222 40.54 2.528 ;
      RECT 40.497 2.219 40.525 2.555 ;
      RECT 40.411 2.211 40.497 2.555 ;
      RECT 40.325 2.2 40.411 2.555 ;
      RECT 40.285 2.185 40.325 2.555 ;
      RECT 40.245 2.159 40.285 2.555 ;
      RECT 40.24 2.141 40.245 2.367 ;
      RECT 40.23 2.137 40.24 2.357 ;
      RECT 40.215 2.127 40.23 2.344 ;
      RECT 40.195 2.111 40.215 2.329 ;
      RECT 40.18 2.096 40.195 2.314 ;
      RECT 40.17 2.085 40.18 2.304 ;
      RECT 40.145 2.069 40.17 2.293 ;
      RECT 40.14 2.056 40.145 2.283 ;
      RECT 40.135 2.052 40.14 2.278 ;
      RECT 40.08 2.038 40.135 2.256 ;
      RECT 40.041 2.019 40.08 2.22 ;
      RECT 39.955 1.993 40.041 2.173 ;
      RECT 39.951 1.975 39.955 2.139 ;
      RECT 39.865 1.956 39.951 2.117 ;
      RECT 39.86 1.938 39.865 2.095 ;
      RECT 39.855 1.936 39.86 2.093 ;
      RECT 39.845 1.935 39.855 2.088 ;
      RECT 39.785 1.922 39.845 2.074 ;
      RECT 39.74 1.9 39.785 2.053 ;
      RECT 39.68 1.877 39.74 2.032 ;
      RECT 39.616 1.852 39.68 2.007 ;
      RECT 39.53 1.822 39.616 1.976 ;
      RECT 39.515 1.802 39.53 1.955 ;
      RECT 39.485 1.797 39.515 1.946 ;
      RECT 39.432 1.795 39.445 1.935 ;
      RECT 39.346 1.795 39.432 1.937 ;
      RECT 39.26 1.795 39.346 1.939 ;
      RECT 39.24 1.795 39.26 1.943 ;
      RECT 39.195 1.797 39.24 1.954 ;
      RECT 39.155 1.807 39.195 1.97 ;
      RECT 39.151 1.816 39.155 1.978 ;
      RECT 39.065 1.836 39.151 1.994 ;
      RECT 39.055 1.855 39.065 2.012 ;
      RECT 39.05 1.857 39.055 2.015 ;
      RECT 39.04 1.861 39.05 2.018 ;
      RECT 39.02 1.866 39.04 2.028 ;
      RECT 38.99 1.876 39.02 2.048 ;
      RECT 38.985 1.883 38.99 2.062 ;
      RECT 38.975 1.887 38.985 2.069 ;
      RECT 38.96 1.895 38.975 2.08 ;
      RECT 38.95 1.905 38.96 2.091 ;
      RECT 38.94 1.912 38.95 2.099 ;
      RECT 38.915 1.925 38.94 2.114 ;
      RECT 38.851 1.961 38.915 2.153 ;
      RECT 38.765 2.024 38.851 2.217 ;
      RECT 38.73 2.075 38.765 2.27 ;
      RECT 38.725 2.092 38.73 2.287 ;
      RECT 38.71 2.101 38.725 2.294 ;
      RECT 38.69 2.116 38.71 2.308 ;
      RECT 38.685 2.127 38.69 2.318 ;
      RECT 38.665 2.14 38.685 2.328 ;
      RECT 38.66 2.15 38.665 2.338 ;
      RECT 38.645 2.155 38.66 2.347 ;
      RECT 38.635 2.165 38.645 2.358 ;
      RECT 38.605 2.182 38.635 2.375 ;
      RECT 38.595 2.2 38.605 2.393 ;
      RECT 38.58 2.211 38.595 2.404 ;
      RECT 38.54 2.235 38.58 2.42 ;
      RECT 38.505 2.269 38.54 2.437 ;
      RECT 38.475 2.292 38.505 2.449 ;
      RECT 38.46 2.302 38.475 2.458 ;
      RECT 38.42 2.312 38.46 2.469 ;
      RECT 38.4 2.323 38.42 2.481 ;
      RECT 38.395 2.327 38.4 2.488 ;
      RECT 38.38 2.331 38.395 2.493 ;
      RECT 38.37 2.336 38.38 2.498 ;
      RECT 38.365 2.339 38.37 2.501 ;
      RECT 38.335 2.345 38.365 2.508 ;
      RECT 38.3 2.355 38.335 2.522 ;
      RECT 38.24 2.37 38.3 2.542 ;
      RECT 38.185 2.39 38.24 2.566 ;
      RECT 38.156 2.405 38.185 2.584 ;
      RECT 38.07 2.425 38.156 2.609 ;
      RECT 38.065 2.44 38.07 2.629 ;
      RECT 38.055 2.443 38.065 2.63 ;
      RECT 38.03 2.45 38.055 2.715 ;
      RECT 40.725 2.943 41.005 3.28 ;
      RECT 40.725 2.953 41.01 3.238 ;
      RECT 40.725 2.962 41.015 3.135 ;
      RECT 40.725 2.977 41.02 3.003 ;
      RECT 40.725 2.805 40.985 3.28 ;
      RECT 31.08 6.66 31.43 7.01 ;
      RECT 39.905 6.615 40.255 6.965 ;
      RECT 31.08 6.69 40.255 6.89 ;
      RECT 38.445 3.685 38.455 3.875 ;
      RECT 36.705 3.56 36.985 3.84 ;
      RECT 39.75 2.5 39.755 2.985 ;
      RECT 39.645 2.5 39.705 2.76 ;
      RECT 39.97 3.47 39.975 3.545 ;
      RECT 39.96 3.337 39.97 3.58 ;
      RECT 39.95 3.172 39.96 3.601 ;
      RECT 39.945 3.042 39.95 3.617 ;
      RECT 39.935 2.932 39.945 3.633 ;
      RECT 39.93 2.831 39.935 3.65 ;
      RECT 39.925 2.813 39.93 3.66 ;
      RECT 39.92 2.795 39.925 3.67 ;
      RECT 39.91 2.77 39.92 3.685 ;
      RECT 39.905 2.75 39.91 3.7 ;
      RECT 39.885 2.5 39.905 3.725 ;
      RECT 39.87 2.5 39.885 3.758 ;
      RECT 39.84 2.5 39.87 3.78 ;
      RECT 39.82 2.5 39.84 3.794 ;
      RECT 39.8 2.5 39.82 3.31 ;
      RECT 39.815 3.377 39.82 3.799 ;
      RECT 39.81 3.407 39.815 3.801 ;
      RECT 39.805 3.42 39.81 3.804 ;
      RECT 39.8 3.43 39.805 3.808 ;
      RECT 39.795 2.5 39.8 3.228 ;
      RECT 39.795 3.44 39.8 3.81 ;
      RECT 39.79 2.5 39.795 3.205 ;
      RECT 39.78 3.462 39.795 3.81 ;
      RECT 39.775 2.5 39.79 3.15 ;
      RECT 39.77 3.487 39.78 3.81 ;
      RECT 39.77 2.5 39.775 3.095 ;
      RECT 39.76 2.5 39.77 3.043 ;
      RECT 39.765 3.5 39.77 3.811 ;
      RECT 39.76 3.512 39.765 3.812 ;
      RECT 39.755 2.5 39.76 3.003 ;
      RECT 39.755 3.525 39.76 3.813 ;
      RECT 39.74 3.54 39.755 3.814 ;
      RECT 39.745 2.5 39.75 2.965 ;
      RECT 39.74 2.5 39.745 2.93 ;
      RECT 39.735 2.5 39.74 2.905 ;
      RECT 39.73 3.567 39.74 3.816 ;
      RECT 39.725 2.5 39.735 2.863 ;
      RECT 39.725 3.585 39.73 3.817 ;
      RECT 39.72 2.5 39.725 2.823 ;
      RECT 39.72 3.592 39.725 3.818 ;
      RECT 39.715 2.5 39.72 2.795 ;
      RECT 39.71 3.61 39.72 3.819 ;
      RECT 39.705 2.5 39.715 2.775 ;
      RECT 39.7 3.63 39.71 3.821 ;
      RECT 39.69 3.647 39.7 3.822 ;
      RECT 39.655 3.67 39.69 3.825 ;
      RECT 39.6 3.688 39.655 3.831 ;
      RECT 39.514 3.696 39.6 3.84 ;
      RECT 39.428 3.707 39.514 3.851 ;
      RECT 39.342 3.717 39.428 3.862 ;
      RECT 39.256 3.727 39.342 3.874 ;
      RECT 39.17 3.737 39.256 3.885 ;
      RECT 39.15 3.743 39.17 3.891 ;
      RECT 39.07 3.745 39.15 3.895 ;
      RECT 39.065 3.744 39.07 3.9 ;
      RECT 39.057 3.743 39.065 3.9 ;
      RECT 38.971 3.739 39.057 3.898 ;
      RECT 38.885 3.731 38.971 3.895 ;
      RECT 38.799 3.722 38.885 3.891 ;
      RECT 38.713 3.714 38.799 3.888 ;
      RECT 38.627 3.706 38.713 3.884 ;
      RECT 38.541 3.697 38.627 3.881 ;
      RECT 38.455 3.689 38.541 3.877 ;
      RECT 38.4 3.682 38.445 3.875 ;
      RECT 38.315 3.675 38.4 3.873 ;
      RECT 38.241 3.667 38.315 3.869 ;
      RECT 38.155 3.659 38.241 3.866 ;
      RECT 38.152 3.655 38.155 3.864 ;
      RECT 38.066 3.651 38.152 3.863 ;
      RECT 37.98 3.643 38.066 3.86 ;
      RECT 37.895 3.638 37.98 3.857 ;
      RECT 37.809 3.635 37.895 3.854 ;
      RECT 37.723 3.633 37.809 3.851 ;
      RECT 37.637 3.63 37.723 3.848 ;
      RECT 37.551 3.627 37.637 3.845 ;
      RECT 37.465 3.624 37.551 3.842 ;
      RECT 37.389 3.622 37.465 3.839 ;
      RECT 37.303 3.619 37.389 3.836 ;
      RECT 37.217 3.616 37.303 3.834 ;
      RECT 37.131 3.614 37.217 3.831 ;
      RECT 37.045 3.611 37.131 3.828 ;
      RECT 36.985 3.602 37.045 3.826 ;
      RECT 39.495 3.22 39.57 3.48 ;
      RECT 39.475 3.2 39.48 3.48 ;
      RECT 38.795 2.985 38.9 3.28 ;
      RECT 33.24 2.96 33.31 3.22 ;
      RECT 39.135 2.835 39.14 3.206 ;
      RECT 39.125 2.89 39.13 3.206 ;
      RECT 39.43 2.06 39.49 2.32 ;
      RECT 39.485 3.215 39.495 3.48 ;
      RECT 39.48 3.205 39.485 3.48 ;
      RECT 39.4 3.152 39.475 3.48 ;
      RECT 39.425 2.06 39.43 2.34 ;
      RECT 39.415 2.06 39.425 2.36 ;
      RECT 39.4 2.06 39.415 2.39 ;
      RECT 39.385 2.06 39.4 2.433 ;
      RECT 39.38 3.095 39.4 3.48 ;
      RECT 39.37 2.06 39.385 2.47 ;
      RECT 39.365 3.075 39.38 3.48 ;
      RECT 39.365 2.06 39.37 2.493 ;
      RECT 39.355 2.06 39.365 2.518 ;
      RECT 39.325 3.042 39.365 3.48 ;
      RECT 39.33 2.06 39.355 2.568 ;
      RECT 39.325 2.06 39.33 2.623 ;
      RECT 39.32 2.06 39.325 2.665 ;
      RECT 39.31 3.005 39.325 3.48 ;
      RECT 39.315 2.06 39.32 2.708 ;
      RECT 39.31 2.06 39.315 2.773 ;
      RECT 39.305 2.06 39.31 2.795 ;
      RECT 39.305 2.993 39.31 3.345 ;
      RECT 39.3 2.06 39.305 2.863 ;
      RECT 39.3 2.985 39.305 3.328 ;
      RECT 39.295 2.06 39.3 2.908 ;
      RECT 39.29 2.967 39.3 3.305 ;
      RECT 39.29 2.06 39.295 2.945 ;
      RECT 39.28 2.06 39.29 3.285 ;
      RECT 39.275 2.06 39.28 3.268 ;
      RECT 39.27 2.06 39.275 3.253 ;
      RECT 39.265 2.06 39.27 3.238 ;
      RECT 39.245 2.06 39.265 3.228 ;
      RECT 39.24 2.06 39.245 3.218 ;
      RECT 39.23 2.06 39.24 3.214 ;
      RECT 39.225 2.337 39.23 3.213 ;
      RECT 39.22 2.36 39.225 3.212 ;
      RECT 39.215 2.39 39.22 3.211 ;
      RECT 39.21 2.417 39.215 3.21 ;
      RECT 39.205 2.445 39.21 3.21 ;
      RECT 39.2 2.472 39.205 3.21 ;
      RECT 39.195 2.492 39.2 3.21 ;
      RECT 39.19 2.52 39.195 3.21 ;
      RECT 39.18 2.562 39.19 3.21 ;
      RECT 39.17 2.607 39.18 3.209 ;
      RECT 39.165 2.66 39.17 3.208 ;
      RECT 39.16 2.692 39.165 3.207 ;
      RECT 39.155 2.712 39.16 3.206 ;
      RECT 39.15 2.75 39.155 3.206 ;
      RECT 39.145 2.772 39.15 3.206 ;
      RECT 39.14 2.797 39.145 3.206 ;
      RECT 39.13 2.862 39.135 3.206 ;
      RECT 39.115 2.922 39.125 3.206 ;
      RECT 39.1 2.932 39.115 3.206 ;
      RECT 39.08 2.942 39.1 3.206 ;
      RECT 39.05 2.947 39.08 3.203 ;
      RECT 38.99 2.957 39.05 3.2 ;
      RECT 38.97 2.966 38.99 3.205 ;
      RECT 38.945 2.972 38.97 3.218 ;
      RECT 38.925 2.977 38.945 3.233 ;
      RECT 38.9 2.982 38.925 3.28 ;
      RECT 38.771 2.984 38.795 3.28 ;
      RECT 38.685 2.979 38.771 3.28 ;
      RECT 38.645 2.976 38.685 3.28 ;
      RECT 38.595 2.978 38.645 3.26 ;
      RECT 38.565 2.982 38.595 3.26 ;
      RECT 38.486 2.992 38.565 3.26 ;
      RECT 38.4 3.007 38.486 3.261 ;
      RECT 38.35 3.017 38.4 3.262 ;
      RECT 38.342 3.02 38.35 3.262 ;
      RECT 38.256 3.022 38.342 3.263 ;
      RECT 38.17 3.026 38.256 3.263 ;
      RECT 38.084 3.03 38.17 3.264 ;
      RECT 37.998 3.033 38.084 3.265 ;
      RECT 37.912 3.037 37.998 3.265 ;
      RECT 37.826 3.041 37.912 3.266 ;
      RECT 37.74 3.044 37.826 3.267 ;
      RECT 37.654 3.048 37.74 3.267 ;
      RECT 37.568 3.052 37.654 3.268 ;
      RECT 37.482 3.056 37.568 3.269 ;
      RECT 37.396 3.059 37.482 3.269 ;
      RECT 37.31 3.063 37.396 3.27 ;
      RECT 37.28 3.065 37.31 3.27 ;
      RECT 37.194 3.068 37.28 3.271 ;
      RECT 37.108 3.072 37.194 3.272 ;
      RECT 37.022 3.076 37.108 3.273 ;
      RECT 36.936 3.079 37.022 3.273 ;
      RECT 36.85 3.083 36.936 3.274 ;
      RECT 36.815 3.088 36.85 3.275 ;
      RECT 36.76 3.098 36.815 3.282 ;
      RECT 36.735 3.11 36.76 3.292 ;
      RECT 36.7 3.123 36.735 3.3 ;
      RECT 36.66 3.14 36.7 3.323 ;
      RECT 36.64 3.153 36.66 3.35 ;
      RECT 36.61 3.165 36.64 3.378 ;
      RECT 36.605 3.173 36.61 3.398 ;
      RECT 36.6 3.176 36.605 3.408 ;
      RECT 36.55 3.188 36.6 3.442 ;
      RECT 36.54 3.203 36.55 3.475 ;
      RECT 36.53 3.209 36.54 3.488 ;
      RECT 36.52 3.216 36.53 3.5 ;
      RECT 36.495 3.229 36.52 3.518 ;
      RECT 36.48 3.244 36.495 3.54 ;
      RECT 36.47 3.252 36.48 3.556 ;
      RECT 36.455 3.261 36.47 3.571 ;
      RECT 36.445 3.271 36.455 3.585 ;
      RECT 36.426 3.284 36.445 3.602 ;
      RECT 36.34 3.329 36.426 3.667 ;
      RECT 36.325 3.374 36.34 3.725 ;
      RECT 36.32 3.383 36.325 3.738 ;
      RECT 36.31 3.39 36.32 3.743 ;
      RECT 36.305 3.395 36.31 3.747 ;
      RECT 36.285 3.405 36.305 3.754 ;
      RECT 36.26 3.425 36.285 3.768 ;
      RECT 36.225 3.45 36.26 3.788 ;
      RECT 36.21 3.473 36.225 3.803 ;
      RECT 36.2 3.483 36.21 3.808 ;
      RECT 36.19 3.491 36.2 3.815 ;
      RECT 36.18 3.5 36.19 3.821 ;
      RECT 36.16 3.512 36.18 3.823 ;
      RECT 36.15 3.525 36.16 3.825 ;
      RECT 36.125 3.54 36.15 3.828 ;
      RECT 36.105 3.557 36.125 3.832 ;
      RECT 36.065 3.585 36.105 3.838 ;
      RECT 36 3.632 36.065 3.847 ;
      RECT 35.985 3.665 36 3.855 ;
      RECT 35.98 3.672 35.985 3.857 ;
      RECT 35.93 3.697 35.98 3.862 ;
      RECT 35.915 3.721 35.93 3.869 ;
      RECT 35.865 3.726 35.915 3.87 ;
      RECT 35.779 3.73 35.865 3.87 ;
      RECT 35.693 3.73 35.779 3.87 ;
      RECT 35.607 3.73 35.693 3.871 ;
      RECT 35.521 3.73 35.607 3.871 ;
      RECT 35.435 3.73 35.521 3.871 ;
      RECT 35.369 3.73 35.435 3.871 ;
      RECT 35.283 3.73 35.369 3.872 ;
      RECT 35.197 3.73 35.283 3.872 ;
      RECT 35.111 3.731 35.197 3.873 ;
      RECT 35.025 3.731 35.111 3.873 ;
      RECT 34.939 3.731 35.025 3.873 ;
      RECT 34.853 3.731 34.939 3.874 ;
      RECT 34.767 3.731 34.853 3.874 ;
      RECT 34.681 3.732 34.767 3.875 ;
      RECT 34.595 3.732 34.681 3.875 ;
      RECT 34.575 3.732 34.595 3.875 ;
      RECT 34.489 3.732 34.575 3.875 ;
      RECT 34.403 3.732 34.489 3.875 ;
      RECT 34.317 3.733 34.403 3.875 ;
      RECT 34.231 3.733 34.317 3.875 ;
      RECT 34.145 3.733 34.231 3.875 ;
      RECT 34.059 3.734 34.145 3.875 ;
      RECT 33.973 3.734 34.059 3.875 ;
      RECT 33.887 3.734 33.973 3.875 ;
      RECT 33.801 3.734 33.887 3.875 ;
      RECT 33.715 3.735 33.801 3.875 ;
      RECT 33.665 3.732 33.715 3.875 ;
      RECT 33.655 3.73 33.665 3.874 ;
      RECT 33.651 3.73 33.655 3.873 ;
      RECT 33.565 3.725 33.651 3.868 ;
      RECT 33.543 3.718 33.565 3.862 ;
      RECT 33.457 3.709 33.543 3.856 ;
      RECT 33.371 3.696 33.457 3.847 ;
      RECT 33.285 3.682 33.371 3.837 ;
      RECT 33.24 3.672 33.285 3.83 ;
      RECT 33.22 2.96 33.24 3.238 ;
      RECT 33.22 3.665 33.24 3.826 ;
      RECT 33.19 2.96 33.22 3.26 ;
      RECT 33.18 3.632 33.22 3.823 ;
      RECT 33.175 2.96 33.19 3.28 ;
      RECT 33.175 3.597 33.18 3.821 ;
      RECT 33.17 2.96 33.175 3.405 ;
      RECT 33.17 3.557 33.175 3.821 ;
      RECT 33.16 2.96 33.17 3.821 ;
      RECT 33.085 2.96 33.16 3.815 ;
      RECT 33.055 2.96 33.085 3.805 ;
      RECT 33.05 2.96 33.055 3.797 ;
      RECT 33.045 3.002 33.05 3.79 ;
      RECT 33.035 3.071 33.045 3.781 ;
      RECT 33.03 3.141 33.035 3.733 ;
      RECT 33.025 3.205 33.03 3.63 ;
      RECT 33.02 3.24 33.025 3.585 ;
      RECT 33.018 3.277 33.02 3.477 ;
      RECT 33.015 3.285 33.018 3.47 ;
      RECT 33.01 3.35 33.015 3.413 ;
      RECT 37.085 2.44 37.365 2.72 ;
      RECT 37.075 2.44 37.365 2.583 ;
      RECT 37.03 2.305 37.29 2.565 ;
      RECT 37.03 2.42 37.345 2.565 ;
      RECT 37.03 2.39 37.34 2.565 ;
      RECT 37.03 2.377 37.33 2.565 ;
      RECT 37.03 2.367 37.325 2.565 ;
      RECT 33.005 2.35 33.265 2.61 ;
      RECT 36.775 1.9 37.035 2.16 ;
      RECT 36.765 1.925 37.035 2.12 ;
      RECT 36.76 1.925 36.765 2.119 ;
      RECT 36.69 1.92 36.76 2.111 ;
      RECT 36.605 1.907 36.69 2.094 ;
      RECT 36.601 1.899 36.605 2.084 ;
      RECT 36.515 1.892 36.601 2.074 ;
      RECT 36.506 1.884 36.515 2.064 ;
      RECT 36.42 1.877 36.506 2.052 ;
      RECT 36.4 1.868 36.42 2.038 ;
      RECT 36.345 1.863 36.4 2.03 ;
      RECT 36.335 1.857 36.345 2.024 ;
      RECT 36.315 1.855 36.335 2.02 ;
      RECT 36.307 1.854 36.315 2.016 ;
      RECT 36.221 1.846 36.307 2.005 ;
      RECT 36.135 1.832 36.221 1.985 ;
      RECT 36.075 1.82 36.135 1.97 ;
      RECT 36.065 1.815 36.075 1.965 ;
      RECT 36.015 1.815 36.065 1.967 ;
      RECT 35.968 1.817 36.015 1.971 ;
      RECT 35.882 1.824 35.968 1.976 ;
      RECT 35.796 1.832 35.882 1.982 ;
      RECT 35.71 1.841 35.796 1.988 ;
      RECT 35.651 1.847 35.71 1.993 ;
      RECT 35.565 1.852 35.651 1.999 ;
      RECT 35.49 1.857 35.565 2.005 ;
      RECT 35.451 1.859 35.49 2.01 ;
      RECT 35.365 1.856 35.451 2.015 ;
      RECT 35.28 1.854 35.365 2.022 ;
      RECT 35.248 1.853 35.28 2.025 ;
      RECT 35.162 1.852 35.248 2.026 ;
      RECT 35.076 1.851 35.162 2.027 ;
      RECT 34.99 1.85 35.076 2.027 ;
      RECT 34.904 1.849 34.99 2.028 ;
      RECT 34.818 1.848 34.904 2.029 ;
      RECT 34.732 1.847 34.818 2.03 ;
      RECT 34.646 1.846 34.732 2.03 ;
      RECT 34.56 1.845 34.646 2.031 ;
      RECT 34.51 1.845 34.56 2.032 ;
      RECT 34.496 1.846 34.51 2.032 ;
      RECT 34.41 1.853 34.496 2.033 ;
      RECT 34.336 1.864 34.41 2.034 ;
      RECT 34.25 1.873 34.336 2.035 ;
      RECT 34.215 1.88 34.25 2.05 ;
      RECT 34.19 1.883 34.215 2.08 ;
      RECT 34.165 1.892 34.19 2.109 ;
      RECT 34.155 1.903 34.165 2.129 ;
      RECT 34.145 1.911 34.155 2.143 ;
      RECT 34.14 1.917 34.145 2.153 ;
      RECT 34.115 1.934 34.14 2.17 ;
      RECT 34.1 1.956 34.115 2.198 ;
      RECT 34.07 1.982 34.1 2.228 ;
      RECT 34.05 2.011 34.07 2.258 ;
      RECT 34.045 2.026 34.05 2.275 ;
      RECT 34.025 2.041 34.045 2.29 ;
      RECT 34.015 2.059 34.025 2.308 ;
      RECT 34.005 2.07 34.015 2.323 ;
      RECT 33.955 2.102 34.005 2.349 ;
      RECT 33.95 2.132 33.955 2.369 ;
      RECT 33.94 2.145 33.95 2.375 ;
      RECT 33.931 2.155 33.94 2.383 ;
      RECT 33.92 2.166 33.931 2.391 ;
      RECT 33.915 2.176 33.92 2.397 ;
      RECT 33.9 2.197 33.915 2.404 ;
      RECT 33.885 2.227 33.9 2.412 ;
      RECT 33.85 2.257 33.885 2.418 ;
      RECT 33.825 2.275 33.85 2.425 ;
      RECT 33.775 2.283 33.825 2.434 ;
      RECT 33.75 2.288 33.775 2.443 ;
      RECT 33.695 2.294 33.75 2.453 ;
      RECT 33.69 2.299 33.695 2.461 ;
      RECT 33.676 2.302 33.69 2.463 ;
      RECT 33.59 2.314 33.676 2.475 ;
      RECT 33.58 2.326 33.59 2.488 ;
      RECT 33.495 2.339 33.58 2.5 ;
      RECT 33.451 2.356 33.495 2.514 ;
      RECT 33.365 2.373 33.451 2.53 ;
      RECT 33.335 2.387 33.365 2.544 ;
      RECT 33.325 2.392 33.335 2.549 ;
      RECT 33.265 2.395 33.325 2.558 ;
      RECT 36.155 2.665 36.415 2.925 ;
      RECT 36.155 2.665 36.435 2.778 ;
      RECT 36.155 2.665 36.46 2.745 ;
      RECT 36.155 2.665 36.465 2.725 ;
      RECT 36.205 2.44 36.485 2.72 ;
      RECT 35.76 3.175 36.02 3.435 ;
      RECT 35.75 3.032 35.945 3.373 ;
      RECT 35.745 3.14 35.96 3.365 ;
      RECT 35.74 3.19 36.02 3.355 ;
      RECT 35.73 3.267 36.02 3.34 ;
      RECT 35.75 3.115 35.96 3.373 ;
      RECT 35.76 2.99 35.945 3.435 ;
      RECT 35.76 2.885 35.925 3.435 ;
      RECT 35.77 2.872 35.925 3.435 ;
      RECT 35.77 2.83 35.915 3.435 ;
      RECT 35.775 2.755 35.915 3.435 ;
      RECT 35.805 2.405 35.915 3.435 ;
      RECT 35.81 2.135 35.935 2.758 ;
      RECT 35.78 2.71 35.935 2.758 ;
      RECT 35.795 2.512 35.915 3.435 ;
      RECT 35.785 2.622 35.935 2.758 ;
      RECT 35.81 2.135 35.95 2.615 ;
      RECT 35.81 2.135 35.97 2.49 ;
      RECT 35.775 2.135 36.035 2.395 ;
      RECT 35.245 2.44 35.525 2.72 ;
      RECT 35.23 2.44 35.525 2.7 ;
      RECT 33.285 3.305 33.545 3.565 ;
      RECT 35.07 3.16 35.33 3.42 ;
      RECT 35.05 3.18 35.33 3.395 ;
      RECT 35.007 3.18 35.05 3.394 ;
      RECT 34.921 3.181 35.007 3.391 ;
      RECT 34.835 3.182 34.921 3.387 ;
      RECT 34.76 3.184 34.835 3.384 ;
      RECT 34.737 3.185 34.76 3.382 ;
      RECT 34.651 3.186 34.737 3.38 ;
      RECT 34.565 3.187 34.651 3.377 ;
      RECT 34.541 3.188 34.565 3.375 ;
      RECT 34.455 3.19 34.541 3.372 ;
      RECT 34.37 3.192 34.455 3.373 ;
      RECT 34.313 3.193 34.37 3.379 ;
      RECT 34.227 3.195 34.313 3.389 ;
      RECT 34.141 3.198 34.227 3.402 ;
      RECT 34.055 3.2 34.141 3.414 ;
      RECT 34.041 3.201 34.055 3.421 ;
      RECT 33.955 3.202 34.041 3.429 ;
      RECT 33.915 3.204 33.955 3.438 ;
      RECT 33.906 3.205 33.915 3.441 ;
      RECT 33.82 3.213 33.906 3.447 ;
      RECT 33.8 3.222 33.82 3.455 ;
      RECT 33.715 3.237 33.8 3.463 ;
      RECT 33.655 3.26 33.715 3.474 ;
      RECT 33.645 3.272 33.655 3.479 ;
      RECT 33.605 3.282 33.645 3.483 ;
      RECT 33.55 3.299 33.605 3.491 ;
      RECT 33.545 3.309 33.55 3.495 ;
      RECT 34.611 2.44 34.67 2.837 ;
      RECT 34.525 2.44 34.73 2.828 ;
      RECT 34.52 2.47 34.73 2.823 ;
      RECT 34.486 2.47 34.73 2.821 ;
      RECT 34.4 2.47 34.73 2.815 ;
      RECT 34.355 2.47 34.75 2.793 ;
      RECT 34.355 2.47 34.77 2.748 ;
      RECT 34.315 2.47 34.77 2.738 ;
      RECT 34.525 2.44 34.805 2.72 ;
      RECT 34.26 2.44 34.52 2.7 ;
      RECT 33.445 1.92 33.705 2.18 ;
      RECT 33.525 1.88 33.805 2.16 ;
      RECT 27.9 6.22 28.22 6.545 ;
      RECT 27.93 5.695 28.1 6.545 ;
      RECT 27.93 5.695 28.105 6.045 ;
      RECT 27.93 5.695 28.905 5.87 ;
      RECT 28.73 1.965 28.905 5.87 ;
      RECT 28.675 1.965 29.025 2.315 ;
      RECT 28.7 6.655 29.025 6.98 ;
      RECT 27.585 6.745 29.025 6.915 ;
      RECT 27.585 2.395 27.745 6.915 ;
      RECT 27.9 2.365 28.22 2.685 ;
      RECT 27.585 2.395 28.22 2.565 ;
      RECT 26.85 5.855 27.2 6.205 ;
      RECT 26.92 2.705 27.095 6.205 ;
      RECT 26.845 2.705 27.195 3.055 ;
      RECT 16.31 3 16.59 3.28 ;
      RECT 16.28 3 16.59 3.265 ;
      RECT 16.275 3 16.59 3.263 ;
      RECT 16.27 1.33 16.44 3.257 ;
      RECT 16.265 2.967 16.535 3.25 ;
      RECT 16.26 3 16.59 3.243 ;
      RECT 16.23 2.97 16.535 3.23 ;
      RECT 16.23 2.997 16.555 3.23 ;
      RECT 16.23 2.987 16.55 3.23 ;
      RECT 16.23 2.972 16.545 3.23 ;
      RECT 16.27 2.962 16.535 3.257 ;
      RECT 16.27 2.957 16.525 3.257 ;
      RECT 16.27 2.956 16.51 3.257 ;
      RECT 26.24 1.34 26.59 1.69 ;
      RECT 26.235 1.34 26.59 1.595 ;
      RECT 16.27 1.33 26.48 1.5 ;
      RECT 25.915 2.85 26.285 3.22 ;
      RECT 26 2.235 26.17 3.22 ;
      RECT 22.02 2.455 22.255 2.715 ;
      RECT 25.165 2.235 25.33 2.495 ;
      RECT 25.07 2.225 25.085 2.495 ;
      RECT 25.165 2.235 26.17 2.415 ;
      RECT 23.67 1.795 23.71 1.935 ;
      RECT 25.085 2.23 25.165 2.495 ;
      RECT 25.03 2.225 25.07 2.461 ;
      RECT 25.016 2.225 25.03 2.461 ;
      RECT 24.93 2.23 25.016 2.463 ;
      RECT 24.885 2.237 24.93 2.465 ;
      RECT 24.855 2.237 24.885 2.467 ;
      RECT 24.83 2.232 24.855 2.469 ;
      RECT 24.8 2.228 24.83 2.478 ;
      RECT 24.79 2.225 24.8 2.49 ;
      RECT 24.785 2.225 24.79 2.498 ;
      RECT 24.78 2.225 24.785 2.503 ;
      RECT 24.77 2.224 24.78 2.513 ;
      RECT 24.765 2.223 24.77 2.523 ;
      RECT 24.75 2.222 24.765 2.528 ;
      RECT 24.722 2.219 24.75 2.555 ;
      RECT 24.636 2.211 24.722 2.555 ;
      RECT 24.55 2.2 24.636 2.555 ;
      RECT 24.51 2.185 24.55 2.555 ;
      RECT 24.47 2.159 24.51 2.555 ;
      RECT 24.465 2.141 24.47 2.367 ;
      RECT 24.455 2.137 24.465 2.357 ;
      RECT 24.44 2.127 24.455 2.344 ;
      RECT 24.42 2.111 24.44 2.329 ;
      RECT 24.405 2.096 24.42 2.314 ;
      RECT 24.395 2.085 24.405 2.304 ;
      RECT 24.37 2.069 24.395 2.293 ;
      RECT 24.365 2.056 24.37 2.283 ;
      RECT 24.36 2.052 24.365 2.278 ;
      RECT 24.305 2.038 24.36 2.256 ;
      RECT 24.266 2.019 24.305 2.22 ;
      RECT 24.18 1.993 24.266 2.173 ;
      RECT 24.176 1.975 24.18 2.139 ;
      RECT 24.09 1.956 24.176 2.117 ;
      RECT 24.085 1.938 24.09 2.095 ;
      RECT 24.08 1.936 24.085 2.093 ;
      RECT 24.07 1.935 24.08 2.088 ;
      RECT 24.01 1.922 24.07 2.074 ;
      RECT 23.965 1.9 24.01 2.053 ;
      RECT 23.905 1.877 23.965 2.032 ;
      RECT 23.841 1.852 23.905 2.007 ;
      RECT 23.755 1.822 23.841 1.976 ;
      RECT 23.74 1.802 23.755 1.955 ;
      RECT 23.71 1.797 23.74 1.946 ;
      RECT 23.657 1.795 23.67 1.935 ;
      RECT 23.571 1.795 23.657 1.937 ;
      RECT 23.485 1.795 23.571 1.939 ;
      RECT 23.465 1.795 23.485 1.943 ;
      RECT 23.42 1.797 23.465 1.954 ;
      RECT 23.38 1.807 23.42 1.97 ;
      RECT 23.376 1.816 23.38 1.978 ;
      RECT 23.29 1.836 23.376 1.994 ;
      RECT 23.28 1.855 23.29 2.012 ;
      RECT 23.275 1.857 23.28 2.015 ;
      RECT 23.265 1.861 23.275 2.018 ;
      RECT 23.245 1.866 23.265 2.028 ;
      RECT 23.215 1.876 23.245 2.048 ;
      RECT 23.21 1.883 23.215 2.062 ;
      RECT 23.2 1.887 23.21 2.069 ;
      RECT 23.185 1.895 23.2 2.08 ;
      RECT 23.175 1.905 23.185 2.091 ;
      RECT 23.165 1.912 23.175 2.099 ;
      RECT 23.14 1.925 23.165 2.114 ;
      RECT 23.076 1.961 23.14 2.153 ;
      RECT 22.99 2.024 23.076 2.217 ;
      RECT 22.955 2.075 22.99 2.27 ;
      RECT 22.95 2.092 22.955 2.287 ;
      RECT 22.935 2.101 22.95 2.294 ;
      RECT 22.915 2.116 22.935 2.308 ;
      RECT 22.91 2.127 22.915 2.318 ;
      RECT 22.89 2.14 22.91 2.328 ;
      RECT 22.885 2.15 22.89 2.338 ;
      RECT 22.87 2.155 22.885 2.347 ;
      RECT 22.86 2.165 22.87 2.358 ;
      RECT 22.83 2.182 22.86 2.375 ;
      RECT 22.82 2.2 22.83 2.393 ;
      RECT 22.805 2.211 22.82 2.404 ;
      RECT 22.765 2.235 22.805 2.42 ;
      RECT 22.73 2.269 22.765 2.437 ;
      RECT 22.7 2.292 22.73 2.449 ;
      RECT 22.685 2.302 22.7 2.458 ;
      RECT 22.645 2.312 22.685 2.469 ;
      RECT 22.625 2.323 22.645 2.481 ;
      RECT 22.62 2.327 22.625 2.488 ;
      RECT 22.605 2.331 22.62 2.493 ;
      RECT 22.595 2.336 22.605 2.498 ;
      RECT 22.59 2.339 22.595 2.501 ;
      RECT 22.56 2.345 22.59 2.508 ;
      RECT 22.525 2.355 22.56 2.522 ;
      RECT 22.465 2.37 22.525 2.542 ;
      RECT 22.41 2.39 22.465 2.566 ;
      RECT 22.381 2.405 22.41 2.584 ;
      RECT 22.295 2.425 22.381 2.609 ;
      RECT 22.29 2.44 22.295 2.629 ;
      RECT 22.28 2.443 22.29 2.63 ;
      RECT 22.255 2.45 22.28 2.715 ;
      RECT 24.95 2.943 25.23 3.28 ;
      RECT 24.95 2.953 25.235 3.238 ;
      RECT 24.95 2.962 25.24 3.135 ;
      RECT 24.95 2.977 25.245 3.003 ;
      RECT 24.95 2.805 25.21 3.28 ;
      RECT 15.3 6.655 15.65 7.005 ;
      RECT 24.125 6.61 24.475 6.96 ;
      RECT 15.3 6.685 24.475 6.885 ;
      RECT 22.67 3.685 22.68 3.875 ;
      RECT 20.93 3.56 21.21 3.84 ;
      RECT 23.975 2.5 23.98 2.985 ;
      RECT 23.87 2.5 23.93 2.76 ;
      RECT 24.195 3.47 24.2 3.545 ;
      RECT 24.185 3.337 24.195 3.58 ;
      RECT 24.175 3.172 24.185 3.601 ;
      RECT 24.17 3.042 24.175 3.617 ;
      RECT 24.16 2.932 24.17 3.633 ;
      RECT 24.155 2.831 24.16 3.65 ;
      RECT 24.15 2.813 24.155 3.66 ;
      RECT 24.145 2.795 24.15 3.67 ;
      RECT 24.135 2.77 24.145 3.685 ;
      RECT 24.13 2.75 24.135 3.7 ;
      RECT 24.11 2.5 24.13 3.725 ;
      RECT 24.095 2.5 24.11 3.758 ;
      RECT 24.065 2.5 24.095 3.78 ;
      RECT 24.045 2.5 24.065 3.794 ;
      RECT 24.025 2.5 24.045 3.31 ;
      RECT 24.04 3.377 24.045 3.799 ;
      RECT 24.035 3.407 24.04 3.801 ;
      RECT 24.03 3.42 24.035 3.804 ;
      RECT 24.025 3.43 24.03 3.808 ;
      RECT 24.02 2.5 24.025 3.228 ;
      RECT 24.02 3.44 24.025 3.81 ;
      RECT 24.015 2.5 24.02 3.205 ;
      RECT 24.005 3.462 24.02 3.81 ;
      RECT 24 2.5 24.015 3.15 ;
      RECT 23.995 3.487 24.005 3.81 ;
      RECT 23.995 2.5 24 3.095 ;
      RECT 23.985 2.5 23.995 3.043 ;
      RECT 23.99 3.5 23.995 3.811 ;
      RECT 23.985 3.512 23.99 3.812 ;
      RECT 23.98 2.5 23.985 3.003 ;
      RECT 23.98 3.525 23.985 3.813 ;
      RECT 23.965 3.54 23.98 3.814 ;
      RECT 23.97 2.5 23.975 2.965 ;
      RECT 23.965 2.5 23.97 2.93 ;
      RECT 23.96 2.5 23.965 2.905 ;
      RECT 23.955 3.567 23.965 3.816 ;
      RECT 23.95 2.5 23.96 2.863 ;
      RECT 23.95 3.585 23.955 3.817 ;
      RECT 23.945 2.5 23.95 2.823 ;
      RECT 23.945 3.592 23.95 3.818 ;
      RECT 23.94 2.5 23.945 2.795 ;
      RECT 23.935 3.61 23.945 3.819 ;
      RECT 23.93 2.5 23.94 2.775 ;
      RECT 23.925 3.63 23.935 3.821 ;
      RECT 23.915 3.647 23.925 3.822 ;
      RECT 23.88 3.67 23.915 3.825 ;
      RECT 23.825 3.688 23.88 3.831 ;
      RECT 23.739 3.696 23.825 3.84 ;
      RECT 23.653 3.707 23.739 3.851 ;
      RECT 23.567 3.717 23.653 3.862 ;
      RECT 23.481 3.727 23.567 3.874 ;
      RECT 23.395 3.737 23.481 3.885 ;
      RECT 23.375 3.743 23.395 3.891 ;
      RECT 23.295 3.745 23.375 3.895 ;
      RECT 23.29 3.744 23.295 3.9 ;
      RECT 23.282 3.743 23.29 3.9 ;
      RECT 23.196 3.739 23.282 3.898 ;
      RECT 23.11 3.731 23.196 3.895 ;
      RECT 23.024 3.722 23.11 3.891 ;
      RECT 22.938 3.714 23.024 3.888 ;
      RECT 22.852 3.706 22.938 3.884 ;
      RECT 22.766 3.697 22.852 3.881 ;
      RECT 22.68 3.689 22.766 3.877 ;
      RECT 22.625 3.682 22.67 3.875 ;
      RECT 22.54 3.675 22.625 3.873 ;
      RECT 22.466 3.667 22.54 3.869 ;
      RECT 22.38 3.659 22.466 3.866 ;
      RECT 22.377 3.655 22.38 3.864 ;
      RECT 22.291 3.651 22.377 3.863 ;
      RECT 22.205 3.643 22.291 3.86 ;
      RECT 22.12 3.638 22.205 3.857 ;
      RECT 22.034 3.635 22.12 3.854 ;
      RECT 21.948 3.633 22.034 3.851 ;
      RECT 21.862 3.63 21.948 3.848 ;
      RECT 21.776 3.627 21.862 3.845 ;
      RECT 21.69 3.624 21.776 3.842 ;
      RECT 21.614 3.622 21.69 3.839 ;
      RECT 21.528 3.619 21.614 3.836 ;
      RECT 21.442 3.616 21.528 3.834 ;
      RECT 21.356 3.614 21.442 3.831 ;
      RECT 21.27 3.611 21.356 3.828 ;
      RECT 21.21 3.602 21.27 3.826 ;
      RECT 23.72 3.22 23.795 3.48 ;
      RECT 23.7 3.2 23.705 3.48 ;
      RECT 23.02 2.985 23.125 3.28 ;
      RECT 17.465 2.96 17.535 3.22 ;
      RECT 23.36 2.835 23.365 3.206 ;
      RECT 23.35 2.89 23.355 3.206 ;
      RECT 23.655 2.06 23.715 2.32 ;
      RECT 23.71 3.215 23.72 3.48 ;
      RECT 23.705 3.205 23.71 3.48 ;
      RECT 23.625 3.152 23.7 3.48 ;
      RECT 23.65 2.06 23.655 2.34 ;
      RECT 23.64 2.06 23.65 2.36 ;
      RECT 23.625 2.06 23.64 2.39 ;
      RECT 23.61 2.06 23.625 2.433 ;
      RECT 23.605 3.095 23.625 3.48 ;
      RECT 23.595 2.06 23.61 2.47 ;
      RECT 23.59 3.075 23.605 3.48 ;
      RECT 23.59 2.06 23.595 2.493 ;
      RECT 23.58 2.06 23.59 2.518 ;
      RECT 23.55 3.042 23.59 3.48 ;
      RECT 23.555 2.06 23.58 2.568 ;
      RECT 23.55 2.06 23.555 2.623 ;
      RECT 23.545 2.06 23.55 2.665 ;
      RECT 23.535 3.005 23.55 3.48 ;
      RECT 23.54 2.06 23.545 2.708 ;
      RECT 23.535 2.06 23.54 2.773 ;
      RECT 23.53 2.06 23.535 2.795 ;
      RECT 23.53 2.993 23.535 3.345 ;
      RECT 23.525 2.06 23.53 2.863 ;
      RECT 23.525 2.985 23.53 3.328 ;
      RECT 23.52 2.06 23.525 2.908 ;
      RECT 23.515 2.967 23.525 3.305 ;
      RECT 23.515 2.06 23.52 2.945 ;
      RECT 23.505 2.06 23.515 3.285 ;
      RECT 23.5 2.06 23.505 3.268 ;
      RECT 23.495 2.06 23.5 3.253 ;
      RECT 23.49 2.06 23.495 3.238 ;
      RECT 23.47 2.06 23.49 3.228 ;
      RECT 23.465 2.06 23.47 3.218 ;
      RECT 23.455 2.06 23.465 3.214 ;
      RECT 23.45 2.337 23.455 3.213 ;
      RECT 23.445 2.36 23.45 3.212 ;
      RECT 23.44 2.39 23.445 3.211 ;
      RECT 23.435 2.417 23.44 3.21 ;
      RECT 23.43 2.445 23.435 3.21 ;
      RECT 23.425 2.472 23.43 3.21 ;
      RECT 23.42 2.492 23.425 3.21 ;
      RECT 23.415 2.52 23.42 3.21 ;
      RECT 23.405 2.562 23.415 3.21 ;
      RECT 23.395 2.607 23.405 3.209 ;
      RECT 23.39 2.66 23.395 3.208 ;
      RECT 23.385 2.692 23.39 3.207 ;
      RECT 23.38 2.712 23.385 3.206 ;
      RECT 23.375 2.75 23.38 3.206 ;
      RECT 23.37 2.772 23.375 3.206 ;
      RECT 23.365 2.797 23.37 3.206 ;
      RECT 23.355 2.862 23.36 3.206 ;
      RECT 23.34 2.922 23.35 3.206 ;
      RECT 23.325 2.932 23.34 3.206 ;
      RECT 23.305 2.942 23.325 3.206 ;
      RECT 23.275 2.947 23.305 3.203 ;
      RECT 23.215 2.957 23.275 3.2 ;
      RECT 23.195 2.966 23.215 3.205 ;
      RECT 23.17 2.972 23.195 3.218 ;
      RECT 23.15 2.977 23.17 3.233 ;
      RECT 23.125 2.982 23.15 3.28 ;
      RECT 22.996 2.984 23.02 3.28 ;
      RECT 22.91 2.979 22.996 3.28 ;
      RECT 22.87 2.976 22.91 3.28 ;
      RECT 22.82 2.978 22.87 3.26 ;
      RECT 22.79 2.982 22.82 3.26 ;
      RECT 22.711 2.992 22.79 3.26 ;
      RECT 22.625 3.007 22.711 3.261 ;
      RECT 22.575 3.017 22.625 3.262 ;
      RECT 22.567 3.02 22.575 3.262 ;
      RECT 22.481 3.022 22.567 3.263 ;
      RECT 22.395 3.026 22.481 3.263 ;
      RECT 22.309 3.03 22.395 3.264 ;
      RECT 22.223 3.033 22.309 3.265 ;
      RECT 22.137 3.037 22.223 3.265 ;
      RECT 22.051 3.041 22.137 3.266 ;
      RECT 21.965 3.044 22.051 3.267 ;
      RECT 21.879 3.048 21.965 3.267 ;
      RECT 21.793 3.052 21.879 3.268 ;
      RECT 21.707 3.056 21.793 3.269 ;
      RECT 21.621 3.059 21.707 3.269 ;
      RECT 21.535 3.063 21.621 3.27 ;
      RECT 21.505 3.065 21.535 3.27 ;
      RECT 21.419 3.068 21.505 3.271 ;
      RECT 21.333 3.072 21.419 3.272 ;
      RECT 21.247 3.076 21.333 3.273 ;
      RECT 21.161 3.079 21.247 3.273 ;
      RECT 21.075 3.083 21.161 3.274 ;
      RECT 21.04 3.088 21.075 3.275 ;
      RECT 20.985 3.098 21.04 3.282 ;
      RECT 20.96 3.11 20.985 3.292 ;
      RECT 20.925 3.123 20.96 3.3 ;
      RECT 20.885 3.14 20.925 3.323 ;
      RECT 20.865 3.153 20.885 3.35 ;
      RECT 20.835 3.165 20.865 3.378 ;
      RECT 20.83 3.173 20.835 3.398 ;
      RECT 20.825 3.176 20.83 3.408 ;
      RECT 20.775 3.188 20.825 3.442 ;
      RECT 20.765 3.203 20.775 3.475 ;
      RECT 20.755 3.209 20.765 3.488 ;
      RECT 20.745 3.216 20.755 3.5 ;
      RECT 20.72 3.229 20.745 3.518 ;
      RECT 20.705 3.244 20.72 3.54 ;
      RECT 20.695 3.252 20.705 3.556 ;
      RECT 20.68 3.261 20.695 3.571 ;
      RECT 20.67 3.271 20.68 3.585 ;
      RECT 20.651 3.284 20.67 3.602 ;
      RECT 20.565 3.329 20.651 3.667 ;
      RECT 20.55 3.374 20.565 3.725 ;
      RECT 20.545 3.383 20.55 3.738 ;
      RECT 20.535 3.39 20.545 3.743 ;
      RECT 20.53 3.395 20.535 3.747 ;
      RECT 20.51 3.405 20.53 3.754 ;
      RECT 20.485 3.425 20.51 3.768 ;
      RECT 20.45 3.45 20.485 3.788 ;
      RECT 20.435 3.473 20.45 3.803 ;
      RECT 20.425 3.483 20.435 3.808 ;
      RECT 20.415 3.491 20.425 3.815 ;
      RECT 20.405 3.5 20.415 3.821 ;
      RECT 20.385 3.512 20.405 3.823 ;
      RECT 20.375 3.525 20.385 3.825 ;
      RECT 20.35 3.54 20.375 3.828 ;
      RECT 20.33 3.557 20.35 3.832 ;
      RECT 20.29 3.585 20.33 3.838 ;
      RECT 20.225 3.632 20.29 3.847 ;
      RECT 20.21 3.665 20.225 3.855 ;
      RECT 20.205 3.672 20.21 3.857 ;
      RECT 20.155 3.697 20.205 3.862 ;
      RECT 20.14 3.721 20.155 3.869 ;
      RECT 20.09 3.726 20.14 3.87 ;
      RECT 20.004 3.73 20.09 3.87 ;
      RECT 19.918 3.73 20.004 3.87 ;
      RECT 19.832 3.73 19.918 3.871 ;
      RECT 19.746 3.73 19.832 3.871 ;
      RECT 19.66 3.73 19.746 3.871 ;
      RECT 19.594 3.73 19.66 3.871 ;
      RECT 19.508 3.73 19.594 3.872 ;
      RECT 19.422 3.73 19.508 3.872 ;
      RECT 19.336 3.731 19.422 3.873 ;
      RECT 19.25 3.731 19.336 3.873 ;
      RECT 19.164 3.731 19.25 3.873 ;
      RECT 19.078 3.731 19.164 3.874 ;
      RECT 18.992 3.731 19.078 3.874 ;
      RECT 18.906 3.732 18.992 3.875 ;
      RECT 18.82 3.732 18.906 3.875 ;
      RECT 18.8 3.732 18.82 3.875 ;
      RECT 18.714 3.732 18.8 3.875 ;
      RECT 18.628 3.732 18.714 3.875 ;
      RECT 18.542 3.733 18.628 3.875 ;
      RECT 18.456 3.733 18.542 3.875 ;
      RECT 18.37 3.733 18.456 3.875 ;
      RECT 18.284 3.734 18.37 3.875 ;
      RECT 18.198 3.734 18.284 3.875 ;
      RECT 18.112 3.734 18.198 3.875 ;
      RECT 18.026 3.734 18.112 3.875 ;
      RECT 17.94 3.735 18.026 3.875 ;
      RECT 17.89 3.732 17.94 3.875 ;
      RECT 17.88 3.73 17.89 3.874 ;
      RECT 17.876 3.73 17.88 3.873 ;
      RECT 17.79 3.725 17.876 3.868 ;
      RECT 17.768 3.718 17.79 3.862 ;
      RECT 17.682 3.709 17.768 3.856 ;
      RECT 17.596 3.696 17.682 3.847 ;
      RECT 17.51 3.682 17.596 3.837 ;
      RECT 17.465 3.672 17.51 3.83 ;
      RECT 17.445 2.96 17.465 3.238 ;
      RECT 17.445 3.665 17.465 3.826 ;
      RECT 17.415 2.96 17.445 3.26 ;
      RECT 17.405 3.632 17.445 3.823 ;
      RECT 17.4 2.96 17.415 3.28 ;
      RECT 17.4 3.597 17.405 3.821 ;
      RECT 17.395 2.96 17.4 3.405 ;
      RECT 17.395 3.557 17.4 3.821 ;
      RECT 17.385 2.96 17.395 3.821 ;
      RECT 17.31 2.96 17.385 3.815 ;
      RECT 17.28 2.96 17.31 3.805 ;
      RECT 17.275 2.96 17.28 3.797 ;
      RECT 17.27 3.002 17.275 3.79 ;
      RECT 17.26 3.071 17.27 3.781 ;
      RECT 17.255 3.141 17.26 3.733 ;
      RECT 17.25 3.205 17.255 3.63 ;
      RECT 17.245 3.24 17.25 3.585 ;
      RECT 17.243 3.277 17.245 3.477 ;
      RECT 17.24 3.285 17.243 3.47 ;
      RECT 17.235 3.35 17.24 3.413 ;
      RECT 21.31 2.44 21.59 2.72 ;
      RECT 21.3 2.44 21.59 2.583 ;
      RECT 21.255 2.305 21.515 2.565 ;
      RECT 21.255 2.42 21.57 2.565 ;
      RECT 21.255 2.39 21.565 2.565 ;
      RECT 21.255 2.377 21.555 2.565 ;
      RECT 21.255 2.367 21.55 2.565 ;
      RECT 17.23 2.35 17.49 2.61 ;
      RECT 21 1.9 21.26 2.16 ;
      RECT 20.99 1.925 21.26 2.12 ;
      RECT 20.985 1.925 20.99 2.119 ;
      RECT 20.915 1.92 20.985 2.111 ;
      RECT 20.83 1.907 20.915 2.094 ;
      RECT 20.826 1.899 20.83 2.084 ;
      RECT 20.74 1.892 20.826 2.074 ;
      RECT 20.731 1.884 20.74 2.064 ;
      RECT 20.645 1.877 20.731 2.052 ;
      RECT 20.625 1.868 20.645 2.038 ;
      RECT 20.57 1.863 20.625 2.03 ;
      RECT 20.56 1.857 20.57 2.024 ;
      RECT 20.54 1.855 20.56 2.02 ;
      RECT 20.532 1.854 20.54 2.016 ;
      RECT 20.446 1.846 20.532 2.005 ;
      RECT 20.36 1.832 20.446 1.985 ;
      RECT 20.3 1.82 20.36 1.97 ;
      RECT 20.29 1.815 20.3 1.965 ;
      RECT 20.24 1.815 20.29 1.967 ;
      RECT 20.193 1.817 20.24 1.971 ;
      RECT 20.107 1.824 20.193 1.976 ;
      RECT 20.021 1.832 20.107 1.982 ;
      RECT 19.935 1.841 20.021 1.988 ;
      RECT 19.876 1.847 19.935 1.993 ;
      RECT 19.79 1.852 19.876 1.999 ;
      RECT 19.715 1.857 19.79 2.005 ;
      RECT 19.676 1.859 19.715 2.01 ;
      RECT 19.59 1.856 19.676 2.015 ;
      RECT 19.505 1.854 19.59 2.022 ;
      RECT 19.473 1.853 19.505 2.025 ;
      RECT 19.387 1.852 19.473 2.026 ;
      RECT 19.301 1.851 19.387 2.027 ;
      RECT 19.215 1.85 19.301 2.027 ;
      RECT 19.129 1.849 19.215 2.028 ;
      RECT 19.043 1.848 19.129 2.029 ;
      RECT 18.957 1.847 19.043 2.03 ;
      RECT 18.871 1.846 18.957 2.03 ;
      RECT 18.785 1.845 18.871 2.031 ;
      RECT 18.735 1.845 18.785 2.032 ;
      RECT 18.721 1.846 18.735 2.032 ;
      RECT 18.635 1.853 18.721 2.033 ;
      RECT 18.561 1.864 18.635 2.034 ;
      RECT 18.475 1.873 18.561 2.035 ;
      RECT 18.44 1.88 18.475 2.05 ;
      RECT 18.415 1.883 18.44 2.08 ;
      RECT 18.39 1.892 18.415 2.109 ;
      RECT 18.38 1.903 18.39 2.129 ;
      RECT 18.37 1.911 18.38 2.143 ;
      RECT 18.365 1.917 18.37 2.153 ;
      RECT 18.34 1.934 18.365 2.17 ;
      RECT 18.325 1.956 18.34 2.198 ;
      RECT 18.295 1.982 18.325 2.228 ;
      RECT 18.275 2.011 18.295 2.258 ;
      RECT 18.27 2.026 18.275 2.275 ;
      RECT 18.25 2.041 18.27 2.29 ;
      RECT 18.24 2.059 18.25 2.308 ;
      RECT 18.23 2.07 18.24 2.323 ;
      RECT 18.18 2.102 18.23 2.349 ;
      RECT 18.175 2.132 18.18 2.369 ;
      RECT 18.165 2.145 18.175 2.375 ;
      RECT 18.156 2.155 18.165 2.383 ;
      RECT 18.145 2.166 18.156 2.391 ;
      RECT 18.14 2.176 18.145 2.397 ;
      RECT 18.125 2.197 18.14 2.404 ;
      RECT 18.11 2.227 18.125 2.412 ;
      RECT 18.075 2.257 18.11 2.418 ;
      RECT 18.05 2.275 18.075 2.425 ;
      RECT 18 2.283 18.05 2.434 ;
      RECT 17.975 2.288 18 2.443 ;
      RECT 17.92 2.294 17.975 2.453 ;
      RECT 17.915 2.299 17.92 2.461 ;
      RECT 17.901 2.302 17.915 2.463 ;
      RECT 17.815 2.314 17.901 2.475 ;
      RECT 17.805 2.326 17.815 2.488 ;
      RECT 17.72 2.339 17.805 2.5 ;
      RECT 17.676 2.356 17.72 2.514 ;
      RECT 17.59 2.373 17.676 2.53 ;
      RECT 17.56 2.387 17.59 2.544 ;
      RECT 17.55 2.392 17.56 2.549 ;
      RECT 17.49 2.395 17.55 2.558 ;
      RECT 20.38 2.665 20.64 2.925 ;
      RECT 20.38 2.665 20.66 2.778 ;
      RECT 20.38 2.665 20.685 2.745 ;
      RECT 20.38 2.665 20.69 2.725 ;
      RECT 20.43 2.44 20.71 2.72 ;
      RECT 19.985 3.175 20.245 3.435 ;
      RECT 19.975 3.032 20.17 3.373 ;
      RECT 19.97 3.14 20.185 3.365 ;
      RECT 19.965 3.19 20.245 3.355 ;
      RECT 19.955 3.267 20.245 3.34 ;
      RECT 19.975 3.115 20.185 3.373 ;
      RECT 19.985 2.99 20.17 3.435 ;
      RECT 19.985 2.885 20.15 3.435 ;
      RECT 19.995 2.872 20.15 3.435 ;
      RECT 19.995 2.83 20.14 3.435 ;
      RECT 20 2.755 20.14 3.435 ;
      RECT 20.03 2.405 20.14 3.435 ;
      RECT 20.035 2.135 20.16 2.758 ;
      RECT 20.005 2.71 20.16 2.758 ;
      RECT 20.02 2.512 20.14 3.435 ;
      RECT 20.01 2.622 20.16 2.758 ;
      RECT 20.035 2.135 20.175 2.615 ;
      RECT 20.035 2.135 20.195 2.49 ;
      RECT 20 2.135 20.26 2.395 ;
      RECT 19.47 2.44 19.75 2.72 ;
      RECT 19.455 2.44 19.75 2.7 ;
      RECT 17.51 3.305 17.77 3.565 ;
      RECT 19.295 3.16 19.555 3.42 ;
      RECT 19.275 3.18 19.555 3.395 ;
      RECT 19.232 3.18 19.275 3.394 ;
      RECT 19.146 3.181 19.232 3.391 ;
      RECT 19.06 3.182 19.146 3.387 ;
      RECT 18.985 3.184 19.06 3.384 ;
      RECT 18.962 3.185 18.985 3.382 ;
      RECT 18.876 3.186 18.962 3.38 ;
      RECT 18.79 3.187 18.876 3.377 ;
      RECT 18.766 3.188 18.79 3.375 ;
      RECT 18.68 3.19 18.766 3.372 ;
      RECT 18.595 3.192 18.68 3.373 ;
      RECT 18.538 3.193 18.595 3.379 ;
      RECT 18.452 3.195 18.538 3.389 ;
      RECT 18.366 3.198 18.452 3.402 ;
      RECT 18.28 3.2 18.366 3.414 ;
      RECT 18.266 3.201 18.28 3.421 ;
      RECT 18.18 3.202 18.266 3.429 ;
      RECT 18.14 3.204 18.18 3.438 ;
      RECT 18.131 3.205 18.14 3.441 ;
      RECT 18.045 3.213 18.131 3.447 ;
      RECT 18.025 3.222 18.045 3.455 ;
      RECT 17.94 3.237 18.025 3.463 ;
      RECT 17.88 3.26 17.94 3.474 ;
      RECT 17.87 3.272 17.88 3.479 ;
      RECT 17.83 3.282 17.87 3.483 ;
      RECT 17.775 3.299 17.83 3.491 ;
      RECT 17.77 3.309 17.775 3.495 ;
      RECT 18.836 2.44 18.895 2.837 ;
      RECT 18.75 2.44 18.955 2.828 ;
      RECT 18.745 2.47 18.955 2.823 ;
      RECT 18.711 2.47 18.955 2.821 ;
      RECT 18.625 2.47 18.955 2.815 ;
      RECT 18.58 2.47 18.975 2.793 ;
      RECT 18.58 2.47 18.995 2.748 ;
      RECT 18.54 2.47 18.995 2.738 ;
      RECT 18.75 2.44 19.03 2.72 ;
      RECT 18.485 2.44 18.745 2.7 ;
      RECT 17.67 1.92 17.93 2.18 ;
      RECT 17.75 1.88 18.03 2.16 ;
      RECT 12.12 6.22 12.44 6.545 ;
      RECT 12.15 5.695 12.32 6.545 ;
      RECT 12.15 5.695 12.325 6.045 ;
      RECT 12.15 5.695 13.125 5.87 ;
      RECT 12.95 1.965 13.125 5.87 ;
      RECT 12.895 1.965 13.245 2.315 ;
      RECT 12.92 6.655 13.245 6.98 ;
      RECT 11.805 6.745 13.245 6.915 ;
      RECT 11.805 2.395 11.965 6.915 ;
      RECT 12.12 2.365 12.44 2.685 ;
      RECT 11.805 2.395 12.44 2.565 ;
      RECT 11.07 5.855 11.42 6.205 ;
      RECT 11.14 2.705 11.315 6.205 ;
      RECT 11.065 2.705 11.415 3.055 ;
      RECT 0.53 3 0.81 3.28 ;
      RECT 0.5 3 0.81 3.265 ;
      RECT 0.495 3 0.81 3.263 ;
      RECT 0.49 1.33 0.66 3.257 ;
      RECT 0.485 2.967 0.755 3.25 ;
      RECT 0.48 3 0.81 3.243 ;
      RECT 0.45 2.97 0.755 3.23 ;
      RECT 0.45 2.997 0.775 3.23 ;
      RECT 0.45 2.987 0.77 3.23 ;
      RECT 0.45 2.972 0.765 3.23 ;
      RECT 0.49 2.962 0.755 3.257 ;
      RECT 0.49 2.957 0.745 3.257 ;
      RECT 0.49 2.956 0.73 3.257 ;
      RECT 10.46 1.34 10.81 1.69 ;
      RECT 10.455 1.34 10.81 1.595 ;
      RECT 0.49 1.33 10.7 1.5 ;
      RECT 10.135 2.85 10.505 3.22 ;
      RECT 10.22 2.235 10.39 3.22 ;
      RECT 6.24 2.455 6.475 2.715 ;
      RECT 9.385 2.235 9.55 2.495 ;
      RECT 9.29 2.225 9.305 2.495 ;
      RECT 9.385 2.235 10.39 2.415 ;
      RECT 7.89 1.795 7.93 1.935 ;
      RECT 9.305 2.23 9.385 2.495 ;
      RECT 9.25 2.225 9.29 2.461 ;
      RECT 9.236 2.225 9.25 2.461 ;
      RECT 9.15 2.23 9.236 2.463 ;
      RECT 9.105 2.237 9.15 2.465 ;
      RECT 9.075 2.237 9.105 2.467 ;
      RECT 9.05 2.232 9.075 2.469 ;
      RECT 9.02 2.228 9.05 2.478 ;
      RECT 9.01 2.225 9.02 2.49 ;
      RECT 9.005 2.225 9.01 2.498 ;
      RECT 9 2.225 9.005 2.503 ;
      RECT 8.99 2.224 9 2.513 ;
      RECT 8.985 2.223 8.99 2.523 ;
      RECT 8.97 2.222 8.985 2.528 ;
      RECT 8.942 2.219 8.97 2.555 ;
      RECT 8.856 2.211 8.942 2.555 ;
      RECT 8.77 2.2 8.856 2.555 ;
      RECT 8.73 2.185 8.77 2.555 ;
      RECT 8.69 2.159 8.73 2.555 ;
      RECT 8.685 2.141 8.69 2.367 ;
      RECT 8.675 2.137 8.685 2.357 ;
      RECT 8.66 2.127 8.675 2.344 ;
      RECT 8.64 2.111 8.66 2.329 ;
      RECT 8.625 2.096 8.64 2.314 ;
      RECT 8.615 2.085 8.625 2.304 ;
      RECT 8.59 2.069 8.615 2.293 ;
      RECT 8.585 2.056 8.59 2.283 ;
      RECT 8.58 2.052 8.585 2.278 ;
      RECT 8.525 2.038 8.58 2.256 ;
      RECT 8.486 2.019 8.525 2.22 ;
      RECT 8.4 1.993 8.486 2.173 ;
      RECT 8.396 1.975 8.4 2.139 ;
      RECT 8.31 1.956 8.396 2.117 ;
      RECT 8.305 1.938 8.31 2.095 ;
      RECT 8.3 1.936 8.305 2.093 ;
      RECT 8.29 1.935 8.3 2.088 ;
      RECT 8.23 1.922 8.29 2.074 ;
      RECT 8.185 1.9 8.23 2.053 ;
      RECT 8.125 1.877 8.185 2.032 ;
      RECT 8.061 1.852 8.125 2.007 ;
      RECT 7.975 1.822 8.061 1.976 ;
      RECT 7.96 1.802 7.975 1.955 ;
      RECT 7.93 1.797 7.96 1.946 ;
      RECT 7.877 1.795 7.89 1.935 ;
      RECT 7.791 1.795 7.877 1.937 ;
      RECT 7.705 1.795 7.791 1.939 ;
      RECT 7.685 1.795 7.705 1.943 ;
      RECT 7.64 1.797 7.685 1.954 ;
      RECT 7.6 1.807 7.64 1.97 ;
      RECT 7.596 1.816 7.6 1.978 ;
      RECT 7.51 1.836 7.596 1.994 ;
      RECT 7.5 1.855 7.51 2.012 ;
      RECT 7.495 1.857 7.5 2.015 ;
      RECT 7.485 1.861 7.495 2.018 ;
      RECT 7.465 1.866 7.485 2.028 ;
      RECT 7.435 1.876 7.465 2.048 ;
      RECT 7.43 1.883 7.435 2.062 ;
      RECT 7.42 1.887 7.43 2.069 ;
      RECT 7.405 1.895 7.42 2.08 ;
      RECT 7.395 1.905 7.405 2.091 ;
      RECT 7.385 1.912 7.395 2.099 ;
      RECT 7.36 1.925 7.385 2.114 ;
      RECT 7.296 1.961 7.36 2.153 ;
      RECT 7.21 2.024 7.296 2.217 ;
      RECT 7.175 2.075 7.21 2.27 ;
      RECT 7.17 2.092 7.175 2.287 ;
      RECT 7.155 2.101 7.17 2.294 ;
      RECT 7.135 2.116 7.155 2.308 ;
      RECT 7.13 2.127 7.135 2.318 ;
      RECT 7.11 2.14 7.13 2.328 ;
      RECT 7.105 2.15 7.11 2.338 ;
      RECT 7.09 2.155 7.105 2.347 ;
      RECT 7.08 2.165 7.09 2.358 ;
      RECT 7.05 2.182 7.08 2.375 ;
      RECT 7.04 2.2 7.05 2.393 ;
      RECT 7.025 2.211 7.04 2.404 ;
      RECT 6.985 2.235 7.025 2.42 ;
      RECT 6.95 2.269 6.985 2.437 ;
      RECT 6.92 2.292 6.95 2.449 ;
      RECT 6.905 2.302 6.92 2.458 ;
      RECT 6.865 2.312 6.905 2.469 ;
      RECT 6.845 2.323 6.865 2.481 ;
      RECT 6.84 2.327 6.845 2.488 ;
      RECT 6.825 2.331 6.84 2.493 ;
      RECT 6.815 2.336 6.825 2.498 ;
      RECT 6.81 2.339 6.815 2.501 ;
      RECT 6.78 2.345 6.81 2.508 ;
      RECT 6.745 2.355 6.78 2.522 ;
      RECT 6.685 2.37 6.745 2.542 ;
      RECT 6.63 2.39 6.685 2.566 ;
      RECT 6.601 2.405 6.63 2.584 ;
      RECT 6.515 2.425 6.601 2.609 ;
      RECT 6.51 2.44 6.515 2.629 ;
      RECT 6.5 2.443 6.51 2.63 ;
      RECT 6.475 2.45 6.5 2.715 ;
      RECT 9.17 2.943 9.45 3.28 ;
      RECT 9.17 2.953 9.455 3.238 ;
      RECT 9.17 2.962 9.46 3.135 ;
      RECT 9.17 2.977 9.465 3.003 ;
      RECT 9.17 2.805 9.43 3.28 ;
      RECT -1.25 6.995 -0.96 7.345 ;
      RECT -1.25 7.055 0.165 7.225 ;
      RECT -0.005 6.685 0.165 7.225 ;
      RECT 8.315 6.605 8.665 6.955 ;
      RECT -0.005 6.685 8.665 6.855 ;
      RECT 6.89 3.685 6.9 3.875 ;
      RECT 5.15 3.56 5.43 3.84 ;
      RECT 8.195 2.5 8.2 2.985 ;
      RECT 8.09 2.5 8.15 2.76 ;
      RECT 8.415 3.47 8.42 3.545 ;
      RECT 8.405 3.337 8.415 3.58 ;
      RECT 8.395 3.172 8.405 3.601 ;
      RECT 8.39 3.042 8.395 3.617 ;
      RECT 8.38 2.932 8.39 3.633 ;
      RECT 8.375 2.831 8.38 3.65 ;
      RECT 8.37 2.813 8.375 3.66 ;
      RECT 8.365 2.795 8.37 3.67 ;
      RECT 8.355 2.77 8.365 3.685 ;
      RECT 8.35 2.75 8.355 3.7 ;
      RECT 8.33 2.5 8.35 3.725 ;
      RECT 8.315 2.5 8.33 3.758 ;
      RECT 8.285 2.5 8.315 3.78 ;
      RECT 8.265 2.5 8.285 3.794 ;
      RECT 8.245 2.5 8.265 3.31 ;
      RECT 8.26 3.377 8.265 3.799 ;
      RECT 8.255 3.407 8.26 3.801 ;
      RECT 8.25 3.42 8.255 3.804 ;
      RECT 8.245 3.43 8.25 3.808 ;
      RECT 8.24 2.5 8.245 3.228 ;
      RECT 8.24 3.44 8.245 3.81 ;
      RECT 8.235 2.5 8.24 3.205 ;
      RECT 8.225 3.462 8.24 3.81 ;
      RECT 8.22 2.5 8.235 3.15 ;
      RECT 8.215 3.487 8.225 3.81 ;
      RECT 8.215 2.5 8.22 3.095 ;
      RECT 8.205 2.5 8.215 3.043 ;
      RECT 8.21 3.5 8.215 3.811 ;
      RECT 8.205 3.512 8.21 3.812 ;
      RECT 8.2 2.5 8.205 3.003 ;
      RECT 8.2 3.525 8.205 3.813 ;
      RECT 8.185 3.54 8.2 3.814 ;
      RECT 8.19 2.5 8.195 2.965 ;
      RECT 8.185 2.5 8.19 2.93 ;
      RECT 8.18 2.5 8.185 2.905 ;
      RECT 8.175 3.567 8.185 3.816 ;
      RECT 8.17 2.5 8.18 2.863 ;
      RECT 8.17 3.585 8.175 3.817 ;
      RECT 8.165 2.5 8.17 2.823 ;
      RECT 8.165 3.592 8.17 3.818 ;
      RECT 8.16 2.5 8.165 2.795 ;
      RECT 8.155 3.61 8.165 3.819 ;
      RECT 8.15 2.5 8.16 2.775 ;
      RECT 8.145 3.63 8.155 3.821 ;
      RECT 8.135 3.647 8.145 3.822 ;
      RECT 8.1 3.67 8.135 3.825 ;
      RECT 8.045 3.688 8.1 3.831 ;
      RECT 7.959 3.696 8.045 3.84 ;
      RECT 7.873 3.707 7.959 3.851 ;
      RECT 7.787 3.717 7.873 3.862 ;
      RECT 7.701 3.727 7.787 3.874 ;
      RECT 7.615 3.737 7.701 3.885 ;
      RECT 7.595 3.743 7.615 3.891 ;
      RECT 7.515 3.745 7.595 3.895 ;
      RECT 7.51 3.744 7.515 3.9 ;
      RECT 7.502 3.743 7.51 3.9 ;
      RECT 7.416 3.739 7.502 3.898 ;
      RECT 7.33 3.731 7.416 3.895 ;
      RECT 7.244 3.722 7.33 3.891 ;
      RECT 7.158 3.714 7.244 3.888 ;
      RECT 7.072 3.706 7.158 3.884 ;
      RECT 6.986 3.697 7.072 3.881 ;
      RECT 6.9 3.689 6.986 3.877 ;
      RECT 6.845 3.682 6.89 3.875 ;
      RECT 6.76 3.675 6.845 3.873 ;
      RECT 6.686 3.667 6.76 3.869 ;
      RECT 6.6 3.659 6.686 3.866 ;
      RECT 6.597 3.655 6.6 3.864 ;
      RECT 6.511 3.651 6.597 3.863 ;
      RECT 6.425 3.643 6.511 3.86 ;
      RECT 6.34 3.638 6.425 3.857 ;
      RECT 6.254 3.635 6.34 3.854 ;
      RECT 6.168 3.633 6.254 3.851 ;
      RECT 6.082 3.63 6.168 3.848 ;
      RECT 5.996 3.627 6.082 3.845 ;
      RECT 5.91 3.624 5.996 3.842 ;
      RECT 5.834 3.622 5.91 3.839 ;
      RECT 5.748 3.619 5.834 3.836 ;
      RECT 5.662 3.616 5.748 3.834 ;
      RECT 5.576 3.614 5.662 3.831 ;
      RECT 5.49 3.611 5.576 3.828 ;
      RECT 5.43 3.602 5.49 3.826 ;
      RECT 7.94 3.22 8.015 3.48 ;
      RECT 7.92 3.2 7.925 3.48 ;
      RECT 7.24 2.985 7.345 3.28 ;
      RECT 1.685 2.96 1.755 3.22 ;
      RECT 7.58 2.835 7.585 3.206 ;
      RECT 7.57 2.89 7.575 3.206 ;
      RECT 7.875 2.06 7.935 2.32 ;
      RECT 7.93 3.215 7.94 3.48 ;
      RECT 7.925 3.205 7.93 3.48 ;
      RECT 7.845 3.152 7.92 3.48 ;
      RECT 7.87 2.06 7.875 2.34 ;
      RECT 7.86 2.06 7.87 2.36 ;
      RECT 7.845 2.06 7.86 2.39 ;
      RECT 7.83 2.06 7.845 2.433 ;
      RECT 7.825 3.095 7.845 3.48 ;
      RECT 7.815 2.06 7.83 2.47 ;
      RECT 7.81 3.075 7.825 3.48 ;
      RECT 7.81 2.06 7.815 2.493 ;
      RECT 7.8 2.06 7.81 2.518 ;
      RECT 7.77 3.042 7.81 3.48 ;
      RECT 7.775 2.06 7.8 2.568 ;
      RECT 7.77 2.06 7.775 2.623 ;
      RECT 7.765 2.06 7.77 2.665 ;
      RECT 7.755 3.005 7.77 3.48 ;
      RECT 7.76 2.06 7.765 2.708 ;
      RECT 7.755 2.06 7.76 2.773 ;
      RECT 7.75 2.06 7.755 2.795 ;
      RECT 7.75 2.993 7.755 3.345 ;
      RECT 7.745 2.06 7.75 2.863 ;
      RECT 7.745 2.985 7.75 3.328 ;
      RECT 7.74 2.06 7.745 2.908 ;
      RECT 7.735 2.967 7.745 3.305 ;
      RECT 7.735 2.06 7.74 2.945 ;
      RECT 7.725 2.06 7.735 3.285 ;
      RECT 7.72 2.06 7.725 3.268 ;
      RECT 7.715 2.06 7.72 3.253 ;
      RECT 7.71 2.06 7.715 3.238 ;
      RECT 7.69 2.06 7.71 3.228 ;
      RECT 7.685 2.06 7.69 3.218 ;
      RECT 7.675 2.06 7.685 3.214 ;
      RECT 7.67 2.337 7.675 3.213 ;
      RECT 7.665 2.36 7.67 3.212 ;
      RECT 7.66 2.39 7.665 3.211 ;
      RECT 7.655 2.417 7.66 3.21 ;
      RECT 7.65 2.445 7.655 3.21 ;
      RECT 7.645 2.472 7.65 3.21 ;
      RECT 7.64 2.492 7.645 3.21 ;
      RECT 7.635 2.52 7.64 3.21 ;
      RECT 7.625 2.562 7.635 3.21 ;
      RECT 7.615 2.607 7.625 3.209 ;
      RECT 7.61 2.66 7.615 3.208 ;
      RECT 7.605 2.692 7.61 3.207 ;
      RECT 7.6 2.712 7.605 3.206 ;
      RECT 7.595 2.75 7.6 3.206 ;
      RECT 7.59 2.772 7.595 3.206 ;
      RECT 7.585 2.797 7.59 3.206 ;
      RECT 7.575 2.862 7.58 3.206 ;
      RECT 7.56 2.922 7.57 3.206 ;
      RECT 7.545 2.932 7.56 3.206 ;
      RECT 7.525 2.942 7.545 3.206 ;
      RECT 7.495 2.947 7.525 3.203 ;
      RECT 7.435 2.957 7.495 3.2 ;
      RECT 7.415 2.966 7.435 3.205 ;
      RECT 7.39 2.972 7.415 3.218 ;
      RECT 7.37 2.977 7.39 3.233 ;
      RECT 7.345 2.982 7.37 3.28 ;
      RECT 7.216 2.984 7.24 3.28 ;
      RECT 7.13 2.979 7.216 3.28 ;
      RECT 7.09 2.976 7.13 3.28 ;
      RECT 7.04 2.978 7.09 3.26 ;
      RECT 7.01 2.982 7.04 3.26 ;
      RECT 6.931 2.992 7.01 3.26 ;
      RECT 6.845 3.007 6.931 3.261 ;
      RECT 6.795 3.017 6.845 3.262 ;
      RECT 6.787 3.02 6.795 3.262 ;
      RECT 6.701 3.022 6.787 3.263 ;
      RECT 6.615 3.026 6.701 3.263 ;
      RECT 6.529 3.03 6.615 3.264 ;
      RECT 6.443 3.033 6.529 3.265 ;
      RECT 6.357 3.037 6.443 3.265 ;
      RECT 6.271 3.041 6.357 3.266 ;
      RECT 6.185 3.044 6.271 3.267 ;
      RECT 6.099 3.048 6.185 3.267 ;
      RECT 6.013 3.052 6.099 3.268 ;
      RECT 5.927 3.056 6.013 3.269 ;
      RECT 5.841 3.059 5.927 3.269 ;
      RECT 5.755 3.063 5.841 3.27 ;
      RECT 5.725 3.065 5.755 3.27 ;
      RECT 5.639 3.068 5.725 3.271 ;
      RECT 5.553 3.072 5.639 3.272 ;
      RECT 5.467 3.076 5.553 3.273 ;
      RECT 5.381 3.079 5.467 3.273 ;
      RECT 5.295 3.083 5.381 3.274 ;
      RECT 5.26 3.088 5.295 3.275 ;
      RECT 5.205 3.098 5.26 3.282 ;
      RECT 5.18 3.11 5.205 3.292 ;
      RECT 5.145 3.123 5.18 3.3 ;
      RECT 5.105 3.14 5.145 3.323 ;
      RECT 5.085 3.153 5.105 3.35 ;
      RECT 5.055 3.165 5.085 3.378 ;
      RECT 5.05 3.173 5.055 3.398 ;
      RECT 5.045 3.176 5.05 3.408 ;
      RECT 4.995 3.188 5.045 3.442 ;
      RECT 4.985 3.203 4.995 3.475 ;
      RECT 4.975 3.209 4.985 3.488 ;
      RECT 4.965 3.216 4.975 3.5 ;
      RECT 4.94 3.229 4.965 3.518 ;
      RECT 4.925 3.244 4.94 3.54 ;
      RECT 4.915 3.252 4.925 3.556 ;
      RECT 4.9 3.261 4.915 3.571 ;
      RECT 4.89 3.271 4.9 3.585 ;
      RECT 4.871 3.284 4.89 3.602 ;
      RECT 4.785 3.329 4.871 3.667 ;
      RECT 4.77 3.374 4.785 3.725 ;
      RECT 4.765 3.383 4.77 3.738 ;
      RECT 4.755 3.39 4.765 3.743 ;
      RECT 4.75 3.395 4.755 3.747 ;
      RECT 4.73 3.405 4.75 3.754 ;
      RECT 4.705 3.425 4.73 3.768 ;
      RECT 4.67 3.45 4.705 3.788 ;
      RECT 4.655 3.473 4.67 3.803 ;
      RECT 4.645 3.483 4.655 3.808 ;
      RECT 4.635 3.491 4.645 3.815 ;
      RECT 4.625 3.5 4.635 3.821 ;
      RECT 4.605 3.512 4.625 3.823 ;
      RECT 4.595 3.525 4.605 3.825 ;
      RECT 4.57 3.54 4.595 3.828 ;
      RECT 4.55 3.557 4.57 3.832 ;
      RECT 4.51 3.585 4.55 3.838 ;
      RECT 4.445 3.632 4.51 3.847 ;
      RECT 4.43 3.665 4.445 3.855 ;
      RECT 4.425 3.672 4.43 3.857 ;
      RECT 4.375 3.697 4.425 3.862 ;
      RECT 4.36 3.721 4.375 3.869 ;
      RECT 4.31 3.726 4.36 3.87 ;
      RECT 4.224 3.73 4.31 3.87 ;
      RECT 4.138 3.73 4.224 3.87 ;
      RECT 4.052 3.73 4.138 3.871 ;
      RECT 3.966 3.73 4.052 3.871 ;
      RECT 3.88 3.73 3.966 3.871 ;
      RECT 3.814 3.73 3.88 3.871 ;
      RECT 3.728 3.73 3.814 3.872 ;
      RECT 3.642 3.73 3.728 3.872 ;
      RECT 3.556 3.731 3.642 3.873 ;
      RECT 3.47 3.731 3.556 3.873 ;
      RECT 3.384 3.731 3.47 3.873 ;
      RECT 3.298 3.731 3.384 3.874 ;
      RECT 3.212 3.731 3.298 3.874 ;
      RECT 3.126 3.732 3.212 3.875 ;
      RECT 3.04 3.732 3.126 3.875 ;
      RECT 3.02 3.732 3.04 3.875 ;
      RECT 2.934 3.732 3.02 3.875 ;
      RECT 2.848 3.732 2.934 3.875 ;
      RECT 2.762 3.733 2.848 3.875 ;
      RECT 2.676 3.733 2.762 3.875 ;
      RECT 2.59 3.733 2.676 3.875 ;
      RECT 2.504 3.734 2.59 3.875 ;
      RECT 2.418 3.734 2.504 3.875 ;
      RECT 2.332 3.734 2.418 3.875 ;
      RECT 2.246 3.734 2.332 3.875 ;
      RECT 2.16 3.735 2.246 3.875 ;
      RECT 2.11 3.732 2.16 3.875 ;
      RECT 2.1 3.73 2.11 3.874 ;
      RECT 2.096 3.73 2.1 3.873 ;
      RECT 2.01 3.725 2.096 3.868 ;
      RECT 1.988 3.718 2.01 3.862 ;
      RECT 1.902 3.709 1.988 3.856 ;
      RECT 1.816 3.696 1.902 3.847 ;
      RECT 1.73 3.682 1.816 3.837 ;
      RECT 1.685 3.672 1.73 3.83 ;
      RECT 1.665 2.96 1.685 3.238 ;
      RECT 1.665 3.665 1.685 3.826 ;
      RECT 1.635 2.96 1.665 3.26 ;
      RECT 1.625 3.632 1.665 3.823 ;
      RECT 1.62 2.96 1.635 3.28 ;
      RECT 1.62 3.597 1.625 3.821 ;
      RECT 1.615 2.96 1.62 3.405 ;
      RECT 1.615 3.557 1.62 3.821 ;
      RECT 1.605 2.96 1.615 3.821 ;
      RECT 1.53 2.96 1.605 3.815 ;
      RECT 1.5 2.96 1.53 3.805 ;
      RECT 1.495 2.96 1.5 3.797 ;
      RECT 1.49 3.002 1.495 3.79 ;
      RECT 1.48 3.071 1.49 3.781 ;
      RECT 1.475 3.141 1.48 3.733 ;
      RECT 1.47 3.205 1.475 3.63 ;
      RECT 1.465 3.24 1.47 3.585 ;
      RECT 1.463 3.277 1.465 3.477 ;
      RECT 1.46 3.285 1.463 3.47 ;
      RECT 1.455 3.35 1.46 3.413 ;
      RECT 5.53 2.44 5.81 2.72 ;
      RECT 5.52 2.44 5.81 2.583 ;
      RECT 5.475 2.305 5.735 2.565 ;
      RECT 5.475 2.42 5.79 2.565 ;
      RECT 5.475 2.39 5.785 2.565 ;
      RECT 5.475 2.377 5.775 2.565 ;
      RECT 5.475 2.367 5.77 2.565 ;
      RECT 1.45 2.35 1.71 2.61 ;
      RECT 5.22 1.9 5.48 2.16 ;
      RECT 5.21 1.925 5.48 2.12 ;
      RECT 5.205 1.925 5.21 2.119 ;
      RECT 5.135 1.92 5.205 2.111 ;
      RECT 5.05 1.907 5.135 2.094 ;
      RECT 5.046 1.899 5.05 2.084 ;
      RECT 4.96 1.892 5.046 2.074 ;
      RECT 4.951 1.884 4.96 2.064 ;
      RECT 4.865 1.877 4.951 2.052 ;
      RECT 4.845 1.868 4.865 2.038 ;
      RECT 4.79 1.863 4.845 2.03 ;
      RECT 4.78 1.857 4.79 2.024 ;
      RECT 4.76 1.855 4.78 2.02 ;
      RECT 4.752 1.854 4.76 2.016 ;
      RECT 4.666 1.846 4.752 2.005 ;
      RECT 4.58 1.832 4.666 1.985 ;
      RECT 4.52 1.82 4.58 1.97 ;
      RECT 4.51 1.815 4.52 1.965 ;
      RECT 4.46 1.815 4.51 1.967 ;
      RECT 4.413 1.817 4.46 1.971 ;
      RECT 4.327 1.824 4.413 1.976 ;
      RECT 4.241 1.832 4.327 1.982 ;
      RECT 4.155 1.841 4.241 1.988 ;
      RECT 4.096 1.847 4.155 1.993 ;
      RECT 4.01 1.852 4.096 1.999 ;
      RECT 3.935 1.857 4.01 2.005 ;
      RECT 3.896 1.859 3.935 2.01 ;
      RECT 3.81 1.856 3.896 2.015 ;
      RECT 3.725 1.854 3.81 2.022 ;
      RECT 3.693 1.853 3.725 2.025 ;
      RECT 3.607 1.852 3.693 2.026 ;
      RECT 3.521 1.851 3.607 2.027 ;
      RECT 3.435 1.85 3.521 2.027 ;
      RECT 3.349 1.849 3.435 2.028 ;
      RECT 3.263 1.848 3.349 2.029 ;
      RECT 3.177 1.847 3.263 2.03 ;
      RECT 3.091 1.846 3.177 2.03 ;
      RECT 3.005 1.845 3.091 2.031 ;
      RECT 2.955 1.845 3.005 2.032 ;
      RECT 2.941 1.846 2.955 2.032 ;
      RECT 2.855 1.853 2.941 2.033 ;
      RECT 2.781 1.864 2.855 2.034 ;
      RECT 2.695 1.873 2.781 2.035 ;
      RECT 2.66 1.88 2.695 2.05 ;
      RECT 2.635 1.883 2.66 2.08 ;
      RECT 2.61 1.892 2.635 2.109 ;
      RECT 2.6 1.903 2.61 2.129 ;
      RECT 2.59 1.911 2.6 2.143 ;
      RECT 2.585 1.917 2.59 2.153 ;
      RECT 2.56 1.934 2.585 2.17 ;
      RECT 2.545 1.956 2.56 2.198 ;
      RECT 2.515 1.982 2.545 2.228 ;
      RECT 2.495 2.011 2.515 2.258 ;
      RECT 2.49 2.026 2.495 2.275 ;
      RECT 2.47 2.041 2.49 2.29 ;
      RECT 2.46 2.059 2.47 2.308 ;
      RECT 2.45 2.07 2.46 2.323 ;
      RECT 2.4 2.102 2.45 2.349 ;
      RECT 2.395 2.132 2.4 2.369 ;
      RECT 2.385 2.145 2.395 2.375 ;
      RECT 2.376 2.155 2.385 2.383 ;
      RECT 2.365 2.166 2.376 2.391 ;
      RECT 2.36 2.176 2.365 2.397 ;
      RECT 2.345 2.197 2.36 2.404 ;
      RECT 2.33 2.227 2.345 2.412 ;
      RECT 2.295 2.257 2.33 2.418 ;
      RECT 2.27 2.275 2.295 2.425 ;
      RECT 2.22 2.283 2.27 2.434 ;
      RECT 2.195 2.288 2.22 2.443 ;
      RECT 2.14 2.294 2.195 2.453 ;
      RECT 2.135 2.299 2.14 2.461 ;
      RECT 2.121 2.302 2.135 2.463 ;
      RECT 2.035 2.314 2.121 2.475 ;
      RECT 2.025 2.326 2.035 2.488 ;
      RECT 1.94 2.339 2.025 2.5 ;
      RECT 1.896 2.356 1.94 2.514 ;
      RECT 1.81 2.373 1.896 2.53 ;
      RECT 1.78 2.387 1.81 2.544 ;
      RECT 1.77 2.392 1.78 2.549 ;
      RECT 1.71 2.395 1.77 2.558 ;
      RECT 4.6 2.665 4.86 2.925 ;
      RECT 4.6 2.665 4.88 2.778 ;
      RECT 4.6 2.665 4.905 2.745 ;
      RECT 4.6 2.665 4.91 2.725 ;
      RECT 4.65 2.44 4.93 2.72 ;
      RECT 4.205 3.175 4.465 3.435 ;
      RECT 4.195 3.032 4.39 3.373 ;
      RECT 4.19 3.14 4.405 3.365 ;
      RECT 4.185 3.19 4.465 3.355 ;
      RECT 4.175 3.267 4.465 3.34 ;
      RECT 4.195 3.115 4.405 3.373 ;
      RECT 4.205 2.99 4.39 3.435 ;
      RECT 4.205 2.885 4.37 3.435 ;
      RECT 4.215 2.872 4.37 3.435 ;
      RECT 4.215 2.83 4.36 3.435 ;
      RECT 4.22 2.755 4.36 3.435 ;
      RECT 4.25 2.405 4.36 3.435 ;
      RECT 4.255 2.135 4.38 2.758 ;
      RECT 4.225 2.71 4.38 2.758 ;
      RECT 4.24 2.512 4.36 3.435 ;
      RECT 4.23 2.622 4.38 2.758 ;
      RECT 4.255 2.135 4.395 2.615 ;
      RECT 4.255 2.135 4.415 2.49 ;
      RECT 4.22 2.135 4.48 2.395 ;
      RECT 3.69 2.44 3.97 2.72 ;
      RECT 3.675 2.44 3.97 2.7 ;
      RECT 1.73 3.305 1.99 3.565 ;
      RECT 3.515 3.16 3.775 3.42 ;
      RECT 3.495 3.18 3.775 3.395 ;
      RECT 3.452 3.18 3.495 3.394 ;
      RECT 3.366 3.181 3.452 3.391 ;
      RECT 3.28 3.182 3.366 3.387 ;
      RECT 3.205 3.184 3.28 3.384 ;
      RECT 3.182 3.185 3.205 3.382 ;
      RECT 3.096 3.186 3.182 3.38 ;
      RECT 3.01 3.187 3.096 3.377 ;
      RECT 2.986 3.188 3.01 3.375 ;
      RECT 2.9 3.19 2.986 3.372 ;
      RECT 2.815 3.192 2.9 3.373 ;
      RECT 2.758 3.193 2.815 3.379 ;
      RECT 2.672 3.195 2.758 3.389 ;
      RECT 2.586 3.198 2.672 3.402 ;
      RECT 2.5 3.2 2.586 3.414 ;
      RECT 2.486 3.201 2.5 3.421 ;
      RECT 2.4 3.202 2.486 3.429 ;
      RECT 2.36 3.204 2.4 3.438 ;
      RECT 2.351 3.205 2.36 3.441 ;
      RECT 2.265 3.213 2.351 3.447 ;
      RECT 2.245 3.222 2.265 3.455 ;
      RECT 2.16 3.237 2.245 3.463 ;
      RECT 2.1 3.26 2.16 3.474 ;
      RECT 2.09 3.272 2.1 3.479 ;
      RECT 2.05 3.282 2.09 3.483 ;
      RECT 1.995 3.299 2.05 3.491 ;
      RECT 1.99 3.309 1.995 3.495 ;
      RECT 3.056 2.44 3.115 2.837 ;
      RECT 2.97 2.44 3.175 2.828 ;
      RECT 2.965 2.47 3.175 2.823 ;
      RECT 2.931 2.47 3.175 2.821 ;
      RECT 2.845 2.47 3.175 2.815 ;
      RECT 2.8 2.47 3.195 2.793 ;
      RECT 2.8 2.47 3.215 2.748 ;
      RECT 2.76 2.47 3.215 2.738 ;
      RECT 2.97 2.44 3.25 2.72 ;
      RECT 2.705 2.44 2.965 2.7 ;
      RECT 1.89 1.92 2.15 2.18 ;
      RECT 1.97 1.88 2.25 2.16 ;
      RECT 72.48 0.815 72.85 1.185 ;
      RECT 70.77 7.04 71.14 7.41 ;
      RECT 56.695 0.815 57.065 1.185 ;
      RECT 54.985 7.04 55.355 7.41 ;
      RECT 40.91 0.815 41.28 1.185 ;
      RECT 39.2 7.04 39.57 7.41 ;
      RECT 25.135 0.815 25.505 1.185 ;
      RECT 23.425 7.04 23.795 7.41 ;
      RECT 9.355 0.815 9.725 1.185 ;
      RECT 7.645 7.04 8.015 7.41 ;
    LAYER via1 ;
      RECT 78.505 7.375 78.655 7.525 ;
      RECT 76.135 6.74 76.285 6.89 ;
      RECT 76.12 2.065 76.27 2.215 ;
      RECT 75.33 2.45 75.48 2.6 ;
      RECT 75.33 6.325 75.48 6.475 ;
      RECT 74.295 5.955 74.445 6.105 ;
      RECT 74.29 2.805 74.44 2.955 ;
      RECT 73.685 1.44 73.835 1.59 ;
      RECT 73.37 2.96 73.52 3.11 ;
      RECT 72.59 0.925 72.74 1.075 ;
      RECT 72.47 2.29 72.62 2.44 ;
      RECT 72.35 2.86 72.5 3.01 ;
      RECT 71.52 6.71 71.67 6.86 ;
      RECT 71.27 2.555 71.42 2.705 ;
      RECT 70.935 3.275 71.085 3.425 ;
      RECT 70.88 7.15 71.03 7.3 ;
      RECT 70.855 2.115 71.005 2.265 ;
      RECT 69.42 2.51 69.57 2.66 ;
      RECT 68.655 2.36 68.805 2.51 ;
      RECT 68.4 1.955 68.55 2.105 ;
      RECT 67.78 2.72 67.93 2.87 ;
      RECT 67.4 2.19 67.55 2.34 ;
      RECT 67.385 3.23 67.535 3.38 ;
      RECT 66.855 2.495 67.005 2.645 ;
      RECT 66.695 3.215 66.845 3.365 ;
      RECT 65.885 2.495 66.035 2.645 ;
      RECT 65.07 1.975 65.22 2.125 ;
      RECT 64.91 3.36 65.06 3.51 ;
      RECT 64.675 3.015 64.825 3.165 ;
      RECT 64.63 2.405 64.78 2.555 ;
      RECT 63.63 3.025 63.78 3.175 ;
      RECT 62.695 6.755 62.845 6.905 ;
      RECT 60.35 6.74 60.5 6.89 ;
      RECT 60.335 2.065 60.485 2.215 ;
      RECT 59.545 2.45 59.695 2.6 ;
      RECT 59.545 6.325 59.695 6.475 ;
      RECT 58.51 5.955 58.66 6.105 ;
      RECT 58.505 2.805 58.655 2.955 ;
      RECT 57.9 1.44 58.05 1.59 ;
      RECT 57.585 2.96 57.735 3.11 ;
      RECT 56.805 0.925 56.955 1.075 ;
      RECT 56.685 2.29 56.835 2.44 ;
      RECT 56.565 2.86 56.715 3.01 ;
      RECT 55.735 6.71 55.885 6.86 ;
      RECT 55.485 2.555 55.635 2.705 ;
      RECT 55.15 3.275 55.3 3.425 ;
      RECT 55.095 7.15 55.245 7.3 ;
      RECT 55.07 2.115 55.22 2.265 ;
      RECT 53.635 2.51 53.785 2.66 ;
      RECT 52.87 2.36 53.02 2.51 ;
      RECT 52.615 1.955 52.765 2.105 ;
      RECT 51.995 2.72 52.145 2.87 ;
      RECT 51.615 2.19 51.765 2.34 ;
      RECT 51.6 3.23 51.75 3.38 ;
      RECT 51.07 2.495 51.22 2.645 ;
      RECT 50.91 3.215 51.06 3.365 ;
      RECT 50.1 2.495 50.25 2.645 ;
      RECT 49.285 1.975 49.435 2.125 ;
      RECT 49.125 3.36 49.275 3.51 ;
      RECT 48.89 3.015 49.04 3.165 ;
      RECT 48.845 2.405 48.995 2.555 ;
      RECT 47.845 3.025 47.995 3.175 ;
      RECT 46.91 6.755 47.06 6.905 ;
      RECT 44.565 6.74 44.715 6.89 ;
      RECT 44.55 2.065 44.7 2.215 ;
      RECT 43.76 2.45 43.91 2.6 ;
      RECT 43.76 6.325 43.91 6.475 ;
      RECT 42.725 5.955 42.875 6.105 ;
      RECT 42.72 2.805 42.87 2.955 ;
      RECT 42.115 1.44 42.265 1.59 ;
      RECT 41.8 2.96 41.95 3.11 ;
      RECT 41.02 0.925 41.17 1.075 ;
      RECT 40.9 2.29 41.05 2.44 ;
      RECT 40.78 2.86 40.93 3.01 ;
      RECT 40.005 6.715 40.155 6.865 ;
      RECT 39.7 2.555 39.85 2.705 ;
      RECT 39.365 3.275 39.515 3.425 ;
      RECT 39.31 7.15 39.46 7.3 ;
      RECT 39.285 2.115 39.435 2.265 ;
      RECT 37.85 2.51 38 2.66 ;
      RECT 37.085 2.36 37.235 2.51 ;
      RECT 36.83 1.955 36.98 2.105 ;
      RECT 36.21 2.72 36.36 2.87 ;
      RECT 35.83 2.19 35.98 2.34 ;
      RECT 35.815 3.23 35.965 3.38 ;
      RECT 35.285 2.495 35.435 2.645 ;
      RECT 35.125 3.215 35.275 3.365 ;
      RECT 34.315 2.495 34.465 2.645 ;
      RECT 33.5 1.975 33.65 2.125 ;
      RECT 33.34 3.36 33.49 3.51 ;
      RECT 33.105 3.015 33.255 3.165 ;
      RECT 33.06 2.405 33.21 2.555 ;
      RECT 32.06 3.025 32.21 3.175 ;
      RECT 31.18 6.76 31.33 6.91 ;
      RECT 28.79 6.74 28.94 6.89 ;
      RECT 28.775 2.065 28.925 2.215 ;
      RECT 27.985 2.45 28.135 2.6 ;
      RECT 27.985 6.325 28.135 6.475 ;
      RECT 26.95 5.955 27.1 6.105 ;
      RECT 26.945 2.805 27.095 2.955 ;
      RECT 26.34 1.44 26.49 1.59 ;
      RECT 26.025 2.96 26.175 3.11 ;
      RECT 25.245 0.925 25.395 1.075 ;
      RECT 25.125 2.29 25.275 2.44 ;
      RECT 25.005 2.86 25.155 3.01 ;
      RECT 24.225 6.71 24.375 6.86 ;
      RECT 23.925 2.555 24.075 2.705 ;
      RECT 23.59 3.275 23.74 3.425 ;
      RECT 23.535 7.15 23.685 7.3 ;
      RECT 23.51 2.115 23.66 2.265 ;
      RECT 22.075 2.51 22.225 2.66 ;
      RECT 21.31 2.36 21.46 2.51 ;
      RECT 21.055 1.955 21.205 2.105 ;
      RECT 20.435 2.72 20.585 2.87 ;
      RECT 20.055 2.19 20.205 2.34 ;
      RECT 20.04 3.23 20.19 3.38 ;
      RECT 19.51 2.495 19.66 2.645 ;
      RECT 19.35 3.215 19.5 3.365 ;
      RECT 18.54 2.495 18.69 2.645 ;
      RECT 17.725 1.975 17.875 2.125 ;
      RECT 17.565 3.36 17.715 3.51 ;
      RECT 17.33 3.015 17.48 3.165 ;
      RECT 17.285 2.405 17.435 2.555 ;
      RECT 16.285 3.025 16.435 3.175 ;
      RECT 15.4 6.755 15.55 6.905 ;
      RECT 13.01 6.74 13.16 6.89 ;
      RECT 12.995 2.065 13.145 2.215 ;
      RECT 12.205 2.45 12.355 2.6 ;
      RECT 12.205 6.325 12.355 6.475 ;
      RECT 11.17 5.955 11.32 6.105 ;
      RECT 11.165 2.805 11.315 2.955 ;
      RECT 10.56 1.44 10.71 1.59 ;
      RECT 10.245 2.96 10.395 3.11 ;
      RECT 9.465 0.925 9.615 1.075 ;
      RECT 9.345 2.29 9.495 2.44 ;
      RECT 9.225 2.86 9.375 3.01 ;
      RECT 8.415 6.705 8.565 6.855 ;
      RECT 8.145 2.555 8.295 2.705 ;
      RECT 7.81 3.275 7.96 3.425 ;
      RECT 7.755 7.15 7.905 7.3 ;
      RECT 7.73 2.115 7.88 2.265 ;
      RECT 6.295 2.51 6.445 2.66 ;
      RECT 5.53 2.36 5.68 2.51 ;
      RECT 5.275 1.955 5.425 2.105 ;
      RECT 4.655 2.72 4.805 2.87 ;
      RECT 4.275 2.19 4.425 2.34 ;
      RECT 4.26 3.23 4.41 3.38 ;
      RECT 3.73 2.495 3.88 2.645 ;
      RECT 3.57 3.215 3.72 3.365 ;
      RECT 2.76 2.495 2.91 2.645 ;
      RECT 1.945 1.975 2.095 2.125 ;
      RECT 1.785 3.36 1.935 3.51 ;
      RECT 1.55 3.015 1.7 3.165 ;
      RECT 1.505 2.405 1.655 2.555 ;
      RECT 0.505 3.025 0.655 3.175 ;
      RECT -1.18 7.095 -1.03 7.245 ;
      RECT -1.555 6.355 -1.405 6.505 ;
    LAYER met1 ;
      RECT 63.38 1.26 73.04 1.74 ;
      RECT 47.595 1.26 57.255 1.74 ;
      RECT 31.81 1.26 41.47 1.74 ;
      RECT 16.035 1.26 25.695 1.74 ;
      RECT 0.255 1.26 9.915 1.74 ;
      RECT 63.38 1.26 73.095 1.59 ;
      RECT 47.595 1.26 57.31 1.59 ;
      RECT 31.81 1.26 41.525 1.59 ;
      RECT 16.035 1.26 25.75 1.59 ;
      RECT 0.255 1.26 9.97 1.59 ;
      RECT 63.495 0 73.21 1.585 ;
      RECT 47.71 0 57.425 1.585 ;
      RECT 31.925 0 41.64 1.585 ;
      RECT 16.15 0 25.865 1.585 ;
      RECT 0.37 0 10.085 1.585 ;
      RECT -2.79 0 78.975 0.305 ;
      RECT 69.065 4.135 78.975 4.745 ;
      RECT 53.28 4.135 68.68 4.745 ;
      RECT 37.495 4.135 52.895 4.745 ;
      RECT 21.72 4.135 37.11 4.745 ;
      RECT 5.94 4.135 21.335 4.745 ;
      RECT -2.79 4.44 5.555 4.745 ;
      RECT 63.38 3.98 73.04 4.74 ;
      RECT 0.005 4.135 78.975 4.74 ;
      RECT 47.595 3.98 57.255 4.74 ;
      RECT 31.81 3.98 41.47 4.74 ;
      RECT 16.035 3.98 25.695 4.74 ;
      RECT 0.255 3.98 9.915 4.74 ;
      RECT -2.79 8.575 78.975 8.88 ;
      RECT 70.065 6.315 70.235 8.88 ;
      RECT 54.28 6.315 54.45 8.88 ;
      RECT 38.495 6.315 38.665 8.88 ;
      RECT 22.72 6.315 22.89 8.88 ;
      RECT 6.94 6.315 7.11 8.88 ;
      RECT 70.435 6.285 70.725 6.515 ;
      RECT 54.65 6.285 54.94 6.515 ;
      RECT 38.865 6.285 39.155 6.515 ;
      RECT 23.09 6.285 23.38 6.515 ;
      RECT 7.31 6.285 7.6 6.515 ;
      RECT 70.065 6.315 70.725 6.485 ;
      RECT 54.28 6.315 54.94 6.485 ;
      RECT 38.495 6.315 39.155 6.485 ;
      RECT 22.72 6.315 23.38 6.485 ;
      RECT 6.94 6.315 7.6 6.485 ;
      RECT 78.375 7.765 78.665 7.995 ;
      RECT 78.435 6.285 78.605 7.995 ;
      RECT 78.405 7.275 78.755 7.625 ;
      RECT 78.375 6.285 78.665 6.515 ;
      RECT 78.375 2.365 78.665 2.595 ;
      RECT 78.435 0.885 78.605 2.595 ;
      RECT 78.375 0.885 78.665 1.115 ;
      RECT 77.965 2.735 78.295 2.965 ;
      RECT 77.965 2.765 78.465 2.935 ;
      RECT 77.965 2.395 78.155 2.965 ;
      RECT 77.385 2.365 77.675 2.595 ;
      RECT 77.385 2.395 78.155 2.565 ;
      RECT 77.445 0.885 77.615 2.595 ;
      RECT 77.385 0.885 77.675 1.115 ;
      RECT 77.385 7.765 77.675 7.995 ;
      RECT 77.445 6.285 77.615 7.995 ;
      RECT 77.385 6.285 77.675 6.515 ;
      RECT 77.385 6.325 78.235 6.485 ;
      RECT 78.065 5.915 78.235 6.485 ;
      RECT 77.385 6.32 77.775 6.485 ;
      RECT 78.005 5.915 78.295 6.145 ;
      RECT 78.005 5.945 78.465 6.115 ;
      RECT 77.015 2.735 77.305 2.965 ;
      RECT 77.015 2.765 77.475 2.935 ;
      RECT 77.075 1.655 77.24 2.965 ;
      RECT 75.59 1.625 75.88 1.855 ;
      RECT 75.59 1.655 77.24 1.825 ;
      RECT 75.65 0.885 75.82 1.855 ;
      RECT 75.59 0.885 75.88 1.115 ;
      RECT 75.59 7.765 75.88 7.995 ;
      RECT 75.65 7.025 75.82 7.995 ;
      RECT 75.65 7.12 77.24 7.29 ;
      RECT 77.07 5.915 77.24 7.29 ;
      RECT 75.59 7.025 75.88 7.255 ;
      RECT 77.015 5.915 77.305 6.145 ;
      RECT 77.015 5.945 77.475 6.115 ;
      RECT 76.02 1.965 76.37 2.315 ;
      RECT 73.685 2.025 76.37 2.195 ;
      RECT 73.685 1.34 73.855 2.195 ;
      RECT 73.585 1.34 73.935 1.69 ;
      RECT 76.045 6.655 76.37 6.98 ;
      RECT 71.42 6.61 71.77 6.96 ;
      RECT 76.02 6.655 76.37 6.885 ;
      RECT 71.24 6.655 71.77 6.885 ;
      RECT 71.07 6.685 76.37 6.855 ;
      RECT 75.245 2.365 75.565 2.685 ;
      RECT 75.215 2.365 75.565 2.595 ;
      RECT 75.045 2.395 75.565 2.565 ;
      RECT 75.245 6.255 75.565 6.545 ;
      RECT 75.215 6.285 75.565 6.515 ;
      RECT 75.045 6.315 75.565 6.485 ;
      RECT 74.19 2.705 74.54 3.055 ;
      RECT 74.19 2.765 74.68 2.935 ;
      RECT 74.195 5.855 74.545 6.205 ;
      RECT 69.44 5.915 69.73 6.145 ;
      RECT 69.44 5.945 74.68 6.115 ;
      RECT 71.88 2.465 72.065 2.675 ;
      RECT 71.87 2.47 72.08 2.668 ;
      RECT 71.87 2.47 72.166 2.645 ;
      RECT 71.87 2.47 72.225 2.62 ;
      RECT 71.87 2.47 72.28 2.6 ;
      RECT 71.87 2.47 72.29 2.588 ;
      RECT 71.87 2.47 72.485 2.527 ;
      RECT 71.87 2.47 72.515 2.51 ;
      RECT 71.87 2.47 72.535 2.5 ;
      RECT 72.415 2.235 72.675 2.495 ;
      RECT 72.4 2.325 72.415 2.542 ;
      RECT 71.935 2.457 72.675 2.495 ;
      RECT 72.386 2.336 72.4 2.548 ;
      RECT 71.975 2.45 72.675 2.495 ;
      RECT 72.3 2.376 72.386 2.567 ;
      RECT 72.225 2.437 72.675 2.495 ;
      RECT 72.295 2.412 72.3 2.584 ;
      RECT 72.28 2.422 72.675 2.495 ;
      RECT 72.29 2.417 72.295 2.586 ;
      RECT 72.585 2.922 72.59 3.014 ;
      RECT 72.58 2.9 72.585 3.031 ;
      RECT 72.575 2.89 72.58 3.043 ;
      RECT 72.565 2.881 72.575 3.053 ;
      RECT 72.56 2.876 72.565 3.061 ;
      RECT 72.555 2.735 72.56 3.064 ;
      RECT 72.521 2.735 72.555 3.075 ;
      RECT 72.435 2.735 72.521 3.11 ;
      RECT 72.355 2.735 72.435 3.158 ;
      RECT 72.326 2.735 72.355 3.182 ;
      RECT 72.24 2.735 72.326 3.188 ;
      RECT 72.235 2.919 72.24 3.193 ;
      RECT 72.2 2.93 72.235 3.196 ;
      RECT 72.175 2.945 72.2 3.2 ;
      RECT 72.161 2.954 72.175 3.202 ;
      RECT 72.075 2.981 72.161 3.208 ;
      RECT 72.01 3.022 72.075 3.217 ;
      RECT 71.995 3.042 72.01 3.222 ;
      RECT 71.965 3.052 71.995 3.225 ;
      RECT 71.96 3.062 71.965 3.228 ;
      RECT 71.93 3.067 71.96 3.23 ;
      RECT 71.91 3.072 71.93 3.234 ;
      RECT 71.825 3.075 71.91 3.241 ;
      RECT 71.81 3.072 71.825 3.247 ;
      RECT 71.8 3.069 71.81 3.249 ;
      RECT 71.78 3.066 71.8 3.251 ;
      RECT 71.76 3.062 71.78 3.252 ;
      RECT 71.745 3.058 71.76 3.254 ;
      RECT 71.735 3.055 71.745 3.255 ;
      RECT 71.695 3.049 71.735 3.253 ;
      RECT 71.685 3.044 71.695 3.251 ;
      RECT 71.67 3.041 71.685 3.247 ;
      RECT 71.645 3.036 71.67 3.24 ;
      RECT 71.595 3.027 71.645 3.228 ;
      RECT 71.525 3.013 71.595 3.21 ;
      RECT 71.467 2.998 71.525 3.192 ;
      RECT 71.381 2.981 71.467 3.172 ;
      RECT 71.295 2.96 71.381 3.147 ;
      RECT 71.245 2.945 71.295 3.128 ;
      RECT 71.241 2.939 71.245 3.12 ;
      RECT 71.155 2.929 71.241 3.107 ;
      RECT 71.12 2.914 71.155 3.09 ;
      RECT 71.105 2.907 71.12 3.083 ;
      RECT 71.045 2.895 71.105 3.071 ;
      RECT 71.025 2.882 71.045 3.059 ;
      RECT 70.985 2.873 71.025 3.051 ;
      RECT 70.98 2.865 70.985 3.044 ;
      RECT 70.9 2.855 70.98 3.03 ;
      RECT 70.885 2.842 70.9 3.015 ;
      RECT 70.88 2.84 70.885 3.013 ;
      RECT 70.801 2.828 70.88 3 ;
      RECT 70.715 2.803 70.801 2.975 ;
      RECT 70.7 2.772 70.715 2.96 ;
      RECT 70.685 2.747 70.7 2.956 ;
      RECT 70.67 2.74 70.685 2.952 ;
      RECT 70.495 2.745 70.5 2.948 ;
      RECT 70.49 2.75 70.495 2.943 ;
      RECT 70.5 2.74 70.67 2.95 ;
      RECT 71.215 2.5 71.32 2.76 ;
      RECT 72.03 2.025 72.035 2.25 ;
      RECT 72.16 2.025 72.215 2.235 ;
      RECT 72.215 2.03 72.225 2.228 ;
      RECT 72.121 2.025 72.16 2.238 ;
      RECT 72.035 2.025 72.121 2.245 ;
      RECT 72.015 2.03 72.03 2.251 ;
      RECT 72.005 2.07 72.015 2.253 ;
      RECT 71.975 2.08 72.005 2.255 ;
      RECT 71.97 2.085 71.975 2.257 ;
      RECT 71.945 2.09 71.97 2.259 ;
      RECT 71.93 2.095 71.945 2.261 ;
      RECT 71.915 2.097 71.93 2.263 ;
      RECT 71.91 2.102 71.915 2.265 ;
      RECT 71.86 2.11 71.91 2.268 ;
      RECT 71.835 2.119 71.86 2.273 ;
      RECT 71.825 2.126 71.835 2.278 ;
      RECT 71.82 2.129 71.825 2.282 ;
      RECT 71.8 2.132 71.82 2.291 ;
      RECT 71.77 2.14 71.8 2.311 ;
      RECT 71.741 2.153 71.77 2.333 ;
      RECT 71.655 2.187 71.741 2.377 ;
      RECT 71.65 2.213 71.655 2.415 ;
      RECT 71.645 2.217 71.65 2.424 ;
      RECT 71.61 2.23 71.645 2.457 ;
      RECT 71.6 2.244 71.61 2.495 ;
      RECT 71.595 2.248 71.6 2.508 ;
      RECT 71.59 2.252 71.595 2.513 ;
      RECT 71.58 2.26 71.59 2.525 ;
      RECT 71.575 2.267 71.58 2.54 ;
      RECT 71.55 2.28 71.575 2.565 ;
      RECT 71.51 2.309 71.55 2.62 ;
      RECT 71.495 2.334 71.51 2.675 ;
      RECT 71.485 2.345 71.495 2.698 ;
      RECT 71.48 2.352 71.485 2.71 ;
      RECT 71.475 2.356 71.48 2.718 ;
      RECT 71.42 2.384 71.475 2.76 ;
      RECT 71.4 2.42 71.42 2.76 ;
      RECT 71.385 2.435 71.4 2.76 ;
      RECT 71.33 2.467 71.385 2.76 ;
      RECT 71.32 2.497 71.33 2.76 ;
      RECT 70.93 2.112 71.115 2.35 ;
      RECT 70.915 2.114 71.125 2.345 ;
      RECT 70.8 2.06 71.06 2.32 ;
      RECT 70.795 2.097 71.06 2.274 ;
      RECT 70.79 2.107 71.06 2.271 ;
      RECT 70.785 2.147 71.125 2.265 ;
      RECT 70.78 2.18 71.125 2.255 ;
      RECT 70.79 2.122 71.14 2.193 ;
      RECT 71.087 3.22 71.1 3.75 ;
      RECT 71.001 3.22 71.1 3.749 ;
      RECT 71.001 3.22 71.105 3.748 ;
      RECT 70.915 3.22 71.105 3.746 ;
      RECT 70.91 3.22 71.105 3.743 ;
      RECT 70.91 3.22 71.115 3.741 ;
      RECT 70.905 3.512 71.115 3.738 ;
      RECT 70.905 3.522 71.12 3.735 ;
      RECT 70.905 3.59 71.125 3.731 ;
      RECT 70.895 3.595 71.125 3.73 ;
      RECT 70.895 3.687 71.13 3.727 ;
      RECT 70.88 3.22 71.14 3.48 ;
      RECT 70.81 7.765 71.1 7.995 ;
      RECT 70.87 7.025 71.04 7.995 ;
      RECT 70.785 7.055 71.125 7.4 ;
      RECT 70.81 7.025 71.1 7.4 ;
      RECT 70.11 2.21 70.155 3.745 ;
      RECT 70.31 2.21 70.34 2.425 ;
      RECT 68.685 1.95 68.805 2.16 ;
      RECT 68.345 1.9 68.605 2.16 ;
      RECT 68.345 1.945 68.64 2.15 ;
      RECT 70.35 2.226 70.355 2.28 ;
      RECT 70.345 2.219 70.35 2.413 ;
      RECT 70.34 2.213 70.345 2.42 ;
      RECT 70.295 2.21 70.31 2.433 ;
      RECT 70.29 2.21 70.295 2.455 ;
      RECT 70.285 2.21 70.29 2.503 ;
      RECT 70.28 2.21 70.285 2.523 ;
      RECT 70.27 2.21 70.28 2.63 ;
      RECT 70.265 2.21 70.27 2.693 ;
      RECT 70.26 2.21 70.265 2.75 ;
      RECT 70.255 2.21 70.26 2.758 ;
      RECT 70.24 2.21 70.255 2.865 ;
      RECT 70.23 2.21 70.24 3 ;
      RECT 70.22 2.21 70.23 3.11 ;
      RECT 70.21 2.21 70.22 3.167 ;
      RECT 70.205 2.21 70.21 3.207 ;
      RECT 70.2 2.21 70.205 3.243 ;
      RECT 70.19 2.21 70.2 3.283 ;
      RECT 70.185 2.21 70.19 3.325 ;
      RECT 70.165 2.21 70.185 3.39 ;
      RECT 70.17 3.535 70.175 3.715 ;
      RECT 70.165 3.517 70.17 3.723 ;
      RECT 70.16 2.21 70.165 3.453 ;
      RECT 70.16 3.497 70.165 3.73 ;
      RECT 70.155 2.21 70.16 3.74 ;
      RECT 70.1 2.21 70.11 2.51 ;
      RECT 70.105 2.757 70.11 3.745 ;
      RECT 70.1 2.822 70.105 3.745 ;
      RECT 70.095 2.211 70.1 2.5 ;
      RECT 70.09 2.887 70.1 3.745 ;
      RECT 70.085 2.212 70.095 2.49 ;
      RECT 70.075 3 70.09 3.745 ;
      RECT 70.08 2.213 70.085 2.48 ;
      RECT 70.06 2.214 70.08 2.458 ;
      RECT 70.065 3.097 70.075 3.745 ;
      RECT 70.06 3.172 70.065 3.745 ;
      RECT 70.05 2.213 70.06 2.435 ;
      RECT 70.055 3.215 70.06 3.745 ;
      RECT 70.05 3.242 70.055 3.745 ;
      RECT 70.04 2.211 70.05 2.423 ;
      RECT 70.045 3.285 70.05 3.745 ;
      RECT 70.04 3.312 70.045 3.745 ;
      RECT 70.03 2.21 70.04 2.41 ;
      RECT 70.035 3.327 70.04 3.745 ;
      RECT 69.995 3.385 70.035 3.745 ;
      RECT 70.025 2.209 70.03 2.395 ;
      RECT 70.02 2.207 70.025 2.388 ;
      RECT 70.01 2.204 70.02 2.378 ;
      RECT 70.005 2.201 70.01 2.363 ;
      RECT 69.99 2.197 70.005 2.356 ;
      RECT 69.985 3.44 69.995 3.745 ;
      RECT 69.985 2.194 69.99 2.351 ;
      RECT 69.97 2.19 69.985 2.345 ;
      RECT 69.98 3.457 69.985 3.745 ;
      RECT 69.97 3.52 69.98 3.745 ;
      RECT 69.89 2.175 69.97 2.325 ;
      RECT 69.965 3.527 69.97 3.74 ;
      RECT 69.96 3.535 69.965 3.73 ;
      RECT 69.88 2.161 69.89 2.309 ;
      RECT 69.865 2.157 69.88 2.307 ;
      RECT 69.855 2.152 69.865 2.303 ;
      RECT 69.83 2.145 69.855 2.295 ;
      RECT 69.825 2.14 69.83 2.29 ;
      RECT 69.815 2.14 69.825 2.288 ;
      RECT 69.805 2.138 69.815 2.286 ;
      RECT 69.775 2.13 69.805 2.28 ;
      RECT 69.76 2.122 69.775 2.273 ;
      RECT 69.74 2.117 69.76 2.266 ;
      RECT 69.735 2.113 69.74 2.261 ;
      RECT 69.705 2.106 69.735 2.255 ;
      RECT 69.68 2.097 69.705 2.245 ;
      RECT 69.65 2.09 69.68 2.237 ;
      RECT 69.625 2.08 69.65 2.228 ;
      RECT 69.61 2.072 69.625 2.222 ;
      RECT 69.585 2.067 69.61 2.217 ;
      RECT 69.575 2.063 69.585 2.212 ;
      RECT 69.555 2.058 69.575 2.207 ;
      RECT 69.52 2.053 69.555 2.2 ;
      RECT 69.46 2.048 69.52 2.193 ;
      RECT 69.447 2.044 69.46 2.191 ;
      RECT 69.361 2.039 69.447 2.188 ;
      RECT 69.275 2.029 69.361 2.184 ;
      RECT 69.234 2.022 69.275 2.181 ;
      RECT 69.148 2.015 69.234 2.178 ;
      RECT 69.062 2.005 69.148 2.174 ;
      RECT 68.976 1.995 69.062 2.169 ;
      RECT 68.89 1.985 68.976 2.165 ;
      RECT 68.88 1.97 68.89 2.163 ;
      RECT 68.87 1.955 68.88 2.163 ;
      RECT 68.805 1.95 68.87 2.162 ;
      RECT 68.64 1.947 68.685 2.155 ;
      RECT 69.885 2.852 69.89 3.043 ;
      RECT 69.88 2.847 69.885 3.05 ;
      RECT 69.866 2.845 69.88 3.056 ;
      RECT 69.78 2.845 69.866 3.058 ;
      RECT 69.776 2.845 69.78 3.061 ;
      RECT 69.69 2.845 69.776 3.079 ;
      RECT 69.68 2.85 69.69 3.098 ;
      RECT 69.67 2.905 69.68 3.102 ;
      RECT 69.645 2.92 69.67 3.109 ;
      RECT 69.605 2.94 69.645 3.122 ;
      RECT 69.6 2.952 69.605 3.132 ;
      RECT 69.585 2.958 69.6 3.137 ;
      RECT 69.58 2.963 69.585 3.141 ;
      RECT 69.56 2.97 69.58 3.146 ;
      RECT 69.49 2.995 69.56 3.163 ;
      RECT 69.45 3.023 69.49 3.183 ;
      RECT 69.445 3.033 69.45 3.191 ;
      RECT 69.425 3.04 69.445 3.193 ;
      RECT 69.42 3.047 69.425 3.196 ;
      RECT 69.39 3.055 69.42 3.199 ;
      RECT 69.385 3.06 69.39 3.203 ;
      RECT 69.311 3.064 69.385 3.211 ;
      RECT 69.225 3.073 69.311 3.227 ;
      RECT 69.221 3.078 69.225 3.236 ;
      RECT 69.135 3.083 69.221 3.246 ;
      RECT 69.095 3.091 69.135 3.258 ;
      RECT 69.045 3.097 69.095 3.265 ;
      RECT 68.96 3.106 69.045 3.28 ;
      RECT 68.885 3.117 68.96 3.298 ;
      RECT 68.85 3.124 68.885 3.308 ;
      RECT 68.775 3.132 68.85 3.313 ;
      RECT 68.72 3.141 68.775 3.313 ;
      RECT 68.695 3.146 68.72 3.311 ;
      RECT 68.685 3.149 68.695 3.309 ;
      RECT 68.65 3.151 68.685 3.307 ;
      RECT 68.62 3.153 68.65 3.303 ;
      RECT 68.575 3.152 68.62 3.299 ;
      RECT 68.555 3.147 68.575 3.296 ;
      RECT 68.505 3.132 68.555 3.293 ;
      RECT 68.495 3.117 68.505 3.288 ;
      RECT 68.445 3.102 68.495 3.278 ;
      RECT 68.395 3.077 68.445 3.258 ;
      RECT 68.385 3.062 68.395 3.24 ;
      RECT 68.38 3.06 68.385 3.234 ;
      RECT 68.36 3.055 68.38 3.229 ;
      RECT 68.355 3.047 68.36 3.223 ;
      RECT 68.34 3.041 68.355 3.216 ;
      RECT 68.335 3.036 68.34 3.208 ;
      RECT 68.315 3.031 68.335 3.2 ;
      RECT 68.3 3.024 68.315 3.193 ;
      RECT 68.285 3.018 68.3 3.184 ;
      RECT 68.28 3.012 68.285 3.177 ;
      RECT 68.235 2.987 68.28 3.163 ;
      RECT 68.22 2.957 68.235 3.145 ;
      RECT 68.205 2.94 68.22 3.136 ;
      RECT 68.18 2.92 68.205 3.124 ;
      RECT 68.14 2.89 68.18 3.104 ;
      RECT 68.13 2.86 68.14 3.089 ;
      RECT 68.115 2.85 68.13 3.082 ;
      RECT 68.06 2.815 68.115 3.061 ;
      RECT 68.045 2.778 68.06 3.04 ;
      RECT 68.035 2.765 68.045 3.032 ;
      RECT 67.985 2.735 68.035 3.014 ;
      RECT 67.97 2.665 67.985 2.995 ;
      RECT 67.925 2.665 67.97 2.978 ;
      RECT 67.9 2.665 67.925 2.96 ;
      RECT 67.89 2.665 67.9 2.953 ;
      RECT 67.811 2.665 67.89 2.946 ;
      RECT 67.725 2.665 67.811 2.938 ;
      RECT 67.71 2.697 67.725 2.933 ;
      RECT 67.635 2.707 67.71 2.929 ;
      RECT 67.615 2.717 67.635 2.924 ;
      RECT 67.59 2.717 67.615 2.921 ;
      RECT 67.58 2.707 67.59 2.92 ;
      RECT 67.57 2.68 67.58 2.919 ;
      RECT 67.53 2.675 67.57 2.917 ;
      RECT 67.485 2.675 67.53 2.913 ;
      RECT 67.46 2.675 67.485 2.908 ;
      RECT 67.41 2.675 67.46 2.895 ;
      RECT 67.37 2.68 67.38 2.88 ;
      RECT 67.38 2.675 67.41 2.885 ;
      RECT 69.365 2.455 69.625 2.715 ;
      RECT 69.36 2.477 69.625 2.673 ;
      RECT 68.6 2.305 68.82 2.67 ;
      RECT 68.582 2.392 68.82 2.669 ;
      RECT 68.565 2.397 68.82 2.666 ;
      RECT 68.565 2.397 68.84 2.665 ;
      RECT 68.535 2.407 68.84 2.663 ;
      RECT 68.53 2.422 68.84 2.659 ;
      RECT 68.53 2.422 68.845 2.658 ;
      RECT 68.525 2.48 68.845 2.656 ;
      RECT 68.525 2.48 68.855 2.653 ;
      RECT 68.52 2.545 68.855 2.648 ;
      RECT 68.6 2.305 68.86 2.565 ;
      RECT 67.345 2.135 67.605 2.395 ;
      RECT 67.345 2.178 67.691 2.369 ;
      RECT 67.345 2.178 67.735 2.368 ;
      RECT 67.345 2.178 67.755 2.366 ;
      RECT 67.345 2.178 67.855 2.365 ;
      RECT 67.345 2.178 67.875 2.363 ;
      RECT 67.345 2.178 67.885 2.358 ;
      RECT 67.755 2.145 67.945 2.355 ;
      RECT 67.755 2.147 67.95 2.353 ;
      RECT 67.745 2.152 67.955 2.345 ;
      RECT 67.691 2.176 67.955 2.345 ;
      RECT 67.735 2.17 67.745 2.367 ;
      RECT 67.745 2.15 67.95 2.353 ;
      RECT 66.7 3.21 66.905 3.44 ;
      RECT 66.64 3.16 66.695 3.42 ;
      RECT 66.7 3.16 66.9 3.44 ;
      RECT 67.67 3.475 67.675 3.502 ;
      RECT 67.66 3.385 67.67 3.507 ;
      RECT 67.655 3.307 67.66 3.513 ;
      RECT 67.645 3.297 67.655 3.52 ;
      RECT 67.64 3.287 67.645 3.526 ;
      RECT 67.63 3.282 67.64 3.528 ;
      RECT 67.615 3.274 67.63 3.536 ;
      RECT 67.6 3.265 67.615 3.548 ;
      RECT 67.59 3.257 67.6 3.558 ;
      RECT 67.555 3.175 67.59 3.576 ;
      RECT 67.52 3.175 67.555 3.595 ;
      RECT 67.505 3.175 67.52 3.603 ;
      RECT 67.45 3.175 67.505 3.603 ;
      RECT 67.416 3.175 67.45 3.594 ;
      RECT 67.33 3.175 67.416 3.57 ;
      RECT 67.32 3.235 67.33 3.552 ;
      RECT 67.28 3.237 67.32 3.543 ;
      RECT 67.275 3.239 67.28 3.533 ;
      RECT 67.255 3.241 67.275 3.528 ;
      RECT 67.245 3.244 67.255 3.523 ;
      RECT 67.235 3.245 67.245 3.518 ;
      RECT 67.211 3.246 67.235 3.51 ;
      RECT 67.125 3.251 67.211 3.488 ;
      RECT 67.07 3.25 67.125 3.461 ;
      RECT 67.055 3.243 67.07 3.448 ;
      RECT 67.02 3.238 67.055 3.444 ;
      RECT 66.965 3.23 67.02 3.443 ;
      RECT 66.905 3.217 66.965 3.441 ;
      RECT 66.695 3.16 66.7 3.428 ;
      RECT 66.77 2.53 66.955 2.74 ;
      RECT 66.76 2.535 66.97 2.733 ;
      RECT 66.8 2.44 67.06 2.7 ;
      RECT 66.755 2.597 67.06 2.623 ;
      RECT 66.1 2.39 66.105 3.19 ;
      RECT 66.045 2.44 66.075 3.19 ;
      RECT 66.035 2.44 66.04 2.75 ;
      RECT 66.02 2.44 66.025 2.745 ;
      RECT 65.565 2.485 65.58 2.7 ;
      RECT 65.495 2.485 65.58 2.695 ;
      RECT 66.76 2.065 66.83 2.275 ;
      RECT 66.83 2.072 66.84 2.27 ;
      RECT 66.726 2.065 66.76 2.282 ;
      RECT 66.64 2.065 66.726 2.306 ;
      RECT 66.63 2.07 66.64 2.325 ;
      RECT 66.625 2.082 66.63 2.328 ;
      RECT 66.61 2.097 66.625 2.332 ;
      RECT 66.605 2.115 66.61 2.336 ;
      RECT 66.565 2.125 66.605 2.345 ;
      RECT 66.55 2.132 66.565 2.357 ;
      RECT 66.535 2.137 66.55 2.362 ;
      RECT 66.52 2.14 66.535 2.367 ;
      RECT 66.51 2.142 66.52 2.371 ;
      RECT 66.475 2.149 66.51 2.379 ;
      RECT 66.44 2.157 66.475 2.393 ;
      RECT 66.43 2.163 66.44 2.402 ;
      RECT 66.425 2.165 66.43 2.404 ;
      RECT 66.405 2.168 66.425 2.41 ;
      RECT 66.375 2.175 66.405 2.421 ;
      RECT 66.365 2.181 66.375 2.428 ;
      RECT 66.34 2.184 66.365 2.435 ;
      RECT 66.33 2.188 66.34 2.443 ;
      RECT 66.325 2.189 66.33 2.465 ;
      RECT 66.32 2.19 66.325 2.48 ;
      RECT 66.315 2.191 66.32 2.495 ;
      RECT 66.31 2.192 66.315 2.51 ;
      RECT 66.305 2.193 66.31 2.54 ;
      RECT 66.295 2.195 66.305 2.573 ;
      RECT 66.28 2.199 66.295 2.62 ;
      RECT 66.27 2.202 66.28 2.665 ;
      RECT 66.265 2.205 66.27 2.693 ;
      RECT 66.255 2.207 66.265 2.72 ;
      RECT 66.25 2.21 66.255 2.755 ;
      RECT 66.22 2.215 66.25 2.813 ;
      RECT 66.215 2.22 66.22 2.898 ;
      RECT 66.21 2.222 66.215 2.933 ;
      RECT 66.205 2.224 66.21 3.015 ;
      RECT 66.2 2.226 66.205 3.103 ;
      RECT 66.19 2.228 66.2 3.185 ;
      RECT 66.175 2.242 66.19 3.19 ;
      RECT 66.14 2.287 66.175 3.19 ;
      RECT 66.13 2.327 66.14 3.19 ;
      RECT 66.115 2.355 66.13 3.19 ;
      RECT 66.11 2.372 66.115 3.19 ;
      RECT 66.105 2.38 66.11 3.19 ;
      RECT 66.095 2.395 66.1 3.19 ;
      RECT 66.09 2.402 66.095 3.19 ;
      RECT 66.08 2.422 66.09 3.19 ;
      RECT 66.075 2.435 66.08 3.19 ;
      RECT 66.04 2.44 66.045 2.775 ;
      RECT 66.025 2.83 66.045 3.19 ;
      RECT 66.025 2.44 66.035 2.748 ;
      RECT 66.02 2.87 66.025 3.19 ;
      RECT 65.97 2.44 66.02 2.743 ;
      RECT 66.015 2.907 66.02 3.19 ;
      RECT 66.005 2.93 66.015 3.19 ;
      RECT 66 2.975 66.005 3.19 ;
      RECT 65.99 2.985 66 3.183 ;
      RECT 65.916 2.44 65.97 2.737 ;
      RECT 65.83 2.44 65.916 2.73 ;
      RECT 65.781 2.487 65.83 2.723 ;
      RECT 65.695 2.495 65.781 2.716 ;
      RECT 65.68 2.492 65.695 2.711 ;
      RECT 65.666 2.485 65.68 2.71 ;
      RECT 65.58 2.485 65.666 2.705 ;
      RECT 65.485 2.49 65.495 2.69 ;
      RECT 65.075 1.92 65.09 2.32 ;
      RECT 65.27 1.92 65.275 2.18 ;
      RECT 65.015 1.92 65.06 2.18 ;
      RECT 65.47 3.225 65.475 3.43 ;
      RECT 65.465 3.215 65.47 3.435 ;
      RECT 65.46 3.202 65.465 3.44 ;
      RECT 65.455 3.182 65.46 3.44 ;
      RECT 65.43 3.135 65.455 3.44 ;
      RECT 65.395 3.05 65.43 3.44 ;
      RECT 65.39 2.987 65.395 3.44 ;
      RECT 65.385 2.972 65.39 3.44 ;
      RECT 65.37 2.932 65.385 3.44 ;
      RECT 65.365 2.907 65.37 3.44 ;
      RECT 65.355 2.89 65.365 3.44 ;
      RECT 65.32 2.812 65.355 3.44 ;
      RECT 65.315 2.755 65.32 3.44 ;
      RECT 65.31 2.742 65.315 3.44 ;
      RECT 65.3 2.72 65.31 3.44 ;
      RECT 65.29 2.685 65.3 3.44 ;
      RECT 65.28 2.655 65.29 3.44 ;
      RECT 65.27 2.57 65.28 3.083 ;
      RECT 65.277 3.215 65.28 3.44 ;
      RECT 65.275 3.225 65.277 3.44 ;
      RECT 65.265 3.235 65.275 3.435 ;
      RECT 65.26 1.92 65.27 2.315 ;
      RECT 65.265 2.447 65.27 3.058 ;
      RECT 65.26 2.345 65.265 3.041 ;
      RECT 65.25 1.92 65.26 3.017 ;
      RECT 65.245 1.92 65.25 2.988 ;
      RECT 65.24 1.92 65.245 2.978 ;
      RECT 65.22 1.92 65.24 2.94 ;
      RECT 65.215 1.92 65.22 2.898 ;
      RECT 65.21 1.92 65.215 2.878 ;
      RECT 65.18 1.92 65.21 2.828 ;
      RECT 65.17 1.92 65.18 2.775 ;
      RECT 65.165 1.92 65.17 2.748 ;
      RECT 65.16 1.92 65.165 2.733 ;
      RECT 65.15 1.92 65.16 2.71 ;
      RECT 65.14 1.92 65.15 2.685 ;
      RECT 65.135 1.92 65.14 2.625 ;
      RECT 65.125 1.92 65.135 2.563 ;
      RECT 65.12 1.92 65.125 2.483 ;
      RECT 65.115 1.92 65.12 2.448 ;
      RECT 65.11 1.92 65.115 2.423 ;
      RECT 65.105 1.92 65.11 2.408 ;
      RECT 65.1 1.92 65.105 2.378 ;
      RECT 65.095 1.92 65.1 2.355 ;
      RECT 65.09 1.92 65.095 2.328 ;
      RECT 65.06 1.92 65.075 2.315 ;
      RECT 64.215 3.455 64.4 3.665 ;
      RECT 64.205 3.46 64.415 3.658 ;
      RECT 64.205 3.46 64.435 3.63 ;
      RECT 64.205 3.46 64.45 3.609 ;
      RECT 64.205 3.46 64.465 3.607 ;
      RECT 64.205 3.46 64.475 3.606 ;
      RECT 64.205 3.46 64.505 3.603 ;
      RECT 64.855 3.305 65.115 3.565 ;
      RECT 64.815 3.352 65.115 3.548 ;
      RECT 64.806 3.36 64.815 3.551 ;
      RECT 64.4 3.453 65.115 3.548 ;
      RECT 64.72 3.378 64.806 3.558 ;
      RECT 64.415 3.45 65.115 3.548 ;
      RECT 64.661 3.4 64.72 3.57 ;
      RECT 64.435 3.446 65.115 3.548 ;
      RECT 64.575 3.412 64.661 3.581 ;
      RECT 64.45 3.442 65.115 3.548 ;
      RECT 64.52 3.425 64.575 3.593 ;
      RECT 64.465 3.44 65.115 3.548 ;
      RECT 64.505 3.431 64.52 3.599 ;
      RECT 64.475 3.436 65.115 3.548 ;
      RECT 64.62 2.96 64.88 3.22 ;
      RECT 64.62 2.98 64.99 3.19 ;
      RECT 64.62 2.985 65 3.185 ;
      RECT 64.811 2.399 64.89 2.63 ;
      RECT 64.725 2.402 64.94 2.625 ;
      RECT 64.72 2.402 64.94 2.62 ;
      RECT 64.72 2.407 64.95 2.618 ;
      RECT 64.695 2.407 64.95 2.615 ;
      RECT 64.695 2.415 64.96 2.613 ;
      RECT 64.575 2.35 64.835 2.61 ;
      RECT 64.575 2.397 64.885 2.61 ;
      RECT 63.83 2.97 63.835 3.23 ;
      RECT 63.66 2.74 63.665 3.23 ;
      RECT 63.545 2.98 63.55 3.205 ;
      RECT 64.255 2.075 64.26 2.285 ;
      RECT 64.26 2.08 64.275 2.28 ;
      RECT 64.195 2.075 64.255 2.293 ;
      RECT 64.18 2.075 64.195 2.303 ;
      RECT 64.13 2.075 64.18 2.32 ;
      RECT 64.11 2.075 64.13 2.343 ;
      RECT 64.095 2.075 64.11 2.355 ;
      RECT 64.075 2.075 64.095 2.365 ;
      RECT 64.065 2.08 64.075 2.374 ;
      RECT 64.06 2.09 64.065 2.379 ;
      RECT 64.055 2.102 64.06 2.383 ;
      RECT 64.045 2.125 64.055 2.388 ;
      RECT 64.04 2.14 64.045 2.392 ;
      RECT 64.035 2.157 64.04 2.395 ;
      RECT 64.03 2.165 64.035 2.398 ;
      RECT 64.02 2.17 64.03 2.402 ;
      RECT 64.015 2.177 64.02 2.407 ;
      RECT 64.005 2.182 64.015 2.411 ;
      RECT 63.98 2.194 64.005 2.422 ;
      RECT 63.96 2.211 63.98 2.438 ;
      RECT 63.935 2.228 63.96 2.46 ;
      RECT 63.9 2.251 63.935 2.518 ;
      RECT 63.88 2.273 63.9 2.58 ;
      RECT 63.875 2.283 63.88 2.615 ;
      RECT 63.865 2.29 63.875 2.653 ;
      RECT 63.86 2.297 63.865 2.673 ;
      RECT 63.855 2.308 63.86 2.71 ;
      RECT 63.85 2.316 63.855 2.775 ;
      RECT 63.84 2.327 63.85 2.828 ;
      RECT 63.835 2.345 63.84 2.898 ;
      RECT 63.83 2.355 63.835 2.935 ;
      RECT 63.825 2.365 63.83 3.23 ;
      RECT 63.82 2.377 63.825 3.23 ;
      RECT 63.815 2.387 63.82 3.23 ;
      RECT 63.805 2.397 63.815 3.23 ;
      RECT 63.795 2.42 63.805 3.23 ;
      RECT 63.78 2.455 63.795 3.23 ;
      RECT 63.74 2.517 63.78 3.23 ;
      RECT 63.735 2.57 63.74 3.23 ;
      RECT 63.71 2.605 63.735 3.23 ;
      RECT 63.695 2.65 63.71 3.23 ;
      RECT 63.69 2.672 63.695 3.23 ;
      RECT 63.68 2.685 63.69 3.23 ;
      RECT 63.67 2.71 63.68 3.23 ;
      RECT 63.665 2.732 63.67 3.23 ;
      RECT 63.64 2.77 63.66 3.23 ;
      RECT 63.6 2.827 63.64 3.23 ;
      RECT 63.595 2.877 63.6 3.23 ;
      RECT 63.59 2.895 63.595 3.23 ;
      RECT 63.585 2.907 63.59 3.23 ;
      RECT 63.575 2.925 63.585 3.23 ;
      RECT 63.565 2.945 63.575 3.205 ;
      RECT 63.56 2.962 63.565 3.205 ;
      RECT 63.55 2.975 63.56 3.205 ;
      RECT 63.52 2.985 63.545 3.205 ;
      RECT 63.51 2.992 63.52 3.205 ;
      RECT 63.495 3.002 63.51 3.2 ;
      RECT 62.59 7.765 62.88 7.995 ;
      RECT 62.65 6.285 62.82 7.995 ;
      RECT 62.595 6.655 62.945 7.005 ;
      RECT 62.59 6.285 62.88 6.515 ;
      RECT 62.59 2.365 62.88 2.595 ;
      RECT 62.65 0.885 62.82 2.595 ;
      RECT 62.59 0.885 62.88 1.115 ;
      RECT 62.18 2.735 62.51 2.965 ;
      RECT 62.18 2.765 62.68 2.935 ;
      RECT 62.18 2.395 62.37 2.965 ;
      RECT 61.6 2.365 61.89 2.595 ;
      RECT 61.6 2.395 62.37 2.565 ;
      RECT 61.66 0.885 61.83 2.595 ;
      RECT 61.6 0.885 61.89 1.115 ;
      RECT 61.6 7.765 61.89 7.995 ;
      RECT 61.66 6.285 61.83 7.995 ;
      RECT 61.6 6.285 61.89 6.515 ;
      RECT 61.6 6.325 62.45 6.485 ;
      RECT 62.28 5.915 62.45 6.485 ;
      RECT 61.6 6.32 61.99 6.485 ;
      RECT 62.22 5.915 62.51 6.145 ;
      RECT 62.22 5.945 62.68 6.115 ;
      RECT 61.23 2.735 61.52 2.965 ;
      RECT 61.23 2.765 61.69 2.935 ;
      RECT 61.29 1.655 61.455 2.965 ;
      RECT 59.805 1.625 60.095 1.855 ;
      RECT 59.805 1.655 61.455 1.825 ;
      RECT 59.865 0.885 60.035 1.855 ;
      RECT 59.805 0.885 60.095 1.115 ;
      RECT 59.805 7.765 60.095 7.995 ;
      RECT 59.865 7.025 60.035 7.995 ;
      RECT 59.865 7.12 61.455 7.29 ;
      RECT 61.285 5.915 61.455 7.29 ;
      RECT 59.805 7.025 60.095 7.255 ;
      RECT 61.23 5.915 61.52 6.145 ;
      RECT 61.23 5.945 61.69 6.115 ;
      RECT 60.235 1.965 60.585 2.315 ;
      RECT 57.9 2.025 60.585 2.195 ;
      RECT 57.9 1.34 58.07 2.195 ;
      RECT 57.8 1.34 58.15 1.69 ;
      RECT 60.26 6.655 60.585 6.98 ;
      RECT 55.635 6.61 55.985 6.96 ;
      RECT 60.235 6.655 60.585 6.885 ;
      RECT 55.455 6.655 55.985 6.885 ;
      RECT 55.285 6.685 60.585 6.855 ;
      RECT 59.46 2.365 59.78 2.685 ;
      RECT 59.43 2.365 59.78 2.595 ;
      RECT 59.26 2.395 59.78 2.565 ;
      RECT 59.46 6.255 59.78 6.545 ;
      RECT 59.43 6.285 59.78 6.515 ;
      RECT 59.26 6.315 59.78 6.485 ;
      RECT 58.405 2.705 58.755 3.055 ;
      RECT 58.405 2.765 58.895 2.935 ;
      RECT 58.41 5.855 58.76 6.205 ;
      RECT 53.655 5.915 53.945 6.145 ;
      RECT 53.655 5.945 58.895 6.115 ;
      RECT 56.095 2.465 56.28 2.675 ;
      RECT 56.085 2.47 56.295 2.668 ;
      RECT 56.085 2.47 56.381 2.645 ;
      RECT 56.085 2.47 56.44 2.62 ;
      RECT 56.085 2.47 56.495 2.6 ;
      RECT 56.085 2.47 56.505 2.588 ;
      RECT 56.085 2.47 56.7 2.527 ;
      RECT 56.085 2.47 56.73 2.51 ;
      RECT 56.085 2.47 56.75 2.5 ;
      RECT 56.63 2.235 56.89 2.495 ;
      RECT 56.615 2.325 56.63 2.542 ;
      RECT 56.15 2.457 56.89 2.495 ;
      RECT 56.601 2.336 56.615 2.548 ;
      RECT 56.19 2.45 56.89 2.495 ;
      RECT 56.515 2.376 56.601 2.567 ;
      RECT 56.44 2.437 56.89 2.495 ;
      RECT 56.51 2.412 56.515 2.584 ;
      RECT 56.495 2.422 56.89 2.495 ;
      RECT 56.505 2.417 56.51 2.586 ;
      RECT 56.8 2.922 56.805 3.014 ;
      RECT 56.795 2.9 56.8 3.031 ;
      RECT 56.79 2.89 56.795 3.043 ;
      RECT 56.78 2.881 56.79 3.053 ;
      RECT 56.775 2.876 56.78 3.061 ;
      RECT 56.77 2.735 56.775 3.064 ;
      RECT 56.736 2.735 56.77 3.075 ;
      RECT 56.65 2.735 56.736 3.11 ;
      RECT 56.57 2.735 56.65 3.158 ;
      RECT 56.541 2.735 56.57 3.182 ;
      RECT 56.455 2.735 56.541 3.188 ;
      RECT 56.45 2.919 56.455 3.193 ;
      RECT 56.415 2.93 56.45 3.196 ;
      RECT 56.39 2.945 56.415 3.2 ;
      RECT 56.376 2.954 56.39 3.202 ;
      RECT 56.29 2.981 56.376 3.208 ;
      RECT 56.225 3.022 56.29 3.217 ;
      RECT 56.21 3.042 56.225 3.222 ;
      RECT 56.18 3.052 56.21 3.225 ;
      RECT 56.175 3.062 56.18 3.228 ;
      RECT 56.145 3.067 56.175 3.23 ;
      RECT 56.125 3.072 56.145 3.234 ;
      RECT 56.04 3.075 56.125 3.241 ;
      RECT 56.025 3.072 56.04 3.247 ;
      RECT 56.015 3.069 56.025 3.249 ;
      RECT 55.995 3.066 56.015 3.251 ;
      RECT 55.975 3.062 55.995 3.252 ;
      RECT 55.96 3.058 55.975 3.254 ;
      RECT 55.95 3.055 55.96 3.255 ;
      RECT 55.91 3.049 55.95 3.253 ;
      RECT 55.9 3.044 55.91 3.251 ;
      RECT 55.885 3.041 55.9 3.247 ;
      RECT 55.86 3.036 55.885 3.24 ;
      RECT 55.81 3.027 55.86 3.228 ;
      RECT 55.74 3.013 55.81 3.21 ;
      RECT 55.682 2.998 55.74 3.192 ;
      RECT 55.596 2.981 55.682 3.172 ;
      RECT 55.51 2.96 55.596 3.147 ;
      RECT 55.46 2.945 55.51 3.128 ;
      RECT 55.456 2.939 55.46 3.12 ;
      RECT 55.37 2.929 55.456 3.107 ;
      RECT 55.335 2.914 55.37 3.09 ;
      RECT 55.32 2.907 55.335 3.083 ;
      RECT 55.26 2.895 55.32 3.071 ;
      RECT 55.24 2.882 55.26 3.059 ;
      RECT 55.2 2.873 55.24 3.051 ;
      RECT 55.195 2.865 55.2 3.044 ;
      RECT 55.115 2.855 55.195 3.03 ;
      RECT 55.1 2.842 55.115 3.015 ;
      RECT 55.095 2.84 55.1 3.013 ;
      RECT 55.016 2.828 55.095 3 ;
      RECT 54.93 2.803 55.016 2.975 ;
      RECT 54.915 2.772 54.93 2.96 ;
      RECT 54.9 2.747 54.915 2.956 ;
      RECT 54.885 2.74 54.9 2.952 ;
      RECT 54.71 2.745 54.715 2.948 ;
      RECT 54.705 2.75 54.71 2.943 ;
      RECT 54.715 2.74 54.885 2.95 ;
      RECT 55.43 2.5 55.535 2.76 ;
      RECT 56.245 2.025 56.25 2.25 ;
      RECT 56.375 2.025 56.43 2.235 ;
      RECT 56.43 2.03 56.44 2.228 ;
      RECT 56.336 2.025 56.375 2.238 ;
      RECT 56.25 2.025 56.336 2.245 ;
      RECT 56.23 2.03 56.245 2.251 ;
      RECT 56.22 2.07 56.23 2.253 ;
      RECT 56.19 2.08 56.22 2.255 ;
      RECT 56.185 2.085 56.19 2.257 ;
      RECT 56.16 2.09 56.185 2.259 ;
      RECT 56.145 2.095 56.16 2.261 ;
      RECT 56.13 2.097 56.145 2.263 ;
      RECT 56.125 2.102 56.13 2.265 ;
      RECT 56.075 2.11 56.125 2.268 ;
      RECT 56.05 2.119 56.075 2.273 ;
      RECT 56.04 2.126 56.05 2.278 ;
      RECT 56.035 2.129 56.04 2.282 ;
      RECT 56.015 2.132 56.035 2.291 ;
      RECT 55.985 2.14 56.015 2.311 ;
      RECT 55.956 2.153 55.985 2.333 ;
      RECT 55.87 2.187 55.956 2.377 ;
      RECT 55.865 2.213 55.87 2.415 ;
      RECT 55.86 2.217 55.865 2.424 ;
      RECT 55.825 2.23 55.86 2.457 ;
      RECT 55.815 2.244 55.825 2.495 ;
      RECT 55.81 2.248 55.815 2.508 ;
      RECT 55.805 2.252 55.81 2.513 ;
      RECT 55.795 2.26 55.805 2.525 ;
      RECT 55.79 2.267 55.795 2.54 ;
      RECT 55.765 2.28 55.79 2.565 ;
      RECT 55.725 2.309 55.765 2.62 ;
      RECT 55.71 2.334 55.725 2.675 ;
      RECT 55.7 2.345 55.71 2.698 ;
      RECT 55.695 2.352 55.7 2.71 ;
      RECT 55.69 2.356 55.695 2.718 ;
      RECT 55.635 2.384 55.69 2.76 ;
      RECT 55.615 2.42 55.635 2.76 ;
      RECT 55.6 2.435 55.615 2.76 ;
      RECT 55.545 2.467 55.6 2.76 ;
      RECT 55.535 2.497 55.545 2.76 ;
      RECT 55.145 2.112 55.33 2.35 ;
      RECT 55.13 2.114 55.34 2.345 ;
      RECT 55.015 2.06 55.275 2.32 ;
      RECT 55.01 2.097 55.275 2.274 ;
      RECT 55.005 2.107 55.275 2.271 ;
      RECT 55 2.147 55.34 2.265 ;
      RECT 54.995 2.18 55.34 2.255 ;
      RECT 55.005 2.122 55.355 2.193 ;
      RECT 55.302 3.22 55.315 3.75 ;
      RECT 55.216 3.22 55.315 3.749 ;
      RECT 55.216 3.22 55.32 3.748 ;
      RECT 55.13 3.22 55.32 3.746 ;
      RECT 55.125 3.22 55.32 3.743 ;
      RECT 55.125 3.22 55.33 3.741 ;
      RECT 55.12 3.512 55.33 3.738 ;
      RECT 55.12 3.522 55.335 3.735 ;
      RECT 55.12 3.59 55.34 3.731 ;
      RECT 55.11 3.595 55.34 3.73 ;
      RECT 55.11 3.687 55.345 3.727 ;
      RECT 55.095 3.22 55.355 3.48 ;
      RECT 55.025 7.765 55.315 7.995 ;
      RECT 55.085 7.025 55.255 7.995 ;
      RECT 55 7.055 55.34 7.4 ;
      RECT 55.025 7.025 55.315 7.4 ;
      RECT 54.325 2.21 54.37 3.745 ;
      RECT 54.525 2.21 54.555 2.425 ;
      RECT 52.9 1.95 53.02 2.16 ;
      RECT 52.56 1.9 52.82 2.16 ;
      RECT 52.56 1.945 52.855 2.15 ;
      RECT 54.565 2.226 54.57 2.28 ;
      RECT 54.56 2.219 54.565 2.413 ;
      RECT 54.555 2.213 54.56 2.42 ;
      RECT 54.51 2.21 54.525 2.433 ;
      RECT 54.505 2.21 54.51 2.455 ;
      RECT 54.5 2.21 54.505 2.503 ;
      RECT 54.495 2.21 54.5 2.523 ;
      RECT 54.485 2.21 54.495 2.63 ;
      RECT 54.48 2.21 54.485 2.693 ;
      RECT 54.475 2.21 54.48 2.75 ;
      RECT 54.47 2.21 54.475 2.758 ;
      RECT 54.455 2.21 54.47 2.865 ;
      RECT 54.445 2.21 54.455 3 ;
      RECT 54.435 2.21 54.445 3.11 ;
      RECT 54.425 2.21 54.435 3.167 ;
      RECT 54.42 2.21 54.425 3.207 ;
      RECT 54.415 2.21 54.42 3.243 ;
      RECT 54.405 2.21 54.415 3.283 ;
      RECT 54.4 2.21 54.405 3.325 ;
      RECT 54.38 2.21 54.4 3.39 ;
      RECT 54.385 3.535 54.39 3.715 ;
      RECT 54.38 3.517 54.385 3.723 ;
      RECT 54.375 2.21 54.38 3.453 ;
      RECT 54.375 3.497 54.38 3.73 ;
      RECT 54.37 2.21 54.375 3.74 ;
      RECT 54.315 2.21 54.325 2.51 ;
      RECT 54.32 2.757 54.325 3.745 ;
      RECT 54.315 2.822 54.32 3.745 ;
      RECT 54.31 2.211 54.315 2.5 ;
      RECT 54.305 2.887 54.315 3.745 ;
      RECT 54.3 2.212 54.31 2.49 ;
      RECT 54.29 3 54.305 3.745 ;
      RECT 54.295 2.213 54.3 2.48 ;
      RECT 54.275 2.214 54.295 2.458 ;
      RECT 54.28 3.097 54.29 3.745 ;
      RECT 54.275 3.172 54.28 3.745 ;
      RECT 54.265 2.213 54.275 2.435 ;
      RECT 54.27 3.215 54.275 3.745 ;
      RECT 54.265 3.242 54.27 3.745 ;
      RECT 54.255 2.211 54.265 2.423 ;
      RECT 54.26 3.285 54.265 3.745 ;
      RECT 54.255 3.312 54.26 3.745 ;
      RECT 54.245 2.21 54.255 2.41 ;
      RECT 54.25 3.327 54.255 3.745 ;
      RECT 54.21 3.385 54.25 3.745 ;
      RECT 54.24 2.209 54.245 2.395 ;
      RECT 54.235 2.207 54.24 2.388 ;
      RECT 54.225 2.204 54.235 2.378 ;
      RECT 54.22 2.201 54.225 2.363 ;
      RECT 54.205 2.197 54.22 2.356 ;
      RECT 54.2 3.44 54.21 3.745 ;
      RECT 54.2 2.194 54.205 2.351 ;
      RECT 54.185 2.19 54.2 2.345 ;
      RECT 54.195 3.457 54.2 3.745 ;
      RECT 54.185 3.52 54.195 3.745 ;
      RECT 54.105 2.175 54.185 2.325 ;
      RECT 54.18 3.527 54.185 3.74 ;
      RECT 54.175 3.535 54.18 3.73 ;
      RECT 54.095 2.161 54.105 2.309 ;
      RECT 54.08 2.157 54.095 2.307 ;
      RECT 54.07 2.152 54.08 2.303 ;
      RECT 54.045 2.145 54.07 2.295 ;
      RECT 54.04 2.14 54.045 2.29 ;
      RECT 54.03 2.14 54.04 2.288 ;
      RECT 54.02 2.138 54.03 2.286 ;
      RECT 53.99 2.13 54.02 2.28 ;
      RECT 53.975 2.122 53.99 2.273 ;
      RECT 53.955 2.117 53.975 2.266 ;
      RECT 53.95 2.113 53.955 2.261 ;
      RECT 53.92 2.106 53.95 2.255 ;
      RECT 53.895 2.097 53.92 2.245 ;
      RECT 53.865 2.09 53.895 2.237 ;
      RECT 53.84 2.08 53.865 2.228 ;
      RECT 53.825 2.072 53.84 2.222 ;
      RECT 53.8 2.067 53.825 2.217 ;
      RECT 53.79 2.063 53.8 2.212 ;
      RECT 53.77 2.058 53.79 2.207 ;
      RECT 53.735 2.053 53.77 2.2 ;
      RECT 53.675 2.048 53.735 2.193 ;
      RECT 53.662 2.044 53.675 2.191 ;
      RECT 53.576 2.039 53.662 2.188 ;
      RECT 53.49 2.029 53.576 2.184 ;
      RECT 53.449 2.022 53.49 2.181 ;
      RECT 53.363 2.015 53.449 2.178 ;
      RECT 53.277 2.005 53.363 2.174 ;
      RECT 53.191 1.995 53.277 2.169 ;
      RECT 53.105 1.985 53.191 2.165 ;
      RECT 53.095 1.97 53.105 2.163 ;
      RECT 53.085 1.955 53.095 2.163 ;
      RECT 53.02 1.95 53.085 2.162 ;
      RECT 52.855 1.947 52.9 2.155 ;
      RECT 54.1 2.852 54.105 3.043 ;
      RECT 54.095 2.847 54.1 3.05 ;
      RECT 54.081 2.845 54.095 3.056 ;
      RECT 53.995 2.845 54.081 3.058 ;
      RECT 53.991 2.845 53.995 3.061 ;
      RECT 53.905 2.845 53.991 3.079 ;
      RECT 53.895 2.85 53.905 3.098 ;
      RECT 53.885 2.905 53.895 3.102 ;
      RECT 53.86 2.92 53.885 3.109 ;
      RECT 53.82 2.94 53.86 3.122 ;
      RECT 53.815 2.952 53.82 3.132 ;
      RECT 53.8 2.958 53.815 3.137 ;
      RECT 53.795 2.963 53.8 3.141 ;
      RECT 53.775 2.97 53.795 3.146 ;
      RECT 53.705 2.995 53.775 3.163 ;
      RECT 53.665 3.023 53.705 3.183 ;
      RECT 53.66 3.033 53.665 3.191 ;
      RECT 53.64 3.04 53.66 3.193 ;
      RECT 53.635 3.047 53.64 3.196 ;
      RECT 53.605 3.055 53.635 3.199 ;
      RECT 53.6 3.06 53.605 3.203 ;
      RECT 53.526 3.064 53.6 3.211 ;
      RECT 53.44 3.073 53.526 3.227 ;
      RECT 53.436 3.078 53.44 3.236 ;
      RECT 53.35 3.083 53.436 3.246 ;
      RECT 53.31 3.091 53.35 3.258 ;
      RECT 53.26 3.097 53.31 3.265 ;
      RECT 53.175 3.106 53.26 3.28 ;
      RECT 53.1 3.117 53.175 3.298 ;
      RECT 53.065 3.124 53.1 3.308 ;
      RECT 52.99 3.132 53.065 3.313 ;
      RECT 52.935 3.141 52.99 3.313 ;
      RECT 52.91 3.146 52.935 3.311 ;
      RECT 52.9 3.149 52.91 3.309 ;
      RECT 52.865 3.151 52.9 3.307 ;
      RECT 52.835 3.153 52.865 3.303 ;
      RECT 52.79 3.152 52.835 3.299 ;
      RECT 52.77 3.147 52.79 3.296 ;
      RECT 52.72 3.132 52.77 3.293 ;
      RECT 52.71 3.117 52.72 3.288 ;
      RECT 52.66 3.102 52.71 3.278 ;
      RECT 52.61 3.077 52.66 3.258 ;
      RECT 52.6 3.062 52.61 3.24 ;
      RECT 52.595 3.06 52.6 3.234 ;
      RECT 52.575 3.055 52.595 3.229 ;
      RECT 52.57 3.047 52.575 3.223 ;
      RECT 52.555 3.041 52.57 3.216 ;
      RECT 52.55 3.036 52.555 3.208 ;
      RECT 52.53 3.031 52.55 3.2 ;
      RECT 52.515 3.024 52.53 3.193 ;
      RECT 52.5 3.018 52.515 3.184 ;
      RECT 52.495 3.012 52.5 3.177 ;
      RECT 52.45 2.987 52.495 3.163 ;
      RECT 52.435 2.957 52.45 3.145 ;
      RECT 52.42 2.94 52.435 3.136 ;
      RECT 52.395 2.92 52.42 3.124 ;
      RECT 52.355 2.89 52.395 3.104 ;
      RECT 52.345 2.86 52.355 3.089 ;
      RECT 52.33 2.85 52.345 3.082 ;
      RECT 52.275 2.815 52.33 3.061 ;
      RECT 52.26 2.778 52.275 3.04 ;
      RECT 52.25 2.765 52.26 3.032 ;
      RECT 52.2 2.735 52.25 3.014 ;
      RECT 52.185 2.665 52.2 2.995 ;
      RECT 52.14 2.665 52.185 2.978 ;
      RECT 52.115 2.665 52.14 2.96 ;
      RECT 52.105 2.665 52.115 2.953 ;
      RECT 52.026 2.665 52.105 2.946 ;
      RECT 51.94 2.665 52.026 2.938 ;
      RECT 51.925 2.697 51.94 2.933 ;
      RECT 51.85 2.707 51.925 2.929 ;
      RECT 51.83 2.717 51.85 2.924 ;
      RECT 51.805 2.717 51.83 2.921 ;
      RECT 51.795 2.707 51.805 2.92 ;
      RECT 51.785 2.68 51.795 2.919 ;
      RECT 51.745 2.675 51.785 2.917 ;
      RECT 51.7 2.675 51.745 2.913 ;
      RECT 51.675 2.675 51.7 2.908 ;
      RECT 51.625 2.675 51.675 2.895 ;
      RECT 51.585 2.68 51.595 2.88 ;
      RECT 51.595 2.675 51.625 2.885 ;
      RECT 53.58 2.455 53.84 2.715 ;
      RECT 53.575 2.477 53.84 2.673 ;
      RECT 52.815 2.305 53.035 2.67 ;
      RECT 52.797 2.392 53.035 2.669 ;
      RECT 52.78 2.397 53.035 2.666 ;
      RECT 52.78 2.397 53.055 2.665 ;
      RECT 52.75 2.407 53.055 2.663 ;
      RECT 52.745 2.422 53.055 2.659 ;
      RECT 52.745 2.422 53.06 2.658 ;
      RECT 52.74 2.48 53.06 2.656 ;
      RECT 52.74 2.48 53.07 2.653 ;
      RECT 52.735 2.545 53.07 2.648 ;
      RECT 52.815 2.305 53.075 2.565 ;
      RECT 51.56 2.135 51.82 2.395 ;
      RECT 51.56 2.178 51.906 2.369 ;
      RECT 51.56 2.178 51.95 2.368 ;
      RECT 51.56 2.178 51.97 2.366 ;
      RECT 51.56 2.178 52.07 2.365 ;
      RECT 51.56 2.178 52.09 2.363 ;
      RECT 51.56 2.178 52.1 2.358 ;
      RECT 51.97 2.145 52.16 2.355 ;
      RECT 51.97 2.147 52.165 2.353 ;
      RECT 51.96 2.152 52.17 2.345 ;
      RECT 51.906 2.176 52.17 2.345 ;
      RECT 51.95 2.17 51.96 2.367 ;
      RECT 51.96 2.15 52.165 2.353 ;
      RECT 50.915 3.21 51.12 3.44 ;
      RECT 50.855 3.16 50.91 3.42 ;
      RECT 50.915 3.16 51.115 3.44 ;
      RECT 51.885 3.475 51.89 3.502 ;
      RECT 51.875 3.385 51.885 3.507 ;
      RECT 51.87 3.307 51.875 3.513 ;
      RECT 51.86 3.297 51.87 3.52 ;
      RECT 51.855 3.287 51.86 3.526 ;
      RECT 51.845 3.282 51.855 3.528 ;
      RECT 51.83 3.274 51.845 3.536 ;
      RECT 51.815 3.265 51.83 3.548 ;
      RECT 51.805 3.257 51.815 3.558 ;
      RECT 51.77 3.175 51.805 3.576 ;
      RECT 51.735 3.175 51.77 3.595 ;
      RECT 51.72 3.175 51.735 3.603 ;
      RECT 51.665 3.175 51.72 3.603 ;
      RECT 51.631 3.175 51.665 3.594 ;
      RECT 51.545 3.175 51.631 3.57 ;
      RECT 51.535 3.235 51.545 3.552 ;
      RECT 51.495 3.237 51.535 3.543 ;
      RECT 51.49 3.239 51.495 3.533 ;
      RECT 51.47 3.241 51.49 3.528 ;
      RECT 51.46 3.244 51.47 3.523 ;
      RECT 51.45 3.245 51.46 3.518 ;
      RECT 51.426 3.246 51.45 3.51 ;
      RECT 51.34 3.251 51.426 3.488 ;
      RECT 51.285 3.25 51.34 3.461 ;
      RECT 51.27 3.243 51.285 3.448 ;
      RECT 51.235 3.238 51.27 3.444 ;
      RECT 51.18 3.23 51.235 3.443 ;
      RECT 51.12 3.217 51.18 3.441 ;
      RECT 50.91 3.16 50.915 3.428 ;
      RECT 50.985 2.53 51.17 2.74 ;
      RECT 50.975 2.535 51.185 2.733 ;
      RECT 51.015 2.44 51.275 2.7 ;
      RECT 50.97 2.597 51.275 2.623 ;
      RECT 50.315 2.39 50.32 3.19 ;
      RECT 50.26 2.44 50.29 3.19 ;
      RECT 50.25 2.44 50.255 2.75 ;
      RECT 50.235 2.44 50.24 2.745 ;
      RECT 49.78 2.485 49.795 2.7 ;
      RECT 49.71 2.485 49.795 2.695 ;
      RECT 50.975 2.065 51.045 2.275 ;
      RECT 51.045 2.072 51.055 2.27 ;
      RECT 50.941 2.065 50.975 2.282 ;
      RECT 50.855 2.065 50.941 2.306 ;
      RECT 50.845 2.07 50.855 2.325 ;
      RECT 50.84 2.082 50.845 2.328 ;
      RECT 50.825 2.097 50.84 2.332 ;
      RECT 50.82 2.115 50.825 2.336 ;
      RECT 50.78 2.125 50.82 2.345 ;
      RECT 50.765 2.132 50.78 2.357 ;
      RECT 50.75 2.137 50.765 2.362 ;
      RECT 50.735 2.14 50.75 2.367 ;
      RECT 50.725 2.142 50.735 2.371 ;
      RECT 50.69 2.149 50.725 2.379 ;
      RECT 50.655 2.157 50.69 2.393 ;
      RECT 50.645 2.163 50.655 2.402 ;
      RECT 50.64 2.165 50.645 2.404 ;
      RECT 50.62 2.168 50.64 2.41 ;
      RECT 50.59 2.175 50.62 2.421 ;
      RECT 50.58 2.181 50.59 2.428 ;
      RECT 50.555 2.184 50.58 2.435 ;
      RECT 50.545 2.188 50.555 2.443 ;
      RECT 50.54 2.189 50.545 2.465 ;
      RECT 50.535 2.19 50.54 2.48 ;
      RECT 50.53 2.191 50.535 2.495 ;
      RECT 50.525 2.192 50.53 2.51 ;
      RECT 50.52 2.193 50.525 2.54 ;
      RECT 50.51 2.195 50.52 2.573 ;
      RECT 50.495 2.199 50.51 2.62 ;
      RECT 50.485 2.202 50.495 2.665 ;
      RECT 50.48 2.205 50.485 2.693 ;
      RECT 50.47 2.207 50.48 2.72 ;
      RECT 50.465 2.21 50.47 2.755 ;
      RECT 50.435 2.215 50.465 2.813 ;
      RECT 50.43 2.22 50.435 2.898 ;
      RECT 50.425 2.222 50.43 2.933 ;
      RECT 50.42 2.224 50.425 3.015 ;
      RECT 50.415 2.226 50.42 3.103 ;
      RECT 50.405 2.228 50.415 3.185 ;
      RECT 50.39 2.242 50.405 3.19 ;
      RECT 50.355 2.287 50.39 3.19 ;
      RECT 50.345 2.327 50.355 3.19 ;
      RECT 50.33 2.355 50.345 3.19 ;
      RECT 50.325 2.372 50.33 3.19 ;
      RECT 50.32 2.38 50.325 3.19 ;
      RECT 50.31 2.395 50.315 3.19 ;
      RECT 50.305 2.402 50.31 3.19 ;
      RECT 50.295 2.422 50.305 3.19 ;
      RECT 50.29 2.435 50.295 3.19 ;
      RECT 50.255 2.44 50.26 2.775 ;
      RECT 50.24 2.83 50.26 3.19 ;
      RECT 50.24 2.44 50.25 2.748 ;
      RECT 50.235 2.87 50.24 3.19 ;
      RECT 50.185 2.44 50.235 2.743 ;
      RECT 50.23 2.907 50.235 3.19 ;
      RECT 50.22 2.93 50.23 3.19 ;
      RECT 50.215 2.975 50.22 3.19 ;
      RECT 50.205 2.985 50.215 3.183 ;
      RECT 50.131 2.44 50.185 2.737 ;
      RECT 50.045 2.44 50.131 2.73 ;
      RECT 49.996 2.487 50.045 2.723 ;
      RECT 49.91 2.495 49.996 2.716 ;
      RECT 49.895 2.492 49.91 2.711 ;
      RECT 49.881 2.485 49.895 2.71 ;
      RECT 49.795 2.485 49.881 2.705 ;
      RECT 49.7 2.49 49.71 2.69 ;
      RECT 49.29 1.92 49.305 2.32 ;
      RECT 49.485 1.92 49.49 2.18 ;
      RECT 49.23 1.92 49.275 2.18 ;
      RECT 49.685 3.225 49.69 3.43 ;
      RECT 49.68 3.215 49.685 3.435 ;
      RECT 49.675 3.202 49.68 3.44 ;
      RECT 49.67 3.182 49.675 3.44 ;
      RECT 49.645 3.135 49.67 3.44 ;
      RECT 49.61 3.05 49.645 3.44 ;
      RECT 49.605 2.987 49.61 3.44 ;
      RECT 49.6 2.972 49.605 3.44 ;
      RECT 49.585 2.932 49.6 3.44 ;
      RECT 49.58 2.907 49.585 3.44 ;
      RECT 49.57 2.89 49.58 3.44 ;
      RECT 49.535 2.812 49.57 3.44 ;
      RECT 49.53 2.755 49.535 3.44 ;
      RECT 49.525 2.742 49.53 3.44 ;
      RECT 49.515 2.72 49.525 3.44 ;
      RECT 49.505 2.685 49.515 3.44 ;
      RECT 49.495 2.655 49.505 3.44 ;
      RECT 49.485 2.57 49.495 3.083 ;
      RECT 49.492 3.215 49.495 3.44 ;
      RECT 49.49 3.225 49.492 3.44 ;
      RECT 49.48 3.235 49.49 3.435 ;
      RECT 49.475 1.92 49.485 2.315 ;
      RECT 49.48 2.447 49.485 3.058 ;
      RECT 49.475 2.345 49.48 3.041 ;
      RECT 49.465 1.92 49.475 3.017 ;
      RECT 49.46 1.92 49.465 2.988 ;
      RECT 49.455 1.92 49.46 2.978 ;
      RECT 49.435 1.92 49.455 2.94 ;
      RECT 49.43 1.92 49.435 2.898 ;
      RECT 49.425 1.92 49.43 2.878 ;
      RECT 49.395 1.92 49.425 2.828 ;
      RECT 49.385 1.92 49.395 2.775 ;
      RECT 49.38 1.92 49.385 2.748 ;
      RECT 49.375 1.92 49.38 2.733 ;
      RECT 49.365 1.92 49.375 2.71 ;
      RECT 49.355 1.92 49.365 2.685 ;
      RECT 49.35 1.92 49.355 2.625 ;
      RECT 49.34 1.92 49.35 2.563 ;
      RECT 49.335 1.92 49.34 2.483 ;
      RECT 49.33 1.92 49.335 2.448 ;
      RECT 49.325 1.92 49.33 2.423 ;
      RECT 49.32 1.92 49.325 2.408 ;
      RECT 49.315 1.92 49.32 2.378 ;
      RECT 49.31 1.92 49.315 2.355 ;
      RECT 49.305 1.92 49.31 2.328 ;
      RECT 49.275 1.92 49.29 2.315 ;
      RECT 48.43 3.455 48.615 3.665 ;
      RECT 48.42 3.46 48.63 3.658 ;
      RECT 48.42 3.46 48.65 3.63 ;
      RECT 48.42 3.46 48.665 3.609 ;
      RECT 48.42 3.46 48.68 3.607 ;
      RECT 48.42 3.46 48.69 3.606 ;
      RECT 48.42 3.46 48.72 3.603 ;
      RECT 49.07 3.305 49.33 3.565 ;
      RECT 49.03 3.352 49.33 3.548 ;
      RECT 49.021 3.36 49.03 3.551 ;
      RECT 48.615 3.453 49.33 3.548 ;
      RECT 48.935 3.378 49.021 3.558 ;
      RECT 48.63 3.45 49.33 3.548 ;
      RECT 48.876 3.4 48.935 3.57 ;
      RECT 48.65 3.446 49.33 3.548 ;
      RECT 48.79 3.412 48.876 3.581 ;
      RECT 48.665 3.442 49.33 3.548 ;
      RECT 48.735 3.425 48.79 3.593 ;
      RECT 48.68 3.44 49.33 3.548 ;
      RECT 48.72 3.431 48.735 3.599 ;
      RECT 48.69 3.436 49.33 3.548 ;
      RECT 48.835 2.96 49.095 3.22 ;
      RECT 48.835 2.98 49.205 3.19 ;
      RECT 48.835 2.985 49.215 3.185 ;
      RECT 49.026 2.399 49.105 2.63 ;
      RECT 48.94 2.402 49.155 2.625 ;
      RECT 48.935 2.402 49.155 2.62 ;
      RECT 48.935 2.407 49.165 2.618 ;
      RECT 48.91 2.407 49.165 2.615 ;
      RECT 48.91 2.415 49.175 2.613 ;
      RECT 48.79 2.35 49.05 2.61 ;
      RECT 48.79 2.397 49.1 2.61 ;
      RECT 48.045 2.97 48.05 3.23 ;
      RECT 47.875 2.74 47.88 3.23 ;
      RECT 47.76 2.98 47.765 3.205 ;
      RECT 48.47 2.075 48.475 2.285 ;
      RECT 48.475 2.08 48.49 2.28 ;
      RECT 48.41 2.075 48.47 2.293 ;
      RECT 48.395 2.075 48.41 2.303 ;
      RECT 48.345 2.075 48.395 2.32 ;
      RECT 48.325 2.075 48.345 2.343 ;
      RECT 48.31 2.075 48.325 2.355 ;
      RECT 48.29 2.075 48.31 2.365 ;
      RECT 48.28 2.08 48.29 2.374 ;
      RECT 48.275 2.09 48.28 2.379 ;
      RECT 48.27 2.102 48.275 2.383 ;
      RECT 48.26 2.125 48.27 2.388 ;
      RECT 48.255 2.14 48.26 2.392 ;
      RECT 48.25 2.157 48.255 2.395 ;
      RECT 48.245 2.165 48.25 2.398 ;
      RECT 48.235 2.17 48.245 2.402 ;
      RECT 48.23 2.177 48.235 2.407 ;
      RECT 48.22 2.182 48.23 2.411 ;
      RECT 48.195 2.194 48.22 2.422 ;
      RECT 48.175 2.211 48.195 2.438 ;
      RECT 48.15 2.228 48.175 2.46 ;
      RECT 48.115 2.251 48.15 2.518 ;
      RECT 48.095 2.273 48.115 2.58 ;
      RECT 48.09 2.283 48.095 2.615 ;
      RECT 48.08 2.29 48.09 2.653 ;
      RECT 48.075 2.297 48.08 2.673 ;
      RECT 48.07 2.308 48.075 2.71 ;
      RECT 48.065 2.316 48.07 2.775 ;
      RECT 48.055 2.327 48.065 2.828 ;
      RECT 48.05 2.345 48.055 2.898 ;
      RECT 48.045 2.355 48.05 2.935 ;
      RECT 48.04 2.365 48.045 3.23 ;
      RECT 48.035 2.377 48.04 3.23 ;
      RECT 48.03 2.387 48.035 3.23 ;
      RECT 48.02 2.397 48.03 3.23 ;
      RECT 48.01 2.42 48.02 3.23 ;
      RECT 47.995 2.455 48.01 3.23 ;
      RECT 47.955 2.517 47.995 3.23 ;
      RECT 47.95 2.57 47.955 3.23 ;
      RECT 47.925 2.605 47.95 3.23 ;
      RECT 47.91 2.65 47.925 3.23 ;
      RECT 47.905 2.672 47.91 3.23 ;
      RECT 47.895 2.685 47.905 3.23 ;
      RECT 47.885 2.71 47.895 3.23 ;
      RECT 47.88 2.732 47.885 3.23 ;
      RECT 47.855 2.77 47.875 3.23 ;
      RECT 47.815 2.827 47.855 3.23 ;
      RECT 47.81 2.877 47.815 3.23 ;
      RECT 47.805 2.895 47.81 3.23 ;
      RECT 47.8 2.907 47.805 3.23 ;
      RECT 47.79 2.925 47.8 3.23 ;
      RECT 47.78 2.945 47.79 3.205 ;
      RECT 47.775 2.962 47.78 3.205 ;
      RECT 47.765 2.975 47.775 3.205 ;
      RECT 47.735 2.985 47.76 3.205 ;
      RECT 47.725 2.992 47.735 3.205 ;
      RECT 47.71 3.002 47.725 3.2 ;
      RECT 46.805 7.765 47.095 7.995 ;
      RECT 46.865 6.285 47.035 7.995 ;
      RECT 46.81 6.655 47.16 7.005 ;
      RECT 46.805 6.285 47.095 6.515 ;
      RECT 46.805 2.365 47.095 2.595 ;
      RECT 46.865 0.885 47.035 2.595 ;
      RECT 46.805 0.885 47.095 1.115 ;
      RECT 46.395 2.735 46.725 2.965 ;
      RECT 46.395 2.765 46.895 2.935 ;
      RECT 46.395 2.395 46.585 2.965 ;
      RECT 45.815 2.365 46.105 2.595 ;
      RECT 45.815 2.395 46.585 2.565 ;
      RECT 45.875 0.885 46.045 2.595 ;
      RECT 45.815 0.885 46.105 1.115 ;
      RECT 45.815 7.765 46.105 7.995 ;
      RECT 45.875 6.285 46.045 7.995 ;
      RECT 45.815 6.285 46.105 6.515 ;
      RECT 45.815 6.325 46.665 6.485 ;
      RECT 46.495 5.915 46.665 6.485 ;
      RECT 45.815 6.32 46.205 6.485 ;
      RECT 46.435 5.915 46.725 6.145 ;
      RECT 46.435 5.945 46.895 6.115 ;
      RECT 45.445 2.735 45.735 2.965 ;
      RECT 45.445 2.765 45.905 2.935 ;
      RECT 45.505 1.655 45.67 2.965 ;
      RECT 44.02 1.625 44.31 1.855 ;
      RECT 44.02 1.655 45.67 1.825 ;
      RECT 44.08 0.885 44.25 1.855 ;
      RECT 44.02 0.885 44.31 1.115 ;
      RECT 44.02 7.765 44.31 7.995 ;
      RECT 44.08 7.025 44.25 7.995 ;
      RECT 44.08 7.12 45.67 7.29 ;
      RECT 45.5 5.915 45.67 7.29 ;
      RECT 44.02 7.025 44.31 7.255 ;
      RECT 45.445 5.915 45.735 6.145 ;
      RECT 45.445 5.945 45.905 6.115 ;
      RECT 44.45 1.965 44.8 2.315 ;
      RECT 42.115 2.025 44.8 2.195 ;
      RECT 42.115 1.34 42.285 2.195 ;
      RECT 42.015 1.34 42.365 1.69 ;
      RECT 44.475 6.655 44.8 6.98 ;
      RECT 39.905 6.615 40.255 6.965 ;
      RECT 44.45 6.655 44.8 6.885 ;
      RECT 39.67 6.655 40.255 6.885 ;
      RECT 39.5 6.685 44.8 6.855 ;
      RECT 43.675 2.365 43.995 2.685 ;
      RECT 43.645 2.365 43.995 2.595 ;
      RECT 43.475 2.395 43.995 2.565 ;
      RECT 43.675 6.255 43.995 6.545 ;
      RECT 43.645 6.285 43.995 6.515 ;
      RECT 43.475 6.315 43.995 6.485 ;
      RECT 42.62 2.705 42.97 3.055 ;
      RECT 42.62 2.765 43.11 2.935 ;
      RECT 42.625 5.855 42.975 6.205 ;
      RECT 37.87 5.915 38.16 6.145 ;
      RECT 37.87 5.945 43.11 6.115 ;
      RECT 40.31 2.465 40.495 2.675 ;
      RECT 40.3 2.47 40.51 2.668 ;
      RECT 40.3 2.47 40.596 2.645 ;
      RECT 40.3 2.47 40.655 2.62 ;
      RECT 40.3 2.47 40.71 2.6 ;
      RECT 40.3 2.47 40.72 2.588 ;
      RECT 40.3 2.47 40.915 2.527 ;
      RECT 40.3 2.47 40.945 2.51 ;
      RECT 40.3 2.47 40.965 2.5 ;
      RECT 40.845 2.235 41.105 2.495 ;
      RECT 40.83 2.325 40.845 2.542 ;
      RECT 40.365 2.457 41.105 2.495 ;
      RECT 40.816 2.336 40.83 2.548 ;
      RECT 40.405 2.45 41.105 2.495 ;
      RECT 40.73 2.376 40.816 2.567 ;
      RECT 40.655 2.437 41.105 2.495 ;
      RECT 40.725 2.412 40.73 2.584 ;
      RECT 40.71 2.422 41.105 2.495 ;
      RECT 40.72 2.417 40.725 2.586 ;
      RECT 41.015 2.922 41.02 3.014 ;
      RECT 41.01 2.9 41.015 3.031 ;
      RECT 41.005 2.89 41.01 3.043 ;
      RECT 40.995 2.881 41.005 3.053 ;
      RECT 40.99 2.876 40.995 3.061 ;
      RECT 40.985 2.735 40.99 3.064 ;
      RECT 40.951 2.735 40.985 3.075 ;
      RECT 40.865 2.735 40.951 3.11 ;
      RECT 40.785 2.735 40.865 3.158 ;
      RECT 40.756 2.735 40.785 3.182 ;
      RECT 40.67 2.735 40.756 3.188 ;
      RECT 40.665 2.919 40.67 3.193 ;
      RECT 40.63 2.93 40.665 3.196 ;
      RECT 40.605 2.945 40.63 3.2 ;
      RECT 40.591 2.954 40.605 3.202 ;
      RECT 40.505 2.981 40.591 3.208 ;
      RECT 40.44 3.022 40.505 3.217 ;
      RECT 40.425 3.042 40.44 3.222 ;
      RECT 40.395 3.052 40.425 3.225 ;
      RECT 40.39 3.062 40.395 3.228 ;
      RECT 40.36 3.067 40.39 3.23 ;
      RECT 40.34 3.072 40.36 3.234 ;
      RECT 40.255 3.075 40.34 3.241 ;
      RECT 40.24 3.072 40.255 3.247 ;
      RECT 40.23 3.069 40.24 3.249 ;
      RECT 40.21 3.066 40.23 3.251 ;
      RECT 40.19 3.062 40.21 3.252 ;
      RECT 40.175 3.058 40.19 3.254 ;
      RECT 40.165 3.055 40.175 3.255 ;
      RECT 40.125 3.049 40.165 3.253 ;
      RECT 40.115 3.044 40.125 3.251 ;
      RECT 40.1 3.041 40.115 3.247 ;
      RECT 40.075 3.036 40.1 3.24 ;
      RECT 40.025 3.027 40.075 3.228 ;
      RECT 39.955 3.013 40.025 3.21 ;
      RECT 39.897 2.998 39.955 3.192 ;
      RECT 39.811 2.981 39.897 3.172 ;
      RECT 39.725 2.96 39.811 3.147 ;
      RECT 39.675 2.945 39.725 3.128 ;
      RECT 39.671 2.939 39.675 3.12 ;
      RECT 39.585 2.929 39.671 3.107 ;
      RECT 39.55 2.914 39.585 3.09 ;
      RECT 39.535 2.907 39.55 3.083 ;
      RECT 39.475 2.895 39.535 3.071 ;
      RECT 39.455 2.882 39.475 3.059 ;
      RECT 39.415 2.873 39.455 3.051 ;
      RECT 39.41 2.865 39.415 3.044 ;
      RECT 39.33 2.855 39.41 3.03 ;
      RECT 39.315 2.842 39.33 3.015 ;
      RECT 39.31 2.84 39.315 3.013 ;
      RECT 39.231 2.828 39.31 3 ;
      RECT 39.145 2.803 39.231 2.975 ;
      RECT 39.13 2.772 39.145 2.96 ;
      RECT 39.115 2.747 39.13 2.956 ;
      RECT 39.1 2.74 39.115 2.952 ;
      RECT 38.925 2.745 38.93 2.948 ;
      RECT 38.92 2.75 38.925 2.943 ;
      RECT 38.93 2.74 39.1 2.95 ;
      RECT 39.645 2.5 39.75 2.76 ;
      RECT 40.46 2.025 40.465 2.25 ;
      RECT 40.59 2.025 40.645 2.235 ;
      RECT 40.645 2.03 40.655 2.228 ;
      RECT 40.551 2.025 40.59 2.238 ;
      RECT 40.465 2.025 40.551 2.245 ;
      RECT 40.445 2.03 40.46 2.251 ;
      RECT 40.435 2.07 40.445 2.253 ;
      RECT 40.405 2.08 40.435 2.255 ;
      RECT 40.4 2.085 40.405 2.257 ;
      RECT 40.375 2.09 40.4 2.259 ;
      RECT 40.36 2.095 40.375 2.261 ;
      RECT 40.345 2.097 40.36 2.263 ;
      RECT 40.34 2.102 40.345 2.265 ;
      RECT 40.29 2.11 40.34 2.268 ;
      RECT 40.265 2.119 40.29 2.273 ;
      RECT 40.255 2.126 40.265 2.278 ;
      RECT 40.25 2.129 40.255 2.282 ;
      RECT 40.23 2.132 40.25 2.291 ;
      RECT 40.2 2.14 40.23 2.311 ;
      RECT 40.171 2.153 40.2 2.333 ;
      RECT 40.085 2.187 40.171 2.377 ;
      RECT 40.08 2.213 40.085 2.415 ;
      RECT 40.075 2.217 40.08 2.424 ;
      RECT 40.04 2.23 40.075 2.457 ;
      RECT 40.03 2.244 40.04 2.495 ;
      RECT 40.025 2.248 40.03 2.508 ;
      RECT 40.02 2.252 40.025 2.513 ;
      RECT 40.01 2.26 40.02 2.525 ;
      RECT 40.005 2.267 40.01 2.54 ;
      RECT 39.98 2.28 40.005 2.565 ;
      RECT 39.94 2.309 39.98 2.62 ;
      RECT 39.925 2.334 39.94 2.675 ;
      RECT 39.915 2.345 39.925 2.698 ;
      RECT 39.91 2.352 39.915 2.71 ;
      RECT 39.905 2.356 39.91 2.718 ;
      RECT 39.85 2.384 39.905 2.76 ;
      RECT 39.83 2.42 39.85 2.76 ;
      RECT 39.815 2.435 39.83 2.76 ;
      RECT 39.76 2.467 39.815 2.76 ;
      RECT 39.75 2.497 39.76 2.76 ;
      RECT 39.36 2.112 39.545 2.35 ;
      RECT 39.345 2.114 39.555 2.345 ;
      RECT 39.23 2.06 39.49 2.32 ;
      RECT 39.225 2.097 39.49 2.274 ;
      RECT 39.22 2.107 39.49 2.271 ;
      RECT 39.215 2.147 39.555 2.265 ;
      RECT 39.21 2.18 39.555 2.255 ;
      RECT 39.22 2.122 39.57 2.193 ;
      RECT 39.517 3.22 39.53 3.75 ;
      RECT 39.431 3.22 39.53 3.749 ;
      RECT 39.431 3.22 39.535 3.748 ;
      RECT 39.345 3.22 39.535 3.746 ;
      RECT 39.34 3.22 39.535 3.743 ;
      RECT 39.34 3.22 39.545 3.741 ;
      RECT 39.335 3.512 39.545 3.738 ;
      RECT 39.335 3.522 39.55 3.735 ;
      RECT 39.335 3.59 39.555 3.731 ;
      RECT 39.325 3.595 39.555 3.73 ;
      RECT 39.325 3.687 39.56 3.727 ;
      RECT 39.31 3.22 39.57 3.48 ;
      RECT 39.24 7.765 39.53 7.995 ;
      RECT 39.3 7.025 39.47 7.995 ;
      RECT 39.215 7.055 39.555 7.4 ;
      RECT 39.24 7.025 39.53 7.4 ;
      RECT 38.54 2.21 38.585 3.745 ;
      RECT 38.74 2.21 38.77 2.425 ;
      RECT 37.115 1.95 37.235 2.16 ;
      RECT 36.775 1.9 37.035 2.16 ;
      RECT 36.775 1.945 37.07 2.15 ;
      RECT 38.78 2.226 38.785 2.28 ;
      RECT 38.775 2.219 38.78 2.413 ;
      RECT 38.77 2.213 38.775 2.42 ;
      RECT 38.725 2.21 38.74 2.433 ;
      RECT 38.72 2.21 38.725 2.455 ;
      RECT 38.715 2.21 38.72 2.503 ;
      RECT 38.71 2.21 38.715 2.523 ;
      RECT 38.7 2.21 38.71 2.63 ;
      RECT 38.695 2.21 38.7 2.693 ;
      RECT 38.69 2.21 38.695 2.75 ;
      RECT 38.685 2.21 38.69 2.758 ;
      RECT 38.67 2.21 38.685 2.865 ;
      RECT 38.66 2.21 38.67 3 ;
      RECT 38.65 2.21 38.66 3.11 ;
      RECT 38.64 2.21 38.65 3.167 ;
      RECT 38.635 2.21 38.64 3.207 ;
      RECT 38.63 2.21 38.635 3.243 ;
      RECT 38.62 2.21 38.63 3.283 ;
      RECT 38.615 2.21 38.62 3.325 ;
      RECT 38.595 2.21 38.615 3.39 ;
      RECT 38.6 3.535 38.605 3.715 ;
      RECT 38.595 3.517 38.6 3.723 ;
      RECT 38.59 2.21 38.595 3.453 ;
      RECT 38.59 3.497 38.595 3.73 ;
      RECT 38.585 2.21 38.59 3.74 ;
      RECT 38.53 2.21 38.54 2.51 ;
      RECT 38.535 2.757 38.54 3.745 ;
      RECT 38.53 2.822 38.535 3.745 ;
      RECT 38.525 2.211 38.53 2.5 ;
      RECT 38.52 2.887 38.53 3.745 ;
      RECT 38.515 2.212 38.525 2.49 ;
      RECT 38.505 3 38.52 3.745 ;
      RECT 38.51 2.213 38.515 2.48 ;
      RECT 38.49 2.214 38.51 2.458 ;
      RECT 38.495 3.097 38.505 3.745 ;
      RECT 38.49 3.172 38.495 3.745 ;
      RECT 38.48 2.213 38.49 2.435 ;
      RECT 38.485 3.215 38.49 3.745 ;
      RECT 38.48 3.242 38.485 3.745 ;
      RECT 38.47 2.211 38.48 2.423 ;
      RECT 38.475 3.285 38.48 3.745 ;
      RECT 38.47 3.312 38.475 3.745 ;
      RECT 38.46 2.21 38.47 2.41 ;
      RECT 38.465 3.327 38.47 3.745 ;
      RECT 38.425 3.385 38.465 3.745 ;
      RECT 38.455 2.209 38.46 2.395 ;
      RECT 38.45 2.207 38.455 2.388 ;
      RECT 38.44 2.204 38.45 2.378 ;
      RECT 38.435 2.201 38.44 2.363 ;
      RECT 38.42 2.197 38.435 2.356 ;
      RECT 38.415 3.44 38.425 3.745 ;
      RECT 38.415 2.194 38.42 2.351 ;
      RECT 38.4 2.19 38.415 2.345 ;
      RECT 38.41 3.457 38.415 3.745 ;
      RECT 38.4 3.52 38.41 3.745 ;
      RECT 38.32 2.175 38.4 2.325 ;
      RECT 38.395 3.527 38.4 3.74 ;
      RECT 38.39 3.535 38.395 3.73 ;
      RECT 38.31 2.161 38.32 2.309 ;
      RECT 38.295 2.157 38.31 2.307 ;
      RECT 38.285 2.152 38.295 2.303 ;
      RECT 38.26 2.145 38.285 2.295 ;
      RECT 38.255 2.14 38.26 2.29 ;
      RECT 38.245 2.14 38.255 2.288 ;
      RECT 38.235 2.138 38.245 2.286 ;
      RECT 38.205 2.13 38.235 2.28 ;
      RECT 38.19 2.122 38.205 2.273 ;
      RECT 38.17 2.117 38.19 2.266 ;
      RECT 38.165 2.113 38.17 2.261 ;
      RECT 38.135 2.106 38.165 2.255 ;
      RECT 38.11 2.097 38.135 2.245 ;
      RECT 38.08 2.09 38.11 2.237 ;
      RECT 38.055 2.08 38.08 2.228 ;
      RECT 38.04 2.072 38.055 2.222 ;
      RECT 38.015 2.067 38.04 2.217 ;
      RECT 38.005 2.063 38.015 2.212 ;
      RECT 37.985 2.058 38.005 2.207 ;
      RECT 37.95 2.053 37.985 2.2 ;
      RECT 37.89 2.048 37.95 2.193 ;
      RECT 37.877 2.044 37.89 2.191 ;
      RECT 37.791 2.039 37.877 2.188 ;
      RECT 37.705 2.029 37.791 2.184 ;
      RECT 37.664 2.022 37.705 2.181 ;
      RECT 37.578 2.015 37.664 2.178 ;
      RECT 37.492 2.005 37.578 2.174 ;
      RECT 37.406 1.995 37.492 2.169 ;
      RECT 37.32 1.985 37.406 2.165 ;
      RECT 37.31 1.97 37.32 2.163 ;
      RECT 37.3 1.955 37.31 2.163 ;
      RECT 37.235 1.95 37.3 2.162 ;
      RECT 37.07 1.947 37.115 2.155 ;
      RECT 38.315 2.852 38.32 3.043 ;
      RECT 38.31 2.847 38.315 3.05 ;
      RECT 38.296 2.845 38.31 3.056 ;
      RECT 38.21 2.845 38.296 3.058 ;
      RECT 38.206 2.845 38.21 3.061 ;
      RECT 38.12 2.845 38.206 3.079 ;
      RECT 38.11 2.85 38.12 3.098 ;
      RECT 38.1 2.905 38.11 3.102 ;
      RECT 38.075 2.92 38.1 3.109 ;
      RECT 38.035 2.94 38.075 3.122 ;
      RECT 38.03 2.952 38.035 3.132 ;
      RECT 38.015 2.958 38.03 3.137 ;
      RECT 38.01 2.963 38.015 3.141 ;
      RECT 37.99 2.97 38.01 3.146 ;
      RECT 37.92 2.995 37.99 3.163 ;
      RECT 37.88 3.023 37.92 3.183 ;
      RECT 37.875 3.033 37.88 3.191 ;
      RECT 37.855 3.04 37.875 3.193 ;
      RECT 37.85 3.047 37.855 3.196 ;
      RECT 37.82 3.055 37.85 3.199 ;
      RECT 37.815 3.06 37.82 3.203 ;
      RECT 37.741 3.064 37.815 3.211 ;
      RECT 37.655 3.073 37.741 3.227 ;
      RECT 37.651 3.078 37.655 3.236 ;
      RECT 37.565 3.083 37.651 3.246 ;
      RECT 37.525 3.091 37.565 3.258 ;
      RECT 37.475 3.097 37.525 3.265 ;
      RECT 37.39 3.106 37.475 3.28 ;
      RECT 37.315 3.117 37.39 3.298 ;
      RECT 37.28 3.124 37.315 3.308 ;
      RECT 37.205 3.132 37.28 3.313 ;
      RECT 37.15 3.141 37.205 3.313 ;
      RECT 37.125 3.146 37.15 3.311 ;
      RECT 37.115 3.149 37.125 3.309 ;
      RECT 37.08 3.151 37.115 3.307 ;
      RECT 37.05 3.153 37.08 3.303 ;
      RECT 37.005 3.152 37.05 3.299 ;
      RECT 36.985 3.147 37.005 3.296 ;
      RECT 36.935 3.132 36.985 3.293 ;
      RECT 36.925 3.117 36.935 3.288 ;
      RECT 36.875 3.102 36.925 3.278 ;
      RECT 36.825 3.077 36.875 3.258 ;
      RECT 36.815 3.062 36.825 3.24 ;
      RECT 36.81 3.06 36.815 3.234 ;
      RECT 36.79 3.055 36.81 3.229 ;
      RECT 36.785 3.047 36.79 3.223 ;
      RECT 36.77 3.041 36.785 3.216 ;
      RECT 36.765 3.036 36.77 3.208 ;
      RECT 36.745 3.031 36.765 3.2 ;
      RECT 36.73 3.024 36.745 3.193 ;
      RECT 36.715 3.018 36.73 3.184 ;
      RECT 36.71 3.012 36.715 3.177 ;
      RECT 36.665 2.987 36.71 3.163 ;
      RECT 36.65 2.957 36.665 3.145 ;
      RECT 36.635 2.94 36.65 3.136 ;
      RECT 36.61 2.92 36.635 3.124 ;
      RECT 36.57 2.89 36.61 3.104 ;
      RECT 36.56 2.86 36.57 3.089 ;
      RECT 36.545 2.85 36.56 3.082 ;
      RECT 36.49 2.815 36.545 3.061 ;
      RECT 36.475 2.778 36.49 3.04 ;
      RECT 36.465 2.765 36.475 3.032 ;
      RECT 36.415 2.735 36.465 3.014 ;
      RECT 36.4 2.665 36.415 2.995 ;
      RECT 36.355 2.665 36.4 2.978 ;
      RECT 36.33 2.665 36.355 2.96 ;
      RECT 36.32 2.665 36.33 2.953 ;
      RECT 36.241 2.665 36.32 2.946 ;
      RECT 36.155 2.665 36.241 2.938 ;
      RECT 36.14 2.697 36.155 2.933 ;
      RECT 36.065 2.707 36.14 2.929 ;
      RECT 36.045 2.717 36.065 2.924 ;
      RECT 36.02 2.717 36.045 2.921 ;
      RECT 36.01 2.707 36.02 2.92 ;
      RECT 36 2.68 36.01 2.919 ;
      RECT 35.96 2.675 36 2.917 ;
      RECT 35.915 2.675 35.96 2.913 ;
      RECT 35.89 2.675 35.915 2.908 ;
      RECT 35.84 2.675 35.89 2.895 ;
      RECT 35.8 2.68 35.81 2.88 ;
      RECT 35.81 2.675 35.84 2.885 ;
      RECT 37.795 2.455 38.055 2.715 ;
      RECT 37.79 2.477 38.055 2.673 ;
      RECT 37.03 2.305 37.25 2.67 ;
      RECT 37.012 2.392 37.25 2.669 ;
      RECT 36.995 2.397 37.25 2.666 ;
      RECT 36.995 2.397 37.27 2.665 ;
      RECT 36.965 2.407 37.27 2.663 ;
      RECT 36.96 2.422 37.27 2.659 ;
      RECT 36.96 2.422 37.275 2.658 ;
      RECT 36.955 2.48 37.275 2.656 ;
      RECT 36.955 2.48 37.285 2.653 ;
      RECT 36.95 2.545 37.285 2.648 ;
      RECT 37.03 2.305 37.29 2.565 ;
      RECT 35.775 2.135 36.035 2.395 ;
      RECT 35.775 2.178 36.121 2.369 ;
      RECT 35.775 2.178 36.165 2.368 ;
      RECT 35.775 2.178 36.185 2.366 ;
      RECT 35.775 2.178 36.285 2.365 ;
      RECT 35.775 2.178 36.305 2.363 ;
      RECT 35.775 2.178 36.315 2.358 ;
      RECT 36.185 2.145 36.375 2.355 ;
      RECT 36.185 2.147 36.38 2.353 ;
      RECT 36.175 2.152 36.385 2.345 ;
      RECT 36.121 2.176 36.385 2.345 ;
      RECT 36.165 2.17 36.175 2.367 ;
      RECT 36.175 2.15 36.38 2.353 ;
      RECT 35.13 3.21 35.335 3.44 ;
      RECT 35.07 3.16 35.125 3.42 ;
      RECT 35.13 3.16 35.33 3.44 ;
      RECT 36.1 3.475 36.105 3.502 ;
      RECT 36.09 3.385 36.1 3.507 ;
      RECT 36.085 3.307 36.09 3.513 ;
      RECT 36.075 3.297 36.085 3.52 ;
      RECT 36.07 3.287 36.075 3.526 ;
      RECT 36.06 3.282 36.07 3.528 ;
      RECT 36.045 3.274 36.06 3.536 ;
      RECT 36.03 3.265 36.045 3.548 ;
      RECT 36.02 3.257 36.03 3.558 ;
      RECT 35.985 3.175 36.02 3.576 ;
      RECT 35.95 3.175 35.985 3.595 ;
      RECT 35.935 3.175 35.95 3.603 ;
      RECT 35.88 3.175 35.935 3.603 ;
      RECT 35.846 3.175 35.88 3.594 ;
      RECT 35.76 3.175 35.846 3.57 ;
      RECT 35.75 3.235 35.76 3.552 ;
      RECT 35.71 3.237 35.75 3.543 ;
      RECT 35.705 3.239 35.71 3.533 ;
      RECT 35.685 3.241 35.705 3.528 ;
      RECT 35.675 3.244 35.685 3.523 ;
      RECT 35.665 3.245 35.675 3.518 ;
      RECT 35.641 3.246 35.665 3.51 ;
      RECT 35.555 3.251 35.641 3.488 ;
      RECT 35.5 3.25 35.555 3.461 ;
      RECT 35.485 3.243 35.5 3.448 ;
      RECT 35.45 3.238 35.485 3.444 ;
      RECT 35.395 3.23 35.45 3.443 ;
      RECT 35.335 3.217 35.395 3.441 ;
      RECT 35.125 3.16 35.13 3.428 ;
      RECT 35.2 2.53 35.385 2.74 ;
      RECT 35.19 2.535 35.4 2.733 ;
      RECT 35.23 2.44 35.49 2.7 ;
      RECT 35.185 2.597 35.49 2.623 ;
      RECT 34.53 2.39 34.535 3.19 ;
      RECT 34.475 2.44 34.505 3.19 ;
      RECT 34.465 2.44 34.47 2.75 ;
      RECT 34.45 2.44 34.455 2.745 ;
      RECT 33.995 2.485 34.01 2.7 ;
      RECT 33.925 2.485 34.01 2.695 ;
      RECT 35.19 2.065 35.26 2.275 ;
      RECT 35.26 2.072 35.27 2.27 ;
      RECT 35.156 2.065 35.19 2.282 ;
      RECT 35.07 2.065 35.156 2.306 ;
      RECT 35.06 2.07 35.07 2.325 ;
      RECT 35.055 2.082 35.06 2.328 ;
      RECT 35.04 2.097 35.055 2.332 ;
      RECT 35.035 2.115 35.04 2.336 ;
      RECT 34.995 2.125 35.035 2.345 ;
      RECT 34.98 2.132 34.995 2.357 ;
      RECT 34.965 2.137 34.98 2.362 ;
      RECT 34.95 2.14 34.965 2.367 ;
      RECT 34.94 2.142 34.95 2.371 ;
      RECT 34.905 2.149 34.94 2.379 ;
      RECT 34.87 2.157 34.905 2.393 ;
      RECT 34.86 2.163 34.87 2.402 ;
      RECT 34.855 2.165 34.86 2.404 ;
      RECT 34.835 2.168 34.855 2.41 ;
      RECT 34.805 2.175 34.835 2.421 ;
      RECT 34.795 2.181 34.805 2.428 ;
      RECT 34.77 2.184 34.795 2.435 ;
      RECT 34.76 2.188 34.77 2.443 ;
      RECT 34.755 2.189 34.76 2.465 ;
      RECT 34.75 2.19 34.755 2.48 ;
      RECT 34.745 2.191 34.75 2.495 ;
      RECT 34.74 2.192 34.745 2.51 ;
      RECT 34.735 2.193 34.74 2.54 ;
      RECT 34.725 2.195 34.735 2.573 ;
      RECT 34.71 2.199 34.725 2.62 ;
      RECT 34.7 2.202 34.71 2.665 ;
      RECT 34.695 2.205 34.7 2.693 ;
      RECT 34.685 2.207 34.695 2.72 ;
      RECT 34.68 2.21 34.685 2.755 ;
      RECT 34.65 2.215 34.68 2.813 ;
      RECT 34.645 2.22 34.65 2.898 ;
      RECT 34.64 2.222 34.645 2.933 ;
      RECT 34.635 2.224 34.64 3.015 ;
      RECT 34.63 2.226 34.635 3.103 ;
      RECT 34.62 2.228 34.63 3.185 ;
      RECT 34.605 2.242 34.62 3.19 ;
      RECT 34.57 2.287 34.605 3.19 ;
      RECT 34.56 2.327 34.57 3.19 ;
      RECT 34.545 2.355 34.56 3.19 ;
      RECT 34.54 2.372 34.545 3.19 ;
      RECT 34.535 2.38 34.54 3.19 ;
      RECT 34.525 2.395 34.53 3.19 ;
      RECT 34.52 2.402 34.525 3.19 ;
      RECT 34.51 2.422 34.52 3.19 ;
      RECT 34.505 2.435 34.51 3.19 ;
      RECT 34.47 2.44 34.475 2.775 ;
      RECT 34.455 2.83 34.475 3.19 ;
      RECT 34.455 2.44 34.465 2.748 ;
      RECT 34.45 2.87 34.455 3.19 ;
      RECT 34.4 2.44 34.45 2.743 ;
      RECT 34.445 2.907 34.45 3.19 ;
      RECT 34.435 2.93 34.445 3.19 ;
      RECT 34.43 2.975 34.435 3.19 ;
      RECT 34.42 2.985 34.43 3.183 ;
      RECT 34.346 2.44 34.4 2.737 ;
      RECT 34.26 2.44 34.346 2.73 ;
      RECT 34.211 2.487 34.26 2.723 ;
      RECT 34.125 2.495 34.211 2.716 ;
      RECT 34.11 2.492 34.125 2.711 ;
      RECT 34.096 2.485 34.11 2.71 ;
      RECT 34.01 2.485 34.096 2.705 ;
      RECT 33.915 2.49 33.925 2.69 ;
      RECT 33.505 1.92 33.52 2.32 ;
      RECT 33.7 1.92 33.705 2.18 ;
      RECT 33.445 1.92 33.49 2.18 ;
      RECT 33.9 3.225 33.905 3.43 ;
      RECT 33.895 3.215 33.9 3.435 ;
      RECT 33.89 3.202 33.895 3.44 ;
      RECT 33.885 3.182 33.89 3.44 ;
      RECT 33.86 3.135 33.885 3.44 ;
      RECT 33.825 3.05 33.86 3.44 ;
      RECT 33.82 2.987 33.825 3.44 ;
      RECT 33.815 2.972 33.82 3.44 ;
      RECT 33.8 2.932 33.815 3.44 ;
      RECT 33.795 2.907 33.8 3.44 ;
      RECT 33.785 2.89 33.795 3.44 ;
      RECT 33.75 2.812 33.785 3.44 ;
      RECT 33.745 2.755 33.75 3.44 ;
      RECT 33.74 2.742 33.745 3.44 ;
      RECT 33.73 2.72 33.74 3.44 ;
      RECT 33.72 2.685 33.73 3.44 ;
      RECT 33.71 2.655 33.72 3.44 ;
      RECT 33.7 2.57 33.71 3.083 ;
      RECT 33.707 3.215 33.71 3.44 ;
      RECT 33.705 3.225 33.707 3.44 ;
      RECT 33.695 3.235 33.705 3.435 ;
      RECT 33.69 1.92 33.7 2.315 ;
      RECT 33.695 2.447 33.7 3.058 ;
      RECT 33.69 2.345 33.695 3.041 ;
      RECT 33.68 1.92 33.69 3.017 ;
      RECT 33.675 1.92 33.68 2.988 ;
      RECT 33.67 1.92 33.675 2.978 ;
      RECT 33.65 1.92 33.67 2.94 ;
      RECT 33.645 1.92 33.65 2.898 ;
      RECT 33.64 1.92 33.645 2.878 ;
      RECT 33.61 1.92 33.64 2.828 ;
      RECT 33.6 1.92 33.61 2.775 ;
      RECT 33.595 1.92 33.6 2.748 ;
      RECT 33.59 1.92 33.595 2.733 ;
      RECT 33.58 1.92 33.59 2.71 ;
      RECT 33.57 1.92 33.58 2.685 ;
      RECT 33.565 1.92 33.57 2.625 ;
      RECT 33.555 1.92 33.565 2.563 ;
      RECT 33.55 1.92 33.555 2.483 ;
      RECT 33.545 1.92 33.55 2.448 ;
      RECT 33.54 1.92 33.545 2.423 ;
      RECT 33.535 1.92 33.54 2.408 ;
      RECT 33.53 1.92 33.535 2.378 ;
      RECT 33.525 1.92 33.53 2.355 ;
      RECT 33.52 1.92 33.525 2.328 ;
      RECT 33.49 1.92 33.505 2.315 ;
      RECT 32.645 3.455 32.83 3.665 ;
      RECT 32.635 3.46 32.845 3.658 ;
      RECT 32.635 3.46 32.865 3.63 ;
      RECT 32.635 3.46 32.88 3.609 ;
      RECT 32.635 3.46 32.895 3.607 ;
      RECT 32.635 3.46 32.905 3.606 ;
      RECT 32.635 3.46 32.935 3.603 ;
      RECT 33.285 3.305 33.545 3.565 ;
      RECT 33.245 3.352 33.545 3.548 ;
      RECT 33.236 3.36 33.245 3.551 ;
      RECT 32.83 3.453 33.545 3.548 ;
      RECT 33.15 3.378 33.236 3.558 ;
      RECT 32.845 3.45 33.545 3.548 ;
      RECT 33.091 3.4 33.15 3.57 ;
      RECT 32.865 3.446 33.545 3.548 ;
      RECT 33.005 3.412 33.091 3.581 ;
      RECT 32.88 3.442 33.545 3.548 ;
      RECT 32.95 3.425 33.005 3.593 ;
      RECT 32.895 3.44 33.545 3.548 ;
      RECT 32.935 3.431 32.95 3.599 ;
      RECT 32.905 3.436 33.545 3.548 ;
      RECT 33.05 2.96 33.31 3.22 ;
      RECT 33.05 2.98 33.42 3.19 ;
      RECT 33.05 2.985 33.43 3.185 ;
      RECT 33.241 2.399 33.32 2.63 ;
      RECT 33.155 2.402 33.37 2.625 ;
      RECT 33.15 2.402 33.37 2.62 ;
      RECT 33.15 2.407 33.38 2.618 ;
      RECT 33.125 2.407 33.38 2.615 ;
      RECT 33.125 2.415 33.39 2.613 ;
      RECT 33.005 2.35 33.265 2.61 ;
      RECT 33.005 2.397 33.315 2.61 ;
      RECT 32.26 2.97 32.265 3.23 ;
      RECT 32.09 2.74 32.095 3.23 ;
      RECT 31.975 2.98 31.98 3.205 ;
      RECT 32.685 2.075 32.69 2.285 ;
      RECT 32.69 2.08 32.705 2.28 ;
      RECT 32.625 2.075 32.685 2.293 ;
      RECT 32.61 2.075 32.625 2.303 ;
      RECT 32.56 2.075 32.61 2.32 ;
      RECT 32.54 2.075 32.56 2.343 ;
      RECT 32.525 2.075 32.54 2.355 ;
      RECT 32.505 2.075 32.525 2.365 ;
      RECT 32.495 2.08 32.505 2.374 ;
      RECT 32.49 2.09 32.495 2.379 ;
      RECT 32.485 2.102 32.49 2.383 ;
      RECT 32.475 2.125 32.485 2.388 ;
      RECT 32.47 2.14 32.475 2.392 ;
      RECT 32.465 2.157 32.47 2.395 ;
      RECT 32.46 2.165 32.465 2.398 ;
      RECT 32.45 2.17 32.46 2.402 ;
      RECT 32.445 2.177 32.45 2.407 ;
      RECT 32.435 2.182 32.445 2.411 ;
      RECT 32.41 2.194 32.435 2.422 ;
      RECT 32.39 2.211 32.41 2.438 ;
      RECT 32.365 2.228 32.39 2.46 ;
      RECT 32.33 2.251 32.365 2.518 ;
      RECT 32.31 2.273 32.33 2.58 ;
      RECT 32.305 2.283 32.31 2.615 ;
      RECT 32.295 2.29 32.305 2.653 ;
      RECT 32.29 2.297 32.295 2.673 ;
      RECT 32.285 2.308 32.29 2.71 ;
      RECT 32.28 2.316 32.285 2.775 ;
      RECT 32.27 2.327 32.28 2.828 ;
      RECT 32.265 2.345 32.27 2.898 ;
      RECT 32.26 2.355 32.265 2.935 ;
      RECT 32.255 2.365 32.26 3.23 ;
      RECT 32.25 2.377 32.255 3.23 ;
      RECT 32.245 2.387 32.25 3.23 ;
      RECT 32.235 2.397 32.245 3.23 ;
      RECT 32.225 2.42 32.235 3.23 ;
      RECT 32.21 2.455 32.225 3.23 ;
      RECT 32.17 2.517 32.21 3.23 ;
      RECT 32.165 2.57 32.17 3.23 ;
      RECT 32.14 2.605 32.165 3.23 ;
      RECT 32.125 2.65 32.14 3.23 ;
      RECT 32.12 2.672 32.125 3.23 ;
      RECT 32.11 2.685 32.12 3.23 ;
      RECT 32.1 2.71 32.11 3.23 ;
      RECT 32.095 2.732 32.1 3.23 ;
      RECT 32.07 2.77 32.09 3.23 ;
      RECT 32.03 2.827 32.07 3.23 ;
      RECT 32.025 2.877 32.03 3.23 ;
      RECT 32.02 2.895 32.025 3.23 ;
      RECT 32.015 2.907 32.02 3.23 ;
      RECT 32.005 2.925 32.015 3.23 ;
      RECT 31.995 2.945 32.005 3.205 ;
      RECT 31.99 2.962 31.995 3.205 ;
      RECT 31.98 2.975 31.99 3.205 ;
      RECT 31.95 2.985 31.975 3.205 ;
      RECT 31.94 2.992 31.95 3.205 ;
      RECT 31.925 3.002 31.94 3.2 ;
      RECT 31.03 7.765 31.32 7.995 ;
      RECT 31.09 6.285 31.26 7.995 ;
      RECT 31.075 6.66 31.43 7.015 ;
      RECT 31.03 6.285 31.32 6.515 ;
      RECT 31.03 2.365 31.32 2.595 ;
      RECT 31.09 0.885 31.26 2.595 ;
      RECT 31.03 0.885 31.32 1.115 ;
      RECT 30.62 2.735 30.95 2.965 ;
      RECT 30.62 2.765 31.12 2.935 ;
      RECT 30.62 2.395 30.81 2.965 ;
      RECT 30.04 2.365 30.33 2.595 ;
      RECT 30.04 2.395 30.81 2.565 ;
      RECT 30.1 0.885 30.27 2.595 ;
      RECT 30.04 0.885 30.33 1.115 ;
      RECT 30.04 7.765 30.33 7.995 ;
      RECT 30.1 6.285 30.27 7.995 ;
      RECT 30.04 6.285 30.33 6.515 ;
      RECT 30.04 6.325 30.89 6.485 ;
      RECT 30.72 5.915 30.89 6.485 ;
      RECT 30.04 6.32 30.43 6.485 ;
      RECT 30.66 5.915 30.95 6.145 ;
      RECT 30.66 5.945 31.12 6.115 ;
      RECT 29.67 2.735 29.96 2.965 ;
      RECT 29.67 2.765 30.13 2.935 ;
      RECT 29.73 1.655 29.895 2.965 ;
      RECT 28.245 1.625 28.535 1.855 ;
      RECT 28.245 1.655 29.895 1.825 ;
      RECT 28.305 0.885 28.475 1.855 ;
      RECT 28.245 0.885 28.535 1.115 ;
      RECT 28.245 7.765 28.535 7.995 ;
      RECT 28.305 7.025 28.475 7.995 ;
      RECT 28.305 7.12 29.895 7.29 ;
      RECT 29.725 5.915 29.895 7.29 ;
      RECT 28.245 7.025 28.535 7.255 ;
      RECT 29.67 5.915 29.96 6.145 ;
      RECT 29.67 5.945 30.13 6.115 ;
      RECT 28.675 1.965 29.025 2.315 ;
      RECT 26.34 2.025 29.025 2.195 ;
      RECT 26.34 1.34 26.51 2.195 ;
      RECT 26.24 1.34 26.59 1.69 ;
      RECT 28.7 6.655 29.025 6.98 ;
      RECT 24.125 6.61 24.475 6.96 ;
      RECT 28.675 6.655 29.025 6.885 ;
      RECT 23.895 6.655 24.475 6.885 ;
      RECT 23.725 6.685 29.025 6.855 ;
      RECT 27.9 2.365 28.22 2.685 ;
      RECT 27.87 2.365 28.22 2.595 ;
      RECT 27.7 2.395 28.22 2.565 ;
      RECT 27.9 6.255 28.22 6.545 ;
      RECT 27.87 6.285 28.22 6.515 ;
      RECT 27.7 6.315 28.22 6.485 ;
      RECT 26.845 2.705 27.195 3.055 ;
      RECT 26.845 2.765 27.335 2.935 ;
      RECT 26.85 5.855 27.2 6.205 ;
      RECT 22.095 5.915 22.385 6.145 ;
      RECT 22.095 5.945 27.335 6.115 ;
      RECT 24.535 2.465 24.72 2.675 ;
      RECT 24.525 2.47 24.735 2.668 ;
      RECT 24.525 2.47 24.821 2.645 ;
      RECT 24.525 2.47 24.88 2.62 ;
      RECT 24.525 2.47 24.935 2.6 ;
      RECT 24.525 2.47 24.945 2.588 ;
      RECT 24.525 2.47 25.14 2.527 ;
      RECT 24.525 2.47 25.17 2.51 ;
      RECT 24.525 2.47 25.19 2.5 ;
      RECT 25.07 2.235 25.33 2.495 ;
      RECT 25.055 2.325 25.07 2.542 ;
      RECT 24.59 2.457 25.33 2.495 ;
      RECT 25.041 2.336 25.055 2.548 ;
      RECT 24.63 2.45 25.33 2.495 ;
      RECT 24.955 2.376 25.041 2.567 ;
      RECT 24.88 2.437 25.33 2.495 ;
      RECT 24.95 2.412 24.955 2.584 ;
      RECT 24.935 2.422 25.33 2.495 ;
      RECT 24.945 2.417 24.95 2.586 ;
      RECT 25.24 2.922 25.245 3.014 ;
      RECT 25.235 2.9 25.24 3.031 ;
      RECT 25.23 2.89 25.235 3.043 ;
      RECT 25.22 2.881 25.23 3.053 ;
      RECT 25.215 2.876 25.22 3.061 ;
      RECT 25.21 2.735 25.215 3.064 ;
      RECT 25.176 2.735 25.21 3.075 ;
      RECT 25.09 2.735 25.176 3.11 ;
      RECT 25.01 2.735 25.09 3.158 ;
      RECT 24.981 2.735 25.01 3.182 ;
      RECT 24.895 2.735 24.981 3.188 ;
      RECT 24.89 2.919 24.895 3.193 ;
      RECT 24.855 2.93 24.89 3.196 ;
      RECT 24.83 2.945 24.855 3.2 ;
      RECT 24.816 2.954 24.83 3.202 ;
      RECT 24.73 2.981 24.816 3.208 ;
      RECT 24.665 3.022 24.73 3.217 ;
      RECT 24.65 3.042 24.665 3.222 ;
      RECT 24.62 3.052 24.65 3.225 ;
      RECT 24.615 3.062 24.62 3.228 ;
      RECT 24.585 3.067 24.615 3.23 ;
      RECT 24.565 3.072 24.585 3.234 ;
      RECT 24.48 3.075 24.565 3.241 ;
      RECT 24.465 3.072 24.48 3.247 ;
      RECT 24.455 3.069 24.465 3.249 ;
      RECT 24.435 3.066 24.455 3.251 ;
      RECT 24.415 3.062 24.435 3.252 ;
      RECT 24.4 3.058 24.415 3.254 ;
      RECT 24.39 3.055 24.4 3.255 ;
      RECT 24.35 3.049 24.39 3.253 ;
      RECT 24.34 3.044 24.35 3.251 ;
      RECT 24.325 3.041 24.34 3.247 ;
      RECT 24.3 3.036 24.325 3.24 ;
      RECT 24.25 3.027 24.3 3.228 ;
      RECT 24.18 3.013 24.25 3.21 ;
      RECT 24.122 2.998 24.18 3.192 ;
      RECT 24.036 2.981 24.122 3.172 ;
      RECT 23.95 2.96 24.036 3.147 ;
      RECT 23.9 2.945 23.95 3.128 ;
      RECT 23.896 2.939 23.9 3.12 ;
      RECT 23.81 2.929 23.896 3.107 ;
      RECT 23.775 2.914 23.81 3.09 ;
      RECT 23.76 2.907 23.775 3.083 ;
      RECT 23.7 2.895 23.76 3.071 ;
      RECT 23.68 2.882 23.7 3.059 ;
      RECT 23.64 2.873 23.68 3.051 ;
      RECT 23.635 2.865 23.64 3.044 ;
      RECT 23.555 2.855 23.635 3.03 ;
      RECT 23.54 2.842 23.555 3.015 ;
      RECT 23.535 2.84 23.54 3.013 ;
      RECT 23.456 2.828 23.535 3 ;
      RECT 23.37 2.803 23.456 2.975 ;
      RECT 23.355 2.772 23.37 2.96 ;
      RECT 23.34 2.747 23.355 2.956 ;
      RECT 23.325 2.74 23.34 2.952 ;
      RECT 23.15 2.745 23.155 2.948 ;
      RECT 23.145 2.75 23.15 2.943 ;
      RECT 23.155 2.74 23.325 2.95 ;
      RECT 23.87 2.5 23.975 2.76 ;
      RECT 24.685 2.025 24.69 2.25 ;
      RECT 24.815 2.025 24.87 2.235 ;
      RECT 24.87 2.03 24.88 2.228 ;
      RECT 24.776 2.025 24.815 2.238 ;
      RECT 24.69 2.025 24.776 2.245 ;
      RECT 24.67 2.03 24.685 2.251 ;
      RECT 24.66 2.07 24.67 2.253 ;
      RECT 24.63 2.08 24.66 2.255 ;
      RECT 24.625 2.085 24.63 2.257 ;
      RECT 24.6 2.09 24.625 2.259 ;
      RECT 24.585 2.095 24.6 2.261 ;
      RECT 24.57 2.097 24.585 2.263 ;
      RECT 24.565 2.102 24.57 2.265 ;
      RECT 24.515 2.11 24.565 2.268 ;
      RECT 24.49 2.119 24.515 2.273 ;
      RECT 24.48 2.126 24.49 2.278 ;
      RECT 24.475 2.129 24.48 2.282 ;
      RECT 24.455 2.132 24.475 2.291 ;
      RECT 24.425 2.14 24.455 2.311 ;
      RECT 24.396 2.153 24.425 2.333 ;
      RECT 24.31 2.187 24.396 2.377 ;
      RECT 24.305 2.213 24.31 2.415 ;
      RECT 24.3 2.217 24.305 2.424 ;
      RECT 24.265 2.23 24.3 2.457 ;
      RECT 24.255 2.244 24.265 2.495 ;
      RECT 24.25 2.248 24.255 2.508 ;
      RECT 24.245 2.252 24.25 2.513 ;
      RECT 24.235 2.26 24.245 2.525 ;
      RECT 24.23 2.267 24.235 2.54 ;
      RECT 24.205 2.28 24.23 2.565 ;
      RECT 24.165 2.309 24.205 2.62 ;
      RECT 24.15 2.334 24.165 2.675 ;
      RECT 24.14 2.345 24.15 2.698 ;
      RECT 24.135 2.352 24.14 2.71 ;
      RECT 24.13 2.356 24.135 2.718 ;
      RECT 24.075 2.384 24.13 2.76 ;
      RECT 24.055 2.42 24.075 2.76 ;
      RECT 24.04 2.435 24.055 2.76 ;
      RECT 23.985 2.467 24.04 2.76 ;
      RECT 23.975 2.497 23.985 2.76 ;
      RECT 23.585 2.112 23.77 2.35 ;
      RECT 23.57 2.114 23.78 2.345 ;
      RECT 23.455 2.06 23.715 2.32 ;
      RECT 23.45 2.097 23.715 2.274 ;
      RECT 23.445 2.107 23.715 2.271 ;
      RECT 23.44 2.147 23.78 2.265 ;
      RECT 23.435 2.18 23.78 2.255 ;
      RECT 23.445 2.122 23.795 2.193 ;
      RECT 23.742 3.22 23.755 3.75 ;
      RECT 23.656 3.22 23.755 3.749 ;
      RECT 23.656 3.22 23.76 3.748 ;
      RECT 23.57 3.22 23.76 3.746 ;
      RECT 23.565 3.22 23.76 3.743 ;
      RECT 23.565 3.22 23.77 3.741 ;
      RECT 23.56 3.512 23.77 3.738 ;
      RECT 23.56 3.522 23.775 3.735 ;
      RECT 23.56 3.59 23.78 3.731 ;
      RECT 23.55 3.595 23.78 3.73 ;
      RECT 23.55 3.687 23.785 3.727 ;
      RECT 23.535 3.22 23.795 3.48 ;
      RECT 23.465 7.765 23.755 7.995 ;
      RECT 23.525 7.025 23.695 7.995 ;
      RECT 23.44 7.055 23.78 7.4 ;
      RECT 23.465 7.025 23.755 7.4 ;
      RECT 22.765 2.21 22.81 3.745 ;
      RECT 22.965 2.21 22.995 2.425 ;
      RECT 21.34 1.95 21.46 2.16 ;
      RECT 21 1.9 21.26 2.16 ;
      RECT 21 1.945 21.295 2.15 ;
      RECT 23.005 2.226 23.01 2.28 ;
      RECT 23 2.219 23.005 2.413 ;
      RECT 22.995 2.213 23 2.42 ;
      RECT 22.95 2.21 22.965 2.433 ;
      RECT 22.945 2.21 22.95 2.455 ;
      RECT 22.94 2.21 22.945 2.503 ;
      RECT 22.935 2.21 22.94 2.523 ;
      RECT 22.925 2.21 22.935 2.63 ;
      RECT 22.92 2.21 22.925 2.693 ;
      RECT 22.915 2.21 22.92 2.75 ;
      RECT 22.91 2.21 22.915 2.758 ;
      RECT 22.895 2.21 22.91 2.865 ;
      RECT 22.885 2.21 22.895 3 ;
      RECT 22.875 2.21 22.885 3.11 ;
      RECT 22.865 2.21 22.875 3.167 ;
      RECT 22.86 2.21 22.865 3.207 ;
      RECT 22.855 2.21 22.86 3.243 ;
      RECT 22.845 2.21 22.855 3.283 ;
      RECT 22.84 2.21 22.845 3.325 ;
      RECT 22.82 2.21 22.84 3.39 ;
      RECT 22.825 3.535 22.83 3.715 ;
      RECT 22.82 3.517 22.825 3.723 ;
      RECT 22.815 2.21 22.82 3.453 ;
      RECT 22.815 3.497 22.82 3.73 ;
      RECT 22.81 2.21 22.815 3.74 ;
      RECT 22.755 2.21 22.765 2.51 ;
      RECT 22.76 2.757 22.765 3.745 ;
      RECT 22.755 2.822 22.76 3.745 ;
      RECT 22.75 2.211 22.755 2.5 ;
      RECT 22.745 2.887 22.755 3.745 ;
      RECT 22.74 2.212 22.75 2.49 ;
      RECT 22.73 3 22.745 3.745 ;
      RECT 22.735 2.213 22.74 2.48 ;
      RECT 22.715 2.214 22.735 2.458 ;
      RECT 22.72 3.097 22.73 3.745 ;
      RECT 22.715 3.172 22.72 3.745 ;
      RECT 22.705 2.213 22.715 2.435 ;
      RECT 22.71 3.215 22.715 3.745 ;
      RECT 22.705 3.242 22.71 3.745 ;
      RECT 22.695 2.211 22.705 2.423 ;
      RECT 22.7 3.285 22.705 3.745 ;
      RECT 22.695 3.312 22.7 3.745 ;
      RECT 22.685 2.21 22.695 2.41 ;
      RECT 22.69 3.327 22.695 3.745 ;
      RECT 22.65 3.385 22.69 3.745 ;
      RECT 22.68 2.209 22.685 2.395 ;
      RECT 22.675 2.207 22.68 2.388 ;
      RECT 22.665 2.204 22.675 2.378 ;
      RECT 22.66 2.201 22.665 2.363 ;
      RECT 22.645 2.197 22.66 2.356 ;
      RECT 22.64 3.44 22.65 3.745 ;
      RECT 22.64 2.194 22.645 2.351 ;
      RECT 22.625 2.19 22.64 2.345 ;
      RECT 22.635 3.457 22.64 3.745 ;
      RECT 22.625 3.52 22.635 3.745 ;
      RECT 22.545 2.175 22.625 2.325 ;
      RECT 22.62 3.527 22.625 3.74 ;
      RECT 22.615 3.535 22.62 3.73 ;
      RECT 22.535 2.161 22.545 2.309 ;
      RECT 22.52 2.157 22.535 2.307 ;
      RECT 22.51 2.152 22.52 2.303 ;
      RECT 22.485 2.145 22.51 2.295 ;
      RECT 22.48 2.14 22.485 2.29 ;
      RECT 22.47 2.14 22.48 2.288 ;
      RECT 22.46 2.138 22.47 2.286 ;
      RECT 22.43 2.13 22.46 2.28 ;
      RECT 22.415 2.122 22.43 2.273 ;
      RECT 22.395 2.117 22.415 2.266 ;
      RECT 22.39 2.113 22.395 2.261 ;
      RECT 22.36 2.106 22.39 2.255 ;
      RECT 22.335 2.097 22.36 2.245 ;
      RECT 22.305 2.09 22.335 2.237 ;
      RECT 22.28 2.08 22.305 2.228 ;
      RECT 22.265 2.072 22.28 2.222 ;
      RECT 22.24 2.067 22.265 2.217 ;
      RECT 22.23 2.063 22.24 2.212 ;
      RECT 22.21 2.058 22.23 2.207 ;
      RECT 22.175 2.053 22.21 2.2 ;
      RECT 22.115 2.048 22.175 2.193 ;
      RECT 22.102 2.044 22.115 2.191 ;
      RECT 22.016 2.039 22.102 2.188 ;
      RECT 21.93 2.029 22.016 2.184 ;
      RECT 21.889 2.022 21.93 2.181 ;
      RECT 21.803 2.015 21.889 2.178 ;
      RECT 21.717 2.005 21.803 2.174 ;
      RECT 21.631 1.995 21.717 2.169 ;
      RECT 21.545 1.985 21.631 2.165 ;
      RECT 21.535 1.97 21.545 2.163 ;
      RECT 21.525 1.955 21.535 2.163 ;
      RECT 21.46 1.95 21.525 2.162 ;
      RECT 21.295 1.947 21.34 2.155 ;
      RECT 22.54 2.852 22.545 3.043 ;
      RECT 22.535 2.847 22.54 3.05 ;
      RECT 22.521 2.845 22.535 3.056 ;
      RECT 22.435 2.845 22.521 3.058 ;
      RECT 22.431 2.845 22.435 3.061 ;
      RECT 22.345 2.845 22.431 3.079 ;
      RECT 22.335 2.85 22.345 3.098 ;
      RECT 22.325 2.905 22.335 3.102 ;
      RECT 22.3 2.92 22.325 3.109 ;
      RECT 22.26 2.94 22.3 3.122 ;
      RECT 22.255 2.952 22.26 3.132 ;
      RECT 22.24 2.958 22.255 3.137 ;
      RECT 22.235 2.963 22.24 3.141 ;
      RECT 22.215 2.97 22.235 3.146 ;
      RECT 22.145 2.995 22.215 3.163 ;
      RECT 22.105 3.023 22.145 3.183 ;
      RECT 22.1 3.033 22.105 3.191 ;
      RECT 22.08 3.04 22.1 3.193 ;
      RECT 22.075 3.047 22.08 3.196 ;
      RECT 22.045 3.055 22.075 3.199 ;
      RECT 22.04 3.06 22.045 3.203 ;
      RECT 21.966 3.064 22.04 3.211 ;
      RECT 21.88 3.073 21.966 3.227 ;
      RECT 21.876 3.078 21.88 3.236 ;
      RECT 21.79 3.083 21.876 3.246 ;
      RECT 21.75 3.091 21.79 3.258 ;
      RECT 21.7 3.097 21.75 3.265 ;
      RECT 21.615 3.106 21.7 3.28 ;
      RECT 21.54 3.117 21.615 3.298 ;
      RECT 21.505 3.124 21.54 3.308 ;
      RECT 21.43 3.132 21.505 3.313 ;
      RECT 21.375 3.141 21.43 3.313 ;
      RECT 21.35 3.146 21.375 3.311 ;
      RECT 21.34 3.149 21.35 3.309 ;
      RECT 21.305 3.151 21.34 3.307 ;
      RECT 21.275 3.153 21.305 3.303 ;
      RECT 21.23 3.152 21.275 3.299 ;
      RECT 21.21 3.147 21.23 3.296 ;
      RECT 21.16 3.132 21.21 3.293 ;
      RECT 21.15 3.117 21.16 3.288 ;
      RECT 21.1 3.102 21.15 3.278 ;
      RECT 21.05 3.077 21.1 3.258 ;
      RECT 21.04 3.062 21.05 3.24 ;
      RECT 21.035 3.06 21.04 3.234 ;
      RECT 21.015 3.055 21.035 3.229 ;
      RECT 21.01 3.047 21.015 3.223 ;
      RECT 20.995 3.041 21.01 3.216 ;
      RECT 20.99 3.036 20.995 3.208 ;
      RECT 20.97 3.031 20.99 3.2 ;
      RECT 20.955 3.024 20.97 3.193 ;
      RECT 20.94 3.018 20.955 3.184 ;
      RECT 20.935 3.012 20.94 3.177 ;
      RECT 20.89 2.987 20.935 3.163 ;
      RECT 20.875 2.957 20.89 3.145 ;
      RECT 20.86 2.94 20.875 3.136 ;
      RECT 20.835 2.92 20.86 3.124 ;
      RECT 20.795 2.89 20.835 3.104 ;
      RECT 20.785 2.86 20.795 3.089 ;
      RECT 20.77 2.85 20.785 3.082 ;
      RECT 20.715 2.815 20.77 3.061 ;
      RECT 20.7 2.778 20.715 3.04 ;
      RECT 20.69 2.765 20.7 3.032 ;
      RECT 20.64 2.735 20.69 3.014 ;
      RECT 20.625 2.665 20.64 2.995 ;
      RECT 20.58 2.665 20.625 2.978 ;
      RECT 20.555 2.665 20.58 2.96 ;
      RECT 20.545 2.665 20.555 2.953 ;
      RECT 20.466 2.665 20.545 2.946 ;
      RECT 20.38 2.665 20.466 2.938 ;
      RECT 20.365 2.697 20.38 2.933 ;
      RECT 20.29 2.707 20.365 2.929 ;
      RECT 20.27 2.717 20.29 2.924 ;
      RECT 20.245 2.717 20.27 2.921 ;
      RECT 20.235 2.707 20.245 2.92 ;
      RECT 20.225 2.68 20.235 2.919 ;
      RECT 20.185 2.675 20.225 2.917 ;
      RECT 20.14 2.675 20.185 2.913 ;
      RECT 20.115 2.675 20.14 2.908 ;
      RECT 20.065 2.675 20.115 2.895 ;
      RECT 20.025 2.68 20.035 2.88 ;
      RECT 20.035 2.675 20.065 2.885 ;
      RECT 22.02 2.455 22.28 2.715 ;
      RECT 22.015 2.477 22.28 2.673 ;
      RECT 21.255 2.305 21.475 2.67 ;
      RECT 21.237 2.392 21.475 2.669 ;
      RECT 21.22 2.397 21.475 2.666 ;
      RECT 21.22 2.397 21.495 2.665 ;
      RECT 21.19 2.407 21.495 2.663 ;
      RECT 21.185 2.422 21.495 2.659 ;
      RECT 21.185 2.422 21.5 2.658 ;
      RECT 21.18 2.48 21.5 2.656 ;
      RECT 21.18 2.48 21.51 2.653 ;
      RECT 21.175 2.545 21.51 2.648 ;
      RECT 21.255 2.305 21.515 2.565 ;
      RECT 20 2.135 20.26 2.395 ;
      RECT 20 2.178 20.346 2.369 ;
      RECT 20 2.178 20.39 2.368 ;
      RECT 20 2.178 20.41 2.366 ;
      RECT 20 2.178 20.51 2.365 ;
      RECT 20 2.178 20.53 2.363 ;
      RECT 20 2.178 20.54 2.358 ;
      RECT 20.41 2.145 20.6 2.355 ;
      RECT 20.41 2.147 20.605 2.353 ;
      RECT 20.4 2.152 20.61 2.345 ;
      RECT 20.346 2.176 20.61 2.345 ;
      RECT 20.39 2.17 20.4 2.367 ;
      RECT 20.4 2.15 20.605 2.353 ;
      RECT 19.355 3.21 19.56 3.44 ;
      RECT 19.295 3.16 19.35 3.42 ;
      RECT 19.355 3.16 19.555 3.44 ;
      RECT 20.325 3.475 20.33 3.502 ;
      RECT 20.315 3.385 20.325 3.507 ;
      RECT 20.31 3.307 20.315 3.513 ;
      RECT 20.3 3.297 20.31 3.52 ;
      RECT 20.295 3.287 20.3 3.526 ;
      RECT 20.285 3.282 20.295 3.528 ;
      RECT 20.27 3.274 20.285 3.536 ;
      RECT 20.255 3.265 20.27 3.548 ;
      RECT 20.245 3.257 20.255 3.558 ;
      RECT 20.21 3.175 20.245 3.576 ;
      RECT 20.175 3.175 20.21 3.595 ;
      RECT 20.16 3.175 20.175 3.603 ;
      RECT 20.105 3.175 20.16 3.603 ;
      RECT 20.071 3.175 20.105 3.594 ;
      RECT 19.985 3.175 20.071 3.57 ;
      RECT 19.975 3.235 19.985 3.552 ;
      RECT 19.935 3.237 19.975 3.543 ;
      RECT 19.93 3.239 19.935 3.533 ;
      RECT 19.91 3.241 19.93 3.528 ;
      RECT 19.9 3.244 19.91 3.523 ;
      RECT 19.89 3.245 19.9 3.518 ;
      RECT 19.866 3.246 19.89 3.51 ;
      RECT 19.78 3.251 19.866 3.488 ;
      RECT 19.725 3.25 19.78 3.461 ;
      RECT 19.71 3.243 19.725 3.448 ;
      RECT 19.675 3.238 19.71 3.444 ;
      RECT 19.62 3.23 19.675 3.443 ;
      RECT 19.56 3.217 19.62 3.441 ;
      RECT 19.35 3.16 19.355 3.428 ;
      RECT 19.425 2.53 19.61 2.74 ;
      RECT 19.415 2.535 19.625 2.733 ;
      RECT 19.455 2.44 19.715 2.7 ;
      RECT 19.41 2.597 19.715 2.623 ;
      RECT 18.755 2.39 18.76 3.19 ;
      RECT 18.7 2.44 18.73 3.19 ;
      RECT 18.69 2.44 18.695 2.75 ;
      RECT 18.675 2.44 18.68 2.745 ;
      RECT 18.22 2.485 18.235 2.7 ;
      RECT 18.15 2.485 18.235 2.695 ;
      RECT 19.415 2.065 19.485 2.275 ;
      RECT 19.485 2.072 19.495 2.27 ;
      RECT 19.381 2.065 19.415 2.282 ;
      RECT 19.295 2.065 19.381 2.306 ;
      RECT 19.285 2.07 19.295 2.325 ;
      RECT 19.28 2.082 19.285 2.328 ;
      RECT 19.265 2.097 19.28 2.332 ;
      RECT 19.26 2.115 19.265 2.336 ;
      RECT 19.22 2.125 19.26 2.345 ;
      RECT 19.205 2.132 19.22 2.357 ;
      RECT 19.19 2.137 19.205 2.362 ;
      RECT 19.175 2.14 19.19 2.367 ;
      RECT 19.165 2.142 19.175 2.371 ;
      RECT 19.13 2.149 19.165 2.379 ;
      RECT 19.095 2.157 19.13 2.393 ;
      RECT 19.085 2.163 19.095 2.402 ;
      RECT 19.08 2.165 19.085 2.404 ;
      RECT 19.06 2.168 19.08 2.41 ;
      RECT 19.03 2.175 19.06 2.421 ;
      RECT 19.02 2.181 19.03 2.428 ;
      RECT 18.995 2.184 19.02 2.435 ;
      RECT 18.985 2.188 18.995 2.443 ;
      RECT 18.98 2.189 18.985 2.465 ;
      RECT 18.975 2.19 18.98 2.48 ;
      RECT 18.97 2.191 18.975 2.495 ;
      RECT 18.965 2.192 18.97 2.51 ;
      RECT 18.96 2.193 18.965 2.54 ;
      RECT 18.95 2.195 18.96 2.573 ;
      RECT 18.935 2.199 18.95 2.62 ;
      RECT 18.925 2.202 18.935 2.665 ;
      RECT 18.92 2.205 18.925 2.693 ;
      RECT 18.91 2.207 18.92 2.72 ;
      RECT 18.905 2.21 18.91 2.755 ;
      RECT 18.875 2.215 18.905 2.813 ;
      RECT 18.87 2.22 18.875 2.898 ;
      RECT 18.865 2.222 18.87 2.933 ;
      RECT 18.86 2.224 18.865 3.015 ;
      RECT 18.855 2.226 18.86 3.103 ;
      RECT 18.845 2.228 18.855 3.185 ;
      RECT 18.83 2.242 18.845 3.19 ;
      RECT 18.795 2.287 18.83 3.19 ;
      RECT 18.785 2.327 18.795 3.19 ;
      RECT 18.77 2.355 18.785 3.19 ;
      RECT 18.765 2.372 18.77 3.19 ;
      RECT 18.76 2.38 18.765 3.19 ;
      RECT 18.75 2.395 18.755 3.19 ;
      RECT 18.745 2.402 18.75 3.19 ;
      RECT 18.735 2.422 18.745 3.19 ;
      RECT 18.73 2.435 18.735 3.19 ;
      RECT 18.695 2.44 18.7 2.775 ;
      RECT 18.68 2.83 18.7 3.19 ;
      RECT 18.68 2.44 18.69 2.748 ;
      RECT 18.675 2.87 18.68 3.19 ;
      RECT 18.625 2.44 18.675 2.743 ;
      RECT 18.67 2.907 18.675 3.19 ;
      RECT 18.66 2.93 18.67 3.19 ;
      RECT 18.655 2.975 18.66 3.19 ;
      RECT 18.645 2.985 18.655 3.183 ;
      RECT 18.571 2.44 18.625 2.737 ;
      RECT 18.485 2.44 18.571 2.73 ;
      RECT 18.436 2.487 18.485 2.723 ;
      RECT 18.35 2.495 18.436 2.716 ;
      RECT 18.335 2.492 18.35 2.711 ;
      RECT 18.321 2.485 18.335 2.71 ;
      RECT 18.235 2.485 18.321 2.705 ;
      RECT 18.14 2.49 18.15 2.69 ;
      RECT 17.73 1.92 17.745 2.32 ;
      RECT 17.925 1.92 17.93 2.18 ;
      RECT 17.67 1.92 17.715 2.18 ;
      RECT 18.125 3.225 18.13 3.43 ;
      RECT 18.12 3.215 18.125 3.435 ;
      RECT 18.115 3.202 18.12 3.44 ;
      RECT 18.11 3.182 18.115 3.44 ;
      RECT 18.085 3.135 18.11 3.44 ;
      RECT 18.05 3.05 18.085 3.44 ;
      RECT 18.045 2.987 18.05 3.44 ;
      RECT 18.04 2.972 18.045 3.44 ;
      RECT 18.025 2.932 18.04 3.44 ;
      RECT 18.02 2.907 18.025 3.44 ;
      RECT 18.01 2.89 18.02 3.44 ;
      RECT 17.975 2.812 18.01 3.44 ;
      RECT 17.97 2.755 17.975 3.44 ;
      RECT 17.965 2.742 17.97 3.44 ;
      RECT 17.955 2.72 17.965 3.44 ;
      RECT 17.945 2.685 17.955 3.44 ;
      RECT 17.935 2.655 17.945 3.44 ;
      RECT 17.925 2.57 17.935 3.083 ;
      RECT 17.932 3.215 17.935 3.44 ;
      RECT 17.93 3.225 17.932 3.44 ;
      RECT 17.92 3.235 17.93 3.435 ;
      RECT 17.915 1.92 17.925 2.315 ;
      RECT 17.92 2.447 17.925 3.058 ;
      RECT 17.915 2.345 17.92 3.041 ;
      RECT 17.905 1.92 17.915 3.017 ;
      RECT 17.9 1.92 17.905 2.988 ;
      RECT 17.895 1.92 17.9 2.978 ;
      RECT 17.875 1.92 17.895 2.94 ;
      RECT 17.87 1.92 17.875 2.898 ;
      RECT 17.865 1.92 17.87 2.878 ;
      RECT 17.835 1.92 17.865 2.828 ;
      RECT 17.825 1.92 17.835 2.775 ;
      RECT 17.82 1.92 17.825 2.748 ;
      RECT 17.815 1.92 17.82 2.733 ;
      RECT 17.805 1.92 17.815 2.71 ;
      RECT 17.795 1.92 17.805 2.685 ;
      RECT 17.79 1.92 17.795 2.625 ;
      RECT 17.78 1.92 17.79 2.563 ;
      RECT 17.775 1.92 17.78 2.483 ;
      RECT 17.77 1.92 17.775 2.448 ;
      RECT 17.765 1.92 17.77 2.423 ;
      RECT 17.76 1.92 17.765 2.408 ;
      RECT 17.755 1.92 17.76 2.378 ;
      RECT 17.75 1.92 17.755 2.355 ;
      RECT 17.745 1.92 17.75 2.328 ;
      RECT 17.715 1.92 17.73 2.315 ;
      RECT 16.87 3.455 17.055 3.665 ;
      RECT 16.86 3.46 17.07 3.658 ;
      RECT 16.86 3.46 17.09 3.63 ;
      RECT 16.86 3.46 17.105 3.609 ;
      RECT 16.86 3.46 17.12 3.607 ;
      RECT 16.86 3.46 17.13 3.606 ;
      RECT 16.86 3.46 17.16 3.603 ;
      RECT 17.51 3.305 17.77 3.565 ;
      RECT 17.47 3.352 17.77 3.548 ;
      RECT 17.461 3.36 17.47 3.551 ;
      RECT 17.055 3.453 17.77 3.548 ;
      RECT 17.375 3.378 17.461 3.558 ;
      RECT 17.07 3.45 17.77 3.548 ;
      RECT 17.316 3.4 17.375 3.57 ;
      RECT 17.09 3.446 17.77 3.548 ;
      RECT 17.23 3.412 17.316 3.581 ;
      RECT 17.105 3.442 17.77 3.548 ;
      RECT 17.175 3.425 17.23 3.593 ;
      RECT 17.12 3.44 17.77 3.548 ;
      RECT 17.16 3.431 17.175 3.599 ;
      RECT 17.13 3.436 17.77 3.548 ;
      RECT 17.275 2.96 17.535 3.22 ;
      RECT 17.275 2.98 17.645 3.19 ;
      RECT 17.275 2.985 17.655 3.185 ;
      RECT 17.466 2.399 17.545 2.63 ;
      RECT 17.38 2.402 17.595 2.625 ;
      RECT 17.375 2.402 17.595 2.62 ;
      RECT 17.375 2.407 17.605 2.618 ;
      RECT 17.35 2.407 17.605 2.615 ;
      RECT 17.35 2.415 17.615 2.613 ;
      RECT 17.23 2.35 17.49 2.61 ;
      RECT 17.23 2.397 17.54 2.61 ;
      RECT 16.485 2.97 16.49 3.23 ;
      RECT 16.315 2.74 16.32 3.23 ;
      RECT 16.2 2.98 16.205 3.205 ;
      RECT 16.91 2.075 16.915 2.285 ;
      RECT 16.915 2.08 16.93 2.28 ;
      RECT 16.85 2.075 16.91 2.293 ;
      RECT 16.835 2.075 16.85 2.303 ;
      RECT 16.785 2.075 16.835 2.32 ;
      RECT 16.765 2.075 16.785 2.343 ;
      RECT 16.75 2.075 16.765 2.355 ;
      RECT 16.73 2.075 16.75 2.365 ;
      RECT 16.72 2.08 16.73 2.374 ;
      RECT 16.715 2.09 16.72 2.379 ;
      RECT 16.71 2.102 16.715 2.383 ;
      RECT 16.7 2.125 16.71 2.388 ;
      RECT 16.695 2.14 16.7 2.392 ;
      RECT 16.69 2.157 16.695 2.395 ;
      RECT 16.685 2.165 16.69 2.398 ;
      RECT 16.675 2.17 16.685 2.402 ;
      RECT 16.67 2.177 16.675 2.407 ;
      RECT 16.66 2.182 16.67 2.411 ;
      RECT 16.635 2.194 16.66 2.422 ;
      RECT 16.615 2.211 16.635 2.438 ;
      RECT 16.59 2.228 16.615 2.46 ;
      RECT 16.555 2.251 16.59 2.518 ;
      RECT 16.535 2.273 16.555 2.58 ;
      RECT 16.53 2.283 16.535 2.615 ;
      RECT 16.52 2.29 16.53 2.653 ;
      RECT 16.515 2.297 16.52 2.673 ;
      RECT 16.51 2.308 16.515 2.71 ;
      RECT 16.505 2.316 16.51 2.775 ;
      RECT 16.495 2.327 16.505 2.828 ;
      RECT 16.49 2.345 16.495 2.898 ;
      RECT 16.485 2.355 16.49 2.935 ;
      RECT 16.48 2.365 16.485 3.23 ;
      RECT 16.475 2.377 16.48 3.23 ;
      RECT 16.47 2.387 16.475 3.23 ;
      RECT 16.46 2.397 16.47 3.23 ;
      RECT 16.45 2.42 16.46 3.23 ;
      RECT 16.435 2.455 16.45 3.23 ;
      RECT 16.395 2.517 16.435 3.23 ;
      RECT 16.39 2.57 16.395 3.23 ;
      RECT 16.365 2.605 16.39 3.23 ;
      RECT 16.35 2.65 16.365 3.23 ;
      RECT 16.345 2.672 16.35 3.23 ;
      RECT 16.335 2.685 16.345 3.23 ;
      RECT 16.325 2.71 16.335 3.23 ;
      RECT 16.32 2.732 16.325 3.23 ;
      RECT 16.295 2.77 16.315 3.23 ;
      RECT 16.255 2.827 16.295 3.23 ;
      RECT 16.25 2.877 16.255 3.23 ;
      RECT 16.245 2.895 16.25 3.23 ;
      RECT 16.24 2.907 16.245 3.23 ;
      RECT 16.23 2.925 16.24 3.23 ;
      RECT 16.22 2.945 16.23 3.205 ;
      RECT 16.215 2.962 16.22 3.205 ;
      RECT 16.205 2.975 16.215 3.205 ;
      RECT 16.175 2.985 16.2 3.205 ;
      RECT 16.165 2.992 16.175 3.205 ;
      RECT 16.15 3.002 16.165 3.2 ;
      RECT 15.25 7.765 15.54 7.995 ;
      RECT 15.31 6.285 15.48 7.995 ;
      RECT 15.3 6.655 15.65 7.005 ;
      RECT 15.25 6.285 15.54 6.515 ;
      RECT 15.25 2.365 15.54 2.595 ;
      RECT 15.31 0.885 15.48 2.595 ;
      RECT 15.25 0.885 15.54 1.115 ;
      RECT 14.84 2.735 15.17 2.965 ;
      RECT 14.84 2.765 15.34 2.935 ;
      RECT 14.84 2.395 15.03 2.965 ;
      RECT 14.26 2.365 14.55 2.595 ;
      RECT 14.26 2.395 15.03 2.565 ;
      RECT 14.32 0.885 14.49 2.595 ;
      RECT 14.26 0.885 14.55 1.115 ;
      RECT 14.26 7.765 14.55 7.995 ;
      RECT 14.32 6.285 14.49 7.995 ;
      RECT 14.26 6.285 14.55 6.515 ;
      RECT 14.26 6.325 15.11 6.485 ;
      RECT 14.94 5.915 15.11 6.485 ;
      RECT 14.26 6.32 14.65 6.485 ;
      RECT 14.88 5.915 15.17 6.145 ;
      RECT 14.88 5.945 15.34 6.115 ;
      RECT 13.89 2.735 14.18 2.965 ;
      RECT 13.89 2.765 14.35 2.935 ;
      RECT 13.95 1.655 14.115 2.965 ;
      RECT 12.465 1.625 12.755 1.855 ;
      RECT 12.465 1.655 14.115 1.825 ;
      RECT 12.525 0.885 12.695 1.855 ;
      RECT 12.465 0.885 12.755 1.115 ;
      RECT 12.465 7.765 12.755 7.995 ;
      RECT 12.525 7.025 12.695 7.995 ;
      RECT 12.525 7.12 14.115 7.29 ;
      RECT 13.945 5.915 14.115 7.29 ;
      RECT 12.465 7.025 12.755 7.255 ;
      RECT 13.89 5.915 14.18 6.145 ;
      RECT 13.89 5.945 14.35 6.115 ;
      RECT 12.895 1.965 13.245 2.315 ;
      RECT 10.56 2.025 13.245 2.195 ;
      RECT 10.56 1.34 10.73 2.195 ;
      RECT 10.46 1.34 10.81 1.69 ;
      RECT 12.92 6.655 13.245 6.98 ;
      RECT 8.315 6.605 8.665 6.955 ;
      RECT 12.895 6.655 13.245 6.885 ;
      RECT 8.115 6.655 8.665 6.885 ;
      RECT 7.945 6.685 13.245 6.855 ;
      RECT 12.12 2.365 12.44 2.685 ;
      RECT 12.09 2.365 12.44 2.595 ;
      RECT 11.92 2.395 12.44 2.565 ;
      RECT 12.12 6.255 12.44 6.545 ;
      RECT 12.09 6.285 12.44 6.515 ;
      RECT 11.92 6.315 12.44 6.485 ;
      RECT 11.065 2.705 11.415 3.055 ;
      RECT 11.065 2.765 11.555 2.935 ;
      RECT 11.07 5.855 11.42 6.205 ;
      RECT 6.315 5.915 6.605 6.145 ;
      RECT 6.315 5.945 11.555 6.115 ;
      RECT 8.755 2.465 8.94 2.675 ;
      RECT 8.745 2.47 8.955 2.668 ;
      RECT 8.745 2.47 9.041 2.645 ;
      RECT 8.745 2.47 9.1 2.62 ;
      RECT 8.745 2.47 9.155 2.6 ;
      RECT 8.745 2.47 9.165 2.588 ;
      RECT 8.745 2.47 9.36 2.527 ;
      RECT 8.745 2.47 9.39 2.51 ;
      RECT 8.745 2.47 9.41 2.5 ;
      RECT 9.29 2.235 9.55 2.495 ;
      RECT 9.275 2.325 9.29 2.542 ;
      RECT 8.81 2.457 9.55 2.495 ;
      RECT 9.261 2.336 9.275 2.548 ;
      RECT 8.85 2.45 9.55 2.495 ;
      RECT 9.175 2.376 9.261 2.567 ;
      RECT 9.1 2.437 9.55 2.495 ;
      RECT 9.17 2.412 9.175 2.584 ;
      RECT 9.155 2.422 9.55 2.495 ;
      RECT 9.165 2.417 9.17 2.586 ;
      RECT 9.46 2.922 9.465 3.014 ;
      RECT 9.455 2.9 9.46 3.031 ;
      RECT 9.45 2.89 9.455 3.043 ;
      RECT 9.44 2.881 9.45 3.053 ;
      RECT 9.435 2.876 9.44 3.061 ;
      RECT 9.43 2.735 9.435 3.064 ;
      RECT 9.396 2.735 9.43 3.075 ;
      RECT 9.31 2.735 9.396 3.11 ;
      RECT 9.23 2.735 9.31 3.158 ;
      RECT 9.201 2.735 9.23 3.182 ;
      RECT 9.115 2.735 9.201 3.188 ;
      RECT 9.11 2.919 9.115 3.193 ;
      RECT 9.075 2.93 9.11 3.196 ;
      RECT 9.05 2.945 9.075 3.2 ;
      RECT 9.036 2.954 9.05 3.202 ;
      RECT 8.95 2.981 9.036 3.208 ;
      RECT 8.885 3.022 8.95 3.217 ;
      RECT 8.87 3.042 8.885 3.222 ;
      RECT 8.84 3.052 8.87 3.225 ;
      RECT 8.835 3.062 8.84 3.228 ;
      RECT 8.805 3.067 8.835 3.23 ;
      RECT 8.785 3.072 8.805 3.234 ;
      RECT 8.7 3.075 8.785 3.241 ;
      RECT 8.685 3.072 8.7 3.247 ;
      RECT 8.675 3.069 8.685 3.249 ;
      RECT 8.655 3.066 8.675 3.251 ;
      RECT 8.635 3.062 8.655 3.252 ;
      RECT 8.62 3.058 8.635 3.254 ;
      RECT 8.61 3.055 8.62 3.255 ;
      RECT 8.57 3.049 8.61 3.253 ;
      RECT 8.56 3.044 8.57 3.251 ;
      RECT 8.545 3.041 8.56 3.247 ;
      RECT 8.52 3.036 8.545 3.24 ;
      RECT 8.47 3.027 8.52 3.228 ;
      RECT 8.4 3.013 8.47 3.21 ;
      RECT 8.342 2.998 8.4 3.192 ;
      RECT 8.256 2.981 8.342 3.172 ;
      RECT 8.17 2.96 8.256 3.147 ;
      RECT 8.12 2.945 8.17 3.128 ;
      RECT 8.116 2.939 8.12 3.12 ;
      RECT 8.03 2.929 8.116 3.107 ;
      RECT 7.995 2.914 8.03 3.09 ;
      RECT 7.98 2.907 7.995 3.083 ;
      RECT 7.92 2.895 7.98 3.071 ;
      RECT 7.9 2.882 7.92 3.059 ;
      RECT 7.86 2.873 7.9 3.051 ;
      RECT 7.855 2.865 7.86 3.044 ;
      RECT 7.775 2.855 7.855 3.03 ;
      RECT 7.76 2.842 7.775 3.015 ;
      RECT 7.755 2.84 7.76 3.013 ;
      RECT 7.676 2.828 7.755 3 ;
      RECT 7.59 2.803 7.676 2.975 ;
      RECT 7.575 2.772 7.59 2.96 ;
      RECT 7.56 2.747 7.575 2.956 ;
      RECT 7.545 2.74 7.56 2.952 ;
      RECT 7.37 2.745 7.375 2.948 ;
      RECT 7.365 2.75 7.37 2.943 ;
      RECT 7.375 2.74 7.545 2.95 ;
      RECT 8.09 2.5 8.195 2.76 ;
      RECT 8.905 2.025 8.91 2.25 ;
      RECT 9.035 2.025 9.09 2.235 ;
      RECT 9.09 2.03 9.1 2.228 ;
      RECT 8.996 2.025 9.035 2.238 ;
      RECT 8.91 2.025 8.996 2.245 ;
      RECT 8.89 2.03 8.905 2.251 ;
      RECT 8.88 2.07 8.89 2.253 ;
      RECT 8.85 2.08 8.88 2.255 ;
      RECT 8.845 2.085 8.85 2.257 ;
      RECT 8.82 2.09 8.845 2.259 ;
      RECT 8.805 2.095 8.82 2.261 ;
      RECT 8.79 2.097 8.805 2.263 ;
      RECT 8.785 2.102 8.79 2.265 ;
      RECT 8.735 2.11 8.785 2.268 ;
      RECT 8.71 2.119 8.735 2.273 ;
      RECT 8.7 2.126 8.71 2.278 ;
      RECT 8.695 2.129 8.7 2.282 ;
      RECT 8.675 2.132 8.695 2.291 ;
      RECT 8.645 2.14 8.675 2.311 ;
      RECT 8.616 2.153 8.645 2.333 ;
      RECT 8.53 2.187 8.616 2.377 ;
      RECT 8.525 2.213 8.53 2.415 ;
      RECT 8.52 2.217 8.525 2.424 ;
      RECT 8.485 2.23 8.52 2.457 ;
      RECT 8.475 2.244 8.485 2.495 ;
      RECT 8.47 2.248 8.475 2.508 ;
      RECT 8.465 2.252 8.47 2.513 ;
      RECT 8.455 2.26 8.465 2.525 ;
      RECT 8.45 2.267 8.455 2.54 ;
      RECT 8.425 2.28 8.45 2.565 ;
      RECT 8.385 2.309 8.425 2.62 ;
      RECT 8.37 2.334 8.385 2.675 ;
      RECT 8.36 2.345 8.37 2.698 ;
      RECT 8.355 2.352 8.36 2.71 ;
      RECT 8.35 2.356 8.355 2.718 ;
      RECT 8.295 2.384 8.35 2.76 ;
      RECT 8.275 2.42 8.295 2.76 ;
      RECT 8.26 2.435 8.275 2.76 ;
      RECT 8.205 2.467 8.26 2.76 ;
      RECT 8.195 2.497 8.205 2.76 ;
      RECT 7.805 2.112 7.99 2.35 ;
      RECT 7.79 2.114 8 2.345 ;
      RECT 7.675 2.06 7.935 2.32 ;
      RECT 7.67 2.097 7.935 2.274 ;
      RECT 7.665 2.107 7.935 2.271 ;
      RECT 7.66 2.147 8 2.265 ;
      RECT 7.655 2.18 8 2.255 ;
      RECT 7.665 2.122 8.015 2.193 ;
      RECT 7.962 3.22 7.975 3.75 ;
      RECT 7.876 3.22 7.975 3.749 ;
      RECT 7.876 3.22 7.98 3.748 ;
      RECT 7.79 3.22 7.98 3.746 ;
      RECT 7.785 3.22 7.98 3.743 ;
      RECT 7.785 3.22 7.99 3.741 ;
      RECT 7.78 3.512 7.99 3.738 ;
      RECT 7.78 3.522 7.995 3.735 ;
      RECT 7.78 3.59 8 3.731 ;
      RECT 7.77 3.595 8 3.73 ;
      RECT 7.77 3.687 8.005 3.727 ;
      RECT 7.755 3.22 8.015 3.48 ;
      RECT 7.685 7.765 7.975 7.995 ;
      RECT 7.745 7.025 7.915 7.995 ;
      RECT 7.66 7.055 8 7.4 ;
      RECT 7.685 7.025 7.975 7.4 ;
      RECT 6.985 2.21 7.03 3.745 ;
      RECT 7.185 2.21 7.215 2.425 ;
      RECT 5.56 1.95 5.68 2.16 ;
      RECT 5.22 1.9 5.48 2.16 ;
      RECT 5.22 1.945 5.515 2.15 ;
      RECT 7.225 2.226 7.23 2.28 ;
      RECT 7.22 2.219 7.225 2.413 ;
      RECT 7.215 2.213 7.22 2.42 ;
      RECT 7.17 2.21 7.185 2.433 ;
      RECT 7.165 2.21 7.17 2.455 ;
      RECT 7.16 2.21 7.165 2.503 ;
      RECT 7.155 2.21 7.16 2.523 ;
      RECT 7.145 2.21 7.155 2.63 ;
      RECT 7.14 2.21 7.145 2.693 ;
      RECT 7.135 2.21 7.14 2.75 ;
      RECT 7.13 2.21 7.135 2.758 ;
      RECT 7.115 2.21 7.13 2.865 ;
      RECT 7.105 2.21 7.115 3 ;
      RECT 7.095 2.21 7.105 3.11 ;
      RECT 7.085 2.21 7.095 3.167 ;
      RECT 7.08 2.21 7.085 3.207 ;
      RECT 7.075 2.21 7.08 3.243 ;
      RECT 7.065 2.21 7.075 3.283 ;
      RECT 7.06 2.21 7.065 3.325 ;
      RECT 7.04 2.21 7.06 3.39 ;
      RECT 7.045 3.535 7.05 3.715 ;
      RECT 7.04 3.517 7.045 3.723 ;
      RECT 7.035 2.21 7.04 3.453 ;
      RECT 7.035 3.497 7.04 3.73 ;
      RECT 7.03 2.21 7.035 3.74 ;
      RECT 6.975 2.21 6.985 2.51 ;
      RECT 6.98 2.757 6.985 3.745 ;
      RECT 6.975 2.822 6.98 3.745 ;
      RECT 6.97 2.211 6.975 2.5 ;
      RECT 6.965 2.887 6.975 3.745 ;
      RECT 6.96 2.212 6.97 2.49 ;
      RECT 6.95 3 6.965 3.745 ;
      RECT 6.955 2.213 6.96 2.48 ;
      RECT 6.935 2.214 6.955 2.458 ;
      RECT 6.94 3.097 6.95 3.745 ;
      RECT 6.935 3.172 6.94 3.745 ;
      RECT 6.925 2.213 6.935 2.435 ;
      RECT 6.93 3.215 6.935 3.745 ;
      RECT 6.925 3.242 6.93 3.745 ;
      RECT 6.915 2.211 6.925 2.423 ;
      RECT 6.92 3.285 6.925 3.745 ;
      RECT 6.915 3.312 6.92 3.745 ;
      RECT 6.905 2.21 6.915 2.41 ;
      RECT 6.91 3.327 6.915 3.745 ;
      RECT 6.87 3.385 6.91 3.745 ;
      RECT 6.9 2.209 6.905 2.395 ;
      RECT 6.895 2.207 6.9 2.388 ;
      RECT 6.885 2.204 6.895 2.378 ;
      RECT 6.88 2.201 6.885 2.363 ;
      RECT 6.865 2.197 6.88 2.356 ;
      RECT 6.86 3.44 6.87 3.745 ;
      RECT 6.86 2.194 6.865 2.351 ;
      RECT 6.845 2.19 6.86 2.345 ;
      RECT 6.855 3.457 6.86 3.745 ;
      RECT 6.845 3.52 6.855 3.745 ;
      RECT 6.765 2.175 6.845 2.325 ;
      RECT 6.84 3.527 6.845 3.74 ;
      RECT 6.835 3.535 6.84 3.73 ;
      RECT 6.755 2.161 6.765 2.309 ;
      RECT 6.74 2.157 6.755 2.307 ;
      RECT 6.73 2.152 6.74 2.303 ;
      RECT 6.705 2.145 6.73 2.295 ;
      RECT 6.7 2.14 6.705 2.29 ;
      RECT 6.69 2.14 6.7 2.288 ;
      RECT 6.68 2.138 6.69 2.286 ;
      RECT 6.65 2.13 6.68 2.28 ;
      RECT 6.635 2.122 6.65 2.273 ;
      RECT 6.615 2.117 6.635 2.266 ;
      RECT 6.61 2.113 6.615 2.261 ;
      RECT 6.58 2.106 6.61 2.255 ;
      RECT 6.555 2.097 6.58 2.245 ;
      RECT 6.525 2.09 6.555 2.237 ;
      RECT 6.5 2.08 6.525 2.228 ;
      RECT 6.485 2.072 6.5 2.222 ;
      RECT 6.46 2.067 6.485 2.217 ;
      RECT 6.45 2.063 6.46 2.212 ;
      RECT 6.43 2.058 6.45 2.207 ;
      RECT 6.395 2.053 6.43 2.2 ;
      RECT 6.335 2.048 6.395 2.193 ;
      RECT 6.322 2.044 6.335 2.191 ;
      RECT 6.236 2.039 6.322 2.188 ;
      RECT 6.15 2.029 6.236 2.184 ;
      RECT 6.109 2.022 6.15 2.181 ;
      RECT 6.023 2.015 6.109 2.178 ;
      RECT 5.937 2.005 6.023 2.174 ;
      RECT 5.851 1.995 5.937 2.169 ;
      RECT 5.765 1.985 5.851 2.165 ;
      RECT 5.755 1.97 5.765 2.163 ;
      RECT 5.745 1.955 5.755 2.163 ;
      RECT 5.68 1.95 5.745 2.162 ;
      RECT 5.515 1.947 5.56 2.155 ;
      RECT 6.76 2.852 6.765 3.043 ;
      RECT 6.755 2.847 6.76 3.05 ;
      RECT 6.741 2.845 6.755 3.056 ;
      RECT 6.655 2.845 6.741 3.058 ;
      RECT 6.651 2.845 6.655 3.061 ;
      RECT 6.565 2.845 6.651 3.079 ;
      RECT 6.555 2.85 6.565 3.098 ;
      RECT 6.545 2.905 6.555 3.102 ;
      RECT 6.52 2.92 6.545 3.109 ;
      RECT 6.48 2.94 6.52 3.122 ;
      RECT 6.475 2.952 6.48 3.132 ;
      RECT 6.46 2.958 6.475 3.137 ;
      RECT 6.455 2.963 6.46 3.141 ;
      RECT 6.435 2.97 6.455 3.146 ;
      RECT 6.365 2.995 6.435 3.163 ;
      RECT 6.325 3.023 6.365 3.183 ;
      RECT 6.32 3.033 6.325 3.191 ;
      RECT 6.3 3.04 6.32 3.193 ;
      RECT 6.295 3.047 6.3 3.196 ;
      RECT 6.265 3.055 6.295 3.199 ;
      RECT 6.26 3.06 6.265 3.203 ;
      RECT 6.186 3.064 6.26 3.211 ;
      RECT 6.1 3.073 6.186 3.227 ;
      RECT 6.096 3.078 6.1 3.236 ;
      RECT 6.01 3.083 6.096 3.246 ;
      RECT 5.97 3.091 6.01 3.258 ;
      RECT 5.92 3.097 5.97 3.265 ;
      RECT 5.835 3.106 5.92 3.28 ;
      RECT 5.76 3.117 5.835 3.298 ;
      RECT 5.725 3.124 5.76 3.308 ;
      RECT 5.65 3.132 5.725 3.313 ;
      RECT 5.595 3.141 5.65 3.313 ;
      RECT 5.57 3.146 5.595 3.311 ;
      RECT 5.56 3.149 5.57 3.309 ;
      RECT 5.525 3.151 5.56 3.307 ;
      RECT 5.495 3.153 5.525 3.303 ;
      RECT 5.45 3.152 5.495 3.299 ;
      RECT 5.43 3.147 5.45 3.296 ;
      RECT 5.38 3.132 5.43 3.293 ;
      RECT 5.37 3.117 5.38 3.288 ;
      RECT 5.32 3.102 5.37 3.278 ;
      RECT 5.27 3.077 5.32 3.258 ;
      RECT 5.26 3.062 5.27 3.24 ;
      RECT 5.255 3.06 5.26 3.234 ;
      RECT 5.235 3.055 5.255 3.229 ;
      RECT 5.23 3.047 5.235 3.223 ;
      RECT 5.215 3.041 5.23 3.216 ;
      RECT 5.21 3.036 5.215 3.208 ;
      RECT 5.19 3.031 5.21 3.2 ;
      RECT 5.175 3.024 5.19 3.193 ;
      RECT 5.16 3.018 5.175 3.184 ;
      RECT 5.155 3.012 5.16 3.177 ;
      RECT 5.11 2.987 5.155 3.163 ;
      RECT 5.095 2.957 5.11 3.145 ;
      RECT 5.08 2.94 5.095 3.136 ;
      RECT 5.055 2.92 5.08 3.124 ;
      RECT 5.015 2.89 5.055 3.104 ;
      RECT 5.005 2.86 5.015 3.089 ;
      RECT 4.99 2.85 5.005 3.082 ;
      RECT 4.935 2.815 4.99 3.061 ;
      RECT 4.92 2.778 4.935 3.04 ;
      RECT 4.91 2.765 4.92 3.032 ;
      RECT 4.86 2.735 4.91 3.014 ;
      RECT 4.845 2.665 4.86 2.995 ;
      RECT 4.8 2.665 4.845 2.978 ;
      RECT 4.775 2.665 4.8 2.96 ;
      RECT 4.765 2.665 4.775 2.953 ;
      RECT 4.686 2.665 4.765 2.946 ;
      RECT 4.6 2.665 4.686 2.938 ;
      RECT 4.585 2.697 4.6 2.933 ;
      RECT 4.51 2.707 4.585 2.929 ;
      RECT 4.49 2.717 4.51 2.924 ;
      RECT 4.465 2.717 4.49 2.921 ;
      RECT 4.455 2.707 4.465 2.92 ;
      RECT 4.445 2.68 4.455 2.919 ;
      RECT 4.405 2.675 4.445 2.917 ;
      RECT 4.36 2.675 4.405 2.913 ;
      RECT 4.335 2.675 4.36 2.908 ;
      RECT 4.285 2.675 4.335 2.895 ;
      RECT 4.245 2.68 4.255 2.88 ;
      RECT 4.255 2.675 4.285 2.885 ;
      RECT 6.24 2.455 6.5 2.715 ;
      RECT 6.235 2.477 6.5 2.673 ;
      RECT 5.475 2.305 5.695 2.67 ;
      RECT 5.457 2.392 5.695 2.669 ;
      RECT 5.44 2.397 5.695 2.666 ;
      RECT 5.44 2.397 5.715 2.665 ;
      RECT 5.41 2.407 5.715 2.663 ;
      RECT 5.405 2.422 5.715 2.659 ;
      RECT 5.405 2.422 5.72 2.658 ;
      RECT 5.4 2.48 5.72 2.656 ;
      RECT 5.4 2.48 5.73 2.653 ;
      RECT 5.395 2.545 5.73 2.648 ;
      RECT 5.475 2.305 5.735 2.565 ;
      RECT 4.22 2.135 4.48 2.395 ;
      RECT 4.22 2.178 4.566 2.369 ;
      RECT 4.22 2.178 4.61 2.368 ;
      RECT 4.22 2.178 4.63 2.366 ;
      RECT 4.22 2.178 4.73 2.365 ;
      RECT 4.22 2.178 4.75 2.363 ;
      RECT 4.22 2.178 4.76 2.358 ;
      RECT 4.63 2.145 4.82 2.355 ;
      RECT 4.63 2.147 4.825 2.353 ;
      RECT 4.62 2.152 4.83 2.345 ;
      RECT 4.566 2.176 4.83 2.345 ;
      RECT 4.61 2.17 4.62 2.367 ;
      RECT 4.62 2.15 4.825 2.353 ;
      RECT 3.575 3.21 3.78 3.44 ;
      RECT 3.515 3.16 3.57 3.42 ;
      RECT 3.575 3.16 3.775 3.44 ;
      RECT 4.545 3.475 4.55 3.502 ;
      RECT 4.535 3.385 4.545 3.507 ;
      RECT 4.53 3.307 4.535 3.513 ;
      RECT 4.52 3.297 4.53 3.52 ;
      RECT 4.515 3.287 4.52 3.526 ;
      RECT 4.505 3.282 4.515 3.528 ;
      RECT 4.49 3.274 4.505 3.536 ;
      RECT 4.475 3.265 4.49 3.548 ;
      RECT 4.465 3.257 4.475 3.558 ;
      RECT 4.43 3.175 4.465 3.576 ;
      RECT 4.395 3.175 4.43 3.595 ;
      RECT 4.38 3.175 4.395 3.603 ;
      RECT 4.325 3.175 4.38 3.603 ;
      RECT 4.291 3.175 4.325 3.594 ;
      RECT 4.205 3.175 4.291 3.57 ;
      RECT 4.195 3.235 4.205 3.552 ;
      RECT 4.155 3.237 4.195 3.543 ;
      RECT 4.15 3.239 4.155 3.533 ;
      RECT 4.13 3.241 4.15 3.528 ;
      RECT 4.12 3.244 4.13 3.523 ;
      RECT 4.11 3.245 4.12 3.518 ;
      RECT 4.086 3.246 4.11 3.51 ;
      RECT 4 3.251 4.086 3.488 ;
      RECT 3.945 3.25 4 3.461 ;
      RECT 3.93 3.243 3.945 3.448 ;
      RECT 3.895 3.238 3.93 3.444 ;
      RECT 3.84 3.23 3.895 3.443 ;
      RECT 3.78 3.217 3.84 3.441 ;
      RECT 3.57 3.16 3.575 3.428 ;
      RECT 3.645 2.53 3.83 2.74 ;
      RECT 3.635 2.535 3.845 2.733 ;
      RECT 3.675 2.44 3.935 2.7 ;
      RECT 3.63 2.597 3.935 2.623 ;
      RECT 2.975 2.39 2.98 3.19 ;
      RECT 2.92 2.44 2.95 3.19 ;
      RECT 2.91 2.44 2.915 2.75 ;
      RECT 2.895 2.44 2.9 2.745 ;
      RECT 2.44 2.485 2.455 2.7 ;
      RECT 2.37 2.485 2.455 2.695 ;
      RECT 3.635 2.065 3.705 2.275 ;
      RECT 3.705 2.072 3.715 2.27 ;
      RECT 3.601 2.065 3.635 2.282 ;
      RECT 3.515 2.065 3.601 2.306 ;
      RECT 3.505 2.07 3.515 2.325 ;
      RECT 3.5 2.082 3.505 2.328 ;
      RECT 3.485 2.097 3.5 2.332 ;
      RECT 3.48 2.115 3.485 2.336 ;
      RECT 3.44 2.125 3.48 2.345 ;
      RECT 3.425 2.132 3.44 2.357 ;
      RECT 3.41 2.137 3.425 2.362 ;
      RECT 3.395 2.14 3.41 2.367 ;
      RECT 3.385 2.142 3.395 2.371 ;
      RECT 3.35 2.149 3.385 2.379 ;
      RECT 3.315 2.157 3.35 2.393 ;
      RECT 3.305 2.163 3.315 2.402 ;
      RECT 3.3 2.165 3.305 2.404 ;
      RECT 3.28 2.168 3.3 2.41 ;
      RECT 3.25 2.175 3.28 2.421 ;
      RECT 3.24 2.181 3.25 2.428 ;
      RECT 3.215 2.184 3.24 2.435 ;
      RECT 3.205 2.188 3.215 2.443 ;
      RECT 3.2 2.189 3.205 2.465 ;
      RECT 3.195 2.19 3.2 2.48 ;
      RECT 3.19 2.191 3.195 2.495 ;
      RECT 3.185 2.192 3.19 2.51 ;
      RECT 3.18 2.193 3.185 2.54 ;
      RECT 3.17 2.195 3.18 2.573 ;
      RECT 3.155 2.199 3.17 2.62 ;
      RECT 3.145 2.202 3.155 2.665 ;
      RECT 3.14 2.205 3.145 2.693 ;
      RECT 3.13 2.207 3.14 2.72 ;
      RECT 3.125 2.21 3.13 2.755 ;
      RECT 3.095 2.215 3.125 2.813 ;
      RECT 3.09 2.22 3.095 2.898 ;
      RECT 3.085 2.222 3.09 2.933 ;
      RECT 3.08 2.224 3.085 3.015 ;
      RECT 3.075 2.226 3.08 3.103 ;
      RECT 3.065 2.228 3.075 3.185 ;
      RECT 3.05 2.242 3.065 3.19 ;
      RECT 3.015 2.287 3.05 3.19 ;
      RECT 3.005 2.327 3.015 3.19 ;
      RECT 2.99 2.355 3.005 3.19 ;
      RECT 2.985 2.372 2.99 3.19 ;
      RECT 2.98 2.38 2.985 3.19 ;
      RECT 2.97 2.395 2.975 3.19 ;
      RECT 2.965 2.402 2.97 3.19 ;
      RECT 2.955 2.422 2.965 3.19 ;
      RECT 2.95 2.435 2.955 3.19 ;
      RECT 2.915 2.44 2.92 2.775 ;
      RECT 2.9 2.83 2.92 3.19 ;
      RECT 2.9 2.44 2.91 2.748 ;
      RECT 2.895 2.87 2.9 3.19 ;
      RECT 2.845 2.44 2.895 2.743 ;
      RECT 2.89 2.907 2.895 3.19 ;
      RECT 2.88 2.93 2.89 3.19 ;
      RECT 2.875 2.975 2.88 3.19 ;
      RECT 2.865 2.985 2.875 3.183 ;
      RECT 2.791 2.44 2.845 2.737 ;
      RECT 2.705 2.44 2.791 2.73 ;
      RECT 2.656 2.487 2.705 2.723 ;
      RECT 2.57 2.495 2.656 2.716 ;
      RECT 2.555 2.492 2.57 2.711 ;
      RECT 2.541 2.485 2.555 2.71 ;
      RECT 2.455 2.485 2.541 2.705 ;
      RECT 2.36 2.49 2.37 2.69 ;
      RECT 1.95 1.92 1.965 2.32 ;
      RECT 2.145 1.92 2.15 2.18 ;
      RECT 1.89 1.92 1.935 2.18 ;
      RECT 2.345 3.225 2.35 3.43 ;
      RECT 2.34 3.215 2.345 3.435 ;
      RECT 2.335 3.202 2.34 3.44 ;
      RECT 2.33 3.182 2.335 3.44 ;
      RECT 2.305 3.135 2.33 3.44 ;
      RECT 2.27 3.05 2.305 3.44 ;
      RECT 2.265 2.987 2.27 3.44 ;
      RECT 2.26 2.972 2.265 3.44 ;
      RECT 2.245 2.932 2.26 3.44 ;
      RECT 2.24 2.907 2.245 3.44 ;
      RECT 2.23 2.89 2.24 3.44 ;
      RECT 2.195 2.812 2.23 3.44 ;
      RECT 2.19 2.755 2.195 3.44 ;
      RECT 2.185 2.742 2.19 3.44 ;
      RECT 2.175 2.72 2.185 3.44 ;
      RECT 2.165 2.685 2.175 3.44 ;
      RECT 2.155 2.655 2.165 3.44 ;
      RECT 2.145 2.57 2.155 3.083 ;
      RECT 2.152 3.215 2.155 3.44 ;
      RECT 2.15 3.225 2.152 3.44 ;
      RECT 2.14 3.235 2.15 3.435 ;
      RECT 2.135 1.92 2.145 2.315 ;
      RECT 2.14 2.447 2.145 3.058 ;
      RECT 2.135 2.345 2.14 3.041 ;
      RECT 2.125 1.92 2.135 3.017 ;
      RECT 2.12 1.92 2.125 2.988 ;
      RECT 2.115 1.92 2.12 2.978 ;
      RECT 2.095 1.92 2.115 2.94 ;
      RECT 2.09 1.92 2.095 2.898 ;
      RECT 2.085 1.92 2.09 2.878 ;
      RECT 2.055 1.92 2.085 2.828 ;
      RECT 2.045 1.92 2.055 2.775 ;
      RECT 2.04 1.92 2.045 2.748 ;
      RECT 2.035 1.92 2.04 2.733 ;
      RECT 2.025 1.92 2.035 2.71 ;
      RECT 2.015 1.92 2.025 2.685 ;
      RECT 2.01 1.92 2.015 2.625 ;
      RECT 2 1.92 2.01 2.563 ;
      RECT 1.995 1.92 2 2.483 ;
      RECT 1.99 1.92 1.995 2.448 ;
      RECT 1.985 1.92 1.99 2.423 ;
      RECT 1.98 1.92 1.985 2.408 ;
      RECT 1.975 1.92 1.98 2.378 ;
      RECT 1.97 1.92 1.975 2.355 ;
      RECT 1.965 1.92 1.97 2.328 ;
      RECT 1.935 1.92 1.95 2.315 ;
      RECT 1.09 3.455 1.275 3.665 ;
      RECT 1.08 3.46 1.29 3.658 ;
      RECT 1.08 3.46 1.31 3.63 ;
      RECT 1.08 3.46 1.325 3.609 ;
      RECT 1.08 3.46 1.34 3.607 ;
      RECT 1.08 3.46 1.35 3.606 ;
      RECT 1.08 3.46 1.38 3.603 ;
      RECT 1.73 3.305 1.99 3.565 ;
      RECT 1.69 3.352 1.99 3.548 ;
      RECT 1.681 3.36 1.69 3.551 ;
      RECT 1.275 3.453 1.99 3.548 ;
      RECT 1.595 3.378 1.681 3.558 ;
      RECT 1.29 3.45 1.99 3.548 ;
      RECT 1.536 3.4 1.595 3.57 ;
      RECT 1.31 3.446 1.99 3.548 ;
      RECT 1.45 3.412 1.536 3.581 ;
      RECT 1.325 3.442 1.99 3.548 ;
      RECT 1.395 3.425 1.45 3.593 ;
      RECT 1.34 3.44 1.99 3.548 ;
      RECT 1.38 3.431 1.395 3.599 ;
      RECT 1.35 3.436 1.99 3.548 ;
      RECT 1.495 2.96 1.755 3.22 ;
      RECT 1.495 2.98 1.865 3.19 ;
      RECT 1.495 2.985 1.875 3.185 ;
      RECT 1.686 2.399 1.765 2.63 ;
      RECT 1.6 2.402 1.815 2.625 ;
      RECT 1.595 2.402 1.815 2.62 ;
      RECT 1.595 2.407 1.825 2.618 ;
      RECT 1.57 2.407 1.825 2.615 ;
      RECT 1.57 2.415 1.835 2.613 ;
      RECT 1.45 2.35 1.71 2.61 ;
      RECT 1.45 2.397 1.76 2.61 ;
      RECT 0.705 2.97 0.71 3.23 ;
      RECT 0.535 2.74 0.54 3.23 ;
      RECT 0.42 2.98 0.425 3.205 ;
      RECT 1.13 2.075 1.135 2.285 ;
      RECT 1.135 2.08 1.15 2.28 ;
      RECT 1.07 2.075 1.13 2.293 ;
      RECT 1.055 2.075 1.07 2.303 ;
      RECT 1.005 2.075 1.055 2.32 ;
      RECT 0.985 2.075 1.005 2.343 ;
      RECT 0.97 2.075 0.985 2.355 ;
      RECT 0.95 2.075 0.97 2.365 ;
      RECT 0.94 2.08 0.95 2.374 ;
      RECT 0.935 2.09 0.94 2.379 ;
      RECT 0.93 2.102 0.935 2.383 ;
      RECT 0.92 2.125 0.93 2.388 ;
      RECT 0.915 2.14 0.92 2.392 ;
      RECT 0.91 2.157 0.915 2.395 ;
      RECT 0.905 2.165 0.91 2.398 ;
      RECT 0.895 2.17 0.905 2.402 ;
      RECT 0.89 2.177 0.895 2.407 ;
      RECT 0.88 2.182 0.89 2.411 ;
      RECT 0.855 2.194 0.88 2.422 ;
      RECT 0.835 2.211 0.855 2.438 ;
      RECT 0.81 2.228 0.835 2.46 ;
      RECT 0.775 2.251 0.81 2.518 ;
      RECT 0.755 2.273 0.775 2.58 ;
      RECT 0.75 2.283 0.755 2.615 ;
      RECT 0.74 2.29 0.75 2.653 ;
      RECT 0.735 2.297 0.74 2.673 ;
      RECT 0.73 2.308 0.735 2.71 ;
      RECT 0.725 2.316 0.73 2.775 ;
      RECT 0.715 2.327 0.725 2.828 ;
      RECT 0.71 2.345 0.715 2.898 ;
      RECT 0.705 2.355 0.71 2.935 ;
      RECT 0.7 2.365 0.705 3.23 ;
      RECT 0.695 2.377 0.7 3.23 ;
      RECT 0.69 2.387 0.695 3.23 ;
      RECT 0.68 2.397 0.69 3.23 ;
      RECT 0.67 2.42 0.68 3.23 ;
      RECT 0.655 2.455 0.67 3.23 ;
      RECT 0.615 2.517 0.655 3.23 ;
      RECT 0.61 2.57 0.615 3.23 ;
      RECT 0.585 2.605 0.61 3.23 ;
      RECT 0.57 2.65 0.585 3.23 ;
      RECT 0.565 2.672 0.57 3.23 ;
      RECT 0.555 2.685 0.565 3.23 ;
      RECT 0.545 2.71 0.555 3.23 ;
      RECT 0.54 2.732 0.545 3.23 ;
      RECT 0.515 2.77 0.535 3.23 ;
      RECT 0.475 2.827 0.515 3.23 ;
      RECT 0.47 2.877 0.475 3.23 ;
      RECT 0.465 2.895 0.47 3.23 ;
      RECT 0.46 2.907 0.465 3.23 ;
      RECT 0.45 2.925 0.46 3.23 ;
      RECT 0.44 2.945 0.45 3.205 ;
      RECT 0.435 2.962 0.44 3.205 ;
      RECT 0.425 2.975 0.435 3.205 ;
      RECT 0.395 2.985 0.42 3.205 ;
      RECT 0.385 2.992 0.395 3.205 ;
      RECT 0.37 3.002 0.385 3.2 ;
      RECT -0.82 6.655 -0.53 6.885 ;
      RECT -0.99 6.685 -0.53 6.855 ;
      RECT -1.25 7.765 -0.96 7.995 ;
      RECT -1.19 7.025 -1.02 7.995 ;
      RECT -1.28 7.025 -0.93 7.315 ;
      RECT -1.655 6.285 -1.305 6.575 ;
      RECT -1.795 6.315 -1.305 6.485 ;
      RECT -2.62 5.915 -2.33 6.145 ;
      RECT -2.62 5.945 -2.16 6.115 ;
      RECT 73.26 2.85 73.63 3.22 ;
      RECT 57.475 2.85 57.845 3.22 ;
      RECT 41.69 2.85 42.06 3.22 ;
      RECT 25.915 2.85 26.285 3.22 ;
      RECT 10.135 2.85 10.505 3.22 ;
    LAYER mcon ;
      RECT 78.435 0.915 78.605 1.085 ;
      RECT 78.435 2.395 78.605 2.565 ;
      RECT 78.435 6.315 78.605 6.485 ;
      RECT 78.435 7.795 78.605 7.965 ;
      RECT 78.085 0.105 78.255 0.275 ;
      RECT 78.085 4.165 78.255 4.335 ;
      RECT 78.085 4.545 78.255 4.715 ;
      RECT 78.085 8.605 78.255 8.775 ;
      RECT 78.065 2.765 78.235 2.935 ;
      RECT 78.065 5.945 78.235 6.115 ;
      RECT 77.445 0.915 77.615 1.085 ;
      RECT 77.445 2.395 77.615 2.565 ;
      RECT 77.445 6.315 77.615 6.485 ;
      RECT 77.445 7.795 77.615 7.965 ;
      RECT 77.095 0.105 77.265 0.275 ;
      RECT 77.095 4.165 77.265 4.335 ;
      RECT 77.095 4.545 77.265 4.715 ;
      RECT 77.095 8.605 77.265 8.775 ;
      RECT 77.075 2.765 77.245 2.935 ;
      RECT 77.075 5.945 77.245 6.115 ;
      RECT 76.39 0.105 76.56 0.275 ;
      RECT 76.39 4.165 76.56 4.335 ;
      RECT 76.39 4.545 76.56 4.715 ;
      RECT 76.39 8.605 76.56 8.775 ;
      RECT 76.08 2.025 76.25 2.195 ;
      RECT 76.08 6.685 76.25 6.855 ;
      RECT 75.71 0.105 75.88 0.275 ;
      RECT 75.71 8.605 75.88 8.775 ;
      RECT 75.65 0.915 75.82 1.085 ;
      RECT 75.65 1.655 75.82 1.825 ;
      RECT 75.65 7.055 75.82 7.225 ;
      RECT 75.65 7.795 75.82 7.965 ;
      RECT 75.275 2.395 75.445 2.565 ;
      RECT 75.275 6.315 75.445 6.485 ;
      RECT 75.03 0.105 75.2 0.275 ;
      RECT 75.03 8.605 75.2 8.775 ;
      RECT 74.35 0.105 74.52 0.275 ;
      RECT 74.35 8.605 74.52 8.775 ;
      RECT 74.28 2.765 74.45 2.935 ;
      RECT 74.28 5.945 74.45 6.115 ;
      RECT 72.725 1.415 72.895 1.585 ;
      RECT 72.725 4.135 72.895 4.305 ;
      RECT 72.355 2.875 72.525 3.045 ;
      RECT 72.265 1.415 72.435 1.585 ;
      RECT 72.265 4.135 72.435 4.305 ;
      RECT 72.035 2.045 72.205 2.215 ;
      RECT 71.89 2.485 72.06 2.655 ;
      RECT 71.805 1.415 71.975 1.585 ;
      RECT 71.805 4.135 71.975 4.305 ;
      RECT 71.61 4.545 71.78 4.715 ;
      RECT 71.61 8.605 71.78 8.775 ;
      RECT 71.345 1.415 71.515 1.585 ;
      RECT 71.345 4.135 71.515 4.305 ;
      RECT 71.3 6.685 71.47 6.855 ;
      RECT 71.28 2.525 71.45 2.695 ;
      RECT 70.935 2.16 71.105 2.33 ;
      RECT 70.93 8.605 71.1 8.775 ;
      RECT 70.925 3.52 71.095 3.69 ;
      RECT 70.885 1.415 71.055 1.585 ;
      RECT 70.885 4.135 71.055 4.305 ;
      RECT 70.87 7.055 71.04 7.225 ;
      RECT 70.87 7.795 71.04 7.965 ;
      RECT 70.51 2.76 70.68 2.93 ;
      RECT 70.495 6.315 70.665 6.485 ;
      RECT 70.425 1.415 70.595 1.585 ;
      RECT 70.425 4.135 70.595 4.305 ;
      RECT 70.25 8.605 70.42 8.775 ;
      RECT 70.16 2.235 70.33 2.405 ;
      RECT 69.98 3.55 70.15 3.72 ;
      RECT 69.965 1.415 70.135 1.585 ;
      RECT 69.965 4.135 70.135 4.305 ;
      RECT 69.7 2.865 69.87 3.035 ;
      RECT 69.57 8.605 69.74 8.775 ;
      RECT 69.505 1.415 69.675 1.585 ;
      RECT 69.505 4.135 69.675 4.305 ;
      RECT 69.5 5.945 69.67 6.115 ;
      RECT 69.38 2.49 69.55 2.66 ;
      RECT 69.045 1.415 69.215 1.585 ;
      RECT 69.045 4.135 69.215 4.305 ;
      RECT 68.69 1.97 68.86 2.14 ;
      RECT 68.615 2.44 68.785 2.61 ;
      RECT 68.585 1.415 68.755 1.585 ;
      RECT 68.585 4.135 68.755 4.305 ;
      RECT 68.125 1.415 68.295 1.585 ;
      RECT 68.125 4.135 68.295 4.305 ;
      RECT 67.765 2.165 67.935 2.335 ;
      RECT 67.665 1.415 67.835 1.585 ;
      RECT 67.665 4.135 67.835 4.305 ;
      RECT 67.425 3.36 67.595 3.53 ;
      RECT 67.39 2.695 67.56 2.865 ;
      RECT 67.205 1.415 67.375 1.585 ;
      RECT 67.205 4.135 67.375 4.305 ;
      RECT 66.78 2.55 66.95 2.72 ;
      RECT 66.745 1.415 66.915 1.585 ;
      RECT 66.745 4.135 66.915 4.305 ;
      RECT 66.71 3.25 66.88 3.42 ;
      RECT 66.65 2.085 66.82 2.255 ;
      RECT 66.285 1.415 66.455 1.585 ;
      RECT 66.285 4.135 66.455 4.305 ;
      RECT 66.01 3 66.18 3.17 ;
      RECT 65.825 1.415 65.995 1.585 ;
      RECT 65.825 4.135 65.995 4.305 ;
      RECT 65.505 2.505 65.675 2.675 ;
      RECT 65.365 1.415 65.535 1.585 ;
      RECT 65.365 4.135 65.535 4.305 ;
      RECT 65.285 3.25 65.455 3.42 ;
      RECT 65.08 2.13 65.25 2.3 ;
      RECT 64.905 1.415 65.075 1.585 ;
      RECT 64.905 4.135 65.075 4.305 ;
      RECT 64.81 3 64.98 3.17 ;
      RECT 64.77 2.43 64.94 2.6 ;
      RECT 64.445 1.415 64.615 1.585 ;
      RECT 64.445 4.135 64.615 4.305 ;
      RECT 64.225 3.475 64.395 3.645 ;
      RECT 64.085 2.095 64.255 2.265 ;
      RECT 63.985 1.415 64.155 1.585 ;
      RECT 63.985 4.135 64.155 4.305 ;
      RECT 63.525 1.415 63.695 1.585 ;
      RECT 63.525 4.135 63.695 4.305 ;
      RECT 63.515 3.015 63.685 3.185 ;
      RECT 62.65 0.915 62.82 1.085 ;
      RECT 62.65 2.395 62.82 2.565 ;
      RECT 62.65 6.315 62.82 6.485 ;
      RECT 62.65 7.795 62.82 7.965 ;
      RECT 62.3 0.105 62.47 0.275 ;
      RECT 62.3 4.165 62.47 4.335 ;
      RECT 62.3 4.545 62.47 4.715 ;
      RECT 62.3 8.605 62.47 8.775 ;
      RECT 62.28 2.765 62.45 2.935 ;
      RECT 62.28 5.945 62.45 6.115 ;
      RECT 61.66 0.915 61.83 1.085 ;
      RECT 61.66 2.395 61.83 2.565 ;
      RECT 61.66 6.315 61.83 6.485 ;
      RECT 61.66 7.795 61.83 7.965 ;
      RECT 61.31 0.105 61.48 0.275 ;
      RECT 61.31 4.165 61.48 4.335 ;
      RECT 61.31 4.545 61.48 4.715 ;
      RECT 61.31 8.605 61.48 8.775 ;
      RECT 61.29 2.765 61.46 2.935 ;
      RECT 61.29 5.945 61.46 6.115 ;
      RECT 60.605 0.105 60.775 0.275 ;
      RECT 60.605 4.165 60.775 4.335 ;
      RECT 60.605 4.545 60.775 4.715 ;
      RECT 60.605 8.605 60.775 8.775 ;
      RECT 60.295 2.025 60.465 2.195 ;
      RECT 60.295 6.685 60.465 6.855 ;
      RECT 59.925 0.105 60.095 0.275 ;
      RECT 59.925 8.605 60.095 8.775 ;
      RECT 59.865 0.915 60.035 1.085 ;
      RECT 59.865 1.655 60.035 1.825 ;
      RECT 59.865 7.055 60.035 7.225 ;
      RECT 59.865 7.795 60.035 7.965 ;
      RECT 59.49 2.395 59.66 2.565 ;
      RECT 59.49 6.315 59.66 6.485 ;
      RECT 59.245 0.105 59.415 0.275 ;
      RECT 59.245 8.605 59.415 8.775 ;
      RECT 58.565 0.105 58.735 0.275 ;
      RECT 58.565 8.605 58.735 8.775 ;
      RECT 58.495 2.765 58.665 2.935 ;
      RECT 58.495 5.945 58.665 6.115 ;
      RECT 56.94 1.415 57.11 1.585 ;
      RECT 56.94 4.135 57.11 4.305 ;
      RECT 56.57 2.875 56.74 3.045 ;
      RECT 56.48 1.415 56.65 1.585 ;
      RECT 56.48 4.135 56.65 4.305 ;
      RECT 56.25 2.045 56.42 2.215 ;
      RECT 56.105 2.485 56.275 2.655 ;
      RECT 56.02 1.415 56.19 1.585 ;
      RECT 56.02 4.135 56.19 4.305 ;
      RECT 55.825 4.545 55.995 4.715 ;
      RECT 55.825 8.605 55.995 8.775 ;
      RECT 55.56 1.415 55.73 1.585 ;
      RECT 55.56 4.135 55.73 4.305 ;
      RECT 55.515 6.685 55.685 6.855 ;
      RECT 55.495 2.525 55.665 2.695 ;
      RECT 55.15 2.16 55.32 2.33 ;
      RECT 55.145 8.605 55.315 8.775 ;
      RECT 55.14 3.52 55.31 3.69 ;
      RECT 55.1 1.415 55.27 1.585 ;
      RECT 55.1 4.135 55.27 4.305 ;
      RECT 55.085 7.055 55.255 7.225 ;
      RECT 55.085 7.795 55.255 7.965 ;
      RECT 54.725 2.76 54.895 2.93 ;
      RECT 54.71 6.315 54.88 6.485 ;
      RECT 54.64 1.415 54.81 1.585 ;
      RECT 54.64 4.135 54.81 4.305 ;
      RECT 54.465 8.605 54.635 8.775 ;
      RECT 54.375 2.235 54.545 2.405 ;
      RECT 54.195 3.55 54.365 3.72 ;
      RECT 54.18 1.415 54.35 1.585 ;
      RECT 54.18 4.135 54.35 4.305 ;
      RECT 53.915 2.865 54.085 3.035 ;
      RECT 53.785 8.605 53.955 8.775 ;
      RECT 53.72 1.415 53.89 1.585 ;
      RECT 53.72 4.135 53.89 4.305 ;
      RECT 53.715 5.945 53.885 6.115 ;
      RECT 53.595 2.49 53.765 2.66 ;
      RECT 53.26 1.415 53.43 1.585 ;
      RECT 53.26 4.135 53.43 4.305 ;
      RECT 52.905 1.97 53.075 2.14 ;
      RECT 52.83 2.44 53 2.61 ;
      RECT 52.8 1.415 52.97 1.585 ;
      RECT 52.8 4.135 52.97 4.305 ;
      RECT 52.34 1.415 52.51 1.585 ;
      RECT 52.34 4.135 52.51 4.305 ;
      RECT 51.98 2.165 52.15 2.335 ;
      RECT 51.88 1.415 52.05 1.585 ;
      RECT 51.88 4.135 52.05 4.305 ;
      RECT 51.64 3.36 51.81 3.53 ;
      RECT 51.605 2.695 51.775 2.865 ;
      RECT 51.42 1.415 51.59 1.585 ;
      RECT 51.42 4.135 51.59 4.305 ;
      RECT 50.995 2.55 51.165 2.72 ;
      RECT 50.96 1.415 51.13 1.585 ;
      RECT 50.96 4.135 51.13 4.305 ;
      RECT 50.925 3.25 51.095 3.42 ;
      RECT 50.865 2.085 51.035 2.255 ;
      RECT 50.5 1.415 50.67 1.585 ;
      RECT 50.5 4.135 50.67 4.305 ;
      RECT 50.225 3 50.395 3.17 ;
      RECT 50.04 1.415 50.21 1.585 ;
      RECT 50.04 4.135 50.21 4.305 ;
      RECT 49.72 2.505 49.89 2.675 ;
      RECT 49.58 1.415 49.75 1.585 ;
      RECT 49.58 4.135 49.75 4.305 ;
      RECT 49.5 3.25 49.67 3.42 ;
      RECT 49.295 2.13 49.465 2.3 ;
      RECT 49.12 1.415 49.29 1.585 ;
      RECT 49.12 4.135 49.29 4.305 ;
      RECT 49.025 3 49.195 3.17 ;
      RECT 48.985 2.43 49.155 2.6 ;
      RECT 48.66 1.415 48.83 1.585 ;
      RECT 48.66 4.135 48.83 4.305 ;
      RECT 48.44 3.475 48.61 3.645 ;
      RECT 48.3 2.095 48.47 2.265 ;
      RECT 48.2 1.415 48.37 1.585 ;
      RECT 48.2 4.135 48.37 4.305 ;
      RECT 47.74 1.415 47.91 1.585 ;
      RECT 47.74 4.135 47.91 4.305 ;
      RECT 47.73 3.015 47.9 3.185 ;
      RECT 46.865 0.915 47.035 1.085 ;
      RECT 46.865 2.395 47.035 2.565 ;
      RECT 46.865 6.315 47.035 6.485 ;
      RECT 46.865 7.795 47.035 7.965 ;
      RECT 46.515 0.105 46.685 0.275 ;
      RECT 46.515 4.165 46.685 4.335 ;
      RECT 46.515 4.545 46.685 4.715 ;
      RECT 46.515 8.605 46.685 8.775 ;
      RECT 46.495 2.765 46.665 2.935 ;
      RECT 46.495 5.945 46.665 6.115 ;
      RECT 45.875 0.915 46.045 1.085 ;
      RECT 45.875 2.395 46.045 2.565 ;
      RECT 45.875 6.315 46.045 6.485 ;
      RECT 45.875 7.795 46.045 7.965 ;
      RECT 45.525 0.105 45.695 0.275 ;
      RECT 45.525 4.165 45.695 4.335 ;
      RECT 45.525 4.545 45.695 4.715 ;
      RECT 45.525 8.605 45.695 8.775 ;
      RECT 45.505 2.765 45.675 2.935 ;
      RECT 45.505 5.945 45.675 6.115 ;
      RECT 44.82 0.105 44.99 0.275 ;
      RECT 44.82 4.165 44.99 4.335 ;
      RECT 44.82 4.545 44.99 4.715 ;
      RECT 44.82 8.605 44.99 8.775 ;
      RECT 44.51 2.025 44.68 2.195 ;
      RECT 44.51 6.685 44.68 6.855 ;
      RECT 44.14 0.105 44.31 0.275 ;
      RECT 44.14 8.605 44.31 8.775 ;
      RECT 44.08 0.915 44.25 1.085 ;
      RECT 44.08 1.655 44.25 1.825 ;
      RECT 44.08 7.055 44.25 7.225 ;
      RECT 44.08 7.795 44.25 7.965 ;
      RECT 43.705 2.395 43.875 2.565 ;
      RECT 43.705 6.315 43.875 6.485 ;
      RECT 43.46 0.105 43.63 0.275 ;
      RECT 43.46 8.605 43.63 8.775 ;
      RECT 42.78 0.105 42.95 0.275 ;
      RECT 42.78 8.605 42.95 8.775 ;
      RECT 42.71 2.765 42.88 2.935 ;
      RECT 42.71 5.945 42.88 6.115 ;
      RECT 41.155 1.415 41.325 1.585 ;
      RECT 41.155 4.135 41.325 4.305 ;
      RECT 40.785 2.875 40.955 3.045 ;
      RECT 40.695 1.415 40.865 1.585 ;
      RECT 40.695 4.135 40.865 4.305 ;
      RECT 40.465 2.045 40.635 2.215 ;
      RECT 40.32 2.485 40.49 2.655 ;
      RECT 40.235 1.415 40.405 1.585 ;
      RECT 40.235 4.135 40.405 4.305 ;
      RECT 40.04 4.545 40.21 4.715 ;
      RECT 40.04 8.605 40.21 8.775 ;
      RECT 39.775 1.415 39.945 1.585 ;
      RECT 39.775 4.135 39.945 4.305 ;
      RECT 39.73 6.685 39.9 6.855 ;
      RECT 39.71 2.525 39.88 2.695 ;
      RECT 39.365 2.16 39.535 2.33 ;
      RECT 39.36 8.605 39.53 8.775 ;
      RECT 39.355 3.52 39.525 3.69 ;
      RECT 39.315 1.415 39.485 1.585 ;
      RECT 39.315 4.135 39.485 4.305 ;
      RECT 39.3 7.055 39.47 7.225 ;
      RECT 39.3 7.795 39.47 7.965 ;
      RECT 38.94 2.76 39.11 2.93 ;
      RECT 38.925 6.315 39.095 6.485 ;
      RECT 38.855 1.415 39.025 1.585 ;
      RECT 38.855 4.135 39.025 4.305 ;
      RECT 38.68 8.605 38.85 8.775 ;
      RECT 38.59 2.235 38.76 2.405 ;
      RECT 38.41 3.55 38.58 3.72 ;
      RECT 38.395 1.415 38.565 1.585 ;
      RECT 38.395 4.135 38.565 4.305 ;
      RECT 38.13 2.865 38.3 3.035 ;
      RECT 38 8.605 38.17 8.775 ;
      RECT 37.935 1.415 38.105 1.585 ;
      RECT 37.935 4.135 38.105 4.305 ;
      RECT 37.93 5.945 38.1 6.115 ;
      RECT 37.81 2.49 37.98 2.66 ;
      RECT 37.475 1.415 37.645 1.585 ;
      RECT 37.475 4.135 37.645 4.305 ;
      RECT 37.12 1.97 37.29 2.14 ;
      RECT 37.045 2.44 37.215 2.61 ;
      RECT 37.015 1.415 37.185 1.585 ;
      RECT 37.015 4.135 37.185 4.305 ;
      RECT 36.555 1.415 36.725 1.585 ;
      RECT 36.555 4.135 36.725 4.305 ;
      RECT 36.195 2.165 36.365 2.335 ;
      RECT 36.095 1.415 36.265 1.585 ;
      RECT 36.095 4.135 36.265 4.305 ;
      RECT 35.855 3.36 36.025 3.53 ;
      RECT 35.82 2.695 35.99 2.865 ;
      RECT 35.635 1.415 35.805 1.585 ;
      RECT 35.635 4.135 35.805 4.305 ;
      RECT 35.21 2.55 35.38 2.72 ;
      RECT 35.175 1.415 35.345 1.585 ;
      RECT 35.175 4.135 35.345 4.305 ;
      RECT 35.14 3.25 35.31 3.42 ;
      RECT 35.08 2.085 35.25 2.255 ;
      RECT 34.715 1.415 34.885 1.585 ;
      RECT 34.715 4.135 34.885 4.305 ;
      RECT 34.44 3 34.61 3.17 ;
      RECT 34.255 1.415 34.425 1.585 ;
      RECT 34.255 4.135 34.425 4.305 ;
      RECT 33.935 2.505 34.105 2.675 ;
      RECT 33.795 1.415 33.965 1.585 ;
      RECT 33.795 4.135 33.965 4.305 ;
      RECT 33.715 3.25 33.885 3.42 ;
      RECT 33.51 2.13 33.68 2.3 ;
      RECT 33.335 1.415 33.505 1.585 ;
      RECT 33.335 4.135 33.505 4.305 ;
      RECT 33.24 3 33.41 3.17 ;
      RECT 33.2 2.43 33.37 2.6 ;
      RECT 32.875 1.415 33.045 1.585 ;
      RECT 32.875 4.135 33.045 4.305 ;
      RECT 32.655 3.475 32.825 3.645 ;
      RECT 32.515 2.095 32.685 2.265 ;
      RECT 32.415 1.415 32.585 1.585 ;
      RECT 32.415 4.135 32.585 4.305 ;
      RECT 31.955 1.415 32.125 1.585 ;
      RECT 31.955 4.135 32.125 4.305 ;
      RECT 31.945 3.015 32.115 3.185 ;
      RECT 31.09 0.915 31.26 1.085 ;
      RECT 31.09 2.395 31.26 2.565 ;
      RECT 31.09 6.315 31.26 6.485 ;
      RECT 31.09 7.795 31.26 7.965 ;
      RECT 30.74 0.105 30.91 0.275 ;
      RECT 30.74 4.165 30.91 4.335 ;
      RECT 30.74 4.545 30.91 4.715 ;
      RECT 30.74 8.605 30.91 8.775 ;
      RECT 30.72 2.765 30.89 2.935 ;
      RECT 30.72 5.945 30.89 6.115 ;
      RECT 30.1 0.915 30.27 1.085 ;
      RECT 30.1 2.395 30.27 2.565 ;
      RECT 30.1 6.315 30.27 6.485 ;
      RECT 30.1 7.795 30.27 7.965 ;
      RECT 29.75 0.105 29.92 0.275 ;
      RECT 29.75 4.165 29.92 4.335 ;
      RECT 29.75 4.545 29.92 4.715 ;
      RECT 29.75 8.605 29.92 8.775 ;
      RECT 29.73 2.765 29.9 2.935 ;
      RECT 29.73 5.945 29.9 6.115 ;
      RECT 29.045 0.105 29.215 0.275 ;
      RECT 29.045 4.165 29.215 4.335 ;
      RECT 29.045 4.545 29.215 4.715 ;
      RECT 29.045 8.605 29.215 8.775 ;
      RECT 28.735 2.025 28.905 2.195 ;
      RECT 28.735 6.685 28.905 6.855 ;
      RECT 28.365 0.105 28.535 0.275 ;
      RECT 28.365 8.605 28.535 8.775 ;
      RECT 28.305 0.915 28.475 1.085 ;
      RECT 28.305 1.655 28.475 1.825 ;
      RECT 28.305 7.055 28.475 7.225 ;
      RECT 28.305 7.795 28.475 7.965 ;
      RECT 27.93 2.395 28.1 2.565 ;
      RECT 27.93 6.315 28.1 6.485 ;
      RECT 27.685 0.105 27.855 0.275 ;
      RECT 27.685 8.605 27.855 8.775 ;
      RECT 27.005 0.105 27.175 0.275 ;
      RECT 27.005 8.605 27.175 8.775 ;
      RECT 26.935 2.765 27.105 2.935 ;
      RECT 26.935 5.945 27.105 6.115 ;
      RECT 25.38 1.415 25.55 1.585 ;
      RECT 25.38 4.135 25.55 4.305 ;
      RECT 25.01 2.875 25.18 3.045 ;
      RECT 24.92 1.415 25.09 1.585 ;
      RECT 24.92 4.135 25.09 4.305 ;
      RECT 24.69 2.045 24.86 2.215 ;
      RECT 24.545 2.485 24.715 2.655 ;
      RECT 24.46 1.415 24.63 1.585 ;
      RECT 24.46 4.135 24.63 4.305 ;
      RECT 24.265 4.545 24.435 4.715 ;
      RECT 24.265 8.605 24.435 8.775 ;
      RECT 24 1.415 24.17 1.585 ;
      RECT 24 4.135 24.17 4.305 ;
      RECT 23.955 6.685 24.125 6.855 ;
      RECT 23.935 2.525 24.105 2.695 ;
      RECT 23.59 2.16 23.76 2.33 ;
      RECT 23.585 8.605 23.755 8.775 ;
      RECT 23.58 3.52 23.75 3.69 ;
      RECT 23.54 1.415 23.71 1.585 ;
      RECT 23.54 4.135 23.71 4.305 ;
      RECT 23.525 7.055 23.695 7.225 ;
      RECT 23.525 7.795 23.695 7.965 ;
      RECT 23.165 2.76 23.335 2.93 ;
      RECT 23.15 6.315 23.32 6.485 ;
      RECT 23.08 1.415 23.25 1.585 ;
      RECT 23.08 4.135 23.25 4.305 ;
      RECT 22.905 8.605 23.075 8.775 ;
      RECT 22.815 2.235 22.985 2.405 ;
      RECT 22.635 3.55 22.805 3.72 ;
      RECT 22.62 1.415 22.79 1.585 ;
      RECT 22.62 4.135 22.79 4.305 ;
      RECT 22.355 2.865 22.525 3.035 ;
      RECT 22.225 8.605 22.395 8.775 ;
      RECT 22.16 1.415 22.33 1.585 ;
      RECT 22.16 4.135 22.33 4.305 ;
      RECT 22.155 5.945 22.325 6.115 ;
      RECT 22.035 2.49 22.205 2.66 ;
      RECT 21.7 1.415 21.87 1.585 ;
      RECT 21.7 4.135 21.87 4.305 ;
      RECT 21.345 1.97 21.515 2.14 ;
      RECT 21.27 2.44 21.44 2.61 ;
      RECT 21.24 1.415 21.41 1.585 ;
      RECT 21.24 4.135 21.41 4.305 ;
      RECT 20.78 1.415 20.95 1.585 ;
      RECT 20.78 4.135 20.95 4.305 ;
      RECT 20.42 2.165 20.59 2.335 ;
      RECT 20.32 1.415 20.49 1.585 ;
      RECT 20.32 4.135 20.49 4.305 ;
      RECT 20.08 3.36 20.25 3.53 ;
      RECT 20.045 2.695 20.215 2.865 ;
      RECT 19.86 1.415 20.03 1.585 ;
      RECT 19.86 4.135 20.03 4.305 ;
      RECT 19.435 2.55 19.605 2.72 ;
      RECT 19.4 1.415 19.57 1.585 ;
      RECT 19.4 4.135 19.57 4.305 ;
      RECT 19.365 3.25 19.535 3.42 ;
      RECT 19.305 2.085 19.475 2.255 ;
      RECT 18.94 1.415 19.11 1.585 ;
      RECT 18.94 4.135 19.11 4.305 ;
      RECT 18.665 3 18.835 3.17 ;
      RECT 18.48 1.415 18.65 1.585 ;
      RECT 18.48 4.135 18.65 4.305 ;
      RECT 18.16 2.505 18.33 2.675 ;
      RECT 18.02 1.415 18.19 1.585 ;
      RECT 18.02 4.135 18.19 4.305 ;
      RECT 17.94 3.25 18.11 3.42 ;
      RECT 17.735 2.13 17.905 2.3 ;
      RECT 17.56 1.415 17.73 1.585 ;
      RECT 17.56 4.135 17.73 4.305 ;
      RECT 17.465 3 17.635 3.17 ;
      RECT 17.425 2.43 17.595 2.6 ;
      RECT 17.1 1.415 17.27 1.585 ;
      RECT 17.1 4.135 17.27 4.305 ;
      RECT 16.88 3.475 17.05 3.645 ;
      RECT 16.74 2.095 16.91 2.265 ;
      RECT 16.64 1.415 16.81 1.585 ;
      RECT 16.64 4.135 16.81 4.305 ;
      RECT 16.18 1.415 16.35 1.585 ;
      RECT 16.18 4.135 16.35 4.305 ;
      RECT 16.17 3.015 16.34 3.185 ;
      RECT 15.31 0.915 15.48 1.085 ;
      RECT 15.31 2.395 15.48 2.565 ;
      RECT 15.31 6.315 15.48 6.485 ;
      RECT 15.31 7.795 15.48 7.965 ;
      RECT 14.96 0.105 15.13 0.275 ;
      RECT 14.96 4.165 15.13 4.335 ;
      RECT 14.96 4.545 15.13 4.715 ;
      RECT 14.96 8.605 15.13 8.775 ;
      RECT 14.94 2.765 15.11 2.935 ;
      RECT 14.94 5.945 15.11 6.115 ;
      RECT 14.32 0.915 14.49 1.085 ;
      RECT 14.32 2.395 14.49 2.565 ;
      RECT 14.32 6.315 14.49 6.485 ;
      RECT 14.32 7.795 14.49 7.965 ;
      RECT 13.97 0.105 14.14 0.275 ;
      RECT 13.97 4.165 14.14 4.335 ;
      RECT 13.97 4.545 14.14 4.715 ;
      RECT 13.97 8.605 14.14 8.775 ;
      RECT 13.95 2.765 14.12 2.935 ;
      RECT 13.95 5.945 14.12 6.115 ;
      RECT 13.265 0.105 13.435 0.275 ;
      RECT 13.265 4.165 13.435 4.335 ;
      RECT 13.265 4.545 13.435 4.715 ;
      RECT 13.265 8.605 13.435 8.775 ;
      RECT 12.955 2.025 13.125 2.195 ;
      RECT 12.955 6.685 13.125 6.855 ;
      RECT 12.585 0.105 12.755 0.275 ;
      RECT 12.585 8.605 12.755 8.775 ;
      RECT 12.525 0.915 12.695 1.085 ;
      RECT 12.525 1.655 12.695 1.825 ;
      RECT 12.525 7.055 12.695 7.225 ;
      RECT 12.525 7.795 12.695 7.965 ;
      RECT 12.15 2.395 12.32 2.565 ;
      RECT 12.15 6.315 12.32 6.485 ;
      RECT 11.905 0.105 12.075 0.275 ;
      RECT 11.905 8.605 12.075 8.775 ;
      RECT 11.225 0.105 11.395 0.275 ;
      RECT 11.225 8.605 11.395 8.775 ;
      RECT 11.155 2.765 11.325 2.935 ;
      RECT 11.155 5.945 11.325 6.115 ;
      RECT 9.6 1.415 9.77 1.585 ;
      RECT 9.6 4.135 9.77 4.305 ;
      RECT 9.23 2.875 9.4 3.045 ;
      RECT 9.14 1.415 9.31 1.585 ;
      RECT 9.14 4.135 9.31 4.305 ;
      RECT 8.91 2.045 9.08 2.215 ;
      RECT 8.765 2.485 8.935 2.655 ;
      RECT 8.68 1.415 8.85 1.585 ;
      RECT 8.68 4.135 8.85 4.305 ;
      RECT 8.485 4.545 8.655 4.715 ;
      RECT 8.485 8.605 8.655 8.775 ;
      RECT 8.22 1.415 8.39 1.585 ;
      RECT 8.22 4.135 8.39 4.305 ;
      RECT 8.175 6.685 8.345 6.855 ;
      RECT 8.155 2.525 8.325 2.695 ;
      RECT 7.81 2.16 7.98 2.33 ;
      RECT 7.805 8.605 7.975 8.775 ;
      RECT 7.8 3.52 7.97 3.69 ;
      RECT 7.76 1.415 7.93 1.585 ;
      RECT 7.76 4.135 7.93 4.305 ;
      RECT 7.745 7.055 7.915 7.225 ;
      RECT 7.745 7.795 7.915 7.965 ;
      RECT 7.385 2.76 7.555 2.93 ;
      RECT 7.37 6.315 7.54 6.485 ;
      RECT 7.3 1.415 7.47 1.585 ;
      RECT 7.3 4.135 7.47 4.305 ;
      RECT 7.125 8.605 7.295 8.775 ;
      RECT 7.035 2.235 7.205 2.405 ;
      RECT 6.855 3.55 7.025 3.72 ;
      RECT 6.84 1.415 7.01 1.585 ;
      RECT 6.84 4.135 7.01 4.305 ;
      RECT 6.575 2.865 6.745 3.035 ;
      RECT 6.445 8.605 6.615 8.775 ;
      RECT 6.38 1.415 6.55 1.585 ;
      RECT 6.38 4.135 6.55 4.305 ;
      RECT 6.375 5.945 6.545 6.115 ;
      RECT 6.255 2.49 6.425 2.66 ;
      RECT 5.92 1.415 6.09 1.585 ;
      RECT 5.92 4.135 6.09 4.305 ;
      RECT 5.565 1.97 5.735 2.14 ;
      RECT 5.49 2.44 5.66 2.61 ;
      RECT 5.46 1.415 5.63 1.585 ;
      RECT 5.46 4.135 5.63 4.305 ;
      RECT 5 1.415 5.17 1.585 ;
      RECT 5 4.135 5.17 4.305 ;
      RECT 4.64 2.165 4.81 2.335 ;
      RECT 4.54 1.415 4.71 1.585 ;
      RECT 4.54 4.135 4.71 4.305 ;
      RECT 4.3 3.36 4.47 3.53 ;
      RECT 4.265 2.695 4.435 2.865 ;
      RECT 4.08 1.415 4.25 1.585 ;
      RECT 4.08 4.135 4.25 4.305 ;
      RECT 3.655 2.55 3.825 2.72 ;
      RECT 3.62 1.415 3.79 1.585 ;
      RECT 3.62 4.135 3.79 4.305 ;
      RECT 3.585 3.25 3.755 3.42 ;
      RECT 3.525 2.085 3.695 2.255 ;
      RECT 3.16 1.415 3.33 1.585 ;
      RECT 3.16 4.135 3.33 4.305 ;
      RECT 2.885 3 3.055 3.17 ;
      RECT 2.7 1.415 2.87 1.585 ;
      RECT 2.7 4.135 2.87 4.305 ;
      RECT 2.38 2.505 2.55 2.675 ;
      RECT 2.24 1.415 2.41 1.585 ;
      RECT 2.24 4.135 2.41 4.305 ;
      RECT 2.16 3.25 2.33 3.42 ;
      RECT 1.955 2.13 2.125 2.3 ;
      RECT 1.78 1.415 1.95 1.585 ;
      RECT 1.78 4.135 1.95 4.305 ;
      RECT 1.685 3 1.855 3.17 ;
      RECT 1.645 2.43 1.815 2.6 ;
      RECT 1.32 1.415 1.49 1.585 ;
      RECT 1.32 4.135 1.49 4.305 ;
      RECT 1.1 3.475 1.27 3.645 ;
      RECT 0.96 2.095 1.13 2.265 ;
      RECT 0.86 1.415 1.03 1.585 ;
      RECT 0.86 4.135 1.03 4.305 ;
      RECT 0.4 1.415 0.57 1.585 ;
      RECT 0.4 4.135 0.57 4.305 ;
      RECT 0.39 3.015 0.56 3.185 ;
      RECT -0.45 4.545 -0.28 4.715 ;
      RECT -0.45 8.605 -0.28 8.775 ;
      RECT -0.76 6.685 -0.59 6.855 ;
      RECT -1.13 8.605 -0.96 8.775 ;
      RECT -1.19 7.055 -1.02 7.225 ;
      RECT -1.19 7.795 -1.02 7.965 ;
      RECT -1.565 6.315 -1.395 6.485 ;
      RECT -1.81 8.605 -1.64 8.775 ;
      RECT -2.49 8.605 -2.32 8.775 ;
      RECT -2.56 5.945 -2.39 6.115 ;
    LAYER li ;
      RECT 71.51 0 71.68 2.085 ;
      RECT 69.55 0 69.72 2.085 ;
      RECT 67.11 0 67.28 2.085 ;
      RECT 66.15 0 66.32 2.085 ;
      RECT 65.63 0 65.8 2.085 ;
      RECT 64.67 0 64.84 2.085 ;
      RECT 63.71 0 63.88 2.085 ;
      RECT 55.725 0 55.895 2.085 ;
      RECT 53.765 0 53.935 2.085 ;
      RECT 51.325 0 51.495 2.085 ;
      RECT 50.365 0 50.535 2.085 ;
      RECT 49.845 0 50.015 2.085 ;
      RECT 48.885 0 49.055 2.085 ;
      RECT 47.925 0 48.095 2.085 ;
      RECT 39.94 0 40.11 2.085 ;
      RECT 37.98 0 38.15 2.085 ;
      RECT 35.54 0 35.71 2.085 ;
      RECT 34.58 0 34.75 2.085 ;
      RECT 34.06 0 34.23 2.085 ;
      RECT 33.1 0 33.27 2.085 ;
      RECT 32.14 0 32.31 2.085 ;
      RECT 24.165 0 24.335 2.085 ;
      RECT 22.205 0 22.375 2.085 ;
      RECT 19.765 0 19.935 2.085 ;
      RECT 18.805 0 18.975 2.085 ;
      RECT 18.285 0 18.455 2.085 ;
      RECT 17.325 0 17.495 2.085 ;
      RECT 16.365 0 16.535 2.085 ;
      RECT 8.385 0 8.555 2.085 ;
      RECT 6.425 0 6.595 2.085 ;
      RECT 3.985 0 4.155 2.085 ;
      RECT 3.025 0 3.195 2.085 ;
      RECT 2.505 0 2.675 2.085 ;
      RECT 1.545 0 1.715 2.085 ;
      RECT 0.585 0 0.755 2.085 ;
      RECT 63.495 0 73.095 1.59 ;
      RECT 47.71 0 57.31 1.59 ;
      RECT 31.925 0 41.525 1.59 ;
      RECT 16.15 0 25.75 1.59 ;
      RECT 0.37 0 9.97 1.59 ;
      RECT 63.38 1.415 73.21 1.585 ;
      RECT 63.495 0 73.21 1.585 ;
      RECT 47.595 1.415 57.425 1.585 ;
      RECT 47.71 0 57.425 1.585 ;
      RECT 31.81 1.415 41.64 1.585 ;
      RECT 31.925 0 41.64 1.585 ;
      RECT 16.035 1.415 25.865 1.585 ;
      RECT 16.15 0 25.865 1.585 ;
      RECT 0.255 1.415 10.085 1.585 ;
      RECT 0.37 0 10.085 1.585 ;
      RECT 78.005 0 78.175 0.935 ;
      RECT 77.015 0 77.185 0.935 ;
      RECT 74.27 0 74.44 0.935 ;
      RECT 62.22 0 62.39 0.935 ;
      RECT 61.23 0 61.4 0.935 ;
      RECT 58.485 0 58.655 0.935 ;
      RECT 46.435 0 46.605 0.935 ;
      RECT 45.445 0 45.615 0.935 ;
      RECT 42.7 0 42.87 0.935 ;
      RECT 30.66 0 30.83 0.935 ;
      RECT 29.67 0 29.84 0.935 ;
      RECT 26.925 0 27.095 0.935 ;
      RECT 14.88 0 15.05 0.935 ;
      RECT 13.89 0 14.06 0.935 ;
      RECT 11.145 0 11.315 0.935 ;
      RECT -2.79 0 78.975 0.305 ;
      RECT -0.76 4.44 -0.59 8.305 ;
      RECT 78.005 3.405 78.175 5.475 ;
      RECT 77.015 3.405 77.185 5.475 ;
      RECT 74.27 3.405 74.44 5.475 ;
      RECT 69.49 4.135 69.66 5.475 ;
      RECT 62.22 3.405 62.39 5.475 ;
      RECT 61.23 3.405 61.4 5.475 ;
      RECT 58.485 3.405 58.655 5.475 ;
      RECT 53.705 4.135 53.875 5.475 ;
      RECT 46.435 3.405 46.605 5.475 ;
      RECT 45.445 3.405 45.615 5.475 ;
      RECT 42.7 3.405 42.87 5.475 ;
      RECT 37.92 4.135 38.09 5.475 ;
      RECT 30.66 3.405 30.83 5.475 ;
      RECT 29.67 3.405 29.84 5.475 ;
      RECT 26.925 3.405 27.095 5.475 ;
      RECT 22.145 4.135 22.315 5.475 ;
      RECT 14.88 3.405 15.05 5.475 ;
      RECT 13.89 3.405 14.06 5.475 ;
      RECT 11.145 3.405 11.315 5.475 ;
      RECT 6.365 4.135 6.535 5.475 ;
      RECT -2.57 4.44 -2.4 5.475 ;
      RECT -2.79 4.44 78.975 4.745 ;
      RECT 0.005 4.135 78.975 4.745 ;
      RECT 72.47 3.635 72.64 4.745 ;
      RECT 71.51 3.635 71.68 4.745 ;
      RECT 69.07 3.635 69.24 4.745 ;
      RECT 68.07 3.635 68.24 4.745 ;
      RECT 67.11 3.635 67.28 4.745 ;
      RECT 64.67 3.635 64.84 4.745 ;
      RECT 56.685 3.635 56.855 4.745 ;
      RECT 55.725 3.635 55.895 4.745 ;
      RECT 53.285 3.635 53.455 4.745 ;
      RECT 52.285 3.635 52.455 4.745 ;
      RECT 51.325 3.635 51.495 4.745 ;
      RECT 48.885 3.635 49.055 4.745 ;
      RECT 40.9 3.635 41.07 4.745 ;
      RECT 39.94 3.635 40.11 4.745 ;
      RECT 37.5 3.635 37.67 4.745 ;
      RECT 36.5 3.635 36.67 4.745 ;
      RECT 35.54 3.635 35.71 4.745 ;
      RECT 33.1 3.635 33.27 4.745 ;
      RECT 25.125 3.635 25.295 4.745 ;
      RECT 24.165 3.635 24.335 4.745 ;
      RECT 21.725 3.635 21.895 4.745 ;
      RECT 20.725 3.635 20.895 4.745 ;
      RECT 19.765 3.635 19.935 4.745 ;
      RECT 17.325 3.635 17.495 4.745 ;
      RECT 9.345 3.635 9.515 4.745 ;
      RECT 8.385 3.635 8.555 4.745 ;
      RECT 5.945 3.635 6.115 4.745 ;
      RECT 4.945 3.635 5.115 4.745 ;
      RECT 3.985 3.635 4.155 4.745 ;
      RECT 1.545 3.635 1.715 4.745 ;
      RECT -2.79 8.575 78.975 8.88 ;
      RECT 78.005 7.945 78.175 8.88 ;
      RECT 77.015 7.945 77.185 8.88 ;
      RECT 74.27 7.945 74.44 8.88 ;
      RECT 69.49 7.945 69.66 8.88 ;
      RECT 62.22 7.945 62.39 8.88 ;
      RECT 61.23 7.945 61.4 8.88 ;
      RECT 58.485 7.945 58.655 8.88 ;
      RECT 53.705 7.945 53.875 8.88 ;
      RECT 46.435 7.945 46.605 8.88 ;
      RECT 45.445 7.945 45.615 8.88 ;
      RECT 42.7 7.945 42.87 8.88 ;
      RECT 37.92 7.945 38.09 8.88 ;
      RECT 30.66 7.945 30.83 8.88 ;
      RECT 29.67 7.945 29.84 8.88 ;
      RECT 26.925 7.945 27.095 8.88 ;
      RECT 22.145 7.945 22.315 8.88 ;
      RECT 14.88 7.945 15.05 8.88 ;
      RECT 13.89 7.945 14.06 8.88 ;
      RECT 11.145 7.945 11.315 8.88 ;
      RECT 6.365 7.945 6.535 8.88 ;
      RECT -2.57 7.945 -2.4 8.88 ;
      RECT 78.065 1.74 78.235 2.935 ;
      RECT 78.065 1.74 78.53 1.91 ;
      RECT 78.065 6.97 78.53 7.14 ;
      RECT 78.065 5.945 78.235 7.14 ;
      RECT 77.075 1.74 77.245 2.935 ;
      RECT 77.075 1.74 77.54 1.91 ;
      RECT 77.075 6.97 77.54 7.14 ;
      RECT 77.075 5.945 77.245 7.14 ;
      RECT 75.22 2.635 75.39 3.865 ;
      RECT 75.275 0.855 75.445 2.805 ;
      RECT 75.22 0.575 75.39 1.025 ;
      RECT 75.22 7.855 75.39 8.305 ;
      RECT 75.275 6.075 75.445 8.025 ;
      RECT 75.22 5.015 75.39 6.245 ;
      RECT 74.7 0.575 74.87 3.865 ;
      RECT 74.7 2.075 75.105 2.405 ;
      RECT 74.7 1.235 75.105 1.565 ;
      RECT 74.7 5.015 74.87 8.305 ;
      RECT 74.7 7.315 75.105 7.645 ;
      RECT 74.7 6.475 75.105 6.805 ;
      RECT 72.035 1.975 72.765 2.215 ;
      RECT 72.577 1.77 72.765 2.215 ;
      RECT 72.405 1.782 72.78 2.209 ;
      RECT 72.32 1.797 72.8 2.194 ;
      RECT 72.32 1.812 72.805 2.184 ;
      RECT 72.275 1.832 72.82 2.176 ;
      RECT 72.252 1.867 72.835 2.13 ;
      RECT 72.166 1.89 72.84 2.09 ;
      RECT 72.166 1.908 72.85 2.06 ;
      RECT 72.035 1.977 72.855 2.023 ;
      RECT 72.08 1.92 72.85 2.06 ;
      RECT 72.166 1.872 72.835 2.13 ;
      RECT 72.252 1.841 72.82 2.176 ;
      RECT 72.275 1.822 72.805 2.184 ;
      RECT 72.32 1.795 72.78 2.209 ;
      RECT 72.405 1.777 72.765 2.215 ;
      RECT 72.491 1.771 72.765 2.215 ;
      RECT 72.577 1.766 72.71 2.215 ;
      RECT 72.663 1.761 72.71 2.215 ;
      RECT 72.355 2.659 72.525 3.045 ;
      RECT 72.35 2.659 72.525 3.04 ;
      RECT 72.325 2.659 72.525 3.005 ;
      RECT 72.325 2.687 72.535 2.995 ;
      RECT 72.305 2.687 72.535 2.955 ;
      RECT 72.3 2.687 72.535 2.928 ;
      RECT 72.3 2.705 72.54 2.92 ;
      RECT 72.245 2.705 72.54 2.855 ;
      RECT 72.245 2.722 72.55 2.838 ;
      RECT 72.235 2.722 72.55 2.778 ;
      RECT 72.235 2.739 72.555 2.775 ;
      RECT 72.23 2.575 72.4 2.753 ;
      RECT 72.23 2.609 72.486 2.753 ;
      RECT 72.225 3.375 72.23 3.388 ;
      RECT 72.22 3.27 72.225 3.393 ;
      RECT 72.195 3.13 72.22 3.408 ;
      RECT 72.16 3.081 72.195 3.44 ;
      RECT 72.155 3.049 72.16 3.46 ;
      RECT 72.15 3.04 72.155 3.46 ;
      RECT 72.07 3.005 72.15 3.46 ;
      RECT 72.007 2.975 72.07 3.46 ;
      RECT 71.921 2.963 72.007 3.46 ;
      RECT 71.835 2.949 71.921 3.46 ;
      RECT 71.755 2.936 71.835 3.446 ;
      RECT 71.72 2.928 71.755 3.426 ;
      RECT 71.71 2.925 71.72 3.417 ;
      RECT 71.68 2.92 71.71 3.404 ;
      RECT 71.63 2.895 71.68 3.38 ;
      RECT 71.616 2.869 71.63 3.362 ;
      RECT 71.53 2.829 71.616 3.338 ;
      RECT 71.485 2.777 71.53 3.307 ;
      RECT 71.475 2.752 71.485 3.294 ;
      RECT 71.47 2.533 71.475 2.555 ;
      RECT 71.465 2.735 71.475 3.29 ;
      RECT 71.465 2.531 71.47 2.645 ;
      RECT 71.455 2.527 71.465 3.286 ;
      RECT 71.411 2.525 71.455 3.274 ;
      RECT 71.325 2.525 71.411 3.245 ;
      RECT 71.295 2.525 71.325 3.218 ;
      RECT 71.28 2.525 71.295 3.206 ;
      RECT 71.24 2.537 71.28 3.191 ;
      RECT 71.22 2.556 71.24 3.17 ;
      RECT 71.21 2.566 71.22 3.154 ;
      RECT 71.2 2.572 71.21 3.143 ;
      RECT 71.18 2.582 71.2 3.126 ;
      RECT 71.175 2.591 71.18 3.113 ;
      RECT 71.17 2.595 71.175 3.063 ;
      RECT 71.16 2.601 71.17 2.98 ;
      RECT 71.155 2.605 71.16 2.894 ;
      RECT 71.15 2.625 71.155 2.831 ;
      RECT 71.145 2.648 71.15 2.778 ;
      RECT 71.14 2.666 71.145 2.723 ;
      RECT 71.75 2.485 71.92 2.745 ;
      RECT 71.92 2.45 71.965 2.731 ;
      RECT 71.881 2.452 71.97 2.714 ;
      RECT 71.77 2.469 72.056 2.685 ;
      RECT 71.77 2.484 72.06 2.657 ;
      RECT 71.77 2.465 71.97 2.714 ;
      RECT 71.795 2.453 71.92 2.745 ;
      RECT 71.881 2.451 71.965 2.731 ;
      RECT 70.935 1.84 71.105 2.33 ;
      RECT 70.935 1.84 71.14 2.31 ;
      RECT 71.07 1.76 71.18 2.27 ;
      RECT 71.051 1.764 71.2 2.24 ;
      RECT 70.965 1.772 71.22 2.223 ;
      RECT 70.965 1.778 71.225 2.213 ;
      RECT 70.965 1.787 71.245 2.201 ;
      RECT 70.94 1.812 71.275 2.179 ;
      RECT 70.94 1.832 71.28 2.159 ;
      RECT 70.935 1.845 71.29 2.139 ;
      RECT 70.935 1.912 71.295 2.12 ;
      RECT 70.935 2.045 71.3 2.107 ;
      RECT 70.93 1.85 71.29 1.94 ;
      RECT 70.94 1.807 71.245 2.201 ;
      RECT 71.051 1.762 71.18 2.27 ;
      RECT 70.925 3.515 71.225 3.77 ;
      RECT 71.01 3.481 71.225 3.77 ;
      RECT 71.01 3.484 71.23 3.63 ;
      RECT 70.945 3.505 71.23 3.63 ;
      RECT 70.98 3.495 71.225 3.77 ;
      RECT 70.975 3.5 71.23 3.63 ;
      RECT 71.01 3.479 71.211 3.77 ;
      RECT 71.096 3.47 71.211 3.77 ;
      RECT 71.096 3.464 71.125 3.77 ;
      RECT 70.585 3.105 70.595 3.595 ;
      RECT 70.245 3.04 70.255 3.34 ;
      RECT 70.76 3.212 70.765 3.431 ;
      RECT 70.75 3.192 70.76 3.448 ;
      RECT 70.74 3.172 70.75 3.478 ;
      RECT 70.735 3.162 70.74 3.493 ;
      RECT 70.73 3.158 70.735 3.498 ;
      RECT 70.715 3.15 70.73 3.505 ;
      RECT 70.675 3.13 70.715 3.53 ;
      RECT 70.65 3.112 70.675 3.563 ;
      RECT 70.645 3.11 70.65 3.576 ;
      RECT 70.625 3.107 70.645 3.58 ;
      RECT 70.595 3.105 70.625 3.59 ;
      RECT 70.525 3.107 70.585 3.591 ;
      RECT 70.505 3.107 70.525 3.585 ;
      RECT 70.48 3.105 70.505 3.582 ;
      RECT 70.445 3.1 70.48 3.578 ;
      RECT 70.425 3.094 70.445 3.565 ;
      RECT 70.415 3.091 70.425 3.553 ;
      RECT 70.395 3.088 70.415 3.538 ;
      RECT 70.375 3.084 70.395 3.52 ;
      RECT 70.37 3.081 70.375 3.51 ;
      RECT 70.365 3.08 70.37 3.508 ;
      RECT 70.355 3.077 70.365 3.5 ;
      RECT 70.345 3.071 70.355 3.483 ;
      RECT 70.335 3.065 70.345 3.465 ;
      RECT 70.325 3.059 70.335 3.453 ;
      RECT 70.315 3.053 70.325 3.433 ;
      RECT 70.31 3.049 70.315 3.418 ;
      RECT 70.305 3.047 70.31 3.41 ;
      RECT 70.3 3.045 70.305 3.403 ;
      RECT 70.295 3.043 70.3 3.393 ;
      RECT 70.29 3.041 70.295 3.387 ;
      RECT 70.28 3.04 70.29 3.377 ;
      RECT 70.27 3.04 70.28 3.368 ;
      RECT 70.255 3.04 70.27 3.353 ;
      RECT 70.215 3.04 70.245 3.337 ;
      RECT 70.195 3.042 70.215 3.332 ;
      RECT 70.19 3.047 70.195 3.33 ;
      RECT 70.16 3.055 70.19 3.328 ;
      RECT 70.13 3.07 70.16 3.327 ;
      RECT 70.085 3.092 70.13 3.332 ;
      RECT 70.08 3.107 70.085 3.336 ;
      RECT 70.065 3.112 70.08 3.338 ;
      RECT 70.06 3.116 70.065 3.34 ;
      RECT 70 3.139 70.06 3.349 ;
      RECT 69.98 3.165 70 3.362 ;
      RECT 69.97 3.172 69.98 3.366 ;
      RECT 69.955 3.179 69.97 3.369 ;
      RECT 69.935 3.189 69.955 3.372 ;
      RECT 69.93 3.197 69.935 3.375 ;
      RECT 69.885 3.202 69.93 3.382 ;
      RECT 69.875 3.205 69.885 3.389 ;
      RECT 69.865 3.205 69.875 3.393 ;
      RECT 69.83 3.207 69.865 3.405 ;
      RECT 69.81 3.21 69.83 3.418 ;
      RECT 69.77 3.213 69.81 3.429 ;
      RECT 69.755 3.215 69.77 3.442 ;
      RECT 69.745 3.215 69.755 3.447 ;
      RECT 69.72 3.216 69.745 3.455 ;
      RECT 69.71 3.218 69.72 3.46 ;
      RECT 69.705 3.219 69.71 3.463 ;
      RECT 69.68 3.217 69.705 3.466 ;
      RECT 69.665 3.215 69.68 3.467 ;
      RECT 69.645 3.212 69.665 3.469 ;
      RECT 69.625 3.207 69.645 3.469 ;
      RECT 69.565 3.202 69.625 3.466 ;
      RECT 69.53 3.177 69.565 3.462 ;
      RECT 69.52 3.154 69.53 3.46 ;
      RECT 69.49 3.131 69.52 3.46 ;
      RECT 69.48 3.11 69.49 3.46 ;
      RECT 69.455 3.092 69.48 3.458 ;
      RECT 69.44 3.07 69.455 3.455 ;
      RECT 69.425 3.052 69.44 3.453 ;
      RECT 69.405 3.042 69.425 3.451 ;
      RECT 69.39 3.037 69.405 3.45 ;
      RECT 69.375 3.035 69.39 3.449 ;
      RECT 69.345 3.036 69.375 3.447 ;
      RECT 69.325 3.039 69.345 3.445 ;
      RECT 69.268 3.043 69.325 3.445 ;
      RECT 69.182 3.052 69.268 3.445 ;
      RECT 69.096 3.063 69.182 3.445 ;
      RECT 69.01 3.074 69.096 3.445 ;
      RECT 68.99 3.081 69.01 3.453 ;
      RECT 68.98 3.084 68.99 3.46 ;
      RECT 68.915 3.089 68.98 3.478 ;
      RECT 68.885 3.096 68.915 3.503 ;
      RECT 68.875 3.099 68.885 3.51 ;
      RECT 68.83 3.103 68.875 3.515 ;
      RECT 68.8 3.108 68.83 3.52 ;
      RECT 68.799 3.11 68.8 3.52 ;
      RECT 68.713 3.116 68.799 3.52 ;
      RECT 68.627 3.127 68.713 3.52 ;
      RECT 68.541 3.139 68.627 3.52 ;
      RECT 68.455 3.15 68.541 3.52 ;
      RECT 68.44 3.157 68.455 3.515 ;
      RECT 68.435 3.159 68.44 3.509 ;
      RECT 68.415 3.17 68.435 3.504 ;
      RECT 68.405 3.188 68.415 3.498 ;
      RECT 68.4 3.2 68.405 3.298 ;
      RECT 70.695 1.953 70.715 2.04 ;
      RECT 70.69 1.888 70.695 2.072 ;
      RECT 70.68 1.855 70.69 2.077 ;
      RECT 70.675 1.835 70.68 2.083 ;
      RECT 70.645 1.835 70.675 2.1 ;
      RECT 70.596 1.835 70.645 2.136 ;
      RECT 70.51 1.835 70.596 2.194 ;
      RECT 70.481 1.845 70.51 2.243 ;
      RECT 70.395 1.887 70.481 2.296 ;
      RECT 70.375 1.925 70.395 2.343 ;
      RECT 70.35 1.942 70.375 2.363 ;
      RECT 70.34 1.956 70.35 2.383 ;
      RECT 70.335 1.962 70.34 2.393 ;
      RECT 70.33 1.966 70.335 2.4 ;
      RECT 70.28 1.986 70.33 2.405 ;
      RECT 70.215 2.03 70.28 2.405 ;
      RECT 70.19 2.08 70.215 2.405 ;
      RECT 70.18 2.11 70.19 2.405 ;
      RECT 70.175 2.137 70.18 2.405 ;
      RECT 70.17 2.155 70.175 2.405 ;
      RECT 70.16 2.197 70.17 2.405 ;
      RECT 70.51 2.755 70.68 2.93 ;
      RECT 70.45 2.583 70.51 2.918 ;
      RECT 70.44 2.576 70.45 2.901 ;
      RECT 70.395 2.755 70.68 2.881 ;
      RECT 70.376 2.755 70.68 2.859 ;
      RECT 70.29 2.755 70.68 2.824 ;
      RECT 70.27 2.575 70.44 2.78 ;
      RECT 70.27 2.722 70.675 2.78 ;
      RECT 70.27 2.67 70.65 2.78 ;
      RECT 70.27 2.625 70.615 2.78 ;
      RECT 70.27 2.607 70.58 2.78 ;
      RECT 70.27 2.597 70.575 2.78 ;
      RECT 70.44 7.855 70.61 8.305 ;
      RECT 70.495 6.075 70.665 8.025 ;
      RECT 70.44 5.015 70.61 6.245 ;
      RECT 69.92 5.015 70.09 8.305 ;
      RECT 69.92 7.315 70.325 7.645 ;
      RECT 69.92 6.475 70.325 6.805 ;
      RECT 69.99 3.555 70.18 3.78 ;
      RECT 69.98 3.556 70.185 3.775 ;
      RECT 69.98 3.558 70.195 3.755 ;
      RECT 69.98 3.562 70.2 3.74 ;
      RECT 69.98 3.549 70.15 3.775 ;
      RECT 69.98 3.552 70.175 3.775 ;
      RECT 69.99 3.548 70.15 3.78 ;
      RECT 70.076 3.546 70.15 3.78 ;
      RECT 69.7 2.797 69.87 3.035 ;
      RECT 69.7 2.797 69.956 2.949 ;
      RECT 69.7 2.797 69.96 2.859 ;
      RECT 69.75 2.57 69.97 2.838 ;
      RECT 69.745 2.587 69.975 2.811 ;
      RECT 69.71 2.745 69.975 2.811 ;
      RECT 69.73 2.595 69.87 3.035 ;
      RECT 69.72 2.677 69.98 2.794 ;
      RECT 69.715 2.725 69.98 2.794 ;
      RECT 69.72 2.635 69.975 2.811 ;
      RECT 69.745 2.572 69.97 2.838 ;
      RECT 69.31 2.547 69.48 2.745 ;
      RECT 69.31 2.547 69.525 2.72 ;
      RECT 69.38 2.49 69.55 2.678 ;
      RECT 69.355 2.505 69.55 2.678 ;
      RECT 68.97 2.551 69 2.745 ;
      RECT 68.965 2.523 68.97 2.745 ;
      RECT 68.935 2.497 68.965 2.747 ;
      RECT 68.91 2.455 68.935 2.75 ;
      RECT 68.9 2.427 68.91 2.752 ;
      RECT 68.865 2.407 68.9 2.754 ;
      RECT 68.8 2.392 68.865 2.76 ;
      RECT 68.75 2.39 68.8 2.766 ;
      RECT 68.727 2.392 68.75 2.771 ;
      RECT 68.641 2.403 68.727 2.777 ;
      RECT 68.555 2.421 68.641 2.787 ;
      RECT 68.54 2.432 68.555 2.793 ;
      RECT 68.47 2.455 68.54 2.799 ;
      RECT 68.415 2.487 68.47 2.807 ;
      RECT 68.375 2.51 68.415 2.813 ;
      RECT 68.361 2.523 68.375 2.816 ;
      RECT 68.275 2.545 68.361 2.822 ;
      RECT 68.26 2.57 68.275 2.828 ;
      RECT 68.22 2.585 68.26 2.832 ;
      RECT 68.17 2.6 68.22 2.837 ;
      RECT 68.145 2.607 68.17 2.841 ;
      RECT 68.085 2.602 68.145 2.845 ;
      RECT 68.07 2.593 68.085 2.849 ;
      RECT 68 2.583 68.07 2.845 ;
      RECT 67.975 2.575 67.995 2.835 ;
      RECT 67.916 2.575 67.975 2.813 ;
      RECT 67.83 2.575 67.916 2.77 ;
      RECT 67.995 2.575 68 2.84 ;
      RECT 68.69 1.806 68.86 2.14 ;
      RECT 68.66 1.806 68.86 2.135 ;
      RECT 68.6 1.773 68.66 2.123 ;
      RECT 68.6 1.829 68.87 2.118 ;
      RECT 68.575 1.829 68.87 2.112 ;
      RECT 68.57 1.77 68.6 2.109 ;
      RECT 68.555 1.776 68.69 2.107 ;
      RECT 68.55 1.784 68.775 2.095 ;
      RECT 68.55 1.836 68.885 2.048 ;
      RECT 68.535 1.792 68.775 2.043 ;
      RECT 68.535 1.862 68.895 1.984 ;
      RECT 68.505 1.812 68.86 1.945 ;
      RECT 68.505 1.902 68.905 1.941 ;
      RECT 68.555 1.781 68.775 2.107 ;
      RECT 67.895 2.111 67.95 2.375 ;
      RECT 67.895 2.111 68.015 2.374 ;
      RECT 67.895 2.111 68.04 2.373 ;
      RECT 67.895 2.111 68.105 2.372 ;
      RECT 68.04 2.077 68.12 2.371 ;
      RECT 67.855 2.121 68.265 2.37 ;
      RECT 67.895 2.118 68.265 2.37 ;
      RECT 67.855 2.126 68.27 2.363 ;
      RECT 67.84 2.128 68.27 2.362 ;
      RECT 67.84 2.135 68.275 2.358 ;
      RECT 67.82 2.134 68.27 2.354 ;
      RECT 67.82 2.142 68.28 2.353 ;
      RECT 67.815 2.139 68.275 2.349 ;
      RECT 67.815 2.152 68.29 2.348 ;
      RECT 67.8 2.142 68.28 2.347 ;
      RECT 67.765 2.155 68.29 2.34 ;
      RECT 67.95 2.11 68.26 2.37 ;
      RECT 67.95 2.095 68.21 2.37 ;
      RECT 68.015 2.082 68.145 2.37 ;
      RECT 67.56 3.171 67.575 3.564 ;
      RECT 67.525 3.176 67.575 3.563 ;
      RECT 67.56 3.175 67.62 3.562 ;
      RECT 67.505 3.186 67.62 3.561 ;
      RECT 67.52 3.182 67.62 3.561 ;
      RECT 67.485 3.192 67.695 3.558 ;
      RECT 67.485 3.211 67.74 3.556 ;
      RECT 67.485 3.218 67.745 3.553 ;
      RECT 67.47 3.195 67.695 3.55 ;
      RECT 67.45 3.2 67.695 3.543 ;
      RECT 67.445 3.204 67.695 3.539 ;
      RECT 67.445 3.221 67.755 3.538 ;
      RECT 67.425 3.215 67.74 3.534 ;
      RECT 67.425 3.224 67.76 3.528 ;
      RECT 67.42 3.23 67.76 3.3 ;
      RECT 67.485 3.19 67.62 3.558 ;
      RECT 67.36 2.553 67.56 2.865 ;
      RECT 67.435 2.531 67.56 2.865 ;
      RECT 67.375 2.55 67.565 2.85 ;
      RECT 67.345 2.561 67.565 2.848 ;
      RECT 67.36 2.556 67.57 2.814 ;
      RECT 67.345 2.66 67.575 2.781 ;
      RECT 67.375 2.532 67.56 2.865 ;
      RECT 67.435 2.51 67.535 2.865 ;
      RECT 67.46 2.507 67.535 2.865 ;
      RECT 67.46 2.502 67.48 2.865 ;
      RECT 66.865 2.57 67.04 2.745 ;
      RECT 66.86 2.57 67.04 2.743 ;
      RECT 66.835 2.57 67.04 2.738 ;
      RECT 66.78 2.55 66.95 2.728 ;
      RECT 66.78 2.557 67.015 2.728 ;
      RECT 66.865 3.237 66.88 3.42 ;
      RECT 66.855 3.215 66.865 3.42 ;
      RECT 66.84 3.195 66.855 3.42 ;
      RECT 66.83 3.17 66.84 3.42 ;
      RECT 66.8 3.135 66.83 3.42 ;
      RECT 66.765 3.075 66.8 3.42 ;
      RECT 66.76 3.037 66.765 3.42 ;
      RECT 66.71 2.988 66.76 3.42 ;
      RECT 66.7 2.938 66.71 3.408 ;
      RECT 66.685 2.917 66.7 3.368 ;
      RECT 66.665 2.885 66.685 3.318 ;
      RECT 66.64 2.841 66.665 3.258 ;
      RECT 66.635 2.813 66.64 3.213 ;
      RECT 66.63 2.804 66.635 3.199 ;
      RECT 66.625 2.797 66.63 3.186 ;
      RECT 66.62 2.792 66.625 3.175 ;
      RECT 66.615 2.777 66.62 3.165 ;
      RECT 66.61 2.755 66.615 3.152 ;
      RECT 66.6 2.715 66.61 3.127 ;
      RECT 66.575 2.645 66.6 3.083 ;
      RECT 66.57 2.585 66.575 3.048 ;
      RECT 66.555 2.565 66.57 3.015 ;
      RECT 66.55 2.565 66.555 2.99 ;
      RECT 66.52 2.565 66.55 2.945 ;
      RECT 66.475 2.565 66.52 2.885 ;
      RECT 66.4 2.565 66.475 2.833 ;
      RECT 66.395 2.565 66.4 2.798 ;
      RECT 66.39 2.565 66.395 2.788 ;
      RECT 66.385 2.565 66.39 2.768 ;
      RECT 66.65 1.785 66.82 2.255 ;
      RECT 66.595 1.778 66.79 2.239 ;
      RECT 66.595 1.792 66.825 2.238 ;
      RECT 66.58 1.793 66.825 2.219 ;
      RECT 66.575 1.811 66.825 2.205 ;
      RECT 66.58 1.794 66.83 2.203 ;
      RECT 66.565 1.825 66.83 2.188 ;
      RECT 66.58 1.8 66.835 2.173 ;
      RECT 66.56 1.84 66.835 2.17 ;
      RECT 66.575 1.812 66.84 2.155 ;
      RECT 66.575 1.824 66.845 2.135 ;
      RECT 66.56 1.84 66.85 2.118 ;
      RECT 66.56 1.85 66.855 1.973 ;
      RECT 66.555 1.85 66.855 1.93 ;
      RECT 66.555 1.865 66.86 1.908 ;
      RECT 66.65 1.775 66.79 2.255 ;
      RECT 66.65 1.773 66.76 2.255 ;
      RECT 66.736 1.77 66.76 2.255 ;
      RECT 66.395 3.437 66.4 3.483 ;
      RECT 66.385 3.285 66.395 3.507 ;
      RECT 66.38 3.13 66.385 3.532 ;
      RECT 66.365 3.092 66.38 3.543 ;
      RECT 66.36 3.075 66.365 3.55 ;
      RECT 66.35 3.063 66.36 3.557 ;
      RECT 66.345 3.054 66.35 3.559 ;
      RECT 66.34 3.052 66.345 3.563 ;
      RECT 66.295 3.043 66.34 3.578 ;
      RECT 66.29 3.035 66.295 3.592 ;
      RECT 66.285 3.032 66.29 3.596 ;
      RECT 66.27 3.027 66.285 3.604 ;
      RECT 66.215 3.017 66.27 3.615 ;
      RECT 66.18 3.005 66.215 3.616 ;
      RECT 66.171 3 66.18 3.61 ;
      RECT 66.085 3 66.171 3.6 ;
      RECT 66.055 3 66.085 3.578 ;
      RECT 66.045 3 66.05 3.558 ;
      RECT 66.04 3 66.045 3.52 ;
      RECT 66.035 3 66.04 3.478 ;
      RECT 66.03 3 66.035 3.438 ;
      RECT 66.025 3 66.03 3.368 ;
      RECT 66.015 3 66.025 3.29 ;
      RECT 66.01 3 66.015 3.19 ;
      RECT 66.05 3 66.055 3.56 ;
      RECT 65.545 3.082 65.635 3.56 ;
      RECT 65.53 3.085 65.65 3.558 ;
      RECT 65.545 3.084 65.65 3.558 ;
      RECT 65.51 3.091 65.675 3.548 ;
      RECT 65.53 3.085 65.675 3.548 ;
      RECT 65.495 3.097 65.675 3.536 ;
      RECT 65.53 3.088 65.725 3.529 ;
      RECT 65.481 3.105 65.725 3.527 ;
      RECT 65.51 3.095 65.735 3.515 ;
      RECT 65.481 3.116 65.765 3.506 ;
      RECT 65.395 3.14 65.765 3.5 ;
      RECT 65.395 3.153 65.805 3.483 ;
      RECT 65.39 3.175 65.805 3.476 ;
      RECT 65.36 3.19 65.805 3.466 ;
      RECT 65.355 3.201 65.805 3.456 ;
      RECT 65.325 3.214 65.805 3.447 ;
      RECT 65.31 3.232 65.805 3.436 ;
      RECT 65.285 3.245 65.805 3.426 ;
      RECT 65.545 3.081 65.555 3.56 ;
      RECT 65.591 2.505 65.63 2.75 ;
      RECT 65.505 2.505 65.64 2.748 ;
      RECT 65.39 2.53 65.64 2.745 ;
      RECT 65.39 2.53 65.645 2.743 ;
      RECT 65.39 2.53 65.66 2.738 ;
      RECT 65.496 2.505 65.675 2.718 ;
      RECT 65.41 2.513 65.675 2.718 ;
      RECT 65.08 1.865 65.25 2.3 ;
      RECT 65.07 1.899 65.25 2.283 ;
      RECT 65.15 1.835 65.32 2.27 ;
      RECT 65.055 1.91 65.32 2.248 ;
      RECT 65.15 1.845 65.325 2.238 ;
      RECT 65.08 1.897 65.355 2.223 ;
      RECT 65.04 1.923 65.355 2.208 ;
      RECT 65.04 1.965 65.365 2.188 ;
      RECT 65.035 1.99 65.37 2.17 ;
      RECT 65.035 2 65.375 2.155 ;
      RECT 65.03 1.937 65.355 2.153 ;
      RECT 65.03 2.01 65.38 2.138 ;
      RECT 65.025 1.947 65.355 2.135 ;
      RECT 65.02 2.031 65.385 2.118 ;
      RECT 65.02 2.063 65.39 2.098 ;
      RECT 65.015 1.977 65.365 2.09 ;
      RECT 65.02 1.962 65.355 2.118 ;
      RECT 65.035 1.932 65.355 2.17 ;
      RECT 64.88 2.519 65.105 2.775 ;
      RECT 64.88 2.552 65.125 2.765 ;
      RECT 64.845 2.552 65.125 2.763 ;
      RECT 64.845 2.565 65.13 2.753 ;
      RECT 64.845 2.585 65.14 2.745 ;
      RECT 64.845 2.682 65.145 2.738 ;
      RECT 64.825 2.43 64.955 2.728 ;
      RECT 64.78 2.585 65.14 2.67 ;
      RECT 64.77 2.43 64.955 2.615 ;
      RECT 64.77 2.462 65.041 2.615 ;
      RECT 64.735 2.992 64.755 3.17 ;
      RECT 64.7 2.945 64.735 3.17 ;
      RECT 64.685 2.885 64.7 3.17 ;
      RECT 64.66 2.832 64.685 3.17 ;
      RECT 64.645 2.785 64.66 3.17 ;
      RECT 64.625 2.762 64.645 3.17 ;
      RECT 64.6 2.727 64.625 3.17 ;
      RECT 64.59 2.573 64.6 3.17 ;
      RECT 64.56 2.568 64.59 3.161 ;
      RECT 64.555 2.565 64.56 3.151 ;
      RECT 64.54 2.565 64.555 3.125 ;
      RECT 64.535 2.565 64.54 3.088 ;
      RECT 64.51 2.565 64.535 3.04 ;
      RECT 64.49 2.565 64.51 2.965 ;
      RECT 64.48 2.565 64.49 2.925 ;
      RECT 64.475 2.565 64.48 2.9 ;
      RECT 64.47 2.565 64.475 2.883 ;
      RECT 64.465 2.565 64.47 2.865 ;
      RECT 64.46 2.566 64.465 2.855 ;
      RECT 64.45 2.568 64.46 2.823 ;
      RECT 64.44 2.57 64.45 2.79 ;
      RECT 64.43 2.573 64.44 2.763 ;
      RECT 64.755 3 64.98 3.17 ;
      RECT 64.085 1.812 64.255 2.265 ;
      RECT 64.085 1.812 64.345 2.231 ;
      RECT 64.085 1.812 64.375 2.215 ;
      RECT 64.085 1.812 64.405 2.188 ;
      RECT 64.341 1.79 64.42 2.17 ;
      RECT 64.12 1.797 64.425 2.155 ;
      RECT 64.12 1.805 64.435 2.118 ;
      RECT 64.08 1.832 64.435 2.09 ;
      RECT 64.065 1.845 64.435 2.055 ;
      RECT 64.085 1.82 64.455 2.045 ;
      RECT 64.06 1.885 64.455 2.015 ;
      RECT 64.06 1.915 64.46 1.998 ;
      RECT 64.055 1.945 64.46 1.985 ;
      RECT 64.12 1.794 64.42 2.17 ;
      RECT 64.255 1.791 64.341 2.249 ;
      RECT 64.206 1.792 64.42 2.17 ;
      RECT 64.35 3.452 64.395 3.645 ;
      RECT 64.34 3.422 64.35 3.645 ;
      RECT 64.335 3.407 64.34 3.645 ;
      RECT 64.295 3.317 64.335 3.645 ;
      RECT 64.29 3.23 64.295 3.645 ;
      RECT 64.28 3.2 64.29 3.645 ;
      RECT 64.275 3.16 64.28 3.645 ;
      RECT 64.265 3.122 64.275 3.645 ;
      RECT 64.26 3.087 64.265 3.645 ;
      RECT 64.24 3.04 64.26 3.645 ;
      RECT 64.225 2.965 64.24 3.645 ;
      RECT 64.22 2.92 64.225 3.64 ;
      RECT 64.215 2.9 64.22 3.613 ;
      RECT 64.21 2.88 64.215 3.598 ;
      RECT 64.205 2.855 64.21 3.578 ;
      RECT 64.2 2.833 64.205 3.563 ;
      RECT 64.195 2.811 64.2 3.545 ;
      RECT 64.19 2.79 64.195 3.535 ;
      RECT 64.18 2.762 64.19 3.505 ;
      RECT 64.17 2.725 64.18 3.473 ;
      RECT 64.16 2.685 64.17 3.44 ;
      RECT 64.15 2.663 64.16 3.41 ;
      RECT 64.12 2.615 64.15 3.342 ;
      RECT 64.105 2.575 64.12 3.269 ;
      RECT 64.095 2.575 64.105 3.235 ;
      RECT 64.09 2.575 64.095 3.21 ;
      RECT 64.085 2.575 64.09 3.195 ;
      RECT 64.08 2.575 64.085 3.173 ;
      RECT 64.075 2.575 64.08 3.16 ;
      RECT 64.06 2.575 64.075 3.125 ;
      RECT 64.04 2.575 64.06 3.065 ;
      RECT 64.03 2.575 64.04 3.015 ;
      RECT 64.01 2.575 64.03 2.963 ;
      RECT 63.99 2.575 64.01 2.92 ;
      RECT 63.98 2.575 63.99 2.908 ;
      RECT 63.95 2.575 63.98 2.895 ;
      RECT 63.92 2.596 63.95 2.875 ;
      RECT 63.91 2.624 63.92 2.855 ;
      RECT 63.895 2.641 63.91 2.823 ;
      RECT 63.89 2.655 63.895 2.79 ;
      RECT 63.885 2.663 63.89 2.763 ;
      RECT 63.88 2.671 63.885 2.725 ;
      RECT 63.885 3.195 63.89 3.53 ;
      RECT 63.85 3.182 63.885 3.529 ;
      RECT 63.78 3.122 63.85 3.528 ;
      RECT 63.7 3.065 63.78 3.527 ;
      RECT 63.565 3.025 63.7 3.526 ;
      RECT 63.565 3.212 63.9 3.515 ;
      RECT 63.525 3.212 63.9 3.505 ;
      RECT 63.525 3.23 63.905 3.5 ;
      RECT 63.525 3.32 63.91 3.49 ;
      RECT 63.52 3.015 63.685 3.47 ;
      RECT 63.515 3.015 63.685 3.213 ;
      RECT 63.515 3.172 63.88 3.213 ;
      RECT 63.515 3.16 63.875 3.213 ;
      RECT 62.28 1.74 62.45 2.935 ;
      RECT 62.28 1.74 62.745 1.91 ;
      RECT 62.28 6.97 62.745 7.14 ;
      RECT 62.28 5.945 62.45 7.14 ;
      RECT 61.29 1.74 61.46 2.935 ;
      RECT 61.29 1.74 61.755 1.91 ;
      RECT 61.29 6.97 61.755 7.14 ;
      RECT 61.29 5.945 61.46 7.14 ;
      RECT 59.435 2.635 59.605 3.865 ;
      RECT 59.49 0.855 59.66 2.805 ;
      RECT 59.435 0.575 59.605 1.025 ;
      RECT 59.435 7.855 59.605 8.305 ;
      RECT 59.49 6.075 59.66 8.025 ;
      RECT 59.435 5.015 59.605 6.245 ;
      RECT 58.915 0.575 59.085 3.865 ;
      RECT 58.915 2.075 59.32 2.405 ;
      RECT 58.915 1.235 59.32 1.565 ;
      RECT 58.915 5.015 59.085 8.305 ;
      RECT 58.915 7.315 59.32 7.645 ;
      RECT 58.915 6.475 59.32 6.805 ;
      RECT 56.25 1.975 56.98 2.215 ;
      RECT 56.792 1.77 56.98 2.215 ;
      RECT 56.62 1.782 56.995 2.209 ;
      RECT 56.535 1.797 57.015 2.194 ;
      RECT 56.535 1.812 57.02 2.184 ;
      RECT 56.49 1.832 57.035 2.176 ;
      RECT 56.467 1.867 57.05 2.13 ;
      RECT 56.381 1.89 57.055 2.09 ;
      RECT 56.381 1.908 57.065 2.06 ;
      RECT 56.25 1.977 57.07 2.023 ;
      RECT 56.295 1.92 57.065 2.06 ;
      RECT 56.381 1.872 57.05 2.13 ;
      RECT 56.467 1.841 57.035 2.176 ;
      RECT 56.49 1.822 57.02 2.184 ;
      RECT 56.535 1.795 56.995 2.209 ;
      RECT 56.62 1.777 56.98 2.215 ;
      RECT 56.706 1.771 56.98 2.215 ;
      RECT 56.792 1.766 56.925 2.215 ;
      RECT 56.878 1.761 56.925 2.215 ;
      RECT 56.57 2.659 56.74 3.045 ;
      RECT 56.565 2.659 56.74 3.04 ;
      RECT 56.54 2.659 56.74 3.005 ;
      RECT 56.54 2.687 56.75 2.995 ;
      RECT 56.52 2.687 56.75 2.955 ;
      RECT 56.515 2.687 56.75 2.928 ;
      RECT 56.515 2.705 56.755 2.92 ;
      RECT 56.46 2.705 56.755 2.855 ;
      RECT 56.46 2.722 56.765 2.838 ;
      RECT 56.45 2.722 56.765 2.778 ;
      RECT 56.45 2.739 56.77 2.775 ;
      RECT 56.445 2.575 56.615 2.753 ;
      RECT 56.445 2.609 56.701 2.753 ;
      RECT 56.44 3.375 56.445 3.388 ;
      RECT 56.435 3.27 56.44 3.393 ;
      RECT 56.41 3.13 56.435 3.408 ;
      RECT 56.375 3.081 56.41 3.44 ;
      RECT 56.37 3.049 56.375 3.46 ;
      RECT 56.365 3.04 56.37 3.46 ;
      RECT 56.285 3.005 56.365 3.46 ;
      RECT 56.222 2.975 56.285 3.46 ;
      RECT 56.136 2.963 56.222 3.46 ;
      RECT 56.05 2.949 56.136 3.46 ;
      RECT 55.97 2.936 56.05 3.446 ;
      RECT 55.935 2.928 55.97 3.426 ;
      RECT 55.925 2.925 55.935 3.417 ;
      RECT 55.895 2.92 55.925 3.404 ;
      RECT 55.845 2.895 55.895 3.38 ;
      RECT 55.831 2.869 55.845 3.362 ;
      RECT 55.745 2.829 55.831 3.338 ;
      RECT 55.7 2.777 55.745 3.307 ;
      RECT 55.69 2.752 55.7 3.294 ;
      RECT 55.685 2.533 55.69 2.555 ;
      RECT 55.68 2.735 55.69 3.29 ;
      RECT 55.68 2.531 55.685 2.645 ;
      RECT 55.67 2.527 55.68 3.286 ;
      RECT 55.626 2.525 55.67 3.274 ;
      RECT 55.54 2.525 55.626 3.245 ;
      RECT 55.51 2.525 55.54 3.218 ;
      RECT 55.495 2.525 55.51 3.206 ;
      RECT 55.455 2.537 55.495 3.191 ;
      RECT 55.435 2.556 55.455 3.17 ;
      RECT 55.425 2.566 55.435 3.154 ;
      RECT 55.415 2.572 55.425 3.143 ;
      RECT 55.395 2.582 55.415 3.126 ;
      RECT 55.39 2.591 55.395 3.113 ;
      RECT 55.385 2.595 55.39 3.063 ;
      RECT 55.375 2.601 55.385 2.98 ;
      RECT 55.37 2.605 55.375 2.894 ;
      RECT 55.365 2.625 55.37 2.831 ;
      RECT 55.36 2.648 55.365 2.778 ;
      RECT 55.355 2.666 55.36 2.723 ;
      RECT 55.965 2.485 56.135 2.745 ;
      RECT 56.135 2.45 56.18 2.731 ;
      RECT 56.096 2.452 56.185 2.714 ;
      RECT 55.985 2.469 56.271 2.685 ;
      RECT 55.985 2.484 56.275 2.657 ;
      RECT 55.985 2.465 56.185 2.714 ;
      RECT 56.01 2.453 56.135 2.745 ;
      RECT 56.096 2.451 56.18 2.731 ;
      RECT 55.15 1.84 55.32 2.33 ;
      RECT 55.15 1.84 55.355 2.31 ;
      RECT 55.285 1.76 55.395 2.27 ;
      RECT 55.266 1.764 55.415 2.24 ;
      RECT 55.18 1.772 55.435 2.223 ;
      RECT 55.18 1.778 55.44 2.213 ;
      RECT 55.18 1.787 55.46 2.201 ;
      RECT 55.155 1.812 55.49 2.179 ;
      RECT 55.155 1.832 55.495 2.159 ;
      RECT 55.15 1.845 55.505 2.139 ;
      RECT 55.15 1.912 55.51 2.12 ;
      RECT 55.15 2.045 55.515 2.107 ;
      RECT 55.145 1.85 55.505 1.94 ;
      RECT 55.155 1.807 55.46 2.201 ;
      RECT 55.266 1.762 55.395 2.27 ;
      RECT 55.14 3.515 55.44 3.77 ;
      RECT 55.225 3.481 55.44 3.77 ;
      RECT 55.225 3.484 55.445 3.63 ;
      RECT 55.16 3.505 55.445 3.63 ;
      RECT 55.195 3.495 55.44 3.77 ;
      RECT 55.19 3.5 55.445 3.63 ;
      RECT 55.225 3.479 55.426 3.77 ;
      RECT 55.311 3.47 55.426 3.77 ;
      RECT 55.311 3.464 55.34 3.77 ;
      RECT 54.8 3.105 54.81 3.595 ;
      RECT 54.46 3.04 54.47 3.34 ;
      RECT 54.975 3.212 54.98 3.431 ;
      RECT 54.965 3.192 54.975 3.448 ;
      RECT 54.955 3.172 54.965 3.478 ;
      RECT 54.95 3.162 54.955 3.493 ;
      RECT 54.945 3.158 54.95 3.498 ;
      RECT 54.93 3.15 54.945 3.505 ;
      RECT 54.89 3.13 54.93 3.53 ;
      RECT 54.865 3.112 54.89 3.563 ;
      RECT 54.86 3.11 54.865 3.576 ;
      RECT 54.84 3.107 54.86 3.58 ;
      RECT 54.81 3.105 54.84 3.59 ;
      RECT 54.74 3.107 54.8 3.591 ;
      RECT 54.72 3.107 54.74 3.585 ;
      RECT 54.695 3.105 54.72 3.582 ;
      RECT 54.66 3.1 54.695 3.578 ;
      RECT 54.64 3.094 54.66 3.565 ;
      RECT 54.63 3.091 54.64 3.553 ;
      RECT 54.61 3.088 54.63 3.538 ;
      RECT 54.59 3.084 54.61 3.52 ;
      RECT 54.585 3.081 54.59 3.51 ;
      RECT 54.58 3.08 54.585 3.508 ;
      RECT 54.57 3.077 54.58 3.5 ;
      RECT 54.56 3.071 54.57 3.483 ;
      RECT 54.55 3.065 54.56 3.465 ;
      RECT 54.54 3.059 54.55 3.453 ;
      RECT 54.53 3.053 54.54 3.433 ;
      RECT 54.525 3.049 54.53 3.418 ;
      RECT 54.52 3.047 54.525 3.41 ;
      RECT 54.515 3.045 54.52 3.403 ;
      RECT 54.51 3.043 54.515 3.393 ;
      RECT 54.505 3.041 54.51 3.387 ;
      RECT 54.495 3.04 54.505 3.377 ;
      RECT 54.485 3.04 54.495 3.368 ;
      RECT 54.47 3.04 54.485 3.353 ;
      RECT 54.43 3.04 54.46 3.337 ;
      RECT 54.41 3.042 54.43 3.332 ;
      RECT 54.405 3.047 54.41 3.33 ;
      RECT 54.375 3.055 54.405 3.328 ;
      RECT 54.345 3.07 54.375 3.327 ;
      RECT 54.3 3.092 54.345 3.332 ;
      RECT 54.295 3.107 54.3 3.336 ;
      RECT 54.28 3.112 54.295 3.338 ;
      RECT 54.275 3.116 54.28 3.34 ;
      RECT 54.215 3.139 54.275 3.349 ;
      RECT 54.195 3.165 54.215 3.362 ;
      RECT 54.185 3.172 54.195 3.366 ;
      RECT 54.17 3.179 54.185 3.369 ;
      RECT 54.15 3.189 54.17 3.372 ;
      RECT 54.145 3.197 54.15 3.375 ;
      RECT 54.1 3.202 54.145 3.382 ;
      RECT 54.09 3.205 54.1 3.389 ;
      RECT 54.08 3.205 54.09 3.393 ;
      RECT 54.045 3.207 54.08 3.405 ;
      RECT 54.025 3.21 54.045 3.418 ;
      RECT 53.985 3.213 54.025 3.429 ;
      RECT 53.97 3.215 53.985 3.442 ;
      RECT 53.96 3.215 53.97 3.447 ;
      RECT 53.935 3.216 53.96 3.455 ;
      RECT 53.925 3.218 53.935 3.46 ;
      RECT 53.92 3.219 53.925 3.463 ;
      RECT 53.895 3.217 53.92 3.466 ;
      RECT 53.88 3.215 53.895 3.467 ;
      RECT 53.86 3.212 53.88 3.469 ;
      RECT 53.84 3.207 53.86 3.469 ;
      RECT 53.78 3.202 53.84 3.466 ;
      RECT 53.745 3.177 53.78 3.462 ;
      RECT 53.735 3.154 53.745 3.46 ;
      RECT 53.705 3.131 53.735 3.46 ;
      RECT 53.695 3.11 53.705 3.46 ;
      RECT 53.67 3.092 53.695 3.458 ;
      RECT 53.655 3.07 53.67 3.455 ;
      RECT 53.64 3.052 53.655 3.453 ;
      RECT 53.62 3.042 53.64 3.451 ;
      RECT 53.605 3.037 53.62 3.45 ;
      RECT 53.59 3.035 53.605 3.449 ;
      RECT 53.56 3.036 53.59 3.447 ;
      RECT 53.54 3.039 53.56 3.445 ;
      RECT 53.483 3.043 53.54 3.445 ;
      RECT 53.397 3.052 53.483 3.445 ;
      RECT 53.311 3.063 53.397 3.445 ;
      RECT 53.225 3.074 53.311 3.445 ;
      RECT 53.205 3.081 53.225 3.453 ;
      RECT 53.195 3.084 53.205 3.46 ;
      RECT 53.13 3.089 53.195 3.478 ;
      RECT 53.1 3.096 53.13 3.503 ;
      RECT 53.09 3.099 53.1 3.51 ;
      RECT 53.045 3.103 53.09 3.515 ;
      RECT 53.015 3.108 53.045 3.52 ;
      RECT 53.014 3.11 53.015 3.52 ;
      RECT 52.928 3.116 53.014 3.52 ;
      RECT 52.842 3.127 52.928 3.52 ;
      RECT 52.756 3.139 52.842 3.52 ;
      RECT 52.67 3.15 52.756 3.52 ;
      RECT 52.655 3.157 52.67 3.515 ;
      RECT 52.65 3.159 52.655 3.509 ;
      RECT 52.63 3.17 52.65 3.504 ;
      RECT 52.62 3.188 52.63 3.498 ;
      RECT 52.615 3.2 52.62 3.298 ;
      RECT 54.91 1.953 54.93 2.04 ;
      RECT 54.905 1.888 54.91 2.072 ;
      RECT 54.895 1.855 54.905 2.077 ;
      RECT 54.89 1.835 54.895 2.083 ;
      RECT 54.86 1.835 54.89 2.1 ;
      RECT 54.811 1.835 54.86 2.136 ;
      RECT 54.725 1.835 54.811 2.194 ;
      RECT 54.696 1.845 54.725 2.243 ;
      RECT 54.61 1.887 54.696 2.296 ;
      RECT 54.59 1.925 54.61 2.343 ;
      RECT 54.565 1.942 54.59 2.363 ;
      RECT 54.555 1.956 54.565 2.383 ;
      RECT 54.55 1.962 54.555 2.393 ;
      RECT 54.545 1.966 54.55 2.4 ;
      RECT 54.495 1.986 54.545 2.405 ;
      RECT 54.43 2.03 54.495 2.405 ;
      RECT 54.405 2.08 54.43 2.405 ;
      RECT 54.395 2.11 54.405 2.405 ;
      RECT 54.39 2.137 54.395 2.405 ;
      RECT 54.385 2.155 54.39 2.405 ;
      RECT 54.375 2.197 54.385 2.405 ;
      RECT 54.725 2.755 54.895 2.93 ;
      RECT 54.665 2.583 54.725 2.918 ;
      RECT 54.655 2.576 54.665 2.901 ;
      RECT 54.61 2.755 54.895 2.881 ;
      RECT 54.591 2.755 54.895 2.859 ;
      RECT 54.505 2.755 54.895 2.824 ;
      RECT 54.485 2.575 54.655 2.78 ;
      RECT 54.485 2.722 54.89 2.78 ;
      RECT 54.485 2.67 54.865 2.78 ;
      RECT 54.485 2.625 54.83 2.78 ;
      RECT 54.485 2.607 54.795 2.78 ;
      RECT 54.485 2.597 54.79 2.78 ;
      RECT 54.655 7.855 54.825 8.305 ;
      RECT 54.71 6.075 54.88 8.025 ;
      RECT 54.655 5.015 54.825 6.245 ;
      RECT 54.135 5.015 54.305 8.305 ;
      RECT 54.135 7.315 54.54 7.645 ;
      RECT 54.135 6.475 54.54 6.805 ;
      RECT 54.205 3.555 54.395 3.78 ;
      RECT 54.195 3.556 54.4 3.775 ;
      RECT 54.195 3.558 54.41 3.755 ;
      RECT 54.195 3.562 54.415 3.74 ;
      RECT 54.195 3.549 54.365 3.775 ;
      RECT 54.195 3.552 54.39 3.775 ;
      RECT 54.205 3.548 54.365 3.78 ;
      RECT 54.291 3.546 54.365 3.78 ;
      RECT 53.915 2.797 54.085 3.035 ;
      RECT 53.915 2.797 54.171 2.949 ;
      RECT 53.915 2.797 54.175 2.859 ;
      RECT 53.965 2.57 54.185 2.838 ;
      RECT 53.96 2.587 54.19 2.811 ;
      RECT 53.925 2.745 54.19 2.811 ;
      RECT 53.945 2.595 54.085 3.035 ;
      RECT 53.935 2.677 54.195 2.794 ;
      RECT 53.93 2.725 54.195 2.794 ;
      RECT 53.935 2.635 54.19 2.811 ;
      RECT 53.96 2.572 54.185 2.838 ;
      RECT 53.525 2.547 53.695 2.745 ;
      RECT 53.525 2.547 53.74 2.72 ;
      RECT 53.595 2.49 53.765 2.678 ;
      RECT 53.57 2.505 53.765 2.678 ;
      RECT 53.185 2.551 53.215 2.745 ;
      RECT 53.18 2.523 53.185 2.745 ;
      RECT 53.15 2.497 53.18 2.747 ;
      RECT 53.125 2.455 53.15 2.75 ;
      RECT 53.115 2.427 53.125 2.752 ;
      RECT 53.08 2.407 53.115 2.754 ;
      RECT 53.015 2.392 53.08 2.76 ;
      RECT 52.965 2.39 53.015 2.766 ;
      RECT 52.942 2.392 52.965 2.771 ;
      RECT 52.856 2.403 52.942 2.777 ;
      RECT 52.77 2.421 52.856 2.787 ;
      RECT 52.755 2.432 52.77 2.793 ;
      RECT 52.685 2.455 52.755 2.799 ;
      RECT 52.63 2.487 52.685 2.807 ;
      RECT 52.59 2.51 52.63 2.813 ;
      RECT 52.576 2.523 52.59 2.816 ;
      RECT 52.49 2.545 52.576 2.822 ;
      RECT 52.475 2.57 52.49 2.828 ;
      RECT 52.435 2.585 52.475 2.832 ;
      RECT 52.385 2.6 52.435 2.837 ;
      RECT 52.36 2.607 52.385 2.841 ;
      RECT 52.3 2.602 52.36 2.845 ;
      RECT 52.285 2.593 52.3 2.849 ;
      RECT 52.215 2.583 52.285 2.845 ;
      RECT 52.19 2.575 52.21 2.835 ;
      RECT 52.131 2.575 52.19 2.813 ;
      RECT 52.045 2.575 52.131 2.77 ;
      RECT 52.21 2.575 52.215 2.84 ;
      RECT 52.905 1.806 53.075 2.14 ;
      RECT 52.875 1.806 53.075 2.135 ;
      RECT 52.815 1.773 52.875 2.123 ;
      RECT 52.815 1.829 53.085 2.118 ;
      RECT 52.79 1.829 53.085 2.112 ;
      RECT 52.785 1.77 52.815 2.109 ;
      RECT 52.77 1.776 52.905 2.107 ;
      RECT 52.765 1.784 52.99 2.095 ;
      RECT 52.765 1.836 53.1 2.048 ;
      RECT 52.75 1.792 52.99 2.043 ;
      RECT 52.75 1.862 53.11 1.984 ;
      RECT 52.72 1.812 53.075 1.945 ;
      RECT 52.72 1.902 53.12 1.941 ;
      RECT 52.77 1.781 52.99 2.107 ;
      RECT 52.11 2.111 52.165 2.375 ;
      RECT 52.11 2.111 52.23 2.374 ;
      RECT 52.11 2.111 52.255 2.373 ;
      RECT 52.11 2.111 52.32 2.372 ;
      RECT 52.255 2.077 52.335 2.371 ;
      RECT 52.07 2.121 52.48 2.37 ;
      RECT 52.11 2.118 52.48 2.37 ;
      RECT 52.07 2.126 52.485 2.363 ;
      RECT 52.055 2.128 52.485 2.362 ;
      RECT 52.055 2.135 52.49 2.358 ;
      RECT 52.035 2.134 52.485 2.354 ;
      RECT 52.035 2.142 52.495 2.353 ;
      RECT 52.03 2.139 52.49 2.349 ;
      RECT 52.03 2.152 52.505 2.348 ;
      RECT 52.015 2.142 52.495 2.347 ;
      RECT 51.98 2.155 52.505 2.34 ;
      RECT 52.165 2.11 52.475 2.37 ;
      RECT 52.165 2.095 52.425 2.37 ;
      RECT 52.23 2.082 52.36 2.37 ;
      RECT 51.775 3.171 51.79 3.564 ;
      RECT 51.74 3.176 51.79 3.563 ;
      RECT 51.775 3.175 51.835 3.562 ;
      RECT 51.72 3.186 51.835 3.561 ;
      RECT 51.735 3.182 51.835 3.561 ;
      RECT 51.7 3.192 51.91 3.558 ;
      RECT 51.7 3.211 51.955 3.556 ;
      RECT 51.7 3.218 51.96 3.553 ;
      RECT 51.685 3.195 51.91 3.55 ;
      RECT 51.665 3.2 51.91 3.543 ;
      RECT 51.66 3.204 51.91 3.539 ;
      RECT 51.66 3.221 51.97 3.538 ;
      RECT 51.64 3.215 51.955 3.534 ;
      RECT 51.64 3.224 51.975 3.528 ;
      RECT 51.635 3.23 51.975 3.3 ;
      RECT 51.7 3.19 51.835 3.558 ;
      RECT 51.575 2.553 51.775 2.865 ;
      RECT 51.65 2.531 51.775 2.865 ;
      RECT 51.59 2.55 51.78 2.85 ;
      RECT 51.56 2.561 51.78 2.848 ;
      RECT 51.575 2.556 51.785 2.814 ;
      RECT 51.56 2.66 51.79 2.781 ;
      RECT 51.59 2.532 51.775 2.865 ;
      RECT 51.65 2.51 51.75 2.865 ;
      RECT 51.675 2.507 51.75 2.865 ;
      RECT 51.675 2.502 51.695 2.865 ;
      RECT 51.08 2.57 51.255 2.745 ;
      RECT 51.075 2.57 51.255 2.743 ;
      RECT 51.05 2.57 51.255 2.738 ;
      RECT 50.995 2.55 51.165 2.728 ;
      RECT 50.995 2.557 51.23 2.728 ;
      RECT 51.08 3.237 51.095 3.42 ;
      RECT 51.07 3.215 51.08 3.42 ;
      RECT 51.055 3.195 51.07 3.42 ;
      RECT 51.045 3.17 51.055 3.42 ;
      RECT 51.015 3.135 51.045 3.42 ;
      RECT 50.98 3.075 51.015 3.42 ;
      RECT 50.975 3.037 50.98 3.42 ;
      RECT 50.925 2.988 50.975 3.42 ;
      RECT 50.915 2.938 50.925 3.408 ;
      RECT 50.9 2.917 50.915 3.368 ;
      RECT 50.88 2.885 50.9 3.318 ;
      RECT 50.855 2.841 50.88 3.258 ;
      RECT 50.85 2.813 50.855 3.213 ;
      RECT 50.845 2.804 50.85 3.199 ;
      RECT 50.84 2.797 50.845 3.186 ;
      RECT 50.835 2.792 50.84 3.175 ;
      RECT 50.83 2.777 50.835 3.165 ;
      RECT 50.825 2.755 50.83 3.152 ;
      RECT 50.815 2.715 50.825 3.127 ;
      RECT 50.79 2.645 50.815 3.083 ;
      RECT 50.785 2.585 50.79 3.048 ;
      RECT 50.77 2.565 50.785 3.015 ;
      RECT 50.765 2.565 50.77 2.99 ;
      RECT 50.735 2.565 50.765 2.945 ;
      RECT 50.69 2.565 50.735 2.885 ;
      RECT 50.615 2.565 50.69 2.833 ;
      RECT 50.61 2.565 50.615 2.798 ;
      RECT 50.605 2.565 50.61 2.788 ;
      RECT 50.6 2.565 50.605 2.768 ;
      RECT 50.865 1.785 51.035 2.255 ;
      RECT 50.81 1.778 51.005 2.239 ;
      RECT 50.81 1.792 51.04 2.238 ;
      RECT 50.795 1.793 51.04 2.219 ;
      RECT 50.79 1.811 51.04 2.205 ;
      RECT 50.795 1.794 51.045 2.203 ;
      RECT 50.78 1.825 51.045 2.188 ;
      RECT 50.795 1.8 51.05 2.173 ;
      RECT 50.775 1.84 51.05 2.17 ;
      RECT 50.79 1.812 51.055 2.155 ;
      RECT 50.79 1.824 51.06 2.135 ;
      RECT 50.775 1.84 51.065 2.118 ;
      RECT 50.775 1.85 51.07 1.973 ;
      RECT 50.77 1.85 51.07 1.93 ;
      RECT 50.77 1.865 51.075 1.908 ;
      RECT 50.865 1.775 51.005 2.255 ;
      RECT 50.865 1.773 50.975 2.255 ;
      RECT 50.951 1.77 50.975 2.255 ;
      RECT 50.61 3.437 50.615 3.483 ;
      RECT 50.6 3.285 50.61 3.507 ;
      RECT 50.595 3.13 50.6 3.532 ;
      RECT 50.58 3.092 50.595 3.543 ;
      RECT 50.575 3.075 50.58 3.55 ;
      RECT 50.565 3.063 50.575 3.557 ;
      RECT 50.56 3.054 50.565 3.559 ;
      RECT 50.555 3.052 50.56 3.563 ;
      RECT 50.51 3.043 50.555 3.578 ;
      RECT 50.505 3.035 50.51 3.592 ;
      RECT 50.5 3.032 50.505 3.596 ;
      RECT 50.485 3.027 50.5 3.604 ;
      RECT 50.43 3.017 50.485 3.615 ;
      RECT 50.395 3.005 50.43 3.616 ;
      RECT 50.386 3 50.395 3.61 ;
      RECT 50.3 3 50.386 3.6 ;
      RECT 50.27 3 50.3 3.578 ;
      RECT 50.26 3 50.265 3.558 ;
      RECT 50.255 3 50.26 3.52 ;
      RECT 50.25 3 50.255 3.478 ;
      RECT 50.245 3 50.25 3.438 ;
      RECT 50.24 3 50.245 3.368 ;
      RECT 50.23 3 50.24 3.29 ;
      RECT 50.225 3 50.23 3.19 ;
      RECT 50.265 3 50.27 3.56 ;
      RECT 49.76 3.082 49.85 3.56 ;
      RECT 49.745 3.085 49.865 3.558 ;
      RECT 49.76 3.084 49.865 3.558 ;
      RECT 49.725 3.091 49.89 3.548 ;
      RECT 49.745 3.085 49.89 3.548 ;
      RECT 49.71 3.097 49.89 3.536 ;
      RECT 49.745 3.088 49.94 3.529 ;
      RECT 49.696 3.105 49.94 3.527 ;
      RECT 49.725 3.095 49.95 3.515 ;
      RECT 49.696 3.116 49.98 3.506 ;
      RECT 49.61 3.14 49.98 3.5 ;
      RECT 49.61 3.153 50.02 3.483 ;
      RECT 49.605 3.175 50.02 3.476 ;
      RECT 49.575 3.19 50.02 3.466 ;
      RECT 49.57 3.201 50.02 3.456 ;
      RECT 49.54 3.214 50.02 3.447 ;
      RECT 49.525 3.232 50.02 3.436 ;
      RECT 49.5 3.245 50.02 3.426 ;
      RECT 49.76 3.081 49.77 3.56 ;
      RECT 49.806 2.505 49.845 2.75 ;
      RECT 49.72 2.505 49.855 2.748 ;
      RECT 49.605 2.53 49.855 2.745 ;
      RECT 49.605 2.53 49.86 2.743 ;
      RECT 49.605 2.53 49.875 2.738 ;
      RECT 49.711 2.505 49.89 2.718 ;
      RECT 49.625 2.513 49.89 2.718 ;
      RECT 49.295 1.865 49.465 2.3 ;
      RECT 49.285 1.899 49.465 2.283 ;
      RECT 49.365 1.835 49.535 2.27 ;
      RECT 49.27 1.91 49.535 2.248 ;
      RECT 49.365 1.845 49.54 2.238 ;
      RECT 49.295 1.897 49.57 2.223 ;
      RECT 49.255 1.923 49.57 2.208 ;
      RECT 49.255 1.965 49.58 2.188 ;
      RECT 49.25 1.99 49.585 2.17 ;
      RECT 49.25 2 49.59 2.155 ;
      RECT 49.245 1.937 49.57 2.153 ;
      RECT 49.245 2.01 49.595 2.138 ;
      RECT 49.24 1.947 49.57 2.135 ;
      RECT 49.235 2.031 49.6 2.118 ;
      RECT 49.235 2.063 49.605 2.098 ;
      RECT 49.23 1.977 49.58 2.09 ;
      RECT 49.235 1.962 49.57 2.118 ;
      RECT 49.25 1.932 49.57 2.17 ;
      RECT 49.095 2.519 49.32 2.775 ;
      RECT 49.095 2.552 49.34 2.765 ;
      RECT 49.06 2.552 49.34 2.763 ;
      RECT 49.06 2.565 49.345 2.753 ;
      RECT 49.06 2.585 49.355 2.745 ;
      RECT 49.06 2.682 49.36 2.738 ;
      RECT 49.04 2.43 49.17 2.728 ;
      RECT 48.995 2.585 49.355 2.67 ;
      RECT 48.985 2.43 49.17 2.615 ;
      RECT 48.985 2.462 49.256 2.615 ;
      RECT 48.95 2.992 48.97 3.17 ;
      RECT 48.915 2.945 48.95 3.17 ;
      RECT 48.9 2.885 48.915 3.17 ;
      RECT 48.875 2.832 48.9 3.17 ;
      RECT 48.86 2.785 48.875 3.17 ;
      RECT 48.84 2.762 48.86 3.17 ;
      RECT 48.815 2.727 48.84 3.17 ;
      RECT 48.805 2.573 48.815 3.17 ;
      RECT 48.775 2.568 48.805 3.161 ;
      RECT 48.77 2.565 48.775 3.151 ;
      RECT 48.755 2.565 48.77 3.125 ;
      RECT 48.75 2.565 48.755 3.088 ;
      RECT 48.725 2.565 48.75 3.04 ;
      RECT 48.705 2.565 48.725 2.965 ;
      RECT 48.695 2.565 48.705 2.925 ;
      RECT 48.69 2.565 48.695 2.9 ;
      RECT 48.685 2.565 48.69 2.883 ;
      RECT 48.68 2.565 48.685 2.865 ;
      RECT 48.675 2.566 48.68 2.855 ;
      RECT 48.665 2.568 48.675 2.823 ;
      RECT 48.655 2.57 48.665 2.79 ;
      RECT 48.645 2.573 48.655 2.763 ;
      RECT 48.97 3 49.195 3.17 ;
      RECT 48.3 1.812 48.47 2.265 ;
      RECT 48.3 1.812 48.56 2.231 ;
      RECT 48.3 1.812 48.59 2.215 ;
      RECT 48.3 1.812 48.62 2.188 ;
      RECT 48.556 1.79 48.635 2.17 ;
      RECT 48.335 1.797 48.64 2.155 ;
      RECT 48.335 1.805 48.65 2.118 ;
      RECT 48.295 1.832 48.65 2.09 ;
      RECT 48.28 1.845 48.65 2.055 ;
      RECT 48.3 1.82 48.67 2.045 ;
      RECT 48.275 1.885 48.67 2.015 ;
      RECT 48.275 1.915 48.675 1.998 ;
      RECT 48.27 1.945 48.675 1.985 ;
      RECT 48.335 1.794 48.635 2.17 ;
      RECT 48.47 1.791 48.556 2.249 ;
      RECT 48.421 1.792 48.635 2.17 ;
      RECT 48.565 3.452 48.61 3.645 ;
      RECT 48.555 3.422 48.565 3.645 ;
      RECT 48.55 3.407 48.555 3.645 ;
      RECT 48.51 3.317 48.55 3.645 ;
      RECT 48.505 3.23 48.51 3.645 ;
      RECT 48.495 3.2 48.505 3.645 ;
      RECT 48.49 3.16 48.495 3.645 ;
      RECT 48.48 3.122 48.49 3.645 ;
      RECT 48.475 3.087 48.48 3.645 ;
      RECT 48.455 3.04 48.475 3.645 ;
      RECT 48.44 2.965 48.455 3.645 ;
      RECT 48.435 2.92 48.44 3.64 ;
      RECT 48.43 2.9 48.435 3.613 ;
      RECT 48.425 2.88 48.43 3.598 ;
      RECT 48.42 2.855 48.425 3.578 ;
      RECT 48.415 2.833 48.42 3.563 ;
      RECT 48.41 2.811 48.415 3.545 ;
      RECT 48.405 2.79 48.41 3.535 ;
      RECT 48.395 2.762 48.405 3.505 ;
      RECT 48.385 2.725 48.395 3.473 ;
      RECT 48.375 2.685 48.385 3.44 ;
      RECT 48.365 2.663 48.375 3.41 ;
      RECT 48.335 2.615 48.365 3.342 ;
      RECT 48.32 2.575 48.335 3.269 ;
      RECT 48.31 2.575 48.32 3.235 ;
      RECT 48.305 2.575 48.31 3.21 ;
      RECT 48.3 2.575 48.305 3.195 ;
      RECT 48.295 2.575 48.3 3.173 ;
      RECT 48.29 2.575 48.295 3.16 ;
      RECT 48.275 2.575 48.29 3.125 ;
      RECT 48.255 2.575 48.275 3.065 ;
      RECT 48.245 2.575 48.255 3.015 ;
      RECT 48.225 2.575 48.245 2.963 ;
      RECT 48.205 2.575 48.225 2.92 ;
      RECT 48.195 2.575 48.205 2.908 ;
      RECT 48.165 2.575 48.195 2.895 ;
      RECT 48.135 2.596 48.165 2.875 ;
      RECT 48.125 2.624 48.135 2.855 ;
      RECT 48.11 2.641 48.125 2.823 ;
      RECT 48.105 2.655 48.11 2.79 ;
      RECT 48.1 2.663 48.105 2.763 ;
      RECT 48.095 2.671 48.1 2.725 ;
      RECT 48.1 3.195 48.105 3.53 ;
      RECT 48.065 3.182 48.1 3.529 ;
      RECT 47.995 3.122 48.065 3.528 ;
      RECT 47.915 3.065 47.995 3.527 ;
      RECT 47.78 3.025 47.915 3.526 ;
      RECT 47.78 3.212 48.115 3.515 ;
      RECT 47.74 3.212 48.115 3.505 ;
      RECT 47.74 3.23 48.12 3.5 ;
      RECT 47.74 3.32 48.125 3.49 ;
      RECT 47.735 3.015 47.9 3.47 ;
      RECT 47.73 3.015 47.9 3.213 ;
      RECT 47.73 3.172 48.095 3.213 ;
      RECT 47.73 3.16 48.09 3.213 ;
      RECT 46.495 1.74 46.665 2.935 ;
      RECT 46.495 1.74 46.96 1.91 ;
      RECT 46.495 6.97 46.96 7.14 ;
      RECT 46.495 5.945 46.665 7.14 ;
      RECT 45.505 1.74 45.675 2.935 ;
      RECT 45.505 1.74 45.97 1.91 ;
      RECT 45.505 6.97 45.97 7.14 ;
      RECT 45.505 5.945 45.675 7.14 ;
      RECT 43.65 2.635 43.82 3.865 ;
      RECT 43.705 0.855 43.875 2.805 ;
      RECT 43.65 0.575 43.82 1.025 ;
      RECT 43.65 7.855 43.82 8.305 ;
      RECT 43.705 6.075 43.875 8.025 ;
      RECT 43.65 5.015 43.82 6.245 ;
      RECT 43.13 0.575 43.3 3.865 ;
      RECT 43.13 2.075 43.535 2.405 ;
      RECT 43.13 1.235 43.535 1.565 ;
      RECT 43.13 5.015 43.3 8.305 ;
      RECT 43.13 7.315 43.535 7.645 ;
      RECT 43.13 6.475 43.535 6.805 ;
      RECT 40.465 1.975 41.195 2.215 ;
      RECT 41.007 1.77 41.195 2.215 ;
      RECT 40.835 1.782 41.21 2.209 ;
      RECT 40.75 1.797 41.23 2.194 ;
      RECT 40.75 1.812 41.235 2.184 ;
      RECT 40.705 1.832 41.25 2.176 ;
      RECT 40.682 1.867 41.265 2.13 ;
      RECT 40.596 1.89 41.27 2.09 ;
      RECT 40.596 1.908 41.28 2.06 ;
      RECT 40.465 1.977 41.285 2.023 ;
      RECT 40.51 1.92 41.28 2.06 ;
      RECT 40.596 1.872 41.265 2.13 ;
      RECT 40.682 1.841 41.25 2.176 ;
      RECT 40.705 1.822 41.235 2.184 ;
      RECT 40.75 1.795 41.21 2.209 ;
      RECT 40.835 1.777 41.195 2.215 ;
      RECT 40.921 1.771 41.195 2.215 ;
      RECT 41.007 1.766 41.14 2.215 ;
      RECT 41.093 1.761 41.14 2.215 ;
      RECT 40.785 2.659 40.955 3.045 ;
      RECT 40.78 2.659 40.955 3.04 ;
      RECT 40.755 2.659 40.955 3.005 ;
      RECT 40.755 2.687 40.965 2.995 ;
      RECT 40.735 2.687 40.965 2.955 ;
      RECT 40.73 2.687 40.965 2.928 ;
      RECT 40.73 2.705 40.97 2.92 ;
      RECT 40.675 2.705 40.97 2.855 ;
      RECT 40.675 2.722 40.98 2.838 ;
      RECT 40.665 2.722 40.98 2.778 ;
      RECT 40.665 2.739 40.985 2.775 ;
      RECT 40.66 2.575 40.83 2.753 ;
      RECT 40.66 2.609 40.916 2.753 ;
      RECT 40.655 3.375 40.66 3.388 ;
      RECT 40.65 3.27 40.655 3.393 ;
      RECT 40.625 3.13 40.65 3.408 ;
      RECT 40.59 3.081 40.625 3.44 ;
      RECT 40.585 3.049 40.59 3.46 ;
      RECT 40.58 3.04 40.585 3.46 ;
      RECT 40.5 3.005 40.58 3.46 ;
      RECT 40.437 2.975 40.5 3.46 ;
      RECT 40.351 2.963 40.437 3.46 ;
      RECT 40.265 2.949 40.351 3.46 ;
      RECT 40.185 2.936 40.265 3.446 ;
      RECT 40.15 2.928 40.185 3.426 ;
      RECT 40.14 2.925 40.15 3.417 ;
      RECT 40.11 2.92 40.14 3.404 ;
      RECT 40.06 2.895 40.11 3.38 ;
      RECT 40.046 2.869 40.06 3.362 ;
      RECT 39.96 2.829 40.046 3.338 ;
      RECT 39.915 2.777 39.96 3.307 ;
      RECT 39.905 2.752 39.915 3.294 ;
      RECT 39.9 2.533 39.905 2.555 ;
      RECT 39.895 2.735 39.905 3.29 ;
      RECT 39.895 2.531 39.9 2.645 ;
      RECT 39.885 2.527 39.895 3.286 ;
      RECT 39.841 2.525 39.885 3.274 ;
      RECT 39.755 2.525 39.841 3.245 ;
      RECT 39.725 2.525 39.755 3.218 ;
      RECT 39.71 2.525 39.725 3.206 ;
      RECT 39.67 2.537 39.71 3.191 ;
      RECT 39.65 2.556 39.67 3.17 ;
      RECT 39.64 2.566 39.65 3.154 ;
      RECT 39.63 2.572 39.64 3.143 ;
      RECT 39.61 2.582 39.63 3.126 ;
      RECT 39.605 2.591 39.61 3.113 ;
      RECT 39.6 2.595 39.605 3.063 ;
      RECT 39.59 2.601 39.6 2.98 ;
      RECT 39.585 2.605 39.59 2.894 ;
      RECT 39.58 2.625 39.585 2.831 ;
      RECT 39.575 2.648 39.58 2.778 ;
      RECT 39.57 2.666 39.575 2.723 ;
      RECT 40.18 2.485 40.35 2.745 ;
      RECT 40.35 2.45 40.395 2.731 ;
      RECT 40.311 2.452 40.4 2.714 ;
      RECT 40.2 2.469 40.486 2.685 ;
      RECT 40.2 2.484 40.49 2.657 ;
      RECT 40.2 2.465 40.4 2.714 ;
      RECT 40.225 2.453 40.35 2.745 ;
      RECT 40.311 2.451 40.395 2.731 ;
      RECT 39.365 1.84 39.535 2.33 ;
      RECT 39.365 1.84 39.57 2.31 ;
      RECT 39.5 1.76 39.61 2.27 ;
      RECT 39.481 1.764 39.63 2.24 ;
      RECT 39.395 1.772 39.65 2.223 ;
      RECT 39.395 1.778 39.655 2.213 ;
      RECT 39.395 1.787 39.675 2.201 ;
      RECT 39.37 1.812 39.705 2.179 ;
      RECT 39.37 1.832 39.71 2.159 ;
      RECT 39.365 1.845 39.72 2.139 ;
      RECT 39.365 1.912 39.725 2.12 ;
      RECT 39.365 2.045 39.73 2.107 ;
      RECT 39.36 1.85 39.72 1.94 ;
      RECT 39.37 1.807 39.675 2.201 ;
      RECT 39.481 1.762 39.61 2.27 ;
      RECT 39.355 3.515 39.655 3.77 ;
      RECT 39.44 3.481 39.655 3.77 ;
      RECT 39.44 3.484 39.66 3.63 ;
      RECT 39.375 3.505 39.66 3.63 ;
      RECT 39.41 3.495 39.655 3.77 ;
      RECT 39.405 3.5 39.66 3.63 ;
      RECT 39.44 3.479 39.641 3.77 ;
      RECT 39.526 3.47 39.641 3.77 ;
      RECT 39.526 3.464 39.555 3.77 ;
      RECT 39.015 3.105 39.025 3.595 ;
      RECT 38.675 3.04 38.685 3.34 ;
      RECT 39.19 3.212 39.195 3.431 ;
      RECT 39.18 3.192 39.19 3.448 ;
      RECT 39.17 3.172 39.18 3.478 ;
      RECT 39.165 3.162 39.17 3.493 ;
      RECT 39.16 3.158 39.165 3.498 ;
      RECT 39.145 3.15 39.16 3.505 ;
      RECT 39.105 3.13 39.145 3.53 ;
      RECT 39.08 3.112 39.105 3.563 ;
      RECT 39.075 3.11 39.08 3.576 ;
      RECT 39.055 3.107 39.075 3.58 ;
      RECT 39.025 3.105 39.055 3.59 ;
      RECT 38.955 3.107 39.015 3.591 ;
      RECT 38.935 3.107 38.955 3.585 ;
      RECT 38.91 3.105 38.935 3.582 ;
      RECT 38.875 3.1 38.91 3.578 ;
      RECT 38.855 3.094 38.875 3.565 ;
      RECT 38.845 3.091 38.855 3.553 ;
      RECT 38.825 3.088 38.845 3.538 ;
      RECT 38.805 3.084 38.825 3.52 ;
      RECT 38.8 3.081 38.805 3.51 ;
      RECT 38.795 3.08 38.8 3.508 ;
      RECT 38.785 3.077 38.795 3.5 ;
      RECT 38.775 3.071 38.785 3.483 ;
      RECT 38.765 3.065 38.775 3.465 ;
      RECT 38.755 3.059 38.765 3.453 ;
      RECT 38.745 3.053 38.755 3.433 ;
      RECT 38.74 3.049 38.745 3.418 ;
      RECT 38.735 3.047 38.74 3.41 ;
      RECT 38.73 3.045 38.735 3.403 ;
      RECT 38.725 3.043 38.73 3.393 ;
      RECT 38.72 3.041 38.725 3.387 ;
      RECT 38.71 3.04 38.72 3.377 ;
      RECT 38.7 3.04 38.71 3.368 ;
      RECT 38.685 3.04 38.7 3.353 ;
      RECT 38.645 3.04 38.675 3.337 ;
      RECT 38.625 3.042 38.645 3.332 ;
      RECT 38.62 3.047 38.625 3.33 ;
      RECT 38.59 3.055 38.62 3.328 ;
      RECT 38.56 3.07 38.59 3.327 ;
      RECT 38.515 3.092 38.56 3.332 ;
      RECT 38.51 3.107 38.515 3.336 ;
      RECT 38.495 3.112 38.51 3.338 ;
      RECT 38.49 3.116 38.495 3.34 ;
      RECT 38.43 3.139 38.49 3.349 ;
      RECT 38.41 3.165 38.43 3.362 ;
      RECT 38.4 3.172 38.41 3.366 ;
      RECT 38.385 3.179 38.4 3.369 ;
      RECT 38.365 3.189 38.385 3.372 ;
      RECT 38.36 3.197 38.365 3.375 ;
      RECT 38.315 3.202 38.36 3.382 ;
      RECT 38.305 3.205 38.315 3.389 ;
      RECT 38.295 3.205 38.305 3.393 ;
      RECT 38.26 3.207 38.295 3.405 ;
      RECT 38.24 3.21 38.26 3.418 ;
      RECT 38.2 3.213 38.24 3.429 ;
      RECT 38.185 3.215 38.2 3.442 ;
      RECT 38.175 3.215 38.185 3.447 ;
      RECT 38.15 3.216 38.175 3.455 ;
      RECT 38.14 3.218 38.15 3.46 ;
      RECT 38.135 3.219 38.14 3.463 ;
      RECT 38.11 3.217 38.135 3.466 ;
      RECT 38.095 3.215 38.11 3.467 ;
      RECT 38.075 3.212 38.095 3.469 ;
      RECT 38.055 3.207 38.075 3.469 ;
      RECT 37.995 3.202 38.055 3.466 ;
      RECT 37.96 3.177 37.995 3.462 ;
      RECT 37.95 3.154 37.96 3.46 ;
      RECT 37.92 3.131 37.95 3.46 ;
      RECT 37.91 3.11 37.92 3.46 ;
      RECT 37.885 3.092 37.91 3.458 ;
      RECT 37.87 3.07 37.885 3.455 ;
      RECT 37.855 3.052 37.87 3.453 ;
      RECT 37.835 3.042 37.855 3.451 ;
      RECT 37.82 3.037 37.835 3.45 ;
      RECT 37.805 3.035 37.82 3.449 ;
      RECT 37.775 3.036 37.805 3.447 ;
      RECT 37.755 3.039 37.775 3.445 ;
      RECT 37.698 3.043 37.755 3.445 ;
      RECT 37.612 3.052 37.698 3.445 ;
      RECT 37.526 3.063 37.612 3.445 ;
      RECT 37.44 3.074 37.526 3.445 ;
      RECT 37.42 3.081 37.44 3.453 ;
      RECT 37.41 3.084 37.42 3.46 ;
      RECT 37.345 3.089 37.41 3.478 ;
      RECT 37.315 3.096 37.345 3.503 ;
      RECT 37.305 3.099 37.315 3.51 ;
      RECT 37.26 3.103 37.305 3.515 ;
      RECT 37.23 3.108 37.26 3.52 ;
      RECT 37.229 3.11 37.23 3.52 ;
      RECT 37.143 3.116 37.229 3.52 ;
      RECT 37.057 3.127 37.143 3.52 ;
      RECT 36.971 3.139 37.057 3.52 ;
      RECT 36.885 3.15 36.971 3.52 ;
      RECT 36.87 3.157 36.885 3.515 ;
      RECT 36.865 3.159 36.87 3.509 ;
      RECT 36.845 3.17 36.865 3.504 ;
      RECT 36.835 3.188 36.845 3.498 ;
      RECT 36.83 3.2 36.835 3.298 ;
      RECT 39.125 1.953 39.145 2.04 ;
      RECT 39.12 1.888 39.125 2.072 ;
      RECT 39.11 1.855 39.12 2.077 ;
      RECT 39.105 1.835 39.11 2.083 ;
      RECT 39.075 1.835 39.105 2.1 ;
      RECT 39.026 1.835 39.075 2.136 ;
      RECT 38.94 1.835 39.026 2.194 ;
      RECT 38.911 1.845 38.94 2.243 ;
      RECT 38.825 1.887 38.911 2.296 ;
      RECT 38.805 1.925 38.825 2.343 ;
      RECT 38.78 1.942 38.805 2.363 ;
      RECT 38.77 1.956 38.78 2.383 ;
      RECT 38.765 1.962 38.77 2.393 ;
      RECT 38.76 1.966 38.765 2.4 ;
      RECT 38.71 1.986 38.76 2.405 ;
      RECT 38.645 2.03 38.71 2.405 ;
      RECT 38.62 2.08 38.645 2.405 ;
      RECT 38.61 2.11 38.62 2.405 ;
      RECT 38.605 2.137 38.61 2.405 ;
      RECT 38.6 2.155 38.605 2.405 ;
      RECT 38.59 2.197 38.6 2.405 ;
      RECT 38.94 2.755 39.11 2.93 ;
      RECT 38.88 2.583 38.94 2.918 ;
      RECT 38.87 2.576 38.88 2.901 ;
      RECT 38.825 2.755 39.11 2.881 ;
      RECT 38.806 2.755 39.11 2.859 ;
      RECT 38.72 2.755 39.11 2.824 ;
      RECT 38.7 2.575 38.87 2.78 ;
      RECT 38.7 2.722 39.105 2.78 ;
      RECT 38.7 2.67 39.08 2.78 ;
      RECT 38.7 2.625 39.045 2.78 ;
      RECT 38.7 2.607 39.01 2.78 ;
      RECT 38.7 2.597 39.005 2.78 ;
      RECT 38.87 7.855 39.04 8.305 ;
      RECT 38.925 6.075 39.095 8.025 ;
      RECT 38.87 5.015 39.04 6.245 ;
      RECT 38.35 5.015 38.52 8.305 ;
      RECT 38.35 7.315 38.755 7.645 ;
      RECT 38.35 6.475 38.755 6.805 ;
      RECT 38.42 3.555 38.61 3.78 ;
      RECT 38.41 3.556 38.615 3.775 ;
      RECT 38.41 3.558 38.625 3.755 ;
      RECT 38.41 3.562 38.63 3.74 ;
      RECT 38.41 3.549 38.58 3.775 ;
      RECT 38.41 3.552 38.605 3.775 ;
      RECT 38.42 3.548 38.58 3.78 ;
      RECT 38.506 3.546 38.58 3.78 ;
      RECT 38.13 2.797 38.3 3.035 ;
      RECT 38.13 2.797 38.386 2.949 ;
      RECT 38.13 2.797 38.39 2.859 ;
      RECT 38.18 2.57 38.4 2.838 ;
      RECT 38.175 2.587 38.405 2.811 ;
      RECT 38.14 2.745 38.405 2.811 ;
      RECT 38.16 2.595 38.3 3.035 ;
      RECT 38.15 2.677 38.41 2.794 ;
      RECT 38.145 2.725 38.41 2.794 ;
      RECT 38.15 2.635 38.405 2.811 ;
      RECT 38.175 2.572 38.4 2.838 ;
      RECT 37.74 2.547 37.91 2.745 ;
      RECT 37.74 2.547 37.955 2.72 ;
      RECT 37.81 2.49 37.98 2.678 ;
      RECT 37.785 2.505 37.98 2.678 ;
      RECT 37.4 2.551 37.43 2.745 ;
      RECT 37.395 2.523 37.4 2.745 ;
      RECT 37.365 2.497 37.395 2.747 ;
      RECT 37.34 2.455 37.365 2.75 ;
      RECT 37.33 2.427 37.34 2.752 ;
      RECT 37.295 2.407 37.33 2.754 ;
      RECT 37.23 2.392 37.295 2.76 ;
      RECT 37.18 2.39 37.23 2.766 ;
      RECT 37.157 2.392 37.18 2.771 ;
      RECT 37.071 2.403 37.157 2.777 ;
      RECT 36.985 2.421 37.071 2.787 ;
      RECT 36.97 2.432 36.985 2.793 ;
      RECT 36.9 2.455 36.97 2.799 ;
      RECT 36.845 2.487 36.9 2.807 ;
      RECT 36.805 2.51 36.845 2.813 ;
      RECT 36.791 2.523 36.805 2.816 ;
      RECT 36.705 2.545 36.791 2.822 ;
      RECT 36.69 2.57 36.705 2.828 ;
      RECT 36.65 2.585 36.69 2.832 ;
      RECT 36.6 2.6 36.65 2.837 ;
      RECT 36.575 2.607 36.6 2.841 ;
      RECT 36.515 2.602 36.575 2.845 ;
      RECT 36.5 2.593 36.515 2.849 ;
      RECT 36.43 2.583 36.5 2.845 ;
      RECT 36.405 2.575 36.425 2.835 ;
      RECT 36.346 2.575 36.405 2.813 ;
      RECT 36.26 2.575 36.346 2.77 ;
      RECT 36.425 2.575 36.43 2.84 ;
      RECT 37.12 1.806 37.29 2.14 ;
      RECT 37.09 1.806 37.29 2.135 ;
      RECT 37.03 1.773 37.09 2.123 ;
      RECT 37.03 1.829 37.3 2.118 ;
      RECT 37.005 1.829 37.3 2.112 ;
      RECT 37 1.77 37.03 2.109 ;
      RECT 36.985 1.776 37.12 2.107 ;
      RECT 36.98 1.784 37.205 2.095 ;
      RECT 36.98 1.836 37.315 2.048 ;
      RECT 36.965 1.792 37.205 2.043 ;
      RECT 36.965 1.862 37.325 1.984 ;
      RECT 36.935 1.812 37.29 1.945 ;
      RECT 36.935 1.902 37.335 1.941 ;
      RECT 36.985 1.781 37.205 2.107 ;
      RECT 36.325 2.111 36.38 2.375 ;
      RECT 36.325 2.111 36.445 2.374 ;
      RECT 36.325 2.111 36.47 2.373 ;
      RECT 36.325 2.111 36.535 2.372 ;
      RECT 36.47 2.077 36.55 2.371 ;
      RECT 36.285 2.121 36.695 2.37 ;
      RECT 36.325 2.118 36.695 2.37 ;
      RECT 36.285 2.126 36.7 2.363 ;
      RECT 36.27 2.128 36.7 2.362 ;
      RECT 36.27 2.135 36.705 2.358 ;
      RECT 36.25 2.134 36.7 2.354 ;
      RECT 36.25 2.142 36.71 2.353 ;
      RECT 36.245 2.139 36.705 2.349 ;
      RECT 36.245 2.152 36.72 2.348 ;
      RECT 36.23 2.142 36.71 2.347 ;
      RECT 36.195 2.155 36.72 2.34 ;
      RECT 36.38 2.11 36.69 2.37 ;
      RECT 36.38 2.095 36.64 2.37 ;
      RECT 36.445 2.082 36.575 2.37 ;
      RECT 35.99 3.171 36.005 3.564 ;
      RECT 35.955 3.176 36.005 3.563 ;
      RECT 35.99 3.175 36.05 3.562 ;
      RECT 35.935 3.186 36.05 3.561 ;
      RECT 35.95 3.182 36.05 3.561 ;
      RECT 35.915 3.192 36.125 3.558 ;
      RECT 35.915 3.211 36.17 3.556 ;
      RECT 35.915 3.218 36.175 3.553 ;
      RECT 35.9 3.195 36.125 3.55 ;
      RECT 35.88 3.2 36.125 3.543 ;
      RECT 35.875 3.204 36.125 3.539 ;
      RECT 35.875 3.221 36.185 3.538 ;
      RECT 35.855 3.215 36.17 3.534 ;
      RECT 35.855 3.224 36.19 3.528 ;
      RECT 35.85 3.23 36.19 3.3 ;
      RECT 35.915 3.19 36.05 3.558 ;
      RECT 35.79 2.553 35.99 2.865 ;
      RECT 35.865 2.531 35.99 2.865 ;
      RECT 35.805 2.55 35.995 2.85 ;
      RECT 35.775 2.561 35.995 2.848 ;
      RECT 35.79 2.556 36 2.814 ;
      RECT 35.775 2.66 36.005 2.781 ;
      RECT 35.805 2.532 35.99 2.865 ;
      RECT 35.865 2.51 35.965 2.865 ;
      RECT 35.89 2.507 35.965 2.865 ;
      RECT 35.89 2.502 35.91 2.865 ;
      RECT 35.295 2.57 35.47 2.745 ;
      RECT 35.29 2.57 35.47 2.743 ;
      RECT 35.265 2.57 35.47 2.738 ;
      RECT 35.21 2.55 35.38 2.728 ;
      RECT 35.21 2.557 35.445 2.728 ;
      RECT 35.295 3.237 35.31 3.42 ;
      RECT 35.285 3.215 35.295 3.42 ;
      RECT 35.27 3.195 35.285 3.42 ;
      RECT 35.26 3.17 35.27 3.42 ;
      RECT 35.23 3.135 35.26 3.42 ;
      RECT 35.195 3.075 35.23 3.42 ;
      RECT 35.19 3.037 35.195 3.42 ;
      RECT 35.14 2.988 35.19 3.42 ;
      RECT 35.13 2.938 35.14 3.408 ;
      RECT 35.115 2.917 35.13 3.368 ;
      RECT 35.095 2.885 35.115 3.318 ;
      RECT 35.07 2.841 35.095 3.258 ;
      RECT 35.065 2.813 35.07 3.213 ;
      RECT 35.06 2.804 35.065 3.199 ;
      RECT 35.055 2.797 35.06 3.186 ;
      RECT 35.05 2.792 35.055 3.175 ;
      RECT 35.045 2.777 35.05 3.165 ;
      RECT 35.04 2.755 35.045 3.152 ;
      RECT 35.03 2.715 35.04 3.127 ;
      RECT 35.005 2.645 35.03 3.083 ;
      RECT 35 2.585 35.005 3.048 ;
      RECT 34.985 2.565 35 3.015 ;
      RECT 34.98 2.565 34.985 2.99 ;
      RECT 34.95 2.565 34.98 2.945 ;
      RECT 34.905 2.565 34.95 2.885 ;
      RECT 34.83 2.565 34.905 2.833 ;
      RECT 34.825 2.565 34.83 2.798 ;
      RECT 34.82 2.565 34.825 2.788 ;
      RECT 34.815 2.565 34.82 2.768 ;
      RECT 35.08 1.785 35.25 2.255 ;
      RECT 35.025 1.778 35.22 2.239 ;
      RECT 35.025 1.792 35.255 2.238 ;
      RECT 35.01 1.793 35.255 2.219 ;
      RECT 35.005 1.811 35.255 2.205 ;
      RECT 35.01 1.794 35.26 2.203 ;
      RECT 34.995 1.825 35.26 2.188 ;
      RECT 35.01 1.8 35.265 2.173 ;
      RECT 34.99 1.84 35.265 2.17 ;
      RECT 35.005 1.812 35.27 2.155 ;
      RECT 35.005 1.824 35.275 2.135 ;
      RECT 34.99 1.84 35.28 2.118 ;
      RECT 34.99 1.85 35.285 1.973 ;
      RECT 34.985 1.85 35.285 1.93 ;
      RECT 34.985 1.865 35.29 1.908 ;
      RECT 35.08 1.775 35.22 2.255 ;
      RECT 35.08 1.773 35.19 2.255 ;
      RECT 35.166 1.77 35.19 2.255 ;
      RECT 34.825 3.437 34.83 3.483 ;
      RECT 34.815 3.285 34.825 3.507 ;
      RECT 34.81 3.13 34.815 3.532 ;
      RECT 34.795 3.092 34.81 3.543 ;
      RECT 34.79 3.075 34.795 3.55 ;
      RECT 34.78 3.063 34.79 3.557 ;
      RECT 34.775 3.054 34.78 3.559 ;
      RECT 34.77 3.052 34.775 3.563 ;
      RECT 34.725 3.043 34.77 3.578 ;
      RECT 34.72 3.035 34.725 3.592 ;
      RECT 34.715 3.032 34.72 3.596 ;
      RECT 34.7 3.027 34.715 3.604 ;
      RECT 34.645 3.017 34.7 3.615 ;
      RECT 34.61 3.005 34.645 3.616 ;
      RECT 34.601 3 34.61 3.61 ;
      RECT 34.515 3 34.601 3.6 ;
      RECT 34.485 3 34.515 3.578 ;
      RECT 34.475 3 34.48 3.558 ;
      RECT 34.47 3 34.475 3.52 ;
      RECT 34.465 3 34.47 3.478 ;
      RECT 34.46 3 34.465 3.438 ;
      RECT 34.455 3 34.46 3.368 ;
      RECT 34.445 3 34.455 3.29 ;
      RECT 34.44 3 34.445 3.19 ;
      RECT 34.48 3 34.485 3.56 ;
      RECT 33.975 3.082 34.065 3.56 ;
      RECT 33.96 3.085 34.08 3.558 ;
      RECT 33.975 3.084 34.08 3.558 ;
      RECT 33.94 3.091 34.105 3.548 ;
      RECT 33.96 3.085 34.105 3.548 ;
      RECT 33.925 3.097 34.105 3.536 ;
      RECT 33.96 3.088 34.155 3.529 ;
      RECT 33.911 3.105 34.155 3.527 ;
      RECT 33.94 3.095 34.165 3.515 ;
      RECT 33.911 3.116 34.195 3.506 ;
      RECT 33.825 3.14 34.195 3.5 ;
      RECT 33.825 3.153 34.235 3.483 ;
      RECT 33.82 3.175 34.235 3.476 ;
      RECT 33.79 3.19 34.235 3.466 ;
      RECT 33.785 3.201 34.235 3.456 ;
      RECT 33.755 3.214 34.235 3.447 ;
      RECT 33.74 3.232 34.235 3.436 ;
      RECT 33.715 3.245 34.235 3.426 ;
      RECT 33.975 3.081 33.985 3.56 ;
      RECT 34.021 2.505 34.06 2.75 ;
      RECT 33.935 2.505 34.07 2.748 ;
      RECT 33.82 2.53 34.07 2.745 ;
      RECT 33.82 2.53 34.075 2.743 ;
      RECT 33.82 2.53 34.09 2.738 ;
      RECT 33.926 2.505 34.105 2.718 ;
      RECT 33.84 2.513 34.105 2.718 ;
      RECT 33.51 1.865 33.68 2.3 ;
      RECT 33.5 1.899 33.68 2.283 ;
      RECT 33.58 1.835 33.75 2.27 ;
      RECT 33.485 1.91 33.75 2.248 ;
      RECT 33.58 1.845 33.755 2.238 ;
      RECT 33.51 1.897 33.785 2.223 ;
      RECT 33.47 1.923 33.785 2.208 ;
      RECT 33.47 1.965 33.795 2.188 ;
      RECT 33.465 1.99 33.8 2.17 ;
      RECT 33.465 2 33.805 2.155 ;
      RECT 33.46 1.937 33.785 2.153 ;
      RECT 33.46 2.01 33.81 2.138 ;
      RECT 33.455 1.947 33.785 2.135 ;
      RECT 33.45 2.031 33.815 2.118 ;
      RECT 33.45 2.063 33.82 2.098 ;
      RECT 33.445 1.977 33.795 2.09 ;
      RECT 33.45 1.962 33.785 2.118 ;
      RECT 33.465 1.932 33.785 2.17 ;
      RECT 33.31 2.519 33.535 2.775 ;
      RECT 33.31 2.552 33.555 2.765 ;
      RECT 33.275 2.552 33.555 2.763 ;
      RECT 33.275 2.565 33.56 2.753 ;
      RECT 33.275 2.585 33.57 2.745 ;
      RECT 33.275 2.682 33.575 2.738 ;
      RECT 33.255 2.43 33.385 2.728 ;
      RECT 33.21 2.585 33.57 2.67 ;
      RECT 33.2 2.43 33.385 2.615 ;
      RECT 33.2 2.462 33.471 2.615 ;
      RECT 33.165 2.992 33.185 3.17 ;
      RECT 33.13 2.945 33.165 3.17 ;
      RECT 33.115 2.885 33.13 3.17 ;
      RECT 33.09 2.832 33.115 3.17 ;
      RECT 33.075 2.785 33.09 3.17 ;
      RECT 33.055 2.762 33.075 3.17 ;
      RECT 33.03 2.727 33.055 3.17 ;
      RECT 33.02 2.573 33.03 3.17 ;
      RECT 32.99 2.568 33.02 3.161 ;
      RECT 32.985 2.565 32.99 3.151 ;
      RECT 32.97 2.565 32.985 3.125 ;
      RECT 32.965 2.565 32.97 3.088 ;
      RECT 32.94 2.565 32.965 3.04 ;
      RECT 32.92 2.565 32.94 2.965 ;
      RECT 32.91 2.565 32.92 2.925 ;
      RECT 32.905 2.565 32.91 2.9 ;
      RECT 32.9 2.565 32.905 2.883 ;
      RECT 32.895 2.565 32.9 2.865 ;
      RECT 32.89 2.566 32.895 2.855 ;
      RECT 32.88 2.568 32.89 2.823 ;
      RECT 32.87 2.57 32.88 2.79 ;
      RECT 32.86 2.573 32.87 2.763 ;
      RECT 33.185 3 33.41 3.17 ;
      RECT 32.515 1.812 32.685 2.265 ;
      RECT 32.515 1.812 32.775 2.231 ;
      RECT 32.515 1.812 32.805 2.215 ;
      RECT 32.515 1.812 32.835 2.188 ;
      RECT 32.771 1.79 32.85 2.17 ;
      RECT 32.55 1.797 32.855 2.155 ;
      RECT 32.55 1.805 32.865 2.118 ;
      RECT 32.51 1.832 32.865 2.09 ;
      RECT 32.495 1.845 32.865 2.055 ;
      RECT 32.515 1.82 32.885 2.045 ;
      RECT 32.49 1.885 32.885 2.015 ;
      RECT 32.49 1.915 32.89 1.998 ;
      RECT 32.485 1.945 32.89 1.985 ;
      RECT 32.55 1.794 32.85 2.17 ;
      RECT 32.685 1.791 32.771 2.249 ;
      RECT 32.636 1.792 32.85 2.17 ;
      RECT 32.78 3.452 32.825 3.645 ;
      RECT 32.77 3.422 32.78 3.645 ;
      RECT 32.765 3.407 32.77 3.645 ;
      RECT 32.725 3.317 32.765 3.645 ;
      RECT 32.72 3.23 32.725 3.645 ;
      RECT 32.71 3.2 32.72 3.645 ;
      RECT 32.705 3.16 32.71 3.645 ;
      RECT 32.695 3.122 32.705 3.645 ;
      RECT 32.69 3.087 32.695 3.645 ;
      RECT 32.67 3.04 32.69 3.645 ;
      RECT 32.655 2.965 32.67 3.645 ;
      RECT 32.65 2.92 32.655 3.64 ;
      RECT 32.645 2.9 32.65 3.613 ;
      RECT 32.64 2.88 32.645 3.598 ;
      RECT 32.635 2.855 32.64 3.578 ;
      RECT 32.63 2.833 32.635 3.563 ;
      RECT 32.625 2.811 32.63 3.545 ;
      RECT 32.62 2.79 32.625 3.535 ;
      RECT 32.61 2.762 32.62 3.505 ;
      RECT 32.6 2.725 32.61 3.473 ;
      RECT 32.59 2.685 32.6 3.44 ;
      RECT 32.58 2.663 32.59 3.41 ;
      RECT 32.55 2.615 32.58 3.342 ;
      RECT 32.535 2.575 32.55 3.269 ;
      RECT 32.525 2.575 32.535 3.235 ;
      RECT 32.52 2.575 32.525 3.21 ;
      RECT 32.515 2.575 32.52 3.195 ;
      RECT 32.51 2.575 32.515 3.173 ;
      RECT 32.505 2.575 32.51 3.16 ;
      RECT 32.49 2.575 32.505 3.125 ;
      RECT 32.47 2.575 32.49 3.065 ;
      RECT 32.46 2.575 32.47 3.015 ;
      RECT 32.44 2.575 32.46 2.963 ;
      RECT 32.42 2.575 32.44 2.92 ;
      RECT 32.41 2.575 32.42 2.908 ;
      RECT 32.38 2.575 32.41 2.895 ;
      RECT 32.35 2.596 32.38 2.875 ;
      RECT 32.34 2.624 32.35 2.855 ;
      RECT 32.325 2.641 32.34 2.823 ;
      RECT 32.32 2.655 32.325 2.79 ;
      RECT 32.315 2.663 32.32 2.763 ;
      RECT 32.31 2.671 32.315 2.725 ;
      RECT 32.315 3.195 32.32 3.53 ;
      RECT 32.28 3.182 32.315 3.529 ;
      RECT 32.21 3.122 32.28 3.528 ;
      RECT 32.13 3.065 32.21 3.527 ;
      RECT 31.995 3.025 32.13 3.526 ;
      RECT 31.995 3.212 32.33 3.515 ;
      RECT 31.955 3.212 32.33 3.505 ;
      RECT 31.955 3.23 32.335 3.5 ;
      RECT 31.955 3.32 32.34 3.49 ;
      RECT 31.95 3.015 32.115 3.47 ;
      RECT 31.945 3.015 32.115 3.213 ;
      RECT 31.945 3.172 32.31 3.213 ;
      RECT 31.945 3.16 32.305 3.213 ;
      RECT 30.72 1.74 30.89 2.935 ;
      RECT 30.72 1.74 31.185 1.91 ;
      RECT 30.72 6.97 31.185 7.14 ;
      RECT 30.72 5.945 30.89 7.14 ;
      RECT 29.73 1.74 29.9 2.935 ;
      RECT 29.73 1.74 30.195 1.91 ;
      RECT 29.73 6.97 30.195 7.14 ;
      RECT 29.73 5.945 29.9 7.14 ;
      RECT 27.875 2.635 28.045 3.865 ;
      RECT 27.93 0.855 28.1 2.805 ;
      RECT 27.875 0.575 28.045 1.025 ;
      RECT 27.875 7.855 28.045 8.305 ;
      RECT 27.93 6.075 28.1 8.025 ;
      RECT 27.875 5.015 28.045 6.245 ;
      RECT 27.355 0.575 27.525 3.865 ;
      RECT 27.355 2.075 27.76 2.405 ;
      RECT 27.355 1.235 27.76 1.565 ;
      RECT 27.355 5.015 27.525 8.305 ;
      RECT 27.355 7.315 27.76 7.645 ;
      RECT 27.355 6.475 27.76 6.805 ;
      RECT 24.69 1.975 25.42 2.215 ;
      RECT 25.232 1.77 25.42 2.215 ;
      RECT 25.06 1.782 25.435 2.209 ;
      RECT 24.975 1.797 25.455 2.194 ;
      RECT 24.975 1.812 25.46 2.184 ;
      RECT 24.93 1.832 25.475 2.176 ;
      RECT 24.907 1.867 25.49 2.13 ;
      RECT 24.821 1.89 25.495 2.09 ;
      RECT 24.821 1.908 25.505 2.06 ;
      RECT 24.69 1.977 25.51 2.023 ;
      RECT 24.735 1.92 25.505 2.06 ;
      RECT 24.821 1.872 25.49 2.13 ;
      RECT 24.907 1.841 25.475 2.176 ;
      RECT 24.93 1.822 25.46 2.184 ;
      RECT 24.975 1.795 25.435 2.209 ;
      RECT 25.06 1.777 25.42 2.215 ;
      RECT 25.146 1.771 25.42 2.215 ;
      RECT 25.232 1.766 25.365 2.215 ;
      RECT 25.318 1.761 25.365 2.215 ;
      RECT 25.01 2.659 25.18 3.045 ;
      RECT 25.005 2.659 25.18 3.04 ;
      RECT 24.98 2.659 25.18 3.005 ;
      RECT 24.98 2.687 25.19 2.995 ;
      RECT 24.96 2.687 25.19 2.955 ;
      RECT 24.955 2.687 25.19 2.928 ;
      RECT 24.955 2.705 25.195 2.92 ;
      RECT 24.9 2.705 25.195 2.855 ;
      RECT 24.9 2.722 25.205 2.838 ;
      RECT 24.89 2.722 25.205 2.778 ;
      RECT 24.89 2.739 25.21 2.775 ;
      RECT 24.885 2.575 25.055 2.753 ;
      RECT 24.885 2.609 25.141 2.753 ;
      RECT 24.88 3.375 24.885 3.388 ;
      RECT 24.875 3.27 24.88 3.393 ;
      RECT 24.85 3.13 24.875 3.408 ;
      RECT 24.815 3.081 24.85 3.44 ;
      RECT 24.81 3.049 24.815 3.46 ;
      RECT 24.805 3.04 24.81 3.46 ;
      RECT 24.725 3.005 24.805 3.46 ;
      RECT 24.662 2.975 24.725 3.46 ;
      RECT 24.576 2.963 24.662 3.46 ;
      RECT 24.49 2.949 24.576 3.46 ;
      RECT 24.41 2.936 24.49 3.446 ;
      RECT 24.375 2.928 24.41 3.426 ;
      RECT 24.365 2.925 24.375 3.417 ;
      RECT 24.335 2.92 24.365 3.404 ;
      RECT 24.285 2.895 24.335 3.38 ;
      RECT 24.271 2.869 24.285 3.362 ;
      RECT 24.185 2.829 24.271 3.338 ;
      RECT 24.14 2.777 24.185 3.307 ;
      RECT 24.13 2.752 24.14 3.294 ;
      RECT 24.125 2.533 24.13 2.555 ;
      RECT 24.12 2.735 24.13 3.29 ;
      RECT 24.12 2.531 24.125 2.645 ;
      RECT 24.11 2.527 24.12 3.286 ;
      RECT 24.066 2.525 24.11 3.274 ;
      RECT 23.98 2.525 24.066 3.245 ;
      RECT 23.95 2.525 23.98 3.218 ;
      RECT 23.935 2.525 23.95 3.206 ;
      RECT 23.895 2.537 23.935 3.191 ;
      RECT 23.875 2.556 23.895 3.17 ;
      RECT 23.865 2.566 23.875 3.154 ;
      RECT 23.855 2.572 23.865 3.143 ;
      RECT 23.835 2.582 23.855 3.126 ;
      RECT 23.83 2.591 23.835 3.113 ;
      RECT 23.825 2.595 23.83 3.063 ;
      RECT 23.815 2.601 23.825 2.98 ;
      RECT 23.81 2.605 23.815 2.894 ;
      RECT 23.805 2.625 23.81 2.831 ;
      RECT 23.8 2.648 23.805 2.778 ;
      RECT 23.795 2.666 23.8 2.723 ;
      RECT 24.405 2.485 24.575 2.745 ;
      RECT 24.575 2.45 24.62 2.731 ;
      RECT 24.536 2.452 24.625 2.714 ;
      RECT 24.425 2.469 24.711 2.685 ;
      RECT 24.425 2.484 24.715 2.657 ;
      RECT 24.425 2.465 24.625 2.714 ;
      RECT 24.45 2.453 24.575 2.745 ;
      RECT 24.536 2.451 24.62 2.731 ;
      RECT 23.59 1.84 23.76 2.33 ;
      RECT 23.59 1.84 23.795 2.31 ;
      RECT 23.725 1.76 23.835 2.27 ;
      RECT 23.706 1.764 23.855 2.24 ;
      RECT 23.62 1.772 23.875 2.223 ;
      RECT 23.62 1.778 23.88 2.213 ;
      RECT 23.62 1.787 23.9 2.201 ;
      RECT 23.595 1.812 23.93 2.179 ;
      RECT 23.595 1.832 23.935 2.159 ;
      RECT 23.59 1.845 23.945 2.139 ;
      RECT 23.59 1.912 23.95 2.12 ;
      RECT 23.59 2.045 23.955 2.107 ;
      RECT 23.585 1.85 23.945 1.94 ;
      RECT 23.595 1.807 23.9 2.201 ;
      RECT 23.706 1.762 23.835 2.27 ;
      RECT 23.58 3.515 23.88 3.77 ;
      RECT 23.665 3.481 23.88 3.77 ;
      RECT 23.665 3.484 23.885 3.63 ;
      RECT 23.6 3.505 23.885 3.63 ;
      RECT 23.635 3.495 23.88 3.77 ;
      RECT 23.63 3.5 23.885 3.63 ;
      RECT 23.665 3.479 23.866 3.77 ;
      RECT 23.751 3.47 23.866 3.77 ;
      RECT 23.751 3.464 23.78 3.77 ;
      RECT 23.24 3.105 23.25 3.595 ;
      RECT 22.9 3.04 22.91 3.34 ;
      RECT 23.415 3.212 23.42 3.431 ;
      RECT 23.405 3.192 23.415 3.448 ;
      RECT 23.395 3.172 23.405 3.478 ;
      RECT 23.39 3.162 23.395 3.493 ;
      RECT 23.385 3.158 23.39 3.498 ;
      RECT 23.37 3.15 23.385 3.505 ;
      RECT 23.33 3.13 23.37 3.53 ;
      RECT 23.305 3.112 23.33 3.563 ;
      RECT 23.3 3.11 23.305 3.576 ;
      RECT 23.28 3.107 23.3 3.58 ;
      RECT 23.25 3.105 23.28 3.59 ;
      RECT 23.18 3.107 23.24 3.591 ;
      RECT 23.16 3.107 23.18 3.585 ;
      RECT 23.135 3.105 23.16 3.582 ;
      RECT 23.1 3.1 23.135 3.578 ;
      RECT 23.08 3.094 23.1 3.565 ;
      RECT 23.07 3.091 23.08 3.553 ;
      RECT 23.05 3.088 23.07 3.538 ;
      RECT 23.03 3.084 23.05 3.52 ;
      RECT 23.025 3.081 23.03 3.51 ;
      RECT 23.02 3.08 23.025 3.508 ;
      RECT 23.01 3.077 23.02 3.5 ;
      RECT 23 3.071 23.01 3.483 ;
      RECT 22.99 3.065 23 3.465 ;
      RECT 22.98 3.059 22.99 3.453 ;
      RECT 22.97 3.053 22.98 3.433 ;
      RECT 22.965 3.049 22.97 3.418 ;
      RECT 22.96 3.047 22.965 3.41 ;
      RECT 22.955 3.045 22.96 3.403 ;
      RECT 22.95 3.043 22.955 3.393 ;
      RECT 22.945 3.041 22.95 3.387 ;
      RECT 22.935 3.04 22.945 3.377 ;
      RECT 22.925 3.04 22.935 3.368 ;
      RECT 22.91 3.04 22.925 3.353 ;
      RECT 22.87 3.04 22.9 3.337 ;
      RECT 22.85 3.042 22.87 3.332 ;
      RECT 22.845 3.047 22.85 3.33 ;
      RECT 22.815 3.055 22.845 3.328 ;
      RECT 22.785 3.07 22.815 3.327 ;
      RECT 22.74 3.092 22.785 3.332 ;
      RECT 22.735 3.107 22.74 3.336 ;
      RECT 22.72 3.112 22.735 3.338 ;
      RECT 22.715 3.116 22.72 3.34 ;
      RECT 22.655 3.139 22.715 3.349 ;
      RECT 22.635 3.165 22.655 3.362 ;
      RECT 22.625 3.172 22.635 3.366 ;
      RECT 22.61 3.179 22.625 3.369 ;
      RECT 22.59 3.189 22.61 3.372 ;
      RECT 22.585 3.197 22.59 3.375 ;
      RECT 22.54 3.202 22.585 3.382 ;
      RECT 22.53 3.205 22.54 3.389 ;
      RECT 22.52 3.205 22.53 3.393 ;
      RECT 22.485 3.207 22.52 3.405 ;
      RECT 22.465 3.21 22.485 3.418 ;
      RECT 22.425 3.213 22.465 3.429 ;
      RECT 22.41 3.215 22.425 3.442 ;
      RECT 22.4 3.215 22.41 3.447 ;
      RECT 22.375 3.216 22.4 3.455 ;
      RECT 22.365 3.218 22.375 3.46 ;
      RECT 22.36 3.219 22.365 3.463 ;
      RECT 22.335 3.217 22.36 3.466 ;
      RECT 22.32 3.215 22.335 3.467 ;
      RECT 22.3 3.212 22.32 3.469 ;
      RECT 22.28 3.207 22.3 3.469 ;
      RECT 22.22 3.202 22.28 3.466 ;
      RECT 22.185 3.177 22.22 3.462 ;
      RECT 22.175 3.154 22.185 3.46 ;
      RECT 22.145 3.131 22.175 3.46 ;
      RECT 22.135 3.11 22.145 3.46 ;
      RECT 22.11 3.092 22.135 3.458 ;
      RECT 22.095 3.07 22.11 3.455 ;
      RECT 22.08 3.052 22.095 3.453 ;
      RECT 22.06 3.042 22.08 3.451 ;
      RECT 22.045 3.037 22.06 3.45 ;
      RECT 22.03 3.035 22.045 3.449 ;
      RECT 22 3.036 22.03 3.447 ;
      RECT 21.98 3.039 22 3.445 ;
      RECT 21.923 3.043 21.98 3.445 ;
      RECT 21.837 3.052 21.923 3.445 ;
      RECT 21.751 3.063 21.837 3.445 ;
      RECT 21.665 3.074 21.751 3.445 ;
      RECT 21.645 3.081 21.665 3.453 ;
      RECT 21.635 3.084 21.645 3.46 ;
      RECT 21.57 3.089 21.635 3.478 ;
      RECT 21.54 3.096 21.57 3.503 ;
      RECT 21.53 3.099 21.54 3.51 ;
      RECT 21.485 3.103 21.53 3.515 ;
      RECT 21.455 3.108 21.485 3.52 ;
      RECT 21.454 3.11 21.455 3.52 ;
      RECT 21.368 3.116 21.454 3.52 ;
      RECT 21.282 3.127 21.368 3.52 ;
      RECT 21.196 3.139 21.282 3.52 ;
      RECT 21.11 3.15 21.196 3.52 ;
      RECT 21.095 3.157 21.11 3.515 ;
      RECT 21.09 3.159 21.095 3.509 ;
      RECT 21.07 3.17 21.09 3.504 ;
      RECT 21.06 3.188 21.07 3.498 ;
      RECT 21.055 3.2 21.06 3.298 ;
      RECT 23.35 1.953 23.37 2.04 ;
      RECT 23.345 1.888 23.35 2.072 ;
      RECT 23.335 1.855 23.345 2.077 ;
      RECT 23.33 1.835 23.335 2.083 ;
      RECT 23.3 1.835 23.33 2.1 ;
      RECT 23.251 1.835 23.3 2.136 ;
      RECT 23.165 1.835 23.251 2.194 ;
      RECT 23.136 1.845 23.165 2.243 ;
      RECT 23.05 1.887 23.136 2.296 ;
      RECT 23.03 1.925 23.05 2.343 ;
      RECT 23.005 1.942 23.03 2.363 ;
      RECT 22.995 1.956 23.005 2.383 ;
      RECT 22.99 1.962 22.995 2.393 ;
      RECT 22.985 1.966 22.99 2.4 ;
      RECT 22.935 1.986 22.985 2.405 ;
      RECT 22.87 2.03 22.935 2.405 ;
      RECT 22.845 2.08 22.87 2.405 ;
      RECT 22.835 2.11 22.845 2.405 ;
      RECT 22.83 2.137 22.835 2.405 ;
      RECT 22.825 2.155 22.83 2.405 ;
      RECT 22.815 2.197 22.825 2.405 ;
      RECT 23.165 2.755 23.335 2.93 ;
      RECT 23.105 2.583 23.165 2.918 ;
      RECT 23.095 2.576 23.105 2.901 ;
      RECT 23.05 2.755 23.335 2.881 ;
      RECT 23.031 2.755 23.335 2.859 ;
      RECT 22.945 2.755 23.335 2.824 ;
      RECT 22.925 2.575 23.095 2.78 ;
      RECT 22.925 2.722 23.33 2.78 ;
      RECT 22.925 2.67 23.305 2.78 ;
      RECT 22.925 2.625 23.27 2.78 ;
      RECT 22.925 2.607 23.235 2.78 ;
      RECT 22.925 2.597 23.23 2.78 ;
      RECT 23.095 7.855 23.265 8.305 ;
      RECT 23.15 6.075 23.32 8.025 ;
      RECT 23.095 5.015 23.265 6.245 ;
      RECT 22.575 5.015 22.745 8.305 ;
      RECT 22.575 7.315 22.98 7.645 ;
      RECT 22.575 6.475 22.98 6.805 ;
      RECT 22.645 3.555 22.835 3.78 ;
      RECT 22.635 3.556 22.84 3.775 ;
      RECT 22.635 3.558 22.85 3.755 ;
      RECT 22.635 3.562 22.855 3.74 ;
      RECT 22.635 3.549 22.805 3.775 ;
      RECT 22.635 3.552 22.83 3.775 ;
      RECT 22.645 3.548 22.805 3.78 ;
      RECT 22.731 3.546 22.805 3.78 ;
      RECT 22.355 2.797 22.525 3.035 ;
      RECT 22.355 2.797 22.611 2.949 ;
      RECT 22.355 2.797 22.615 2.859 ;
      RECT 22.405 2.57 22.625 2.838 ;
      RECT 22.4 2.587 22.63 2.811 ;
      RECT 22.365 2.745 22.63 2.811 ;
      RECT 22.385 2.595 22.525 3.035 ;
      RECT 22.375 2.677 22.635 2.794 ;
      RECT 22.37 2.725 22.635 2.794 ;
      RECT 22.375 2.635 22.63 2.811 ;
      RECT 22.4 2.572 22.625 2.838 ;
      RECT 21.965 2.547 22.135 2.745 ;
      RECT 21.965 2.547 22.18 2.72 ;
      RECT 22.035 2.49 22.205 2.678 ;
      RECT 22.01 2.505 22.205 2.678 ;
      RECT 21.625 2.551 21.655 2.745 ;
      RECT 21.62 2.523 21.625 2.745 ;
      RECT 21.59 2.497 21.62 2.747 ;
      RECT 21.565 2.455 21.59 2.75 ;
      RECT 21.555 2.427 21.565 2.752 ;
      RECT 21.52 2.407 21.555 2.754 ;
      RECT 21.455 2.392 21.52 2.76 ;
      RECT 21.405 2.39 21.455 2.766 ;
      RECT 21.382 2.392 21.405 2.771 ;
      RECT 21.296 2.403 21.382 2.777 ;
      RECT 21.21 2.421 21.296 2.787 ;
      RECT 21.195 2.432 21.21 2.793 ;
      RECT 21.125 2.455 21.195 2.799 ;
      RECT 21.07 2.487 21.125 2.807 ;
      RECT 21.03 2.51 21.07 2.813 ;
      RECT 21.016 2.523 21.03 2.816 ;
      RECT 20.93 2.545 21.016 2.822 ;
      RECT 20.915 2.57 20.93 2.828 ;
      RECT 20.875 2.585 20.915 2.832 ;
      RECT 20.825 2.6 20.875 2.837 ;
      RECT 20.8 2.607 20.825 2.841 ;
      RECT 20.74 2.602 20.8 2.845 ;
      RECT 20.725 2.593 20.74 2.849 ;
      RECT 20.655 2.583 20.725 2.845 ;
      RECT 20.63 2.575 20.65 2.835 ;
      RECT 20.571 2.575 20.63 2.813 ;
      RECT 20.485 2.575 20.571 2.77 ;
      RECT 20.65 2.575 20.655 2.84 ;
      RECT 21.345 1.806 21.515 2.14 ;
      RECT 21.315 1.806 21.515 2.135 ;
      RECT 21.255 1.773 21.315 2.123 ;
      RECT 21.255 1.829 21.525 2.118 ;
      RECT 21.23 1.829 21.525 2.112 ;
      RECT 21.225 1.77 21.255 2.109 ;
      RECT 21.21 1.776 21.345 2.107 ;
      RECT 21.205 1.784 21.43 2.095 ;
      RECT 21.205 1.836 21.54 2.048 ;
      RECT 21.19 1.792 21.43 2.043 ;
      RECT 21.19 1.862 21.55 1.984 ;
      RECT 21.16 1.812 21.515 1.945 ;
      RECT 21.16 1.902 21.56 1.941 ;
      RECT 21.21 1.781 21.43 2.107 ;
      RECT 20.55 2.111 20.605 2.375 ;
      RECT 20.55 2.111 20.67 2.374 ;
      RECT 20.55 2.111 20.695 2.373 ;
      RECT 20.55 2.111 20.76 2.372 ;
      RECT 20.695 2.077 20.775 2.371 ;
      RECT 20.51 2.121 20.92 2.37 ;
      RECT 20.55 2.118 20.92 2.37 ;
      RECT 20.51 2.126 20.925 2.363 ;
      RECT 20.495 2.128 20.925 2.362 ;
      RECT 20.495 2.135 20.93 2.358 ;
      RECT 20.475 2.134 20.925 2.354 ;
      RECT 20.475 2.142 20.935 2.353 ;
      RECT 20.47 2.139 20.93 2.349 ;
      RECT 20.47 2.152 20.945 2.348 ;
      RECT 20.455 2.142 20.935 2.347 ;
      RECT 20.42 2.155 20.945 2.34 ;
      RECT 20.605 2.11 20.915 2.37 ;
      RECT 20.605 2.095 20.865 2.37 ;
      RECT 20.67 2.082 20.8 2.37 ;
      RECT 20.215 3.171 20.23 3.564 ;
      RECT 20.18 3.176 20.23 3.563 ;
      RECT 20.215 3.175 20.275 3.562 ;
      RECT 20.16 3.186 20.275 3.561 ;
      RECT 20.175 3.182 20.275 3.561 ;
      RECT 20.14 3.192 20.35 3.558 ;
      RECT 20.14 3.211 20.395 3.556 ;
      RECT 20.14 3.218 20.4 3.553 ;
      RECT 20.125 3.195 20.35 3.55 ;
      RECT 20.105 3.2 20.35 3.543 ;
      RECT 20.1 3.204 20.35 3.539 ;
      RECT 20.1 3.221 20.41 3.538 ;
      RECT 20.08 3.215 20.395 3.534 ;
      RECT 20.08 3.224 20.415 3.528 ;
      RECT 20.075 3.23 20.415 3.3 ;
      RECT 20.14 3.19 20.275 3.558 ;
      RECT 20.015 2.553 20.215 2.865 ;
      RECT 20.09 2.531 20.215 2.865 ;
      RECT 20.03 2.55 20.22 2.85 ;
      RECT 20 2.561 20.22 2.848 ;
      RECT 20.015 2.556 20.225 2.814 ;
      RECT 20 2.66 20.23 2.781 ;
      RECT 20.03 2.532 20.215 2.865 ;
      RECT 20.09 2.51 20.19 2.865 ;
      RECT 20.115 2.507 20.19 2.865 ;
      RECT 20.115 2.502 20.135 2.865 ;
      RECT 19.52 2.57 19.695 2.745 ;
      RECT 19.515 2.57 19.695 2.743 ;
      RECT 19.49 2.57 19.695 2.738 ;
      RECT 19.435 2.55 19.605 2.728 ;
      RECT 19.435 2.557 19.67 2.728 ;
      RECT 19.52 3.237 19.535 3.42 ;
      RECT 19.51 3.215 19.52 3.42 ;
      RECT 19.495 3.195 19.51 3.42 ;
      RECT 19.485 3.17 19.495 3.42 ;
      RECT 19.455 3.135 19.485 3.42 ;
      RECT 19.42 3.075 19.455 3.42 ;
      RECT 19.415 3.037 19.42 3.42 ;
      RECT 19.365 2.988 19.415 3.42 ;
      RECT 19.355 2.938 19.365 3.408 ;
      RECT 19.34 2.917 19.355 3.368 ;
      RECT 19.32 2.885 19.34 3.318 ;
      RECT 19.295 2.841 19.32 3.258 ;
      RECT 19.29 2.813 19.295 3.213 ;
      RECT 19.285 2.804 19.29 3.199 ;
      RECT 19.28 2.797 19.285 3.186 ;
      RECT 19.275 2.792 19.28 3.175 ;
      RECT 19.27 2.777 19.275 3.165 ;
      RECT 19.265 2.755 19.27 3.152 ;
      RECT 19.255 2.715 19.265 3.127 ;
      RECT 19.23 2.645 19.255 3.083 ;
      RECT 19.225 2.585 19.23 3.048 ;
      RECT 19.21 2.565 19.225 3.015 ;
      RECT 19.205 2.565 19.21 2.99 ;
      RECT 19.175 2.565 19.205 2.945 ;
      RECT 19.13 2.565 19.175 2.885 ;
      RECT 19.055 2.565 19.13 2.833 ;
      RECT 19.05 2.565 19.055 2.798 ;
      RECT 19.045 2.565 19.05 2.788 ;
      RECT 19.04 2.565 19.045 2.768 ;
      RECT 19.305 1.785 19.475 2.255 ;
      RECT 19.25 1.778 19.445 2.239 ;
      RECT 19.25 1.792 19.48 2.238 ;
      RECT 19.235 1.793 19.48 2.219 ;
      RECT 19.23 1.811 19.48 2.205 ;
      RECT 19.235 1.794 19.485 2.203 ;
      RECT 19.22 1.825 19.485 2.188 ;
      RECT 19.235 1.8 19.49 2.173 ;
      RECT 19.215 1.84 19.49 2.17 ;
      RECT 19.23 1.812 19.495 2.155 ;
      RECT 19.23 1.824 19.5 2.135 ;
      RECT 19.215 1.84 19.505 2.118 ;
      RECT 19.215 1.85 19.51 1.973 ;
      RECT 19.21 1.85 19.51 1.93 ;
      RECT 19.21 1.865 19.515 1.908 ;
      RECT 19.305 1.775 19.445 2.255 ;
      RECT 19.305 1.773 19.415 2.255 ;
      RECT 19.391 1.77 19.415 2.255 ;
      RECT 19.05 3.437 19.055 3.483 ;
      RECT 19.04 3.285 19.05 3.507 ;
      RECT 19.035 3.13 19.04 3.532 ;
      RECT 19.02 3.092 19.035 3.543 ;
      RECT 19.015 3.075 19.02 3.55 ;
      RECT 19.005 3.063 19.015 3.557 ;
      RECT 19 3.054 19.005 3.559 ;
      RECT 18.995 3.052 19 3.563 ;
      RECT 18.95 3.043 18.995 3.578 ;
      RECT 18.945 3.035 18.95 3.592 ;
      RECT 18.94 3.032 18.945 3.596 ;
      RECT 18.925 3.027 18.94 3.604 ;
      RECT 18.87 3.017 18.925 3.615 ;
      RECT 18.835 3.005 18.87 3.616 ;
      RECT 18.826 3 18.835 3.61 ;
      RECT 18.74 3 18.826 3.6 ;
      RECT 18.71 3 18.74 3.578 ;
      RECT 18.7 3 18.705 3.558 ;
      RECT 18.695 3 18.7 3.52 ;
      RECT 18.69 3 18.695 3.478 ;
      RECT 18.685 3 18.69 3.438 ;
      RECT 18.68 3 18.685 3.368 ;
      RECT 18.67 3 18.68 3.29 ;
      RECT 18.665 3 18.67 3.19 ;
      RECT 18.705 3 18.71 3.56 ;
      RECT 18.2 3.082 18.29 3.56 ;
      RECT 18.185 3.085 18.305 3.558 ;
      RECT 18.2 3.084 18.305 3.558 ;
      RECT 18.165 3.091 18.33 3.548 ;
      RECT 18.185 3.085 18.33 3.548 ;
      RECT 18.15 3.097 18.33 3.536 ;
      RECT 18.185 3.088 18.38 3.529 ;
      RECT 18.136 3.105 18.38 3.527 ;
      RECT 18.165 3.095 18.39 3.515 ;
      RECT 18.136 3.116 18.42 3.506 ;
      RECT 18.05 3.14 18.42 3.5 ;
      RECT 18.05 3.153 18.46 3.483 ;
      RECT 18.045 3.175 18.46 3.476 ;
      RECT 18.015 3.19 18.46 3.466 ;
      RECT 18.01 3.201 18.46 3.456 ;
      RECT 17.98 3.214 18.46 3.447 ;
      RECT 17.965 3.232 18.46 3.436 ;
      RECT 17.94 3.245 18.46 3.426 ;
      RECT 18.2 3.081 18.21 3.56 ;
      RECT 18.246 2.505 18.285 2.75 ;
      RECT 18.16 2.505 18.295 2.748 ;
      RECT 18.045 2.53 18.295 2.745 ;
      RECT 18.045 2.53 18.3 2.743 ;
      RECT 18.045 2.53 18.315 2.738 ;
      RECT 18.151 2.505 18.33 2.718 ;
      RECT 18.065 2.513 18.33 2.718 ;
      RECT 17.735 1.865 17.905 2.3 ;
      RECT 17.725 1.899 17.905 2.283 ;
      RECT 17.805 1.835 17.975 2.27 ;
      RECT 17.71 1.91 17.975 2.248 ;
      RECT 17.805 1.845 17.98 2.238 ;
      RECT 17.735 1.897 18.01 2.223 ;
      RECT 17.695 1.923 18.01 2.208 ;
      RECT 17.695 1.965 18.02 2.188 ;
      RECT 17.69 1.99 18.025 2.17 ;
      RECT 17.69 2 18.03 2.155 ;
      RECT 17.685 1.937 18.01 2.153 ;
      RECT 17.685 2.01 18.035 2.138 ;
      RECT 17.68 1.947 18.01 2.135 ;
      RECT 17.675 2.031 18.04 2.118 ;
      RECT 17.675 2.063 18.045 2.098 ;
      RECT 17.67 1.977 18.02 2.09 ;
      RECT 17.675 1.962 18.01 2.118 ;
      RECT 17.69 1.932 18.01 2.17 ;
      RECT 17.535 2.519 17.76 2.775 ;
      RECT 17.535 2.552 17.78 2.765 ;
      RECT 17.5 2.552 17.78 2.763 ;
      RECT 17.5 2.565 17.785 2.753 ;
      RECT 17.5 2.585 17.795 2.745 ;
      RECT 17.5 2.682 17.8 2.738 ;
      RECT 17.48 2.43 17.61 2.728 ;
      RECT 17.435 2.585 17.795 2.67 ;
      RECT 17.425 2.43 17.61 2.615 ;
      RECT 17.425 2.462 17.696 2.615 ;
      RECT 17.39 2.992 17.41 3.17 ;
      RECT 17.355 2.945 17.39 3.17 ;
      RECT 17.34 2.885 17.355 3.17 ;
      RECT 17.315 2.832 17.34 3.17 ;
      RECT 17.3 2.785 17.315 3.17 ;
      RECT 17.28 2.762 17.3 3.17 ;
      RECT 17.255 2.727 17.28 3.17 ;
      RECT 17.245 2.573 17.255 3.17 ;
      RECT 17.215 2.568 17.245 3.161 ;
      RECT 17.21 2.565 17.215 3.151 ;
      RECT 17.195 2.565 17.21 3.125 ;
      RECT 17.19 2.565 17.195 3.088 ;
      RECT 17.165 2.565 17.19 3.04 ;
      RECT 17.145 2.565 17.165 2.965 ;
      RECT 17.135 2.565 17.145 2.925 ;
      RECT 17.13 2.565 17.135 2.9 ;
      RECT 17.125 2.565 17.13 2.883 ;
      RECT 17.12 2.565 17.125 2.865 ;
      RECT 17.115 2.566 17.12 2.855 ;
      RECT 17.105 2.568 17.115 2.823 ;
      RECT 17.095 2.57 17.105 2.79 ;
      RECT 17.085 2.573 17.095 2.763 ;
      RECT 17.41 3 17.635 3.17 ;
      RECT 16.74 1.812 16.91 2.265 ;
      RECT 16.74 1.812 17 2.231 ;
      RECT 16.74 1.812 17.03 2.215 ;
      RECT 16.74 1.812 17.06 2.188 ;
      RECT 16.996 1.79 17.075 2.17 ;
      RECT 16.775 1.797 17.08 2.155 ;
      RECT 16.775 1.805 17.09 2.118 ;
      RECT 16.735 1.832 17.09 2.09 ;
      RECT 16.72 1.845 17.09 2.055 ;
      RECT 16.74 1.82 17.11 2.045 ;
      RECT 16.715 1.885 17.11 2.015 ;
      RECT 16.715 1.915 17.115 1.998 ;
      RECT 16.71 1.945 17.115 1.985 ;
      RECT 16.775 1.794 17.075 2.17 ;
      RECT 16.91 1.791 16.996 2.249 ;
      RECT 16.861 1.792 17.075 2.17 ;
      RECT 17.005 3.452 17.05 3.645 ;
      RECT 16.995 3.422 17.005 3.645 ;
      RECT 16.99 3.407 16.995 3.645 ;
      RECT 16.95 3.317 16.99 3.645 ;
      RECT 16.945 3.23 16.95 3.645 ;
      RECT 16.935 3.2 16.945 3.645 ;
      RECT 16.93 3.16 16.935 3.645 ;
      RECT 16.92 3.122 16.93 3.645 ;
      RECT 16.915 3.087 16.92 3.645 ;
      RECT 16.895 3.04 16.915 3.645 ;
      RECT 16.88 2.965 16.895 3.645 ;
      RECT 16.875 2.92 16.88 3.64 ;
      RECT 16.87 2.9 16.875 3.613 ;
      RECT 16.865 2.88 16.87 3.598 ;
      RECT 16.86 2.855 16.865 3.578 ;
      RECT 16.855 2.833 16.86 3.563 ;
      RECT 16.85 2.811 16.855 3.545 ;
      RECT 16.845 2.79 16.85 3.535 ;
      RECT 16.835 2.762 16.845 3.505 ;
      RECT 16.825 2.725 16.835 3.473 ;
      RECT 16.815 2.685 16.825 3.44 ;
      RECT 16.805 2.663 16.815 3.41 ;
      RECT 16.775 2.615 16.805 3.342 ;
      RECT 16.76 2.575 16.775 3.269 ;
      RECT 16.75 2.575 16.76 3.235 ;
      RECT 16.745 2.575 16.75 3.21 ;
      RECT 16.74 2.575 16.745 3.195 ;
      RECT 16.735 2.575 16.74 3.173 ;
      RECT 16.73 2.575 16.735 3.16 ;
      RECT 16.715 2.575 16.73 3.125 ;
      RECT 16.695 2.575 16.715 3.065 ;
      RECT 16.685 2.575 16.695 3.015 ;
      RECT 16.665 2.575 16.685 2.963 ;
      RECT 16.645 2.575 16.665 2.92 ;
      RECT 16.635 2.575 16.645 2.908 ;
      RECT 16.605 2.575 16.635 2.895 ;
      RECT 16.575 2.596 16.605 2.875 ;
      RECT 16.565 2.624 16.575 2.855 ;
      RECT 16.55 2.641 16.565 2.823 ;
      RECT 16.545 2.655 16.55 2.79 ;
      RECT 16.54 2.663 16.545 2.763 ;
      RECT 16.535 2.671 16.54 2.725 ;
      RECT 16.54 3.195 16.545 3.53 ;
      RECT 16.505 3.182 16.54 3.529 ;
      RECT 16.435 3.122 16.505 3.528 ;
      RECT 16.355 3.065 16.435 3.527 ;
      RECT 16.22 3.025 16.355 3.526 ;
      RECT 16.22 3.212 16.555 3.515 ;
      RECT 16.18 3.212 16.555 3.505 ;
      RECT 16.18 3.23 16.56 3.5 ;
      RECT 16.18 3.32 16.565 3.49 ;
      RECT 16.175 3.015 16.34 3.47 ;
      RECT 16.17 3.015 16.34 3.213 ;
      RECT 16.17 3.172 16.535 3.213 ;
      RECT 16.17 3.16 16.53 3.213 ;
      RECT 14.94 1.74 15.11 2.935 ;
      RECT 14.94 1.74 15.405 1.91 ;
      RECT 14.94 6.97 15.405 7.14 ;
      RECT 14.94 5.945 15.11 7.14 ;
      RECT 13.95 1.74 14.12 2.935 ;
      RECT 13.95 1.74 14.415 1.91 ;
      RECT 13.95 6.97 14.415 7.14 ;
      RECT 13.95 5.945 14.12 7.14 ;
      RECT 12.095 2.635 12.265 3.865 ;
      RECT 12.15 0.855 12.32 2.805 ;
      RECT 12.095 0.575 12.265 1.025 ;
      RECT 12.095 7.855 12.265 8.305 ;
      RECT 12.15 6.075 12.32 8.025 ;
      RECT 12.095 5.015 12.265 6.245 ;
      RECT 11.575 0.575 11.745 3.865 ;
      RECT 11.575 2.075 11.98 2.405 ;
      RECT 11.575 1.235 11.98 1.565 ;
      RECT 11.575 5.015 11.745 8.305 ;
      RECT 11.575 7.315 11.98 7.645 ;
      RECT 11.575 6.475 11.98 6.805 ;
      RECT 8.91 1.975 9.64 2.215 ;
      RECT 9.452 1.77 9.64 2.215 ;
      RECT 9.28 1.782 9.655 2.209 ;
      RECT 9.195 1.797 9.675 2.194 ;
      RECT 9.195 1.812 9.68 2.184 ;
      RECT 9.15 1.832 9.695 2.176 ;
      RECT 9.127 1.867 9.71 2.13 ;
      RECT 9.041 1.89 9.715 2.09 ;
      RECT 9.041 1.908 9.725 2.06 ;
      RECT 8.91 1.977 9.73 2.023 ;
      RECT 8.955 1.92 9.725 2.06 ;
      RECT 9.041 1.872 9.71 2.13 ;
      RECT 9.127 1.841 9.695 2.176 ;
      RECT 9.15 1.822 9.68 2.184 ;
      RECT 9.195 1.795 9.655 2.209 ;
      RECT 9.28 1.777 9.64 2.215 ;
      RECT 9.366 1.771 9.64 2.215 ;
      RECT 9.452 1.766 9.585 2.215 ;
      RECT 9.538 1.761 9.585 2.215 ;
      RECT 9.23 2.659 9.4 3.045 ;
      RECT 9.225 2.659 9.4 3.04 ;
      RECT 9.2 2.659 9.4 3.005 ;
      RECT 9.2 2.687 9.41 2.995 ;
      RECT 9.18 2.687 9.41 2.955 ;
      RECT 9.175 2.687 9.41 2.928 ;
      RECT 9.175 2.705 9.415 2.92 ;
      RECT 9.12 2.705 9.415 2.855 ;
      RECT 9.12 2.722 9.425 2.838 ;
      RECT 9.11 2.722 9.425 2.778 ;
      RECT 9.11 2.739 9.43 2.775 ;
      RECT 9.105 2.575 9.275 2.753 ;
      RECT 9.105 2.609 9.361 2.753 ;
      RECT 9.1 3.375 9.105 3.388 ;
      RECT 9.095 3.27 9.1 3.393 ;
      RECT 9.07 3.13 9.095 3.408 ;
      RECT 9.035 3.081 9.07 3.44 ;
      RECT 9.03 3.049 9.035 3.46 ;
      RECT 9.025 3.04 9.03 3.46 ;
      RECT 8.945 3.005 9.025 3.46 ;
      RECT 8.882 2.975 8.945 3.46 ;
      RECT 8.796 2.963 8.882 3.46 ;
      RECT 8.71 2.949 8.796 3.46 ;
      RECT 8.63 2.936 8.71 3.446 ;
      RECT 8.595 2.928 8.63 3.426 ;
      RECT 8.585 2.925 8.595 3.417 ;
      RECT 8.555 2.92 8.585 3.404 ;
      RECT 8.505 2.895 8.555 3.38 ;
      RECT 8.491 2.869 8.505 3.362 ;
      RECT 8.405 2.829 8.491 3.338 ;
      RECT 8.36 2.777 8.405 3.307 ;
      RECT 8.35 2.752 8.36 3.294 ;
      RECT 8.345 2.533 8.35 2.555 ;
      RECT 8.34 2.735 8.35 3.29 ;
      RECT 8.34 2.531 8.345 2.645 ;
      RECT 8.33 2.527 8.34 3.286 ;
      RECT 8.286 2.525 8.33 3.274 ;
      RECT 8.2 2.525 8.286 3.245 ;
      RECT 8.17 2.525 8.2 3.218 ;
      RECT 8.155 2.525 8.17 3.206 ;
      RECT 8.115 2.537 8.155 3.191 ;
      RECT 8.095 2.556 8.115 3.17 ;
      RECT 8.085 2.566 8.095 3.154 ;
      RECT 8.075 2.572 8.085 3.143 ;
      RECT 8.055 2.582 8.075 3.126 ;
      RECT 8.05 2.591 8.055 3.113 ;
      RECT 8.045 2.595 8.05 3.063 ;
      RECT 8.035 2.601 8.045 2.98 ;
      RECT 8.03 2.605 8.035 2.894 ;
      RECT 8.025 2.625 8.03 2.831 ;
      RECT 8.02 2.648 8.025 2.778 ;
      RECT 8.015 2.666 8.02 2.723 ;
      RECT 8.625 2.485 8.795 2.745 ;
      RECT 8.795 2.45 8.84 2.731 ;
      RECT 8.756 2.452 8.845 2.714 ;
      RECT 8.645 2.469 8.931 2.685 ;
      RECT 8.645 2.484 8.935 2.657 ;
      RECT 8.645 2.465 8.845 2.714 ;
      RECT 8.67 2.453 8.795 2.745 ;
      RECT 8.756 2.451 8.84 2.731 ;
      RECT 7.81 1.84 7.98 2.33 ;
      RECT 7.81 1.84 8.015 2.31 ;
      RECT 7.945 1.76 8.055 2.27 ;
      RECT 7.926 1.764 8.075 2.24 ;
      RECT 7.84 1.772 8.095 2.223 ;
      RECT 7.84 1.778 8.1 2.213 ;
      RECT 7.84 1.787 8.12 2.201 ;
      RECT 7.815 1.812 8.15 2.179 ;
      RECT 7.815 1.832 8.155 2.159 ;
      RECT 7.81 1.845 8.165 2.139 ;
      RECT 7.81 1.912 8.17 2.12 ;
      RECT 7.81 2.045 8.175 2.107 ;
      RECT 7.805 1.85 8.165 1.94 ;
      RECT 7.815 1.807 8.12 2.201 ;
      RECT 7.926 1.762 8.055 2.27 ;
      RECT 7.8 3.515 8.1 3.77 ;
      RECT 7.885 3.481 8.1 3.77 ;
      RECT 7.885 3.484 8.105 3.63 ;
      RECT 7.82 3.505 8.105 3.63 ;
      RECT 7.855 3.495 8.1 3.77 ;
      RECT 7.85 3.5 8.105 3.63 ;
      RECT 7.885 3.479 8.086 3.77 ;
      RECT 7.971 3.47 8.086 3.77 ;
      RECT 7.971 3.464 8 3.77 ;
      RECT 7.46 3.105 7.47 3.595 ;
      RECT 7.12 3.04 7.13 3.34 ;
      RECT 7.635 3.212 7.64 3.431 ;
      RECT 7.625 3.192 7.635 3.448 ;
      RECT 7.615 3.172 7.625 3.478 ;
      RECT 7.61 3.162 7.615 3.493 ;
      RECT 7.605 3.158 7.61 3.498 ;
      RECT 7.59 3.15 7.605 3.505 ;
      RECT 7.55 3.13 7.59 3.53 ;
      RECT 7.525 3.112 7.55 3.563 ;
      RECT 7.52 3.11 7.525 3.576 ;
      RECT 7.5 3.107 7.52 3.58 ;
      RECT 7.47 3.105 7.5 3.59 ;
      RECT 7.4 3.107 7.46 3.591 ;
      RECT 7.38 3.107 7.4 3.585 ;
      RECT 7.355 3.105 7.38 3.582 ;
      RECT 7.32 3.1 7.355 3.578 ;
      RECT 7.3 3.094 7.32 3.565 ;
      RECT 7.29 3.091 7.3 3.553 ;
      RECT 7.27 3.088 7.29 3.538 ;
      RECT 7.25 3.084 7.27 3.52 ;
      RECT 7.245 3.081 7.25 3.51 ;
      RECT 7.24 3.08 7.245 3.508 ;
      RECT 7.23 3.077 7.24 3.5 ;
      RECT 7.22 3.071 7.23 3.483 ;
      RECT 7.21 3.065 7.22 3.465 ;
      RECT 7.2 3.059 7.21 3.453 ;
      RECT 7.19 3.053 7.2 3.433 ;
      RECT 7.185 3.049 7.19 3.418 ;
      RECT 7.18 3.047 7.185 3.41 ;
      RECT 7.175 3.045 7.18 3.403 ;
      RECT 7.17 3.043 7.175 3.393 ;
      RECT 7.165 3.041 7.17 3.387 ;
      RECT 7.155 3.04 7.165 3.377 ;
      RECT 7.145 3.04 7.155 3.368 ;
      RECT 7.13 3.04 7.145 3.353 ;
      RECT 7.09 3.04 7.12 3.337 ;
      RECT 7.07 3.042 7.09 3.332 ;
      RECT 7.065 3.047 7.07 3.33 ;
      RECT 7.035 3.055 7.065 3.328 ;
      RECT 7.005 3.07 7.035 3.327 ;
      RECT 6.96 3.092 7.005 3.332 ;
      RECT 6.955 3.107 6.96 3.336 ;
      RECT 6.94 3.112 6.955 3.338 ;
      RECT 6.935 3.116 6.94 3.34 ;
      RECT 6.875 3.139 6.935 3.349 ;
      RECT 6.855 3.165 6.875 3.362 ;
      RECT 6.845 3.172 6.855 3.366 ;
      RECT 6.83 3.179 6.845 3.369 ;
      RECT 6.81 3.189 6.83 3.372 ;
      RECT 6.805 3.197 6.81 3.375 ;
      RECT 6.76 3.202 6.805 3.382 ;
      RECT 6.75 3.205 6.76 3.389 ;
      RECT 6.74 3.205 6.75 3.393 ;
      RECT 6.705 3.207 6.74 3.405 ;
      RECT 6.685 3.21 6.705 3.418 ;
      RECT 6.645 3.213 6.685 3.429 ;
      RECT 6.63 3.215 6.645 3.442 ;
      RECT 6.62 3.215 6.63 3.447 ;
      RECT 6.595 3.216 6.62 3.455 ;
      RECT 6.585 3.218 6.595 3.46 ;
      RECT 6.58 3.219 6.585 3.463 ;
      RECT 6.555 3.217 6.58 3.466 ;
      RECT 6.54 3.215 6.555 3.467 ;
      RECT 6.52 3.212 6.54 3.469 ;
      RECT 6.5 3.207 6.52 3.469 ;
      RECT 6.44 3.202 6.5 3.466 ;
      RECT 6.405 3.177 6.44 3.462 ;
      RECT 6.395 3.154 6.405 3.46 ;
      RECT 6.365 3.131 6.395 3.46 ;
      RECT 6.355 3.11 6.365 3.46 ;
      RECT 6.33 3.092 6.355 3.458 ;
      RECT 6.315 3.07 6.33 3.455 ;
      RECT 6.3 3.052 6.315 3.453 ;
      RECT 6.28 3.042 6.3 3.451 ;
      RECT 6.265 3.037 6.28 3.45 ;
      RECT 6.25 3.035 6.265 3.449 ;
      RECT 6.22 3.036 6.25 3.447 ;
      RECT 6.2 3.039 6.22 3.445 ;
      RECT 6.143 3.043 6.2 3.445 ;
      RECT 6.057 3.052 6.143 3.445 ;
      RECT 5.971 3.063 6.057 3.445 ;
      RECT 5.885 3.074 5.971 3.445 ;
      RECT 5.865 3.081 5.885 3.453 ;
      RECT 5.855 3.084 5.865 3.46 ;
      RECT 5.79 3.089 5.855 3.478 ;
      RECT 5.76 3.096 5.79 3.503 ;
      RECT 5.75 3.099 5.76 3.51 ;
      RECT 5.705 3.103 5.75 3.515 ;
      RECT 5.675 3.108 5.705 3.52 ;
      RECT 5.674 3.11 5.675 3.52 ;
      RECT 5.588 3.116 5.674 3.52 ;
      RECT 5.502 3.127 5.588 3.52 ;
      RECT 5.416 3.139 5.502 3.52 ;
      RECT 5.33 3.15 5.416 3.52 ;
      RECT 5.315 3.157 5.33 3.515 ;
      RECT 5.31 3.159 5.315 3.509 ;
      RECT 5.29 3.17 5.31 3.504 ;
      RECT 5.28 3.188 5.29 3.498 ;
      RECT 5.275 3.2 5.28 3.298 ;
      RECT 7.57 1.953 7.59 2.04 ;
      RECT 7.565 1.888 7.57 2.072 ;
      RECT 7.555 1.855 7.565 2.077 ;
      RECT 7.55 1.835 7.555 2.083 ;
      RECT 7.52 1.835 7.55 2.1 ;
      RECT 7.471 1.835 7.52 2.136 ;
      RECT 7.385 1.835 7.471 2.194 ;
      RECT 7.356 1.845 7.385 2.243 ;
      RECT 7.27 1.887 7.356 2.296 ;
      RECT 7.25 1.925 7.27 2.343 ;
      RECT 7.225 1.942 7.25 2.363 ;
      RECT 7.215 1.956 7.225 2.383 ;
      RECT 7.21 1.962 7.215 2.393 ;
      RECT 7.205 1.966 7.21 2.4 ;
      RECT 7.155 1.986 7.205 2.405 ;
      RECT 7.09 2.03 7.155 2.405 ;
      RECT 7.065 2.08 7.09 2.405 ;
      RECT 7.055 2.11 7.065 2.405 ;
      RECT 7.05 2.137 7.055 2.405 ;
      RECT 7.045 2.155 7.05 2.405 ;
      RECT 7.035 2.197 7.045 2.405 ;
      RECT 7.385 2.755 7.555 2.93 ;
      RECT 7.325 2.583 7.385 2.918 ;
      RECT 7.315 2.576 7.325 2.901 ;
      RECT 7.27 2.755 7.555 2.881 ;
      RECT 7.251 2.755 7.555 2.859 ;
      RECT 7.165 2.755 7.555 2.824 ;
      RECT 7.145 2.575 7.315 2.78 ;
      RECT 7.145 2.722 7.55 2.78 ;
      RECT 7.145 2.67 7.525 2.78 ;
      RECT 7.145 2.625 7.49 2.78 ;
      RECT 7.145 2.607 7.455 2.78 ;
      RECT 7.145 2.597 7.45 2.78 ;
      RECT 7.315 7.855 7.485 8.305 ;
      RECT 7.37 6.075 7.54 8.025 ;
      RECT 7.315 5.015 7.485 6.245 ;
      RECT 6.795 5.015 6.965 8.305 ;
      RECT 6.795 7.315 7.2 7.645 ;
      RECT 6.795 6.475 7.2 6.805 ;
      RECT 6.865 3.555 7.055 3.78 ;
      RECT 6.855 3.556 7.06 3.775 ;
      RECT 6.855 3.558 7.07 3.755 ;
      RECT 6.855 3.562 7.075 3.74 ;
      RECT 6.855 3.549 7.025 3.775 ;
      RECT 6.855 3.552 7.05 3.775 ;
      RECT 6.865 3.548 7.025 3.78 ;
      RECT 6.951 3.546 7.025 3.78 ;
      RECT 6.575 2.797 6.745 3.035 ;
      RECT 6.575 2.797 6.831 2.949 ;
      RECT 6.575 2.797 6.835 2.859 ;
      RECT 6.625 2.57 6.845 2.838 ;
      RECT 6.62 2.587 6.85 2.811 ;
      RECT 6.585 2.745 6.85 2.811 ;
      RECT 6.605 2.595 6.745 3.035 ;
      RECT 6.595 2.677 6.855 2.794 ;
      RECT 6.59 2.725 6.855 2.794 ;
      RECT 6.595 2.635 6.85 2.811 ;
      RECT 6.62 2.572 6.845 2.838 ;
      RECT 6.185 2.547 6.355 2.745 ;
      RECT 6.185 2.547 6.4 2.72 ;
      RECT 6.255 2.49 6.425 2.678 ;
      RECT 6.23 2.505 6.425 2.678 ;
      RECT 5.845 2.551 5.875 2.745 ;
      RECT 5.84 2.523 5.845 2.745 ;
      RECT 5.81 2.497 5.84 2.747 ;
      RECT 5.785 2.455 5.81 2.75 ;
      RECT 5.775 2.427 5.785 2.752 ;
      RECT 5.74 2.407 5.775 2.754 ;
      RECT 5.675 2.392 5.74 2.76 ;
      RECT 5.625 2.39 5.675 2.766 ;
      RECT 5.602 2.392 5.625 2.771 ;
      RECT 5.516 2.403 5.602 2.777 ;
      RECT 5.43 2.421 5.516 2.787 ;
      RECT 5.415 2.432 5.43 2.793 ;
      RECT 5.345 2.455 5.415 2.799 ;
      RECT 5.29 2.487 5.345 2.807 ;
      RECT 5.25 2.51 5.29 2.813 ;
      RECT 5.236 2.523 5.25 2.816 ;
      RECT 5.15 2.545 5.236 2.822 ;
      RECT 5.135 2.57 5.15 2.828 ;
      RECT 5.095 2.585 5.135 2.832 ;
      RECT 5.045 2.6 5.095 2.837 ;
      RECT 5.02 2.607 5.045 2.841 ;
      RECT 4.96 2.602 5.02 2.845 ;
      RECT 4.945 2.593 4.96 2.849 ;
      RECT 4.875 2.583 4.945 2.845 ;
      RECT 4.85 2.575 4.87 2.835 ;
      RECT 4.791 2.575 4.85 2.813 ;
      RECT 4.705 2.575 4.791 2.77 ;
      RECT 4.87 2.575 4.875 2.84 ;
      RECT 5.565 1.806 5.735 2.14 ;
      RECT 5.535 1.806 5.735 2.135 ;
      RECT 5.475 1.773 5.535 2.123 ;
      RECT 5.475 1.829 5.745 2.118 ;
      RECT 5.45 1.829 5.745 2.112 ;
      RECT 5.445 1.77 5.475 2.109 ;
      RECT 5.43 1.776 5.565 2.107 ;
      RECT 5.425 1.784 5.65 2.095 ;
      RECT 5.425 1.836 5.76 2.048 ;
      RECT 5.41 1.792 5.65 2.043 ;
      RECT 5.41 1.862 5.77 1.984 ;
      RECT 5.38 1.812 5.735 1.945 ;
      RECT 5.38 1.902 5.78 1.941 ;
      RECT 5.43 1.781 5.65 2.107 ;
      RECT 4.77 2.111 4.825 2.375 ;
      RECT 4.77 2.111 4.89 2.374 ;
      RECT 4.77 2.111 4.915 2.373 ;
      RECT 4.77 2.111 4.98 2.372 ;
      RECT 4.915 2.077 4.995 2.371 ;
      RECT 4.73 2.121 5.14 2.37 ;
      RECT 4.77 2.118 5.14 2.37 ;
      RECT 4.73 2.126 5.145 2.363 ;
      RECT 4.715 2.128 5.145 2.362 ;
      RECT 4.715 2.135 5.15 2.358 ;
      RECT 4.695 2.134 5.145 2.354 ;
      RECT 4.695 2.142 5.155 2.353 ;
      RECT 4.69 2.139 5.15 2.349 ;
      RECT 4.69 2.152 5.165 2.348 ;
      RECT 4.675 2.142 5.155 2.347 ;
      RECT 4.64 2.155 5.165 2.34 ;
      RECT 4.825 2.11 5.135 2.37 ;
      RECT 4.825 2.095 5.085 2.37 ;
      RECT 4.89 2.082 5.02 2.37 ;
      RECT 4.435 3.171 4.45 3.564 ;
      RECT 4.4 3.176 4.45 3.563 ;
      RECT 4.435 3.175 4.495 3.562 ;
      RECT 4.38 3.186 4.495 3.561 ;
      RECT 4.395 3.182 4.495 3.561 ;
      RECT 4.36 3.192 4.57 3.558 ;
      RECT 4.36 3.211 4.615 3.556 ;
      RECT 4.36 3.218 4.62 3.553 ;
      RECT 4.345 3.195 4.57 3.55 ;
      RECT 4.325 3.2 4.57 3.543 ;
      RECT 4.32 3.204 4.57 3.539 ;
      RECT 4.32 3.221 4.63 3.538 ;
      RECT 4.3 3.215 4.615 3.534 ;
      RECT 4.3 3.224 4.635 3.528 ;
      RECT 4.295 3.23 4.635 3.3 ;
      RECT 4.36 3.19 4.495 3.558 ;
      RECT 4.235 2.553 4.435 2.865 ;
      RECT 4.31 2.531 4.435 2.865 ;
      RECT 4.25 2.55 4.44 2.85 ;
      RECT 4.22 2.561 4.44 2.848 ;
      RECT 4.235 2.556 4.445 2.814 ;
      RECT 4.22 2.66 4.45 2.781 ;
      RECT 4.25 2.532 4.435 2.865 ;
      RECT 4.31 2.51 4.41 2.865 ;
      RECT 4.335 2.507 4.41 2.865 ;
      RECT 4.335 2.502 4.355 2.865 ;
      RECT 3.74 2.57 3.915 2.745 ;
      RECT 3.735 2.57 3.915 2.743 ;
      RECT 3.71 2.57 3.915 2.738 ;
      RECT 3.655 2.55 3.825 2.728 ;
      RECT 3.655 2.557 3.89 2.728 ;
      RECT 3.74 3.237 3.755 3.42 ;
      RECT 3.73 3.215 3.74 3.42 ;
      RECT 3.715 3.195 3.73 3.42 ;
      RECT 3.705 3.17 3.715 3.42 ;
      RECT 3.675 3.135 3.705 3.42 ;
      RECT 3.64 3.075 3.675 3.42 ;
      RECT 3.635 3.037 3.64 3.42 ;
      RECT 3.585 2.988 3.635 3.42 ;
      RECT 3.575 2.938 3.585 3.408 ;
      RECT 3.56 2.917 3.575 3.368 ;
      RECT 3.54 2.885 3.56 3.318 ;
      RECT 3.515 2.841 3.54 3.258 ;
      RECT 3.51 2.813 3.515 3.213 ;
      RECT 3.505 2.804 3.51 3.199 ;
      RECT 3.5 2.797 3.505 3.186 ;
      RECT 3.495 2.792 3.5 3.175 ;
      RECT 3.49 2.777 3.495 3.165 ;
      RECT 3.485 2.755 3.49 3.152 ;
      RECT 3.475 2.715 3.485 3.127 ;
      RECT 3.45 2.645 3.475 3.083 ;
      RECT 3.445 2.585 3.45 3.048 ;
      RECT 3.43 2.565 3.445 3.015 ;
      RECT 3.425 2.565 3.43 2.99 ;
      RECT 3.395 2.565 3.425 2.945 ;
      RECT 3.35 2.565 3.395 2.885 ;
      RECT 3.275 2.565 3.35 2.833 ;
      RECT 3.27 2.565 3.275 2.798 ;
      RECT 3.265 2.565 3.27 2.788 ;
      RECT 3.26 2.565 3.265 2.768 ;
      RECT 3.525 1.785 3.695 2.255 ;
      RECT 3.47 1.778 3.665 2.239 ;
      RECT 3.47 1.792 3.7 2.238 ;
      RECT 3.455 1.793 3.7 2.219 ;
      RECT 3.45 1.811 3.7 2.205 ;
      RECT 3.455 1.794 3.705 2.203 ;
      RECT 3.44 1.825 3.705 2.188 ;
      RECT 3.455 1.8 3.71 2.173 ;
      RECT 3.435 1.84 3.71 2.17 ;
      RECT 3.45 1.812 3.715 2.155 ;
      RECT 3.45 1.824 3.72 2.135 ;
      RECT 3.435 1.84 3.725 2.118 ;
      RECT 3.435 1.85 3.73 1.973 ;
      RECT 3.43 1.85 3.73 1.93 ;
      RECT 3.43 1.865 3.735 1.908 ;
      RECT 3.525 1.775 3.665 2.255 ;
      RECT 3.525 1.773 3.635 2.255 ;
      RECT 3.611 1.77 3.635 2.255 ;
      RECT 3.27 3.437 3.275 3.483 ;
      RECT 3.26 3.285 3.27 3.507 ;
      RECT 3.255 3.13 3.26 3.532 ;
      RECT 3.24 3.092 3.255 3.543 ;
      RECT 3.235 3.075 3.24 3.55 ;
      RECT 3.225 3.063 3.235 3.557 ;
      RECT 3.22 3.054 3.225 3.559 ;
      RECT 3.215 3.052 3.22 3.563 ;
      RECT 3.17 3.043 3.215 3.578 ;
      RECT 3.165 3.035 3.17 3.592 ;
      RECT 3.16 3.032 3.165 3.596 ;
      RECT 3.145 3.027 3.16 3.604 ;
      RECT 3.09 3.017 3.145 3.615 ;
      RECT 3.055 3.005 3.09 3.616 ;
      RECT 3.046 3 3.055 3.61 ;
      RECT 2.96 3 3.046 3.6 ;
      RECT 2.93 3 2.96 3.578 ;
      RECT 2.92 3 2.925 3.558 ;
      RECT 2.915 3 2.92 3.52 ;
      RECT 2.91 3 2.915 3.478 ;
      RECT 2.905 3 2.91 3.438 ;
      RECT 2.9 3 2.905 3.368 ;
      RECT 2.89 3 2.9 3.29 ;
      RECT 2.885 3 2.89 3.19 ;
      RECT 2.925 3 2.93 3.56 ;
      RECT 2.42 3.082 2.51 3.56 ;
      RECT 2.405 3.085 2.525 3.558 ;
      RECT 2.42 3.084 2.525 3.558 ;
      RECT 2.385 3.091 2.55 3.548 ;
      RECT 2.405 3.085 2.55 3.548 ;
      RECT 2.37 3.097 2.55 3.536 ;
      RECT 2.405 3.088 2.6 3.529 ;
      RECT 2.356 3.105 2.6 3.527 ;
      RECT 2.385 3.095 2.61 3.515 ;
      RECT 2.356 3.116 2.64 3.506 ;
      RECT 2.27 3.14 2.64 3.5 ;
      RECT 2.27 3.153 2.68 3.483 ;
      RECT 2.265 3.175 2.68 3.476 ;
      RECT 2.235 3.19 2.68 3.466 ;
      RECT 2.23 3.201 2.68 3.456 ;
      RECT 2.2 3.214 2.68 3.447 ;
      RECT 2.185 3.232 2.68 3.436 ;
      RECT 2.16 3.245 2.68 3.426 ;
      RECT 2.42 3.081 2.43 3.56 ;
      RECT 2.466 2.505 2.505 2.75 ;
      RECT 2.38 2.505 2.515 2.748 ;
      RECT 2.265 2.53 2.515 2.745 ;
      RECT 2.265 2.53 2.52 2.743 ;
      RECT 2.265 2.53 2.535 2.738 ;
      RECT 2.371 2.505 2.55 2.718 ;
      RECT 2.285 2.513 2.55 2.718 ;
      RECT 1.955 1.865 2.125 2.3 ;
      RECT 1.945 1.899 2.125 2.283 ;
      RECT 2.025 1.835 2.195 2.27 ;
      RECT 1.93 1.91 2.195 2.248 ;
      RECT 2.025 1.845 2.2 2.238 ;
      RECT 1.955 1.897 2.23 2.223 ;
      RECT 1.915 1.923 2.23 2.208 ;
      RECT 1.915 1.965 2.24 2.188 ;
      RECT 1.91 1.99 2.245 2.17 ;
      RECT 1.91 2 2.25 2.155 ;
      RECT 1.905 1.937 2.23 2.153 ;
      RECT 1.905 2.01 2.255 2.138 ;
      RECT 1.9 1.947 2.23 2.135 ;
      RECT 1.895 2.031 2.26 2.118 ;
      RECT 1.895 2.063 2.265 2.098 ;
      RECT 1.89 1.977 2.24 2.09 ;
      RECT 1.895 1.962 2.23 2.118 ;
      RECT 1.91 1.932 2.23 2.17 ;
      RECT 1.755 2.519 1.98 2.775 ;
      RECT 1.755 2.552 2 2.765 ;
      RECT 1.72 2.552 2 2.763 ;
      RECT 1.72 2.565 2.005 2.753 ;
      RECT 1.72 2.585 2.015 2.745 ;
      RECT 1.72 2.682 2.02 2.738 ;
      RECT 1.7 2.43 1.83 2.728 ;
      RECT 1.655 2.585 2.015 2.67 ;
      RECT 1.645 2.43 1.83 2.615 ;
      RECT 1.645 2.462 1.916 2.615 ;
      RECT 1.61 2.992 1.63 3.17 ;
      RECT 1.575 2.945 1.61 3.17 ;
      RECT 1.56 2.885 1.575 3.17 ;
      RECT 1.535 2.832 1.56 3.17 ;
      RECT 1.52 2.785 1.535 3.17 ;
      RECT 1.5 2.762 1.52 3.17 ;
      RECT 1.475 2.727 1.5 3.17 ;
      RECT 1.465 2.573 1.475 3.17 ;
      RECT 1.435 2.568 1.465 3.161 ;
      RECT 1.43 2.565 1.435 3.151 ;
      RECT 1.415 2.565 1.43 3.125 ;
      RECT 1.41 2.565 1.415 3.088 ;
      RECT 1.385 2.565 1.41 3.04 ;
      RECT 1.365 2.565 1.385 2.965 ;
      RECT 1.355 2.565 1.365 2.925 ;
      RECT 1.35 2.565 1.355 2.9 ;
      RECT 1.345 2.565 1.35 2.883 ;
      RECT 1.34 2.565 1.345 2.865 ;
      RECT 1.335 2.566 1.34 2.855 ;
      RECT 1.325 2.568 1.335 2.823 ;
      RECT 1.315 2.57 1.325 2.79 ;
      RECT 1.305 2.573 1.315 2.763 ;
      RECT 1.63 3 1.855 3.17 ;
      RECT 0.96 1.812 1.13 2.265 ;
      RECT 0.96 1.812 1.22 2.231 ;
      RECT 0.96 1.812 1.25 2.215 ;
      RECT 0.96 1.812 1.28 2.188 ;
      RECT 1.216 1.79 1.295 2.17 ;
      RECT 0.995 1.797 1.3 2.155 ;
      RECT 0.995 1.805 1.31 2.118 ;
      RECT 0.955 1.832 1.31 2.09 ;
      RECT 0.94 1.845 1.31 2.055 ;
      RECT 0.96 1.82 1.33 2.045 ;
      RECT 0.935 1.885 1.33 2.015 ;
      RECT 0.935 1.915 1.335 1.998 ;
      RECT 0.93 1.945 1.335 1.985 ;
      RECT 0.995 1.794 1.295 2.17 ;
      RECT 1.13 1.791 1.216 2.249 ;
      RECT 1.081 1.792 1.295 2.17 ;
      RECT 1.225 3.452 1.27 3.645 ;
      RECT 1.215 3.422 1.225 3.645 ;
      RECT 1.21 3.407 1.215 3.645 ;
      RECT 1.17 3.317 1.21 3.645 ;
      RECT 1.165 3.23 1.17 3.645 ;
      RECT 1.155 3.2 1.165 3.645 ;
      RECT 1.15 3.16 1.155 3.645 ;
      RECT 1.14 3.122 1.15 3.645 ;
      RECT 1.135 3.087 1.14 3.645 ;
      RECT 1.115 3.04 1.135 3.645 ;
      RECT 1.1 2.965 1.115 3.645 ;
      RECT 1.095 2.92 1.1 3.64 ;
      RECT 1.09 2.9 1.095 3.613 ;
      RECT 1.085 2.88 1.09 3.598 ;
      RECT 1.08 2.855 1.085 3.578 ;
      RECT 1.075 2.833 1.08 3.563 ;
      RECT 1.07 2.811 1.075 3.545 ;
      RECT 1.065 2.79 1.07 3.535 ;
      RECT 1.055 2.762 1.065 3.505 ;
      RECT 1.045 2.725 1.055 3.473 ;
      RECT 1.035 2.685 1.045 3.44 ;
      RECT 1.025 2.663 1.035 3.41 ;
      RECT 0.995 2.615 1.025 3.342 ;
      RECT 0.98 2.575 0.995 3.269 ;
      RECT 0.97 2.575 0.98 3.235 ;
      RECT 0.965 2.575 0.97 3.21 ;
      RECT 0.96 2.575 0.965 3.195 ;
      RECT 0.955 2.575 0.96 3.173 ;
      RECT 0.95 2.575 0.955 3.16 ;
      RECT 0.935 2.575 0.95 3.125 ;
      RECT 0.915 2.575 0.935 3.065 ;
      RECT 0.905 2.575 0.915 3.015 ;
      RECT 0.885 2.575 0.905 2.963 ;
      RECT 0.865 2.575 0.885 2.92 ;
      RECT 0.855 2.575 0.865 2.908 ;
      RECT 0.825 2.575 0.855 2.895 ;
      RECT 0.795 2.596 0.825 2.875 ;
      RECT 0.785 2.624 0.795 2.855 ;
      RECT 0.77 2.641 0.785 2.823 ;
      RECT 0.765 2.655 0.77 2.79 ;
      RECT 0.76 2.663 0.765 2.763 ;
      RECT 0.755 2.671 0.76 2.725 ;
      RECT 0.76 3.195 0.765 3.53 ;
      RECT 0.725 3.182 0.76 3.529 ;
      RECT 0.655 3.122 0.725 3.528 ;
      RECT 0.575 3.065 0.655 3.527 ;
      RECT 0.44 3.025 0.575 3.526 ;
      RECT 0.44 3.212 0.775 3.515 ;
      RECT 0.4 3.212 0.775 3.505 ;
      RECT 0.4 3.23 0.78 3.5 ;
      RECT 0.4 3.32 0.785 3.49 ;
      RECT 0.395 3.015 0.56 3.47 ;
      RECT 0.39 3.015 0.56 3.213 ;
      RECT 0.39 3.172 0.755 3.213 ;
      RECT 0.39 3.16 0.75 3.213 ;
      RECT -1.62 7.855 -1.45 8.305 ;
      RECT -1.565 6.075 -1.395 8.025 ;
      RECT -1.62 5.015 -1.45 6.245 ;
      RECT -2.14 5.015 -1.97 8.305 ;
      RECT -2.14 7.315 -1.735 7.645 ;
      RECT -2.14 6.475 -1.735 6.805 ;
      RECT 78.435 0.575 78.605 1.085 ;
      RECT 78.435 2.395 78.605 3.865 ;
      RECT 78.435 5.015 78.605 6.485 ;
      RECT 78.435 7.795 78.605 8.305 ;
      RECT 77.445 0.575 77.615 1.085 ;
      RECT 77.445 2.395 77.615 3.865 ;
      RECT 77.445 5.015 77.615 6.485 ;
      RECT 77.445 7.795 77.615 8.305 ;
      RECT 76.08 0.575 76.25 3.865 ;
      RECT 76.08 5.015 76.25 8.305 ;
      RECT 75.65 0.575 75.82 1.085 ;
      RECT 75.65 1.655 75.82 3.865 ;
      RECT 75.65 5.015 75.82 7.225 ;
      RECT 75.65 7.795 75.82 8.305 ;
      RECT 74.28 1.66 74.45 2.935 ;
      RECT 74.28 5.945 74.45 7.22 ;
      RECT 73.26 2.85 73.63 3.22 ;
      RECT 71.3 5.015 71.47 8.305 ;
      RECT 70.87 5.015 71.04 7.225 ;
      RECT 70.87 7.795 71.04 8.305 ;
      RECT 69.5 5.945 69.67 7.22 ;
      RECT 62.65 0.575 62.82 1.085 ;
      RECT 62.65 2.395 62.82 3.865 ;
      RECT 62.65 5.015 62.82 6.485 ;
      RECT 62.65 7.795 62.82 8.305 ;
      RECT 61.66 0.575 61.83 1.085 ;
      RECT 61.66 2.395 61.83 3.865 ;
      RECT 61.66 5.015 61.83 6.485 ;
      RECT 61.66 7.795 61.83 8.305 ;
      RECT 60.295 0.575 60.465 3.865 ;
      RECT 60.295 5.015 60.465 8.305 ;
      RECT 59.865 0.575 60.035 1.085 ;
      RECT 59.865 1.655 60.035 3.865 ;
      RECT 59.865 5.015 60.035 7.225 ;
      RECT 59.865 7.795 60.035 8.305 ;
      RECT 58.495 1.66 58.665 2.935 ;
      RECT 58.495 5.945 58.665 7.22 ;
      RECT 57.475 2.85 57.845 3.22 ;
      RECT 55.515 5.015 55.685 8.305 ;
      RECT 55.085 5.015 55.255 7.225 ;
      RECT 55.085 7.795 55.255 8.305 ;
      RECT 53.715 5.945 53.885 7.22 ;
      RECT 46.865 0.575 47.035 1.085 ;
      RECT 46.865 2.395 47.035 3.865 ;
      RECT 46.865 5.015 47.035 6.485 ;
      RECT 46.865 7.795 47.035 8.305 ;
      RECT 45.875 0.575 46.045 1.085 ;
      RECT 45.875 2.395 46.045 3.865 ;
      RECT 45.875 5.015 46.045 6.485 ;
      RECT 45.875 7.795 46.045 8.305 ;
      RECT 44.51 0.575 44.68 3.865 ;
      RECT 44.51 5.015 44.68 8.305 ;
      RECT 44.08 0.575 44.25 1.085 ;
      RECT 44.08 1.655 44.25 3.865 ;
      RECT 44.08 5.015 44.25 7.225 ;
      RECT 44.08 7.795 44.25 8.305 ;
      RECT 42.71 1.66 42.88 2.935 ;
      RECT 42.71 5.945 42.88 7.22 ;
      RECT 41.69 2.85 42.06 3.22 ;
      RECT 39.73 5.015 39.9 8.305 ;
      RECT 39.3 5.015 39.47 7.225 ;
      RECT 39.3 7.795 39.47 8.305 ;
      RECT 37.93 5.945 38.1 7.22 ;
      RECT 31.09 0.575 31.26 1.085 ;
      RECT 31.09 2.395 31.26 3.865 ;
      RECT 31.09 5.015 31.26 6.485 ;
      RECT 31.09 7.795 31.26 8.305 ;
      RECT 30.1 0.575 30.27 1.085 ;
      RECT 30.1 2.395 30.27 3.865 ;
      RECT 30.1 5.015 30.27 6.485 ;
      RECT 30.1 7.795 30.27 8.305 ;
      RECT 28.735 0.575 28.905 3.865 ;
      RECT 28.735 5.015 28.905 8.305 ;
      RECT 28.305 0.575 28.475 1.085 ;
      RECT 28.305 1.655 28.475 3.865 ;
      RECT 28.305 5.015 28.475 7.225 ;
      RECT 28.305 7.795 28.475 8.305 ;
      RECT 26.935 1.66 27.105 2.935 ;
      RECT 26.935 5.945 27.105 7.22 ;
      RECT 25.915 2.85 26.285 3.22 ;
      RECT 23.955 5.015 24.125 8.305 ;
      RECT 23.525 5.015 23.695 7.225 ;
      RECT 23.525 7.795 23.695 8.305 ;
      RECT 22.155 5.945 22.325 7.22 ;
      RECT 15.31 0.575 15.48 1.085 ;
      RECT 15.31 2.395 15.48 3.865 ;
      RECT 15.31 5.015 15.48 6.485 ;
      RECT 15.31 7.795 15.48 8.305 ;
      RECT 14.32 0.575 14.49 1.085 ;
      RECT 14.32 2.395 14.49 3.865 ;
      RECT 14.32 5.015 14.49 6.485 ;
      RECT 14.32 7.795 14.49 8.305 ;
      RECT 12.955 0.575 13.125 3.865 ;
      RECT 12.955 5.015 13.125 8.305 ;
      RECT 12.525 0.575 12.695 1.085 ;
      RECT 12.525 1.655 12.695 3.865 ;
      RECT 12.525 5.015 12.695 7.225 ;
      RECT 12.525 7.795 12.695 8.305 ;
      RECT 11.155 1.66 11.325 2.935 ;
      RECT 11.155 5.945 11.325 7.22 ;
      RECT 10.135 2.85 10.505 3.22 ;
      RECT 8.175 5.015 8.345 8.305 ;
      RECT 7.745 5.015 7.915 7.225 ;
      RECT 7.745 7.795 7.915 8.305 ;
      RECT 6.375 5.945 6.545 7.22 ;
      RECT -1.19 5.015 -1.02 7.225 ;
      RECT -1.19 7.795 -1.02 8.305 ;
      RECT -2.56 5.945 -2.39 7.22 ;
  END
END sky130_osu_ring_oscillator_mpr2aa_8_b0r2

MACRO sky130_osu_ring_oscillator_mpr2at_8_b0r1
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 4.885 0 ;
  SIZE 92.435 BY 8.88 ;
  SYMMETRY X Y R90 ;
  SITE CoreSite ;
  OBS
    LAYER met3 ;
      RECT 79.355 7.055 79.73 7.425 ;
      RECT 79.39 4.925 79.7 7.425 ;
      RECT 79.39 4.925 82.485 5.235 ;
      RECT 82.175 1.125 82.485 5.235 ;
      RECT 82.175 1.14 82.55 1.51 ;
      RECT 79.305 3.685 79.86 4.015 ;
      RECT 79.305 2.02 79.605 4.015 ;
      RECT 75.37 3.125 75.925 3.455 ;
      RECT 75.625 2.02 75.925 3.455 ;
      RECT 76.42 1.885 76.57 2.535 ;
      RECT 75.625 2.02 79.605 2.32 ;
      RECT 74.14 0.96 74.44 3.91 ;
      RECT 74.13 2.565 74.86 2.895 ;
      RECT 74.095 0.96 74.47 1.33 ;
      RECT 72.69 3.125 73.42 3.455 ;
      RECT 72.705 0.96 73.005 3.455 ;
      RECT 70.58 2.565 71.31 2.895 ;
      RECT 70.735 0.93 71.035 2.895 ;
      RECT 72.66 0.96 73.035 1.33 ;
      RECT 70.69 0.93 71.065 1.3 ;
      RECT 70.69 0.97 73.035 1.27 ;
      RECT 61.43 7.055 61.805 7.425 ;
      RECT 61.465 4.925 61.775 7.425 ;
      RECT 61.465 4.925 64.56 5.235 ;
      RECT 64.25 1.125 64.56 5.235 ;
      RECT 64.25 1.14 64.625 1.51 ;
      RECT 61.38 3.685 61.935 4.015 ;
      RECT 61.38 2.02 61.68 4.015 ;
      RECT 57.445 3.125 58 3.455 ;
      RECT 57.7 2.02 58 3.455 ;
      RECT 58.495 1.885 58.645 2.535 ;
      RECT 57.7 2.02 61.68 2.32 ;
      RECT 56.215 0.96 56.515 3.91 ;
      RECT 56.205 2.565 56.935 2.895 ;
      RECT 56.17 0.96 56.545 1.33 ;
      RECT 54.765 3.125 55.495 3.455 ;
      RECT 54.78 0.96 55.08 3.455 ;
      RECT 52.655 2.565 53.385 2.895 ;
      RECT 52.81 0.93 53.11 2.895 ;
      RECT 54.735 0.96 55.11 1.33 ;
      RECT 52.765 0.93 53.14 1.3 ;
      RECT 52.765 0.97 55.11 1.27 ;
      RECT 43.505 7.055 43.88 7.425 ;
      RECT 43.54 4.925 43.85 7.425 ;
      RECT 43.54 4.925 46.635 5.235 ;
      RECT 46.325 1.125 46.635 5.235 ;
      RECT 46.325 1.14 46.7 1.51 ;
      RECT 43.455 3.685 44.01 4.015 ;
      RECT 43.455 2.02 43.755 4.015 ;
      RECT 39.52 3.125 40.075 3.455 ;
      RECT 39.775 2.02 40.075 3.455 ;
      RECT 40.57 1.885 40.72 2.535 ;
      RECT 39.775 2.02 43.755 2.32 ;
      RECT 38.29 0.96 38.59 3.91 ;
      RECT 38.28 2.565 39.01 2.895 ;
      RECT 38.245 0.96 38.62 1.33 ;
      RECT 36.84 3.125 37.57 3.455 ;
      RECT 36.855 0.96 37.155 3.455 ;
      RECT 34.73 2.565 35.46 2.895 ;
      RECT 34.885 0.93 35.185 2.895 ;
      RECT 36.81 0.96 37.185 1.33 ;
      RECT 34.84 0.93 35.215 1.3 ;
      RECT 34.84 0.97 37.185 1.27 ;
      RECT 25.58 7.055 25.955 7.425 ;
      RECT 25.615 4.925 25.925 7.425 ;
      RECT 25.615 4.925 28.71 5.235 ;
      RECT 28.4 1.125 28.71 5.235 ;
      RECT 28.4 1.14 28.775 1.51 ;
      RECT 25.53 3.685 26.085 4.015 ;
      RECT 25.53 2.02 25.83 4.015 ;
      RECT 21.595 3.125 22.15 3.455 ;
      RECT 21.85 2.02 22.15 3.455 ;
      RECT 22.645 1.885 22.795 2.535 ;
      RECT 21.85 2.02 25.83 2.32 ;
      RECT 20.365 0.96 20.665 3.91 ;
      RECT 20.355 2.565 21.085 2.895 ;
      RECT 20.32 0.96 20.695 1.33 ;
      RECT 18.915 3.125 19.645 3.455 ;
      RECT 18.93 0.96 19.23 3.455 ;
      RECT 16.805 2.565 17.535 2.895 ;
      RECT 16.96 0.93 17.26 2.895 ;
      RECT 18.885 0.96 19.26 1.33 ;
      RECT 16.915 0.93 17.29 1.3 ;
      RECT 16.915 0.97 19.26 1.27 ;
      RECT 7.655 7.055 8.03 7.425 ;
      RECT 7.69 4.925 8 7.425 ;
      RECT 7.69 4.925 10.785 5.235 ;
      RECT 10.475 1.125 10.785 5.235 ;
      RECT 10.475 1.14 10.85 1.51 ;
      RECT 7.605 3.685 8.16 4.015 ;
      RECT 7.605 2.02 7.905 4.015 ;
      RECT 3.67 3.125 4.225 3.455 ;
      RECT 3.925 2.02 4.225 3.455 ;
      RECT 4.72 1.885 4.87 2.535 ;
      RECT 3.925 2.02 7.905 2.32 ;
      RECT 2.44 0.96 2.74 3.91 ;
      RECT 2.43 2.565 3.16 2.895 ;
      RECT 2.395 0.96 2.77 1.33 ;
      RECT 0.99 3.125 1.72 3.455 ;
      RECT 1.005 0.96 1.305 3.455 ;
      RECT -1.12 2.565 -0.39 2.895 ;
      RECT -0.965 0.93 -0.665 2.895 ;
      RECT 0.96 0.96 1.335 1.33 ;
      RECT -1.01 0.93 -0.635 1.3 ;
      RECT -1.01 0.97 1.335 1.27 ;
      RECT 80.49 2.005 81.22 2.335 ;
      RECT 78.27 3.685 79 4.015 ;
      RECT 76.57 3.685 77.3 4.015 ;
      RECT 71.615 2.565 72.345 2.895 ;
      RECT 70.25 3.685 70.98 4.015 ;
      RECT 62.565 2.005 63.295 2.335 ;
      RECT 60.345 3.685 61.075 4.015 ;
      RECT 58.645 3.685 59.375 4.015 ;
      RECT 53.69 2.565 54.42 2.895 ;
      RECT 52.325 3.685 53.055 4.015 ;
      RECT 44.64 2.005 45.37 2.335 ;
      RECT 42.42 3.685 43.15 4.015 ;
      RECT 40.72 3.685 41.45 4.015 ;
      RECT 35.765 2.565 36.495 2.895 ;
      RECT 34.4 3.685 35.13 4.015 ;
      RECT 26.715 2.005 27.445 2.335 ;
      RECT 24.495 3.685 25.225 4.015 ;
      RECT 22.795 3.685 23.525 4.015 ;
      RECT 17.84 2.565 18.57 2.895 ;
      RECT 16.475 3.685 17.205 4.015 ;
      RECT 8.79 2.005 9.52 2.335 ;
      RECT 6.57 3.685 7.3 4.015 ;
      RECT 4.87 3.685 5.6 4.015 ;
      RECT -0.085 2.565 0.645 2.895 ;
      RECT -1.45 3.685 -0.72 4.015 ;
    LAYER via2 ;
      RECT 82.265 1.225 82.465 1.425 ;
      RECT 80.555 2.07 80.755 2.27 ;
      RECT 79.595 3.75 79.795 3.95 ;
      RECT 79.445 7.14 79.645 7.34 ;
      RECT 78.595 3.75 78.795 3.95 ;
      RECT 76.635 3.75 76.835 3.95 ;
      RECT 75.435 3.19 75.635 3.39 ;
      RECT 74.195 2.63 74.395 2.83 ;
      RECT 74.185 1.045 74.385 1.245 ;
      RECT 72.755 3.19 72.955 3.39 ;
      RECT 72.75 1.04 72.95 1.24 ;
      RECT 72.015 2.63 72.215 2.83 ;
      RECT 70.795 2.63 70.995 2.83 ;
      RECT 70.78 1.015 70.98 1.215 ;
      RECT 70.315 3.75 70.515 3.95 ;
      RECT 64.34 1.225 64.54 1.425 ;
      RECT 62.63 2.07 62.83 2.27 ;
      RECT 61.67 3.75 61.87 3.95 ;
      RECT 61.52 7.14 61.72 7.34 ;
      RECT 60.67 3.75 60.87 3.95 ;
      RECT 58.71 3.75 58.91 3.95 ;
      RECT 57.51 3.19 57.71 3.39 ;
      RECT 56.27 2.63 56.47 2.83 ;
      RECT 56.26 1.045 56.46 1.245 ;
      RECT 54.83 3.19 55.03 3.39 ;
      RECT 54.825 1.04 55.025 1.24 ;
      RECT 54.09 2.63 54.29 2.83 ;
      RECT 52.87 2.63 53.07 2.83 ;
      RECT 52.855 1.015 53.055 1.215 ;
      RECT 52.39 3.75 52.59 3.95 ;
      RECT 46.415 1.225 46.615 1.425 ;
      RECT 44.705 2.07 44.905 2.27 ;
      RECT 43.745 3.75 43.945 3.95 ;
      RECT 43.595 7.14 43.795 7.34 ;
      RECT 42.745 3.75 42.945 3.95 ;
      RECT 40.785 3.75 40.985 3.95 ;
      RECT 39.585 3.19 39.785 3.39 ;
      RECT 38.345 2.63 38.545 2.83 ;
      RECT 38.335 1.045 38.535 1.245 ;
      RECT 36.905 3.19 37.105 3.39 ;
      RECT 36.9 1.04 37.1 1.24 ;
      RECT 36.165 2.63 36.365 2.83 ;
      RECT 34.945 2.63 35.145 2.83 ;
      RECT 34.93 1.015 35.13 1.215 ;
      RECT 34.465 3.75 34.665 3.95 ;
      RECT 28.49 1.225 28.69 1.425 ;
      RECT 26.78 2.07 26.98 2.27 ;
      RECT 25.82 3.75 26.02 3.95 ;
      RECT 25.67 7.14 25.87 7.34 ;
      RECT 24.82 3.75 25.02 3.95 ;
      RECT 22.86 3.75 23.06 3.95 ;
      RECT 21.66 3.19 21.86 3.39 ;
      RECT 20.42 2.63 20.62 2.83 ;
      RECT 20.41 1.045 20.61 1.245 ;
      RECT 18.98 3.19 19.18 3.39 ;
      RECT 18.975 1.04 19.175 1.24 ;
      RECT 18.24 2.63 18.44 2.83 ;
      RECT 17.02 2.63 17.22 2.83 ;
      RECT 17.005 1.015 17.205 1.215 ;
      RECT 16.54 3.75 16.74 3.95 ;
      RECT 10.565 1.225 10.765 1.425 ;
      RECT 8.855 2.07 9.055 2.27 ;
      RECT 7.895 3.75 8.095 3.95 ;
      RECT 7.745 7.14 7.945 7.34 ;
      RECT 6.895 3.75 7.095 3.95 ;
      RECT 4.935 3.75 5.135 3.95 ;
      RECT 3.735 3.19 3.935 3.39 ;
      RECT 2.495 2.63 2.695 2.83 ;
      RECT 2.485 1.045 2.685 1.245 ;
      RECT 1.055 3.19 1.255 3.39 ;
      RECT 1.05 1.04 1.25 1.24 ;
      RECT 0.315 2.63 0.515 2.83 ;
      RECT -0.905 2.63 -0.705 2.83 ;
      RECT -0.92 1.015 -0.72 1.215 ;
      RECT -1.385 3.75 -1.185 3.95 ;
    LAYER met2 ;
      RECT -3.645 8.4 87.175 8.57 ;
      RECT 87.005 7.275 87.175 8.57 ;
      RECT -3.645 6.255 -3.475 8.57 ;
      RECT 86.975 7.275 87.325 7.625 ;
      RECT -3.7 6.255 -3.41 6.605 ;
      RECT 83.82 6.225 84.14 6.545 ;
      RECT 83.85 5.695 84.02 6.545 ;
      RECT 83.85 5.695 84.025 6.045 ;
      RECT 83.85 5.695 84.825 5.87 ;
      RECT 84.65 1.965 84.825 5.87 ;
      RECT 84.595 1.965 84.945 2.315 ;
      RECT 84.62 6.655 84.945 6.98 ;
      RECT 83.505 6.745 84.945 6.915 ;
      RECT 83.505 2.395 83.665 6.915 ;
      RECT 83.82 2.365 84.14 2.685 ;
      RECT 83.505 2.395 84.14 2.565 ;
      RECT 82.765 5.84 83.115 6.19 ;
      RECT 82.84 2.705 83.015 6.19 ;
      RECT 82.775 2.705 83.125 3.055 ;
      RECT 82.175 1.14 82.55 1.51 ;
      RECT 74.095 0.96 74.47 1.33 ;
      RECT 72.66 0.96 73.035 1.33 ;
      RECT 72.66 1.08 82.48 1.25 ;
      RECT 78.605 4.36 82.46 4.53 ;
      RECT 82.29 3.425 82.46 4.53 ;
      RECT 78.605 3.67 78.775 4.53 ;
      RECT 78.555 3.71 78.835 3.99 ;
      RECT 78.575 3.67 78.835 3.99 ;
      RECT 78.215 3.625 78.32 3.885 ;
      RECT 82.2 3.43 82.55 3.78 ;
      RECT 78.07 2.115 78.16 2.375 ;
      RECT 78.61 3.18 78.615 3.22 ;
      RECT 78.605 3.17 78.61 3.305 ;
      RECT 78.6 3.16 78.605 3.398 ;
      RECT 78.59 3.14 78.6 3.454 ;
      RECT 78.51 3.068 78.59 3.534 ;
      RECT 78.545 3.712 78.555 3.937 ;
      RECT 78.54 3.709 78.545 3.932 ;
      RECT 78.525 3.706 78.54 3.925 ;
      RECT 78.49 3.7 78.525 3.907 ;
      RECT 78.505 3.003 78.51 3.608 ;
      RECT 78.485 2.954 78.505 3.623 ;
      RECT 78.475 3.687 78.49 3.89 ;
      RECT 78.48 2.896 78.485 3.638 ;
      RECT 78.475 2.874 78.48 3.648 ;
      RECT 78.44 2.784 78.475 3.885 ;
      RECT 78.425 2.662 78.44 3.885 ;
      RECT 78.42 2.615 78.425 3.885 ;
      RECT 78.395 2.54 78.42 3.885 ;
      RECT 78.38 2.455 78.395 3.885 ;
      RECT 78.375 2.402 78.38 3.885 ;
      RECT 78.37 2.382 78.375 3.885 ;
      RECT 78.365 2.357 78.37 3.119 ;
      RECT 78.35 3.317 78.37 3.885 ;
      RECT 78.36 2.335 78.365 3.096 ;
      RECT 78.35 2.287 78.36 3.061 ;
      RECT 78.345 2.25 78.35 3.027 ;
      RECT 78.345 3.397 78.35 3.885 ;
      RECT 78.33 2.227 78.345 2.982 ;
      RECT 78.325 3.495 78.345 3.885 ;
      RECT 78.275 2.115 78.33 2.824 ;
      RECT 78.32 3.617 78.325 3.885 ;
      RECT 78.26 2.115 78.275 2.663 ;
      RECT 78.255 2.115 78.26 2.615 ;
      RECT 78.25 2.115 78.255 2.603 ;
      RECT 78.205 2.115 78.25 2.54 ;
      RECT 78.18 2.115 78.205 2.458 ;
      RECT 78.165 2.115 78.18 2.41 ;
      RECT 78.16 2.115 78.165 2.38 ;
      RECT 80.55 2.16 80.81 2.42 ;
      RECT 80.545 2.16 80.81 2.368 ;
      RECT 80.54 2.16 80.81 2.338 ;
      RECT 80.515 2.03 80.795 2.31 ;
      RECT 69.03 6.655 69.38 7.005 ;
      RECT 80.275 6.61 80.625 6.96 ;
      RECT 69.03 6.685 80.625 6.885 ;
      RECT 79.555 3.71 79.835 3.99 ;
      RECT 79.595 3.665 79.86 3.925 ;
      RECT 79.585 3.7 79.86 3.925 ;
      RECT 79.59 3.685 79.835 3.99 ;
      RECT 79.595 3.662 79.805 3.99 ;
      RECT 79.595 3.66 79.79 3.99 ;
      RECT 79.635 3.65 79.79 3.99 ;
      RECT 79.605 3.655 79.79 3.99 ;
      RECT 79.635 3.647 79.735 3.99 ;
      RECT 79.66 3.64 79.735 3.99 ;
      RECT 79.64 3.642 79.735 3.99 ;
      RECT 78.97 3.155 79.23 3.415 ;
      RECT 79.02 3.147 79.21 3.415 ;
      RECT 79.025 3.067 79.21 3.415 ;
      RECT 79.145 2.455 79.21 3.415 ;
      RECT 79.05 2.852 79.21 3.415 ;
      RECT 79.125 2.54 79.21 3.415 ;
      RECT 79.16 2.165 79.296 2.893 ;
      RECT 79.105 2.662 79.296 2.893 ;
      RECT 79.12 2.602 79.21 3.415 ;
      RECT 79.16 2.165 79.32 2.558 ;
      RECT 79.16 2.165 79.33 2.455 ;
      RECT 79.15 2.165 79.41 2.425 ;
      RECT 77.485 3.565 77.53 3.825 ;
      RECT 77.39 2.1 77.535 2.36 ;
      RECT 77.895 2.722 77.905 2.813 ;
      RECT 77.88 2.66 77.895 2.869 ;
      RECT 77.875 2.607 77.88 2.915 ;
      RECT 77.825 2.554 77.875 3.041 ;
      RECT 77.82 2.509 77.825 3.188 ;
      RECT 77.81 2.497 77.82 3.23 ;
      RECT 77.775 2.461 77.81 3.335 ;
      RECT 77.77 2.429 77.775 3.441 ;
      RECT 77.755 2.411 77.77 3.486 ;
      RECT 77.75 2.394 77.755 2.72 ;
      RECT 77.745 2.775 77.755 3.543 ;
      RECT 77.74 2.38 77.75 2.693 ;
      RECT 77.735 2.83 77.745 3.825 ;
      RECT 77.73 2.366 77.74 2.678 ;
      RECT 77.73 2.88 77.735 3.825 ;
      RECT 77.715 2.343 77.73 2.658 ;
      RECT 77.695 3.002 77.73 3.825 ;
      RECT 77.71 2.325 77.715 2.64 ;
      RECT 77.705 2.317 77.71 2.63 ;
      RECT 77.675 2.285 77.705 2.594 ;
      RECT 77.685 3.13 77.695 3.825 ;
      RECT 77.68 3.157 77.685 3.825 ;
      RECT 77.675 3.207 77.68 3.825 ;
      RECT 77.665 2.251 77.675 2.559 ;
      RECT 77.625 3.275 77.675 3.825 ;
      RECT 77.65 2.228 77.665 2.535 ;
      RECT 77.625 2.1 77.65 2.498 ;
      RECT 77.62 2.1 77.625 2.47 ;
      RECT 77.59 3.375 77.625 3.825 ;
      RECT 77.615 2.1 77.62 2.463 ;
      RECT 77.61 2.1 77.615 2.453 ;
      RECT 77.595 2.1 77.61 2.438 ;
      RECT 77.58 2.1 77.595 2.41 ;
      RECT 77.545 3.48 77.59 3.825 ;
      RECT 77.565 2.1 77.58 2.383 ;
      RECT 77.535 2.1 77.565 2.368 ;
      RECT 77.53 3.552 77.545 3.825 ;
      RECT 77.455 2.635 77.495 2.895 ;
      RECT 77.23 2.582 77.235 2.84 ;
      RECT 73.185 2.06 73.445 2.32 ;
      RECT 73.185 2.085 73.46 2.3 ;
      RECT 75.575 1.91 75.58 2.055 ;
      RECT 77.445 2.63 77.455 2.895 ;
      RECT 77.425 2.622 77.445 2.895 ;
      RECT 77.407 2.618 77.425 2.895 ;
      RECT 77.321 2.607 77.407 2.895 ;
      RECT 77.235 2.59 77.321 2.895 ;
      RECT 77.18 2.577 77.23 2.825 ;
      RECT 77.146 2.569 77.18 2.8 ;
      RECT 77.06 2.558 77.146 2.765 ;
      RECT 77.025 2.535 77.06 2.73 ;
      RECT 77.015 2.497 77.025 2.716 ;
      RECT 77.01 2.47 77.015 2.712 ;
      RECT 77.005 2.457 77.01 2.709 ;
      RECT 76.995 2.437 77.005 2.705 ;
      RECT 76.99 2.412 76.995 2.701 ;
      RECT 76.965 2.367 76.99 2.695 ;
      RECT 76.955 2.308 76.965 2.687 ;
      RECT 76.945 2.276 76.955 2.678 ;
      RECT 76.925 2.228 76.945 2.658 ;
      RECT 76.92 2.188 76.925 2.628 ;
      RECT 76.905 2.162 76.92 2.602 ;
      RECT 76.9 2.14 76.905 2.578 ;
      RECT 76.885 2.112 76.9 2.554 ;
      RECT 76.87 2.085 76.885 2.518 ;
      RECT 76.855 2.062 76.87 2.48 ;
      RECT 76.85 2.052 76.855 2.455 ;
      RECT 76.84 2.045 76.85 2.438 ;
      RECT 76.825 2.032 76.84 2.408 ;
      RECT 76.82 2.022 76.825 2.383 ;
      RECT 76.815 2.017 76.82 2.37 ;
      RECT 76.805 2.01 76.815 2.35 ;
      RECT 76.8 2.003 76.805 2.335 ;
      RECT 76.775 1.996 76.8 2.293 ;
      RECT 76.76 1.986 76.775 2.243 ;
      RECT 76.75 1.981 76.76 2.213 ;
      RECT 76.74 1.977 76.75 2.188 ;
      RECT 76.725 1.974 76.74 2.178 ;
      RECT 76.675 1.971 76.725 2.163 ;
      RECT 76.655 1.969 76.675 2.148 ;
      RECT 76.606 1.967 76.655 2.143 ;
      RECT 76.52 1.963 76.606 2.138 ;
      RECT 76.481 1.96 76.52 2.134 ;
      RECT 76.395 1.956 76.481 2.129 ;
      RECT 76.345 1.953 76.395 2.123 ;
      RECT 76.296 1.95 76.345 2.118 ;
      RECT 76.21 1.947 76.296 2.113 ;
      RECT 76.206 1.945 76.21 2.11 ;
      RECT 76.12 1.942 76.206 2.105 ;
      RECT 76.071 1.938 76.12 2.098 ;
      RECT 75.985 1.935 76.071 2.093 ;
      RECT 75.961 1.932 75.985 2.089 ;
      RECT 75.875 1.93 75.961 2.084 ;
      RECT 75.81 1.926 75.875 2.077 ;
      RECT 75.807 1.925 75.81 2.074 ;
      RECT 75.721 1.922 75.807 2.071 ;
      RECT 75.635 1.916 75.721 2.064 ;
      RECT 75.605 1.912 75.635 2.06 ;
      RECT 75.58 1.91 75.605 2.058 ;
      RECT 75.525 1.907 75.575 2.055 ;
      RECT 75.445 1.906 75.525 2.055 ;
      RECT 75.39 1.908 75.445 2.058 ;
      RECT 75.375 1.909 75.39 2.062 ;
      RECT 75.32 1.917 75.375 2.072 ;
      RECT 75.29 1.925 75.32 2.085 ;
      RECT 75.271 1.926 75.29 2.091 ;
      RECT 75.185 1.929 75.271 2.096 ;
      RECT 75.115 1.934 75.185 2.105 ;
      RECT 75.096 1.937 75.115 2.111 ;
      RECT 75.01 1.941 75.096 2.116 ;
      RECT 74.97 1.945 75.01 2.123 ;
      RECT 74.961 1.947 74.97 2.126 ;
      RECT 74.875 1.951 74.961 2.131 ;
      RECT 74.872 1.954 74.875 2.135 ;
      RECT 74.786 1.957 74.872 2.139 ;
      RECT 74.7 1.963 74.786 2.147 ;
      RECT 74.676 1.967 74.7 2.151 ;
      RECT 74.59 1.971 74.676 2.156 ;
      RECT 74.545 1.976 74.59 2.163 ;
      RECT 74.465 1.981 74.545 2.17 ;
      RECT 74.385 1.987 74.465 2.185 ;
      RECT 74.36 1.991 74.385 2.198 ;
      RECT 74.295 1.994 74.36 2.21 ;
      RECT 74.24 1.999 74.295 2.225 ;
      RECT 74.21 2.002 74.24 2.243 ;
      RECT 74.2 2.004 74.21 2.256 ;
      RECT 74.14 2.019 74.2 2.266 ;
      RECT 74.125 2.036 74.14 2.275 ;
      RECT 74.12 2.045 74.125 2.275 ;
      RECT 74.11 2.055 74.12 2.275 ;
      RECT 74.1 2.072 74.11 2.275 ;
      RECT 74.08 2.082 74.1 2.276 ;
      RECT 74.035 2.092 74.08 2.277 ;
      RECT 74 2.101 74.035 2.279 ;
      RECT 73.935 2.106 74 2.281 ;
      RECT 73.855 2.107 73.935 2.284 ;
      RECT 73.851 2.105 73.855 2.285 ;
      RECT 73.765 2.102 73.851 2.287 ;
      RECT 73.718 2.099 73.765 2.289 ;
      RECT 73.632 2.095 73.718 2.292 ;
      RECT 73.546 2.091 73.632 2.295 ;
      RECT 73.46 2.087 73.546 2.299 ;
      RECT 76.845 3.71 76.875 3.99 ;
      RECT 76.595 3.6 76.615 3.99 ;
      RECT 76.55 3.6 76.615 3.86 ;
      RECT 76.38 2.225 76.415 2.485 ;
      RECT 76.155 2.225 76.215 2.485 ;
      RECT 76.835 3.69 76.845 3.99 ;
      RECT 76.83 3.65 76.835 3.99 ;
      RECT 76.815 3.605 76.83 3.99 ;
      RECT 76.81 3.57 76.815 3.99 ;
      RECT 76.805 3.55 76.81 3.99 ;
      RECT 76.775 3.477 76.805 3.99 ;
      RECT 76.755 3.375 76.775 3.99 ;
      RECT 76.745 3.305 76.755 3.99 ;
      RECT 76.7 3.245 76.745 3.99 ;
      RECT 76.615 3.206 76.7 3.99 ;
      RECT 76.61 3.197 76.615 3.57 ;
      RECT 76.6 3.196 76.61 3.553 ;
      RECT 76.575 3.177 76.6 3.523 ;
      RECT 76.57 3.152 76.575 3.502 ;
      RECT 76.56 3.13 76.57 3.493 ;
      RECT 76.555 3.101 76.56 3.483 ;
      RECT 76.515 3.027 76.555 3.455 ;
      RECT 76.495 2.928 76.515 3.42 ;
      RECT 76.48 2.864 76.495 3.403 ;
      RECT 76.45 2.788 76.48 3.375 ;
      RECT 76.43 2.703 76.45 3.348 ;
      RECT 76.39 2.599 76.43 3.255 ;
      RECT 76.385 2.52 76.39 3.163 ;
      RECT 76.38 2.503 76.385 3.14 ;
      RECT 76.375 2.225 76.38 3.12 ;
      RECT 76.345 2.225 76.375 3.058 ;
      RECT 76.34 2.225 76.345 2.99 ;
      RECT 76.33 2.225 76.34 2.955 ;
      RECT 76.32 2.225 76.33 2.92 ;
      RECT 76.255 2.225 76.32 2.775 ;
      RECT 76.25 2.225 76.255 2.645 ;
      RECT 76.22 2.225 76.25 2.578 ;
      RECT 76.215 2.225 76.22 2.503 ;
      RECT 75.395 3.15 75.675 3.43 ;
      RECT 75.435 3.13 75.695 3.39 ;
      RECT 75.425 3.14 75.695 3.39 ;
      RECT 75.435 3.067 75.65 3.43 ;
      RECT 75.49 2.99 75.645 3.43 ;
      RECT 75.495 2.775 75.645 3.43 ;
      RECT 75.485 2.577 75.635 2.828 ;
      RECT 75.475 2.577 75.635 2.695 ;
      RECT 75.47 2.455 75.63 2.598 ;
      RECT 75.455 2.455 75.63 2.503 ;
      RECT 75.45 2.165 75.625 2.48 ;
      RECT 75.435 2.165 75.625 2.45 ;
      RECT 75.395 2.165 75.655 2.425 ;
      RECT 75.305 3.635 75.385 3.895 ;
      RECT 74.71 2.355 74.715 2.62 ;
      RECT 74.59 2.355 74.715 2.615 ;
      RECT 75.265 3.6 75.305 3.895 ;
      RECT 75.22 3.522 75.265 3.895 ;
      RECT 75.2 3.45 75.22 3.895 ;
      RECT 75.19 3.402 75.2 3.895 ;
      RECT 75.155 3.335 75.19 3.895 ;
      RECT 75.125 3.235 75.155 3.895 ;
      RECT 75.105 3.16 75.125 3.695 ;
      RECT 75.095 3.11 75.105 3.65 ;
      RECT 75.09 3.087 75.095 3.623 ;
      RECT 75.085 3.072 75.09 3.61 ;
      RECT 75.08 3.057 75.085 3.588 ;
      RECT 75.075 3.042 75.08 3.57 ;
      RECT 75.05 2.997 75.075 3.525 ;
      RECT 75.04 2.945 75.05 3.468 ;
      RECT 75.03 2.915 75.04 3.435 ;
      RECT 75.02 2.88 75.03 3.403 ;
      RECT 74.985 2.812 75.02 3.335 ;
      RECT 74.98 2.751 74.985 3.27 ;
      RECT 74.97 2.739 74.98 3.25 ;
      RECT 74.965 2.727 74.97 3.23 ;
      RECT 74.96 2.719 74.965 3.218 ;
      RECT 74.955 2.711 74.96 3.198 ;
      RECT 74.945 2.699 74.955 3.17 ;
      RECT 74.935 2.683 74.945 3.14 ;
      RECT 74.91 2.655 74.935 3.078 ;
      RECT 74.9 2.626 74.91 3.023 ;
      RECT 74.885 2.605 74.9 2.983 ;
      RECT 74.88 2.589 74.885 2.955 ;
      RECT 74.875 2.577 74.88 2.945 ;
      RECT 74.87 2.572 74.875 2.918 ;
      RECT 74.865 2.565 74.87 2.905 ;
      RECT 74.85 2.548 74.865 2.878 ;
      RECT 74.84 2.355 74.85 2.838 ;
      RECT 74.83 2.355 74.84 2.805 ;
      RECT 74.82 2.355 74.83 2.78 ;
      RECT 74.75 2.355 74.82 2.715 ;
      RECT 74.74 2.355 74.75 2.663 ;
      RECT 74.725 2.355 74.74 2.645 ;
      RECT 74.715 2.355 74.725 2.63 ;
      RECT 74.545 3.225 74.805 3.485 ;
      RECT 73.08 3.26 73.085 3.467 ;
      RECT 72.715 3.15 72.79 3.465 ;
      RECT 72.53 3.205 72.685 3.465 ;
      RECT 72.715 3.15 72.82 3.43 ;
      RECT 74.53 3.322 74.545 3.483 ;
      RECT 74.505 3.33 74.53 3.488 ;
      RECT 74.48 3.337 74.505 3.493 ;
      RECT 74.417 3.348 74.48 3.502 ;
      RECT 74.331 3.367 74.417 3.519 ;
      RECT 74.245 3.389 74.331 3.538 ;
      RECT 74.23 3.402 74.245 3.549 ;
      RECT 74.19 3.41 74.23 3.556 ;
      RECT 74.17 3.415 74.19 3.563 ;
      RECT 74.132 3.416 74.17 3.566 ;
      RECT 74.046 3.419 74.132 3.567 ;
      RECT 73.96 3.423 74.046 3.568 ;
      RECT 73.911 3.425 73.96 3.57 ;
      RECT 73.825 3.425 73.911 3.572 ;
      RECT 73.785 3.42 73.825 3.574 ;
      RECT 73.775 3.414 73.785 3.575 ;
      RECT 73.735 3.409 73.775 3.572 ;
      RECT 73.725 3.402 73.735 3.568 ;
      RECT 73.71 3.398 73.725 3.566 ;
      RECT 73.693 3.394 73.71 3.564 ;
      RECT 73.607 3.384 73.693 3.556 ;
      RECT 73.521 3.366 73.607 3.542 ;
      RECT 73.435 3.349 73.521 3.528 ;
      RECT 73.41 3.337 73.435 3.519 ;
      RECT 73.34 3.327 73.41 3.512 ;
      RECT 73.295 3.315 73.34 3.503 ;
      RECT 73.235 3.302 73.295 3.495 ;
      RECT 73.23 3.294 73.235 3.49 ;
      RECT 73.195 3.289 73.23 3.488 ;
      RECT 73.14 3.28 73.195 3.481 ;
      RECT 73.1 3.269 73.14 3.473 ;
      RECT 73.085 3.262 73.1 3.469 ;
      RECT 73.065 3.255 73.08 3.466 ;
      RECT 73.05 3.245 73.065 3.464 ;
      RECT 73.035 3.232 73.05 3.461 ;
      RECT 73.01 3.215 73.035 3.457 ;
      RECT 72.995 3.197 73.01 3.454 ;
      RECT 72.97 3.15 72.995 3.452 ;
      RECT 72.946 3.15 72.97 3.449 ;
      RECT 72.86 3.15 72.946 3.441 ;
      RECT 72.82 3.15 72.86 3.433 ;
      RECT 72.685 3.197 72.715 3.465 ;
      RECT 74.365 2.78 74.625 3.04 ;
      RECT 74.325 2.78 74.625 2.918 ;
      RECT 74.29 2.78 74.625 2.903 ;
      RECT 74.235 2.78 74.625 2.883 ;
      RECT 74.155 2.59 74.435 2.87 ;
      RECT 74.155 2.772 74.505 2.87 ;
      RECT 74.155 2.715 74.49 2.87 ;
      RECT 74.155 2.662 74.44 2.87 ;
      RECT 71.985 2.59 72.18 3.375 ;
      RECT 72.065 1.205 72.18 3.375 ;
      RECT 71.92 3.115 71.98 3.375 ;
      RECT 73.29 2.635 73.55 2.895 ;
      RECT 71.975 2.59 72.18 2.87 ;
      RECT 73.285 2.645 73.55 2.83 ;
      RECT 73 2.62 73.01 2.77 ;
      RECT 72.235 1.205 72.315 1.55 ;
      RECT 71.97 1.205 72.18 1.55 ;
      RECT 73.275 2.645 73.285 2.829 ;
      RECT 73.265 2.644 73.275 2.826 ;
      RECT 73.256 2.643 73.265 2.824 ;
      RECT 73.17 2.639 73.256 2.814 ;
      RECT 73.096 2.631 73.17 2.796 ;
      RECT 73.01 2.624 73.096 2.779 ;
      RECT 72.95 2.62 73 2.769 ;
      RECT 72.915 2.619 72.95 2.766 ;
      RECT 72.86 2.619 72.915 2.768 ;
      RECT 72.825 2.619 72.86 2.772 ;
      RECT 72.739 2.618 72.825 2.779 ;
      RECT 72.653 2.617 72.739 2.789 ;
      RECT 72.567 2.616 72.653 2.8 ;
      RECT 72.481 2.616 72.567 2.81 ;
      RECT 72.395 2.615 72.481 2.82 ;
      RECT 72.36 2.615 72.395 2.86 ;
      RECT 72.355 2.615 72.36 2.903 ;
      RECT 72.33 2.615 72.355 2.92 ;
      RECT 72.255 2.615 72.33 2.935 ;
      RECT 72.235 2.59 72.255 2.948 ;
      RECT 72.23 1.205 72.235 2.958 ;
      RECT 72.205 1.205 72.23 3 ;
      RECT 72.18 1.205 72.205 3.078 ;
      RECT 71.98 2.997 71.985 3.375 ;
      RECT 71.315 2.949 71.33 3.405 ;
      RECT 71.31 3.021 71.416 3.403 ;
      RECT 71.33 2.115 71.465 3.401 ;
      RECT 71.315 2.965 71.47 3.4 ;
      RECT 71.315 3.015 71.475 3.398 ;
      RECT 71.3 3.08 71.475 3.397 ;
      RECT 71.31 3.072 71.48 3.394 ;
      RECT 71.29 3.12 71.48 3.389 ;
      RECT 71.29 3.12 71.495 3.386 ;
      RECT 71.285 3.12 71.495 3.383 ;
      RECT 71.26 3.12 71.52 3.38 ;
      RECT 71.33 2.115 71.49 2.768 ;
      RECT 71.325 2.115 71.49 2.74 ;
      RECT 71.32 2.115 71.49 2.568 ;
      RECT 71.32 2.115 71.51 2.508 ;
      RECT 71.275 2.115 71.535 2.375 ;
      RECT 70.755 2.59 71.035 2.87 ;
      RECT 70.745 2.605 71.035 2.865 ;
      RECT 70.7 2.667 71.035 2.863 ;
      RECT 70.775 2.582 70.94 2.87 ;
      RECT 70.775 2.567 70.896 2.87 ;
      RECT 70.81 2.56 70.896 2.87 ;
      RECT 70.275 3.71 70.555 3.99 ;
      RECT 70.235 3.672 70.53 3.783 ;
      RECT 70.22 3.622 70.51 3.678 ;
      RECT 70.165 3.385 70.425 3.645 ;
      RECT 70.165 3.587 70.505 3.645 ;
      RECT 70.165 3.527 70.5 3.645 ;
      RECT 70.165 3.477 70.48 3.645 ;
      RECT 70.165 3.457 70.475 3.645 ;
      RECT 70.165 3.435 70.47 3.645 ;
      RECT 70.165 3.42 70.44 3.645 ;
      RECT 65.895 6.225 66.215 6.545 ;
      RECT 65.925 5.695 66.095 6.545 ;
      RECT 65.925 5.695 66.1 6.045 ;
      RECT 65.925 5.695 66.9 5.87 ;
      RECT 66.725 1.965 66.9 5.87 ;
      RECT 66.67 1.965 67.02 2.315 ;
      RECT 66.695 6.655 67.02 6.98 ;
      RECT 65.58 6.745 67.02 6.915 ;
      RECT 65.58 2.395 65.74 6.915 ;
      RECT 65.895 2.365 66.215 2.685 ;
      RECT 65.58 2.395 66.215 2.565 ;
      RECT 64.84 5.84 65.19 6.19 ;
      RECT 64.915 2.705 65.09 6.19 ;
      RECT 64.85 2.705 65.2 3.055 ;
      RECT 64.25 1.14 64.625 1.51 ;
      RECT 56.17 0.96 56.545 1.33 ;
      RECT 54.735 0.96 55.11 1.33 ;
      RECT 54.735 1.08 64.555 1.25 ;
      RECT 60.68 4.36 64.535 4.53 ;
      RECT 64.365 3.425 64.535 4.53 ;
      RECT 60.68 3.67 60.85 4.53 ;
      RECT 60.63 3.71 60.91 3.99 ;
      RECT 60.65 3.67 60.91 3.99 ;
      RECT 60.29 3.625 60.395 3.885 ;
      RECT 64.275 3.43 64.625 3.78 ;
      RECT 60.145 2.115 60.235 2.375 ;
      RECT 60.685 3.18 60.69 3.22 ;
      RECT 60.68 3.17 60.685 3.305 ;
      RECT 60.675 3.16 60.68 3.398 ;
      RECT 60.665 3.14 60.675 3.454 ;
      RECT 60.585 3.068 60.665 3.534 ;
      RECT 60.62 3.712 60.63 3.937 ;
      RECT 60.615 3.709 60.62 3.932 ;
      RECT 60.6 3.706 60.615 3.925 ;
      RECT 60.565 3.7 60.6 3.907 ;
      RECT 60.58 3.003 60.585 3.608 ;
      RECT 60.56 2.954 60.58 3.623 ;
      RECT 60.55 3.687 60.565 3.89 ;
      RECT 60.555 2.896 60.56 3.638 ;
      RECT 60.55 2.874 60.555 3.648 ;
      RECT 60.515 2.784 60.55 3.885 ;
      RECT 60.5 2.662 60.515 3.885 ;
      RECT 60.495 2.615 60.5 3.885 ;
      RECT 60.47 2.54 60.495 3.885 ;
      RECT 60.455 2.455 60.47 3.885 ;
      RECT 60.45 2.402 60.455 3.885 ;
      RECT 60.445 2.382 60.45 3.885 ;
      RECT 60.44 2.357 60.445 3.119 ;
      RECT 60.425 3.317 60.445 3.885 ;
      RECT 60.435 2.335 60.44 3.096 ;
      RECT 60.425 2.287 60.435 3.061 ;
      RECT 60.42 2.25 60.425 3.027 ;
      RECT 60.42 3.397 60.425 3.885 ;
      RECT 60.405 2.227 60.42 2.982 ;
      RECT 60.4 3.495 60.42 3.885 ;
      RECT 60.35 2.115 60.405 2.824 ;
      RECT 60.395 3.617 60.4 3.885 ;
      RECT 60.335 2.115 60.35 2.663 ;
      RECT 60.33 2.115 60.335 2.615 ;
      RECT 60.325 2.115 60.33 2.603 ;
      RECT 60.28 2.115 60.325 2.54 ;
      RECT 60.255 2.115 60.28 2.458 ;
      RECT 60.24 2.115 60.255 2.41 ;
      RECT 60.235 2.115 60.24 2.38 ;
      RECT 62.625 2.16 62.885 2.42 ;
      RECT 62.62 2.16 62.885 2.368 ;
      RECT 62.615 2.16 62.885 2.338 ;
      RECT 62.59 2.03 62.87 2.31 ;
      RECT 51.105 6.655 51.455 7.005 ;
      RECT 62.07 6.61 62.42 6.96 ;
      RECT 51.105 6.685 62.42 6.885 ;
      RECT 61.63 3.71 61.91 3.99 ;
      RECT 61.67 3.665 61.935 3.925 ;
      RECT 61.66 3.7 61.935 3.925 ;
      RECT 61.665 3.685 61.91 3.99 ;
      RECT 61.67 3.662 61.88 3.99 ;
      RECT 61.67 3.66 61.865 3.99 ;
      RECT 61.71 3.65 61.865 3.99 ;
      RECT 61.68 3.655 61.865 3.99 ;
      RECT 61.71 3.647 61.81 3.99 ;
      RECT 61.735 3.64 61.81 3.99 ;
      RECT 61.715 3.642 61.81 3.99 ;
      RECT 61.045 3.155 61.305 3.415 ;
      RECT 61.095 3.147 61.285 3.415 ;
      RECT 61.1 3.067 61.285 3.415 ;
      RECT 61.22 2.455 61.285 3.415 ;
      RECT 61.125 2.852 61.285 3.415 ;
      RECT 61.2 2.54 61.285 3.415 ;
      RECT 61.235 2.165 61.371 2.893 ;
      RECT 61.18 2.662 61.371 2.893 ;
      RECT 61.195 2.602 61.285 3.415 ;
      RECT 61.235 2.165 61.395 2.558 ;
      RECT 61.235 2.165 61.405 2.455 ;
      RECT 61.225 2.165 61.485 2.425 ;
      RECT 59.56 3.565 59.605 3.825 ;
      RECT 59.465 2.1 59.61 2.36 ;
      RECT 59.97 2.722 59.98 2.813 ;
      RECT 59.955 2.66 59.97 2.869 ;
      RECT 59.95 2.607 59.955 2.915 ;
      RECT 59.9 2.554 59.95 3.041 ;
      RECT 59.895 2.509 59.9 3.188 ;
      RECT 59.885 2.497 59.895 3.23 ;
      RECT 59.85 2.461 59.885 3.335 ;
      RECT 59.845 2.429 59.85 3.441 ;
      RECT 59.83 2.411 59.845 3.486 ;
      RECT 59.825 2.394 59.83 2.72 ;
      RECT 59.82 2.775 59.83 3.543 ;
      RECT 59.815 2.38 59.825 2.693 ;
      RECT 59.81 2.83 59.82 3.825 ;
      RECT 59.805 2.366 59.815 2.678 ;
      RECT 59.805 2.88 59.81 3.825 ;
      RECT 59.79 2.343 59.805 2.658 ;
      RECT 59.77 3.002 59.805 3.825 ;
      RECT 59.785 2.325 59.79 2.64 ;
      RECT 59.78 2.317 59.785 2.63 ;
      RECT 59.75 2.285 59.78 2.594 ;
      RECT 59.76 3.13 59.77 3.825 ;
      RECT 59.755 3.157 59.76 3.825 ;
      RECT 59.75 3.207 59.755 3.825 ;
      RECT 59.74 2.251 59.75 2.559 ;
      RECT 59.7 3.275 59.75 3.825 ;
      RECT 59.725 2.228 59.74 2.535 ;
      RECT 59.7 2.1 59.725 2.498 ;
      RECT 59.695 2.1 59.7 2.47 ;
      RECT 59.665 3.375 59.7 3.825 ;
      RECT 59.69 2.1 59.695 2.463 ;
      RECT 59.685 2.1 59.69 2.453 ;
      RECT 59.67 2.1 59.685 2.438 ;
      RECT 59.655 2.1 59.67 2.41 ;
      RECT 59.62 3.48 59.665 3.825 ;
      RECT 59.64 2.1 59.655 2.383 ;
      RECT 59.61 2.1 59.64 2.368 ;
      RECT 59.605 3.552 59.62 3.825 ;
      RECT 59.53 2.635 59.57 2.895 ;
      RECT 59.305 2.582 59.31 2.84 ;
      RECT 55.26 2.06 55.52 2.32 ;
      RECT 55.26 2.085 55.535 2.3 ;
      RECT 57.65 1.91 57.655 2.055 ;
      RECT 59.52 2.63 59.53 2.895 ;
      RECT 59.5 2.622 59.52 2.895 ;
      RECT 59.482 2.618 59.5 2.895 ;
      RECT 59.396 2.607 59.482 2.895 ;
      RECT 59.31 2.59 59.396 2.895 ;
      RECT 59.255 2.577 59.305 2.825 ;
      RECT 59.221 2.569 59.255 2.8 ;
      RECT 59.135 2.558 59.221 2.765 ;
      RECT 59.1 2.535 59.135 2.73 ;
      RECT 59.09 2.497 59.1 2.716 ;
      RECT 59.085 2.47 59.09 2.712 ;
      RECT 59.08 2.457 59.085 2.709 ;
      RECT 59.07 2.437 59.08 2.705 ;
      RECT 59.065 2.412 59.07 2.701 ;
      RECT 59.04 2.367 59.065 2.695 ;
      RECT 59.03 2.308 59.04 2.687 ;
      RECT 59.02 2.276 59.03 2.678 ;
      RECT 59 2.228 59.02 2.658 ;
      RECT 58.995 2.188 59 2.628 ;
      RECT 58.98 2.162 58.995 2.602 ;
      RECT 58.975 2.14 58.98 2.578 ;
      RECT 58.96 2.112 58.975 2.554 ;
      RECT 58.945 2.085 58.96 2.518 ;
      RECT 58.93 2.062 58.945 2.48 ;
      RECT 58.925 2.052 58.93 2.455 ;
      RECT 58.915 2.045 58.925 2.438 ;
      RECT 58.9 2.032 58.915 2.408 ;
      RECT 58.895 2.022 58.9 2.383 ;
      RECT 58.89 2.017 58.895 2.37 ;
      RECT 58.88 2.01 58.89 2.35 ;
      RECT 58.875 2.003 58.88 2.335 ;
      RECT 58.85 1.996 58.875 2.293 ;
      RECT 58.835 1.986 58.85 2.243 ;
      RECT 58.825 1.981 58.835 2.213 ;
      RECT 58.815 1.977 58.825 2.188 ;
      RECT 58.8 1.974 58.815 2.178 ;
      RECT 58.75 1.971 58.8 2.163 ;
      RECT 58.73 1.969 58.75 2.148 ;
      RECT 58.681 1.967 58.73 2.143 ;
      RECT 58.595 1.963 58.681 2.138 ;
      RECT 58.556 1.96 58.595 2.134 ;
      RECT 58.47 1.956 58.556 2.129 ;
      RECT 58.42 1.953 58.47 2.123 ;
      RECT 58.371 1.95 58.42 2.118 ;
      RECT 58.285 1.947 58.371 2.113 ;
      RECT 58.281 1.945 58.285 2.11 ;
      RECT 58.195 1.942 58.281 2.105 ;
      RECT 58.146 1.938 58.195 2.098 ;
      RECT 58.06 1.935 58.146 2.093 ;
      RECT 58.036 1.932 58.06 2.089 ;
      RECT 57.95 1.93 58.036 2.084 ;
      RECT 57.885 1.926 57.95 2.077 ;
      RECT 57.882 1.925 57.885 2.074 ;
      RECT 57.796 1.922 57.882 2.071 ;
      RECT 57.71 1.916 57.796 2.064 ;
      RECT 57.68 1.912 57.71 2.06 ;
      RECT 57.655 1.91 57.68 2.058 ;
      RECT 57.6 1.907 57.65 2.055 ;
      RECT 57.52 1.906 57.6 2.055 ;
      RECT 57.465 1.908 57.52 2.058 ;
      RECT 57.45 1.909 57.465 2.062 ;
      RECT 57.395 1.917 57.45 2.072 ;
      RECT 57.365 1.925 57.395 2.085 ;
      RECT 57.346 1.926 57.365 2.091 ;
      RECT 57.26 1.929 57.346 2.096 ;
      RECT 57.19 1.934 57.26 2.105 ;
      RECT 57.171 1.937 57.19 2.111 ;
      RECT 57.085 1.941 57.171 2.116 ;
      RECT 57.045 1.945 57.085 2.123 ;
      RECT 57.036 1.947 57.045 2.126 ;
      RECT 56.95 1.951 57.036 2.131 ;
      RECT 56.947 1.954 56.95 2.135 ;
      RECT 56.861 1.957 56.947 2.139 ;
      RECT 56.775 1.963 56.861 2.147 ;
      RECT 56.751 1.967 56.775 2.151 ;
      RECT 56.665 1.971 56.751 2.156 ;
      RECT 56.62 1.976 56.665 2.163 ;
      RECT 56.54 1.981 56.62 2.17 ;
      RECT 56.46 1.987 56.54 2.185 ;
      RECT 56.435 1.991 56.46 2.198 ;
      RECT 56.37 1.994 56.435 2.21 ;
      RECT 56.315 1.999 56.37 2.225 ;
      RECT 56.285 2.002 56.315 2.243 ;
      RECT 56.275 2.004 56.285 2.256 ;
      RECT 56.215 2.019 56.275 2.266 ;
      RECT 56.2 2.036 56.215 2.275 ;
      RECT 56.195 2.045 56.2 2.275 ;
      RECT 56.185 2.055 56.195 2.275 ;
      RECT 56.175 2.072 56.185 2.275 ;
      RECT 56.155 2.082 56.175 2.276 ;
      RECT 56.11 2.092 56.155 2.277 ;
      RECT 56.075 2.101 56.11 2.279 ;
      RECT 56.01 2.106 56.075 2.281 ;
      RECT 55.93 2.107 56.01 2.284 ;
      RECT 55.926 2.105 55.93 2.285 ;
      RECT 55.84 2.102 55.926 2.287 ;
      RECT 55.793 2.099 55.84 2.289 ;
      RECT 55.707 2.095 55.793 2.292 ;
      RECT 55.621 2.091 55.707 2.295 ;
      RECT 55.535 2.087 55.621 2.299 ;
      RECT 58.92 3.71 58.95 3.99 ;
      RECT 58.67 3.6 58.69 3.99 ;
      RECT 58.625 3.6 58.69 3.86 ;
      RECT 58.455 2.225 58.49 2.485 ;
      RECT 58.23 2.225 58.29 2.485 ;
      RECT 58.91 3.69 58.92 3.99 ;
      RECT 58.905 3.65 58.91 3.99 ;
      RECT 58.89 3.605 58.905 3.99 ;
      RECT 58.885 3.57 58.89 3.99 ;
      RECT 58.88 3.55 58.885 3.99 ;
      RECT 58.85 3.477 58.88 3.99 ;
      RECT 58.83 3.375 58.85 3.99 ;
      RECT 58.82 3.305 58.83 3.99 ;
      RECT 58.775 3.245 58.82 3.99 ;
      RECT 58.69 3.206 58.775 3.99 ;
      RECT 58.685 3.197 58.69 3.57 ;
      RECT 58.675 3.196 58.685 3.553 ;
      RECT 58.65 3.177 58.675 3.523 ;
      RECT 58.645 3.152 58.65 3.502 ;
      RECT 58.635 3.13 58.645 3.493 ;
      RECT 58.63 3.101 58.635 3.483 ;
      RECT 58.59 3.027 58.63 3.455 ;
      RECT 58.57 2.928 58.59 3.42 ;
      RECT 58.555 2.864 58.57 3.403 ;
      RECT 58.525 2.788 58.555 3.375 ;
      RECT 58.505 2.703 58.525 3.348 ;
      RECT 58.465 2.599 58.505 3.255 ;
      RECT 58.46 2.52 58.465 3.163 ;
      RECT 58.455 2.503 58.46 3.14 ;
      RECT 58.45 2.225 58.455 3.12 ;
      RECT 58.42 2.225 58.45 3.058 ;
      RECT 58.415 2.225 58.42 2.99 ;
      RECT 58.405 2.225 58.415 2.955 ;
      RECT 58.395 2.225 58.405 2.92 ;
      RECT 58.33 2.225 58.395 2.775 ;
      RECT 58.325 2.225 58.33 2.645 ;
      RECT 58.295 2.225 58.325 2.578 ;
      RECT 58.29 2.225 58.295 2.503 ;
      RECT 57.47 3.15 57.75 3.43 ;
      RECT 57.51 3.13 57.77 3.39 ;
      RECT 57.5 3.14 57.77 3.39 ;
      RECT 57.51 3.067 57.725 3.43 ;
      RECT 57.565 2.99 57.72 3.43 ;
      RECT 57.57 2.775 57.72 3.43 ;
      RECT 57.56 2.577 57.71 2.828 ;
      RECT 57.55 2.577 57.71 2.695 ;
      RECT 57.545 2.455 57.705 2.598 ;
      RECT 57.53 2.455 57.705 2.503 ;
      RECT 57.525 2.165 57.7 2.48 ;
      RECT 57.51 2.165 57.7 2.45 ;
      RECT 57.47 2.165 57.73 2.425 ;
      RECT 57.38 3.635 57.46 3.895 ;
      RECT 56.785 2.355 56.79 2.62 ;
      RECT 56.665 2.355 56.79 2.615 ;
      RECT 57.34 3.6 57.38 3.895 ;
      RECT 57.295 3.522 57.34 3.895 ;
      RECT 57.275 3.45 57.295 3.895 ;
      RECT 57.265 3.402 57.275 3.895 ;
      RECT 57.23 3.335 57.265 3.895 ;
      RECT 57.2 3.235 57.23 3.895 ;
      RECT 57.18 3.16 57.2 3.695 ;
      RECT 57.17 3.11 57.18 3.65 ;
      RECT 57.165 3.087 57.17 3.623 ;
      RECT 57.16 3.072 57.165 3.61 ;
      RECT 57.155 3.057 57.16 3.588 ;
      RECT 57.15 3.042 57.155 3.57 ;
      RECT 57.125 2.997 57.15 3.525 ;
      RECT 57.115 2.945 57.125 3.468 ;
      RECT 57.105 2.915 57.115 3.435 ;
      RECT 57.095 2.88 57.105 3.403 ;
      RECT 57.06 2.812 57.095 3.335 ;
      RECT 57.055 2.751 57.06 3.27 ;
      RECT 57.045 2.739 57.055 3.25 ;
      RECT 57.04 2.727 57.045 3.23 ;
      RECT 57.035 2.719 57.04 3.218 ;
      RECT 57.03 2.711 57.035 3.198 ;
      RECT 57.02 2.699 57.03 3.17 ;
      RECT 57.01 2.683 57.02 3.14 ;
      RECT 56.985 2.655 57.01 3.078 ;
      RECT 56.975 2.626 56.985 3.023 ;
      RECT 56.96 2.605 56.975 2.983 ;
      RECT 56.955 2.589 56.96 2.955 ;
      RECT 56.95 2.577 56.955 2.945 ;
      RECT 56.945 2.572 56.95 2.918 ;
      RECT 56.94 2.565 56.945 2.905 ;
      RECT 56.925 2.548 56.94 2.878 ;
      RECT 56.915 2.355 56.925 2.838 ;
      RECT 56.905 2.355 56.915 2.805 ;
      RECT 56.895 2.355 56.905 2.78 ;
      RECT 56.825 2.355 56.895 2.715 ;
      RECT 56.815 2.355 56.825 2.663 ;
      RECT 56.8 2.355 56.815 2.645 ;
      RECT 56.79 2.355 56.8 2.63 ;
      RECT 56.62 3.225 56.88 3.485 ;
      RECT 55.155 3.26 55.16 3.467 ;
      RECT 54.79 3.15 54.865 3.465 ;
      RECT 54.605 3.205 54.76 3.465 ;
      RECT 54.79 3.15 54.895 3.43 ;
      RECT 56.605 3.322 56.62 3.483 ;
      RECT 56.58 3.33 56.605 3.488 ;
      RECT 56.555 3.337 56.58 3.493 ;
      RECT 56.492 3.348 56.555 3.502 ;
      RECT 56.406 3.367 56.492 3.519 ;
      RECT 56.32 3.389 56.406 3.538 ;
      RECT 56.305 3.402 56.32 3.549 ;
      RECT 56.265 3.41 56.305 3.556 ;
      RECT 56.245 3.415 56.265 3.563 ;
      RECT 56.207 3.416 56.245 3.566 ;
      RECT 56.121 3.419 56.207 3.567 ;
      RECT 56.035 3.423 56.121 3.568 ;
      RECT 55.986 3.425 56.035 3.57 ;
      RECT 55.9 3.425 55.986 3.572 ;
      RECT 55.86 3.42 55.9 3.574 ;
      RECT 55.85 3.414 55.86 3.575 ;
      RECT 55.81 3.409 55.85 3.572 ;
      RECT 55.8 3.402 55.81 3.568 ;
      RECT 55.785 3.398 55.8 3.566 ;
      RECT 55.768 3.394 55.785 3.564 ;
      RECT 55.682 3.384 55.768 3.556 ;
      RECT 55.596 3.366 55.682 3.542 ;
      RECT 55.51 3.349 55.596 3.528 ;
      RECT 55.485 3.337 55.51 3.519 ;
      RECT 55.415 3.327 55.485 3.512 ;
      RECT 55.37 3.315 55.415 3.503 ;
      RECT 55.31 3.302 55.37 3.495 ;
      RECT 55.305 3.294 55.31 3.49 ;
      RECT 55.27 3.289 55.305 3.488 ;
      RECT 55.215 3.28 55.27 3.481 ;
      RECT 55.175 3.269 55.215 3.473 ;
      RECT 55.16 3.262 55.175 3.469 ;
      RECT 55.14 3.255 55.155 3.466 ;
      RECT 55.125 3.245 55.14 3.464 ;
      RECT 55.11 3.232 55.125 3.461 ;
      RECT 55.085 3.215 55.11 3.457 ;
      RECT 55.07 3.197 55.085 3.454 ;
      RECT 55.045 3.15 55.07 3.452 ;
      RECT 55.021 3.15 55.045 3.449 ;
      RECT 54.935 3.15 55.021 3.441 ;
      RECT 54.895 3.15 54.935 3.433 ;
      RECT 54.76 3.197 54.79 3.465 ;
      RECT 56.44 2.78 56.7 3.04 ;
      RECT 56.4 2.78 56.7 2.918 ;
      RECT 56.365 2.78 56.7 2.903 ;
      RECT 56.31 2.78 56.7 2.883 ;
      RECT 56.23 2.59 56.51 2.87 ;
      RECT 56.23 2.772 56.58 2.87 ;
      RECT 56.23 2.715 56.565 2.87 ;
      RECT 56.23 2.662 56.515 2.87 ;
      RECT 54.06 2.59 54.255 3.375 ;
      RECT 54.14 1.205 54.255 3.375 ;
      RECT 53.995 3.115 54.055 3.375 ;
      RECT 55.365 2.635 55.625 2.895 ;
      RECT 54.05 2.59 54.255 2.87 ;
      RECT 55.36 2.645 55.625 2.83 ;
      RECT 55.075 2.62 55.085 2.77 ;
      RECT 54.31 1.205 54.39 1.55 ;
      RECT 54.045 1.205 54.255 1.55 ;
      RECT 55.35 2.645 55.36 2.829 ;
      RECT 55.34 2.644 55.35 2.826 ;
      RECT 55.331 2.643 55.34 2.824 ;
      RECT 55.245 2.639 55.331 2.814 ;
      RECT 55.171 2.631 55.245 2.796 ;
      RECT 55.085 2.624 55.171 2.779 ;
      RECT 55.025 2.62 55.075 2.769 ;
      RECT 54.99 2.619 55.025 2.766 ;
      RECT 54.935 2.619 54.99 2.768 ;
      RECT 54.9 2.619 54.935 2.772 ;
      RECT 54.814 2.618 54.9 2.779 ;
      RECT 54.728 2.617 54.814 2.789 ;
      RECT 54.642 2.616 54.728 2.8 ;
      RECT 54.556 2.616 54.642 2.81 ;
      RECT 54.47 2.615 54.556 2.82 ;
      RECT 54.435 2.615 54.47 2.86 ;
      RECT 54.43 2.615 54.435 2.903 ;
      RECT 54.405 2.615 54.43 2.92 ;
      RECT 54.33 2.615 54.405 2.935 ;
      RECT 54.31 2.59 54.33 2.948 ;
      RECT 54.305 1.205 54.31 2.958 ;
      RECT 54.28 1.205 54.305 3 ;
      RECT 54.255 1.205 54.28 3.078 ;
      RECT 54.055 2.997 54.06 3.375 ;
      RECT 53.39 2.949 53.405 3.405 ;
      RECT 53.385 3.021 53.491 3.403 ;
      RECT 53.405 2.115 53.54 3.401 ;
      RECT 53.39 2.965 53.545 3.4 ;
      RECT 53.39 3.015 53.55 3.398 ;
      RECT 53.375 3.08 53.55 3.397 ;
      RECT 53.385 3.072 53.555 3.394 ;
      RECT 53.365 3.12 53.555 3.389 ;
      RECT 53.365 3.12 53.57 3.386 ;
      RECT 53.36 3.12 53.57 3.383 ;
      RECT 53.335 3.12 53.595 3.38 ;
      RECT 53.405 2.115 53.565 2.768 ;
      RECT 53.4 2.115 53.565 2.74 ;
      RECT 53.395 2.115 53.565 2.568 ;
      RECT 53.395 2.115 53.585 2.508 ;
      RECT 53.35 2.115 53.61 2.375 ;
      RECT 52.83 2.59 53.11 2.87 ;
      RECT 52.82 2.605 53.11 2.865 ;
      RECT 52.775 2.667 53.11 2.863 ;
      RECT 52.85 2.582 53.015 2.87 ;
      RECT 52.85 2.567 52.971 2.87 ;
      RECT 52.885 2.56 52.971 2.87 ;
      RECT 52.35 3.71 52.63 3.99 ;
      RECT 52.31 3.672 52.605 3.783 ;
      RECT 52.295 3.622 52.585 3.678 ;
      RECT 52.24 3.385 52.5 3.645 ;
      RECT 52.24 3.587 52.58 3.645 ;
      RECT 52.24 3.527 52.575 3.645 ;
      RECT 52.24 3.477 52.555 3.645 ;
      RECT 52.24 3.457 52.55 3.645 ;
      RECT 52.24 3.435 52.545 3.645 ;
      RECT 52.24 3.42 52.515 3.645 ;
      RECT 47.97 6.225 48.29 6.545 ;
      RECT 48 5.695 48.17 6.545 ;
      RECT 48 5.695 48.175 6.045 ;
      RECT 48 5.695 48.975 5.87 ;
      RECT 48.8 1.965 48.975 5.87 ;
      RECT 48.745 1.965 49.095 2.315 ;
      RECT 48.77 6.655 49.095 6.98 ;
      RECT 47.655 6.745 49.095 6.915 ;
      RECT 47.655 2.395 47.815 6.915 ;
      RECT 47.97 2.365 48.29 2.685 ;
      RECT 47.655 2.395 48.29 2.565 ;
      RECT 46.915 5.84 47.265 6.19 ;
      RECT 46.99 2.705 47.165 6.19 ;
      RECT 46.925 2.705 47.275 3.055 ;
      RECT 46.325 1.14 46.7 1.51 ;
      RECT 38.245 0.96 38.62 1.33 ;
      RECT 36.81 0.96 37.185 1.33 ;
      RECT 36.81 1.08 46.63 1.25 ;
      RECT 42.755 4.36 46.61 4.53 ;
      RECT 46.44 3.425 46.61 4.53 ;
      RECT 42.755 3.67 42.925 4.53 ;
      RECT 42.705 3.71 42.985 3.99 ;
      RECT 42.725 3.67 42.985 3.99 ;
      RECT 42.365 3.625 42.47 3.885 ;
      RECT 46.35 3.43 46.7 3.78 ;
      RECT 42.22 2.115 42.31 2.375 ;
      RECT 42.76 3.18 42.765 3.22 ;
      RECT 42.755 3.17 42.76 3.305 ;
      RECT 42.75 3.16 42.755 3.398 ;
      RECT 42.74 3.14 42.75 3.454 ;
      RECT 42.66 3.068 42.74 3.534 ;
      RECT 42.695 3.712 42.705 3.937 ;
      RECT 42.69 3.709 42.695 3.932 ;
      RECT 42.675 3.706 42.69 3.925 ;
      RECT 42.64 3.7 42.675 3.907 ;
      RECT 42.655 3.003 42.66 3.608 ;
      RECT 42.635 2.954 42.655 3.623 ;
      RECT 42.625 3.687 42.64 3.89 ;
      RECT 42.63 2.896 42.635 3.638 ;
      RECT 42.625 2.874 42.63 3.648 ;
      RECT 42.59 2.784 42.625 3.885 ;
      RECT 42.575 2.662 42.59 3.885 ;
      RECT 42.57 2.615 42.575 3.885 ;
      RECT 42.545 2.54 42.57 3.885 ;
      RECT 42.53 2.455 42.545 3.885 ;
      RECT 42.525 2.402 42.53 3.885 ;
      RECT 42.52 2.382 42.525 3.885 ;
      RECT 42.515 2.357 42.52 3.119 ;
      RECT 42.5 3.317 42.52 3.885 ;
      RECT 42.51 2.335 42.515 3.096 ;
      RECT 42.5 2.287 42.51 3.061 ;
      RECT 42.495 2.25 42.5 3.027 ;
      RECT 42.495 3.397 42.5 3.885 ;
      RECT 42.48 2.227 42.495 2.982 ;
      RECT 42.475 3.495 42.495 3.885 ;
      RECT 42.425 2.115 42.48 2.824 ;
      RECT 42.47 3.617 42.475 3.885 ;
      RECT 42.41 2.115 42.425 2.663 ;
      RECT 42.405 2.115 42.41 2.615 ;
      RECT 42.4 2.115 42.405 2.603 ;
      RECT 42.355 2.115 42.4 2.54 ;
      RECT 42.33 2.115 42.355 2.458 ;
      RECT 42.315 2.115 42.33 2.41 ;
      RECT 42.31 2.115 42.315 2.38 ;
      RECT 44.7 2.16 44.96 2.42 ;
      RECT 44.695 2.16 44.96 2.368 ;
      RECT 44.69 2.16 44.96 2.338 ;
      RECT 44.665 2.03 44.945 2.31 ;
      RECT 33.225 6.66 33.575 7.01 ;
      RECT 44.2 6.615 44.55 6.965 ;
      RECT 33.225 6.69 44.55 6.89 ;
      RECT 43.705 3.71 43.985 3.99 ;
      RECT 43.745 3.665 44.01 3.925 ;
      RECT 43.735 3.7 44.01 3.925 ;
      RECT 43.74 3.685 43.985 3.99 ;
      RECT 43.745 3.662 43.955 3.99 ;
      RECT 43.745 3.66 43.94 3.99 ;
      RECT 43.785 3.65 43.94 3.99 ;
      RECT 43.755 3.655 43.94 3.99 ;
      RECT 43.785 3.647 43.885 3.99 ;
      RECT 43.81 3.64 43.885 3.99 ;
      RECT 43.79 3.642 43.885 3.99 ;
      RECT 43.12 3.155 43.38 3.415 ;
      RECT 43.17 3.147 43.36 3.415 ;
      RECT 43.175 3.067 43.36 3.415 ;
      RECT 43.295 2.455 43.36 3.415 ;
      RECT 43.2 2.852 43.36 3.415 ;
      RECT 43.275 2.54 43.36 3.415 ;
      RECT 43.31 2.165 43.446 2.893 ;
      RECT 43.255 2.662 43.446 2.893 ;
      RECT 43.27 2.602 43.36 3.415 ;
      RECT 43.31 2.165 43.47 2.558 ;
      RECT 43.31 2.165 43.48 2.455 ;
      RECT 43.3 2.165 43.56 2.425 ;
      RECT 41.635 3.565 41.68 3.825 ;
      RECT 41.54 2.1 41.685 2.36 ;
      RECT 42.045 2.722 42.055 2.813 ;
      RECT 42.03 2.66 42.045 2.869 ;
      RECT 42.025 2.607 42.03 2.915 ;
      RECT 41.975 2.554 42.025 3.041 ;
      RECT 41.97 2.509 41.975 3.188 ;
      RECT 41.96 2.497 41.97 3.23 ;
      RECT 41.925 2.461 41.96 3.335 ;
      RECT 41.92 2.429 41.925 3.441 ;
      RECT 41.905 2.411 41.92 3.486 ;
      RECT 41.9 2.394 41.905 2.72 ;
      RECT 41.895 2.775 41.905 3.543 ;
      RECT 41.89 2.38 41.9 2.693 ;
      RECT 41.885 2.83 41.895 3.825 ;
      RECT 41.88 2.366 41.89 2.678 ;
      RECT 41.88 2.88 41.885 3.825 ;
      RECT 41.865 2.343 41.88 2.658 ;
      RECT 41.845 3.002 41.88 3.825 ;
      RECT 41.86 2.325 41.865 2.64 ;
      RECT 41.855 2.317 41.86 2.63 ;
      RECT 41.825 2.285 41.855 2.594 ;
      RECT 41.835 3.13 41.845 3.825 ;
      RECT 41.83 3.157 41.835 3.825 ;
      RECT 41.825 3.207 41.83 3.825 ;
      RECT 41.815 2.251 41.825 2.559 ;
      RECT 41.775 3.275 41.825 3.825 ;
      RECT 41.8 2.228 41.815 2.535 ;
      RECT 41.775 2.1 41.8 2.498 ;
      RECT 41.77 2.1 41.775 2.47 ;
      RECT 41.74 3.375 41.775 3.825 ;
      RECT 41.765 2.1 41.77 2.463 ;
      RECT 41.76 2.1 41.765 2.453 ;
      RECT 41.745 2.1 41.76 2.438 ;
      RECT 41.73 2.1 41.745 2.41 ;
      RECT 41.695 3.48 41.74 3.825 ;
      RECT 41.715 2.1 41.73 2.383 ;
      RECT 41.685 2.1 41.715 2.368 ;
      RECT 41.68 3.552 41.695 3.825 ;
      RECT 41.605 2.635 41.645 2.895 ;
      RECT 41.38 2.582 41.385 2.84 ;
      RECT 37.335 2.06 37.595 2.32 ;
      RECT 37.335 2.085 37.61 2.3 ;
      RECT 39.725 1.91 39.73 2.055 ;
      RECT 41.595 2.63 41.605 2.895 ;
      RECT 41.575 2.622 41.595 2.895 ;
      RECT 41.557 2.618 41.575 2.895 ;
      RECT 41.471 2.607 41.557 2.895 ;
      RECT 41.385 2.59 41.471 2.895 ;
      RECT 41.33 2.577 41.38 2.825 ;
      RECT 41.296 2.569 41.33 2.8 ;
      RECT 41.21 2.558 41.296 2.765 ;
      RECT 41.175 2.535 41.21 2.73 ;
      RECT 41.165 2.497 41.175 2.716 ;
      RECT 41.16 2.47 41.165 2.712 ;
      RECT 41.155 2.457 41.16 2.709 ;
      RECT 41.145 2.437 41.155 2.705 ;
      RECT 41.14 2.412 41.145 2.701 ;
      RECT 41.115 2.367 41.14 2.695 ;
      RECT 41.105 2.308 41.115 2.687 ;
      RECT 41.095 2.276 41.105 2.678 ;
      RECT 41.075 2.228 41.095 2.658 ;
      RECT 41.07 2.188 41.075 2.628 ;
      RECT 41.055 2.162 41.07 2.602 ;
      RECT 41.05 2.14 41.055 2.578 ;
      RECT 41.035 2.112 41.05 2.554 ;
      RECT 41.02 2.085 41.035 2.518 ;
      RECT 41.005 2.062 41.02 2.48 ;
      RECT 41 2.052 41.005 2.455 ;
      RECT 40.99 2.045 41 2.438 ;
      RECT 40.975 2.032 40.99 2.408 ;
      RECT 40.97 2.022 40.975 2.383 ;
      RECT 40.965 2.017 40.97 2.37 ;
      RECT 40.955 2.01 40.965 2.35 ;
      RECT 40.95 2.003 40.955 2.335 ;
      RECT 40.925 1.996 40.95 2.293 ;
      RECT 40.91 1.986 40.925 2.243 ;
      RECT 40.9 1.981 40.91 2.213 ;
      RECT 40.89 1.977 40.9 2.188 ;
      RECT 40.875 1.974 40.89 2.178 ;
      RECT 40.825 1.971 40.875 2.163 ;
      RECT 40.805 1.969 40.825 2.148 ;
      RECT 40.756 1.967 40.805 2.143 ;
      RECT 40.67 1.963 40.756 2.138 ;
      RECT 40.631 1.96 40.67 2.134 ;
      RECT 40.545 1.956 40.631 2.129 ;
      RECT 40.495 1.953 40.545 2.123 ;
      RECT 40.446 1.95 40.495 2.118 ;
      RECT 40.36 1.947 40.446 2.113 ;
      RECT 40.356 1.945 40.36 2.11 ;
      RECT 40.27 1.942 40.356 2.105 ;
      RECT 40.221 1.938 40.27 2.098 ;
      RECT 40.135 1.935 40.221 2.093 ;
      RECT 40.111 1.932 40.135 2.089 ;
      RECT 40.025 1.93 40.111 2.084 ;
      RECT 39.96 1.926 40.025 2.077 ;
      RECT 39.957 1.925 39.96 2.074 ;
      RECT 39.871 1.922 39.957 2.071 ;
      RECT 39.785 1.916 39.871 2.064 ;
      RECT 39.755 1.912 39.785 2.06 ;
      RECT 39.73 1.91 39.755 2.058 ;
      RECT 39.675 1.907 39.725 2.055 ;
      RECT 39.595 1.906 39.675 2.055 ;
      RECT 39.54 1.908 39.595 2.058 ;
      RECT 39.525 1.909 39.54 2.062 ;
      RECT 39.47 1.917 39.525 2.072 ;
      RECT 39.44 1.925 39.47 2.085 ;
      RECT 39.421 1.926 39.44 2.091 ;
      RECT 39.335 1.929 39.421 2.096 ;
      RECT 39.265 1.934 39.335 2.105 ;
      RECT 39.246 1.937 39.265 2.111 ;
      RECT 39.16 1.941 39.246 2.116 ;
      RECT 39.12 1.945 39.16 2.123 ;
      RECT 39.111 1.947 39.12 2.126 ;
      RECT 39.025 1.951 39.111 2.131 ;
      RECT 39.022 1.954 39.025 2.135 ;
      RECT 38.936 1.957 39.022 2.139 ;
      RECT 38.85 1.963 38.936 2.147 ;
      RECT 38.826 1.967 38.85 2.151 ;
      RECT 38.74 1.971 38.826 2.156 ;
      RECT 38.695 1.976 38.74 2.163 ;
      RECT 38.615 1.981 38.695 2.17 ;
      RECT 38.535 1.987 38.615 2.185 ;
      RECT 38.51 1.991 38.535 2.198 ;
      RECT 38.445 1.994 38.51 2.21 ;
      RECT 38.39 1.999 38.445 2.225 ;
      RECT 38.36 2.002 38.39 2.243 ;
      RECT 38.35 2.004 38.36 2.256 ;
      RECT 38.29 2.019 38.35 2.266 ;
      RECT 38.275 2.036 38.29 2.275 ;
      RECT 38.27 2.045 38.275 2.275 ;
      RECT 38.26 2.055 38.27 2.275 ;
      RECT 38.25 2.072 38.26 2.275 ;
      RECT 38.23 2.082 38.25 2.276 ;
      RECT 38.185 2.092 38.23 2.277 ;
      RECT 38.15 2.101 38.185 2.279 ;
      RECT 38.085 2.106 38.15 2.281 ;
      RECT 38.005 2.107 38.085 2.284 ;
      RECT 38.001 2.105 38.005 2.285 ;
      RECT 37.915 2.102 38.001 2.287 ;
      RECT 37.868 2.099 37.915 2.289 ;
      RECT 37.782 2.095 37.868 2.292 ;
      RECT 37.696 2.091 37.782 2.295 ;
      RECT 37.61 2.087 37.696 2.299 ;
      RECT 40.995 3.71 41.025 3.99 ;
      RECT 40.745 3.6 40.765 3.99 ;
      RECT 40.7 3.6 40.765 3.86 ;
      RECT 40.53 2.225 40.565 2.485 ;
      RECT 40.305 2.225 40.365 2.485 ;
      RECT 40.985 3.69 40.995 3.99 ;
      RECT 40.98 3.65 40.985 3.99 ;
      RECT 40.965 3.605 40.98 3.99 ;
      RECT 40.96 3.57 40.965 3.99 ;
      RECT 40.955 3.55 40.96 3.99 ;
      RECT 40.925 3.477 40.955 3.99 ;
      RECT 40.905 3.375 40.925 3.99 ;
      RECT 40.895 3.305 40.905 3.99 ;
      RECT 40.85 3.245 40.895 3.99 ;
      RECT 40.765 3.206 40.85 3.99 ;
      RECT 40.76 3.197 40.765 3.57 ;
      RECT 40.75 3.196 40.76 3.553 ;
      RECT 40.725 3.177 40.75 3.523 ;
      RECT 40.72 3.152 40.725 3.502 ;
      RECT 40.71 3.13 40.72 3.493 ;
      RECT 40.705 3.101 40.71 3.483 ;
      RECT 40.665 3.027 40.705 3.455 ;
      RECT 40.645 2.928 40.665 3.42 ;
      RECT 40.63 2.864 40.645 3.403 ;
      RECT 40.6 2.788 40.63 3.375 ;
      RECT 40.58 2.703 40.6 3.348 ;
      RECT 40.54 2.599 40.58 3.255 ;
      RECT 40.535 2.52 40.54 3.163 ;
      RECT 40.53 2.503 40.535 3.14 ;
      RECT 40.525 2.225 40.53 3.12 ;
      RECT 40.495 2.225 40.525 3.058 ;
      RECT 40.49 2.225 40.495 2.99 ;
      RECT 40.48 2.225 40.49 2.955 ;
      RECT 40.47 2.225 40.48 2.92 ;
      RECT 40.405 2.225 40.47 2.775 ;
      RECT 40.4 2.225 40.405 2.645 ;
      RECT 40.37 2.225 40.4 2.578 ;
      RECT 40.365 2.225 40.37 2.503 ;
      RECT 39.545 3.15 39.825 3.43 ;
      RECT 39.585 3.13 39.845 3.39 ;
      RECT 39.575 3.14 39.845 3.39 ;
      RECT 39.585 3.067 39.8 3.43 ;
      RECT 39.64 2.99 39.795 3.43 ;
      RECT 39.645 2.775 39.795 3.43 ;
      RECT 39.635 2.577 39.785 2.828 ;
      RECT 39.625 2.577 39.785 2.695 ;
      RECT 39.62 2.455 39.78 2.598 ;
      RECT 39.605 2.455 39.78 2.503 ;
      RECT 39.6 2.165 39.775 2.48 ;
      RECT 39.585 2.165 39.775 2.45 ;
      RECT 39.545 2.165 39.805 2.425 ;
      RECT 39.455 3.635 39.535 3.895 ;
      RECT 38.86 2.355 38.865 2.62 ;
      RECT 38.74 2.355 38.865 2.615 ;
      RECT 39.415 3.6 39.455 3.895 ;
      RECT 39.37 3.522 39.415 3.895 ;
      RECT 39.35 3.45 39.37 3.895 ;
      RECT 39.34 3.402 39.35 3.895 ;
      RECT 39.305 3.335 39.34 3.895 ;
      RECT 39.275 3.235 39.305 3.895 ;
      RECT 39.255 3.16 39.275 3.695 ;
      RECT 39.245 3.11 39.255 3.65 ;
      RECT 39.24 3.087 39.245 3.623 ;
      RECT 39.235 3.072 39.24 3.61 ;
      RECT 39.23 3.057 39.235 3.588 ;
      RECT 39.225 3.042 39.23 3.57 ;
      RECT 39.2 2.997 39.225 3.525 ;
      RECT 39.19 2.945 39.2 3.468 ;
      RECT 39.18 2.915 39.19 3.435 ;
      RECT 39.17 2.88 39.18 3.403 ;
      RECT 39.135 2.812 39.17 3.335 ;
      RECT 39.13 2.751 39.135 3.27 ;
      RECT 39.12 2.739 39.13 3.25 ;
      RECT 39.115 2.727 39.12 3.23 ;
      RECT 39.11 2.719 39.115 3.218 ;
      RECT 39.105 2.711 39.11 3.198 ;
      RECT 39.095 2.699 39.105 3.17 ;
      RECT 39.085 2.683 39.095 3.14 ;
      RECT 39.06 2.655 39.085 3.078 ;
      RECT 39.05 2.626 39.06 3.023 ;
      RECT 39.035 2.605 39.05 2.983 ;
      RECT 39.03 2.589 39.035 2.955 ;
      RECT 39.025 2.577 39.03 2.945 ;
      RECT 39.02 2.572 39.025 2.918 ;
      RECT 39.015 2.565 39.02 2.905 ;
      RECT 39 2.548 39.015 2.878 ;
      RECT 38.99 2.355 39 2.838 ;
      RECT 38.98 2.355 38.99 2.805 ;
      RECT 38.97 2.355 38.98 2.78 ;
      RECT 38.9 2.355 38.97 2.715 ;
      RECT 38.89 2.355 38.9 2.663 ;
      RECT 38.875 2.355 38.89 2.645 ;
      RECT 38.865 2.355 38.875 2.63 ;
      RECT 38.695 3.225 38.955 3.485 ;
      RECT 37.23 3.26 37.235 3.467 ;
      RECT 36.865 3.15 36.94 3.465 ;
      RECT 36.68 3.205 36.835 3.465 ;
      RECT 36.865 3.15 36.97 3.43 ;
      RECT 38.68 3.322 38.695 3.483 ;
      RECT 38.655 3.33 38.68 3.488 ;
      RECT 38.63 3.337 38.655 3.493 ;
      RECT 38.567 3.348 38.63 3.502 ;
      RECT 38.481 3.367 38.567 3.519 ;
      RECT 38.395 3.389 38.481 3.538 ;
      RECT 38.38 3.402 38.395 3.549 ;
      RECT 38.34 3.41 38.38 3.556 ;
      RECT 38.32 3.415 38.34 3.563 ;
      RECT 38.282 3.416 38.32 3.566 ;
      RECT 38.196 3.419 38.282 3.567 ;
      RECT 38.11 3.423 38.196 3.568 ;
      RECT 38.061 3.425 38.11 3.57 ;
      RECT 37.975 3.425 38.061 3.572 ;
      RECT 37.935 3.42 37.975 3.574 ;
      RECT 37.925 3.414 37.935 3.575 ;
      RECT 37.885 3.409 37.925 3.572 ;
      RECT 37.875 3.402 37.885 3.568 ;
      RECT 37.86 3.398 37.875 3.566 ;
      RECT 37.843 3.394 37.86 3.564 ;
      RECT 37.757 3.384 37.843 3.556 ;
      RECT 37.671 3.366 37.757 3.542 ;
      RECT 37.585 3.349 37.671 3.528 ;
      RECT 37.56 3.337 37.585 3.519 ;
      RECT 37.49 3.327 37.56 3.512 ;
      RECT 37.445 3.315 37.49 3.503 ;
      RECT 37.385 3.302 37.445 3.495 ;
      RECT 37.38 3.294 37.385 3.49 ;
      RECT 37.345 3.289 37.38 3.488 ;
      RECT 37.29 3.28 37.345 3.481 ;
      RECT 37.25 3.269 37.29 3.473 ;
      RECT 37.235 3.262 37.25 3.469 ;
      RECT 37.215 3.255 37.23 3.466 ;
      RECT 37.2 3.245 37.215 3.464 ;
      RECT 37.185 3.232 37.2 3.461 ;
      RECT 37.16 3.215 37.185 3.457 ;
      RECT 37.145 3.197 37.16 3.454 ;
      RECT 37.12 3.15 37.145 3.452 ;
      RECT 37.096 3.15 37.12 3.449 ;
      RECT 37.01 3.15 37.096 3.441 ;
      RECT 36.97 3.15 37.01 3.433 ;
      RECT 36.835 3.197 36.865 3.465 ;
      RECT 38.515 2.78 38.775 3.04 ;
      RECT 38.475 2.78 38.775 2.918 ;
      RECT 38.44 2.78 38.775 2.903 ;
      RECT 38.385 2.78 38.775 2.883 ;
      RECT 38.305 2.59 38.585 2.87 ;
      RECT 38.305 2.772 38.655 2.87 ;
      RECT 38.305 2.715 38.64 2.87 ;
      RECT 38.305 2.662 38.59 2.87 ;
      RECT 36.135 2.59 36.33 3.375 ;
      RECT 36.215 1.205 36.33 3.375 ;
      RECT 36.07 3.115 36.13 3.375 ;
      RECT 37.44 2.635 37.7 2.895 ;
      RECT 36.125 2.59 36.33 2.87 ;
      RECT 37.435 2.645 37.7 2.83 ;
      RECT 37.15 2.62 37.16 2.77 ;
      RECT 36.385 1.205 36.465 1.55 ;
      RECT 36.12 1.205 36.33 1.55 ;
      RECT 37.425 2.645 37.435 2.829 ;
      RECT 37.415 2.644 37.425 2.826 ;
      RECT 37.406 2.643 37.415 2.824 ;
      RECT 37.32 2.639 37.406 2.814 ;
      RECT 37.246 2.631 37.32 2.796 ;
      RECT 37.16 2.624 37.246 2.779 ;
      RECT 37.1 2.62 37.15 2.769 ;
      RECT 37.065 2.619 37.1 2.766 ;
      RECT 37.01 2.619 37.065 2.768 ;
      RECT 36.975 2.619 37.01 2.772 ;
      RECT 36.889 2.618 36.975 2.779 ;
      RECT 36.803 2.617 36.889 2.789 ;
      RECT 36.717 2.616 36.803 2.8 ;
      RECT 36.631 2.616 36.717 2.81 ;
      RECT 36.545 2.615 36.631 2.82 ;
      RECT 36.51 2.615 36.545 2.86 ;
      RECT 36.505 2.615 36.51 2.903 ;
      RECT 36.48 2.615 36.505 2.92 ;
      RECT 36.405 2.615 36.48 2.935 ;
      RECT 36.385 2.59 36.405 2.948 ;
      RECT 36.38 1.205 36.385 2.958 ;
      RECT 36.355 1.205 36.38 3 ;
      RECT 36.33 1.205 36.355 3.078 ;
      RECT 36.13 2.997 36.135 3.375 ;
      RECT 35.465 2.949 35.48 3.405 ;
      RECT 35.46 3.021 35.566 3.403 ;
      RECT 35.48 2.115 35.615 3.401 ;
      RECT 35.465 2.965 35.62 3.4 ;
      RECT 35.465 3.015 35.625 3.398 ;
      RECT 35.45 3.08 35.625 3.397 ;
      RECT 35.46 3.072 35.63 3.394 ;
      RECT 35.44 3.12 35.63 3.389 ;
      RECT 35.44 3.12 35.645 3.386 ;
      RECT 35.435 3.12 35.645 3.383 ;
      RECT 35.41 3.12 35.67 3.38 ;
      RECT 35.48 2.115 35.64 2.768 ;
      RECT 35.475 2.115 35.64 2.74 ;
      RECT 35.47 2.115 35.64 2.568 ;
      RECT 35.47 2.115 35.66 2.508 ;
      RECT 35.425 2.115 35.685 2.375 ;
      RECT 34.905 2.59 35.185 2.87 ;
      RECT 34.895 2.605 35.185 2.865 ;
      RECT 34.85 2.667 35.185 2.863 ;
      RECT 34.925 2.582 35.09 2.87 ;
      RECT 34.925 2.567 35.046 2.87 ;
      RECT 34.96 2.56 35.046 2.87 ;
      RECT 34.425 3.71 34.705 3.99 ;
      RECT 34.385 3.672 34.68 3.783 ;
      RECT 34.37 3.622 34.66 3.678 ;
      RECT 34.315 3.385 34.575 3.645 ;
      RECT 34.315 3.587 34.655 3.645 ;
      RECT 34.315 3.527 34.65 3.645 ;
      RECT 34.315 3.477 34.63 3.645 ;
      RECT 34.315 3.457 34.625 3.645 ;
      RECT 34.315 3.435 34.62 3.645 ;
      RECT 34.315 3.42 34.59 3.645 ;
      RECT 30.045 6.225 30.365 6.545 ;
      RECT 30.075 5.695 30.245 6.545 ;
      RECT 30.075 5.695 30.25 6.045 ;
      RECT 30.075 5.695 31.05 5.87 ;
      RECT 30.875 1.965 31.05 5.87 ;
      RECT 30.82 1.965 31.17 2.315 ;
      RECT 30.845 6.655 31.17 6.98 ;
      RECT 29.73 6.745 31.17 6.915 ;
      RECT 29.73 2.395 29.89 6.915 ;
      RECT 30.045 2.365 30.365 2.685 ;
      RECT 29.73 2.395 30.365 2.565 ;
      RECT 28.99 5.84 29.34 6.19 ;
      RECT 29.065 2.705 29.24 6.19 ;
      RECT 29 2.705 29.35 3.055 ;
      RECT 28.4 1.14 28.775 1.51 ;
      RECT 20.32 0.96 20.695 1.33 ;
      RECT 18.885 0.96 19.26 1.33 ;
      RECT 18.885 1.08 28.705 1.25 ;
      RECT 24.83 4.36 28.685 4.53 ;
      RECT 28.515 3.425 28.685 4.53 ;
      RECT 24.83 3.67 25 4.53 ;
      RECT 24.78 3.71 25.06 3.99 ;
      RECT 24.8 3.67 25.06 3.99 ;
      RECT 24.44 3.625 24.545 3.885 ;
      RECT 28.425 3.43 28.775 3.78 ;
      RECT 24.295 2.115 24.385 2.375 ;
      RECT 24.835 3.18 24.84 3.22 ;
      RECT 24.83 3.17 24.835 3.305 ;
      RECT 24.825 3.16 24.83 3.398 ;
      RECT 24.815 3.14 24.825 3.454 ;
      RECT 24.735 3.068 24.815 3.534 ;
      RECT 24.77 3.712 24.78 3.937 ;
      RECT 24.765 3.709 24.77 3.932 ;
      RECT 24.75 3.706 24.765 3.925 ;
      RECT 24.715 3.7 24.75 3.907 ;
      RECT 24.73 3.003 24.735 3.608 ;
      RECT 24.71 2.954 24.73 3.623 ;
      RECT 24.7 3.687 24.715 3.89 ;
      RECT 24.705 2.896 24.71 3.638 ;
      RECT 24.7 2.874 24.705 3.648 ;
      RECT 24.665 2.784 24.7 3.885 ;
      RECT 24.65 2.662 24.665 3.885 ;
      RECT 24.645 2.615 24.65 3.885 ;
      RECT 24.62 2.54 24.645 3.885 ;
      RECT 24.605 2.455 24.62 3.885 ;
      RECT 24.6 2.402 24.605 3.885 ;
      RECT 24.595 2.382 24.6 3.885 ;
      RECT 24.59 2.357 24.595 3.119 ;
      RECT 24.575 3.317 24.595 3.885 ;
      RECT 24.585 2.335 24.59 3.096 ;
      RECT 24.575 2.287 24.585 3.061 ;
      RECT 24.57 2.25 24.575 3.027 ;
      RECT 24.57 3.397 24.575 3.885 ;
      RECT 24.555 2.227 24.57 2.982 ;
      RECT 24.55 3.495 24.57 3.885 ;
      RECT 24.5 2.115 24.555 2.824 ;
      RECT 24.545 3.617 24.55 3.885 ;
      RECT 24.485 2.115 24.5 2.663 ;
      RECT 24.48 2.115 24.485 2.615 ;
      RECT 24.475 2.115 24.48 2.603 ;
      RECT 24.43 2.115 24.475 2.54 ;
      RECT 24.405 2.115 24.43 2.458 ;
      RECT 24.39 2.115 24.405 2.41 ;
      RECT 24.385 2.115 24.39 2.38 ;
      RECT 26.775 2.16 27.035 2.42 ;
      RECT 26.77 2.16 27.035 2.368 ;
      RECT 26.765 2.16 27.035 2.338 ;
      RECT 26.74 2.03 27.02 2.31 ;
      RECT 15.3 6.655 15.65 7.005 ;
      RECT 26.27 6.61 26.62 6.96 ;
      RECT 15.3 6.685 26.62 6.885 ;
      RECT 25.78 3.71 26.06 3.99 ;
      RECT 25.82 3.665 26.085 3.925 ;
      RECT 25.81 3.7 26.085 3.925 ;
      RECT 25.815 3.685 26.06 3.99 ;
      RECT 25.82 3.662 26.03 3.99 ;
      RECT 25.82 3.66 26.015 3.99 ;
      RECT 25.86 3.65 26.015 3.99 ;
      RECT 25.83 3.655 26.015 3.99 ;
      RECT 25.86 3.647 25.96 3.99 ;
      RECT 25.885 3.64 25.96 3.99 ;
      RECT 25.865 3.642 25.96 3.99 ;
      RECT 25.195 3.155 25.455 3.415 ;
      RECT 25.245 3.147 25.435 3.415 ;
      RECT 25.25 3.067 25.435 3.415 ;
      RECT 25.37 2.455 25.435 3.415 ;
      RECT 25.275 2.852 25.435 3.415 ;
      RECT 25.35 2.54 25.435 3.415 ;
      RECT 25.385 2.165 25.521 2.893 ;
      RECT 25.33 2.662 25.521 2.893 ;
      RECT 25.345 2.602 25.435 3.415 ;
      RECT 25.385 2.165 25.545 2.558 ;
      RECT 25.385 2.165 25.555 2.455 ;
      RECT 25.375 2.165 25.635 2.425 ;
      RECT 23.71 3.565 23.755 3.825 ;
      RECT 23.615 2.1 23.76 2.36 ;
      RECT 24.12 2.722 24.13 2.813 ;
      RECT 24.105 2.66 24.12 2.869 ;
      RECT 24.1 2.607 24.105 2.915 ;
      RECT 24.05 2.554 24.1 3.041 ;
      RECT 24.045 2.509 24.05 3.188 ;
      RECT 24.035 2.497 24.045 3.23 ;
      RECT 24 2.461 24.035 3.335 ;
      RECT 23.995 2.429 24 3.441 ;
      RECT 23.98 2.411 23.995 3.486 ;
      RECT 23.975 2.394 23.98 2.72 ;
      RECT 23.97 2.775 23.98 3.543 ;
      RECT 23.965 2.38 23.975 2.693 ;
      RECT 23.96 2.83 23.97 3.825 ;
      RECT 23.955 2.366 23.965 2.678 ;
      RECT 23.955 2.88 23.96 3.825 ;
      RECT 23.94 2.343 23.955 2.658 ;
      RECT 23.92 3.002 23.955 3.825 ;
      RECT 23.935 2.325 23.94 2.64 ;
      RECT 23.93 2.317 23.935 2.63 ;
      RECT 23.9 2.285 23.93 2.594 ;
      RECT 23.91 3.13 23.92 3.825 ;
      RECT 23.905 3.157 23.91 3.825 ;
      RECT 23.9 3.207 23.905 3.825 ;
      RECT 23.89 2.251 23.9 2.559 ;
      RECT 23.85 3.275 23.9 3.825 ;
      RECT 23.875 2.228 23.89 2.535 ;
      RECT 23.85 2.1 23.875 2.498 ;
      RECT 23.845 2.1 23.85 2.47 ;
      RECT 23.815 3.375 23.85 3.825 ;
      RECT 23.84 2.1 23.845 2.463 ;
      RECT 23.835 2.1 23.84 2.453 ;
      RECT 23.82 2.1 23.835 2.438 ;
      RECT 23.805 2.1 23.82 2.41 ;
      RECT 23.77 3.48 23.815 3.825 ;
      RECT 23.79 2.1 23.805 2.383 ;
      RECT 23.76 2.1 23.79 2.368 ;
      RECT 23.755 3.552 23.77 3.825 ;
      RECT 23.68 2.635 23.72 2.895 ;
      RECT 23.455 2.582 23.46 2.84 ;
      RECT 19.41 2.06 19.67 2.32 ;
      RECT 19.41 2.085 19.685 2.3 ;
      RECT 21.8 1.91 21.805 2.055 ;
      RECT 23.67 2.63 23.68 2.895 ;
      RECT 23.65 2.622 23.67 2.895 ;
      RECT 23.632 2.618 23.65 2.895 ;
      RECT 23.546 2.607 23.632 2.895 ;
      RECT 23.46 2.59 23.546 2.895 ;
      RECT 23.405 2.577 23.455 2.825 ;
      RECT 23.371 2.569 23.405 2.8 ;
      RECT 23.285 2.558 23.371 2.765 ;
      RECT 23.25 2.535 23.285 2.73 ;
      RECT 23.24 2.497 23.25 2.716 ;
      RECT 23.235 2.47 23.24 2.712 ;
      RECT 23.23 2.457 23.235 2.709 ;
      RECT 23.22 2.437 23.23 2.705 ;
      RECT 23.215 2.412 23.22 2.701 ;
      RECT 23.19 2.367 23.215 2.695 ;
      RECT 23.18 2.308 23.19 2.687 ;
      RECT 23.17 2.276 23.18 2.678 ;
      RECT 23.15 2.228 23.17 2.658 ;
      RECT 23.145 2.188 23.15 2.628 ;
      RECT 23.13 2.162 23.145 2.602 ;
      RECT 23.125 2.14 23.13 2.578 ;
      RECT 23.11 2.112 23.125 2.554 ;
      RECT 23.095 2.085 23.11 2.518 ;
      RECT 23.08 2.062 23.095 2.48 ;
      RECT 23.075 2.052 23.08 2.455 ;
      RECT 23.065 2.045 23.075 2.438 ;
      RECT 23.05 2.032 23.065 2.408 ;
      RECT 23.045 2.022 23.05 2.383 ;
      RECT 23.04 2.017 23.045 2.37 ;
      RECT 23.03 2.01 23.04 2.35 ;
      RECT 23.025 2.003 23.03 2.335 ;
      RECT 23 1.996 23.025 2.293 ;
      RECT 22.985 1.986 23 2.243 ;
      RECT 22.975 1.981 22.985 2.213 ;
      RECT 22.965 1.977 22.975 2.188 ;
      RECT 22.95 1.974 22.965 2.178 ;
      RECT 22.9 1.971 22.95 2.163 ;
      RECT 22.88 1.969 22.9 2.148 ;
      RECT 22.831 1.967 22.88 2.143 ;
      RECT 22.745 1.963 22.831 2.138 ;
      RECT 22.706 1.96 22.745 2.134 ;
      RECT 22.62 1.956 22.706 2.129 ;
      RECT 22.57 1.953 22.62 2.123 ;
      RECT 22.521 1.95 22.57 2.118 ;
      RECT 22.435 1.947 22.521 2.113 ;
      RECT 22.431 1.945 22.435 2.11 ;
      RECT 22.345 1.942 22.431 2.105 ;
      RECT 22.296 1.938 22.345 2.098 ;
      RECT 22.21 1.935 22.296 2.093 ;
      RECT 22.186 1.932 22.21 2.089 ;
      RECT 22.1 1.93 22.186 2.084 ;
      RECT 22.035 1.926 22.1 2.077 ;
      RECT 22.032 1.925 22.035 2.074 ;
      RECT 21.946 1.922 22.032 2.071 ;
      RECT 21.86 1.916 21.946 2.064 ;
      RECT 21.83 1.912 21.86 2.06 ;
      RECT 21.805 1.91 21.83 2.058 ;
      RECT 21.75 1.907 21.8 2.055 ;
      RECT 21.67 1.906 21.75 2.055 ;
      RECT 21.615 1.908 21.67 2.058 ;
      RECT 21.6 1.909 21.615 2.062 ;
      RECT 21.545 1.917 21.6 2.072 ;
      RECT 21.515 1.925 21.545 2.085 ;
      RECT 21.496 1.926 21.515 2.091 ;
      RECT 21.41 1.929 21.496 2.096 ;
      RECT 21.34 1.934 21.41 2.105 ;
      RECT 21.321 1.937 21.34 2.111 ;
      RECT 21.235 1.941 21.321 2.116 ;
      RECT 21.195 1.945 21.235 2.123 ;
      RECT 21.186 1.947 21.195 2.126 ;
      RECT 21.1 1.951 21.186 2.131 ;
      RECT 21.097 1.954 21.1 2.135 ;
      RECT 21.011 1.957 21.097 2.139 ;
      RECT 20.925 1.963 21.011 2.147 ;
      RECT 20.901 1.967 20.925 2.151 ;
      RECT 20.815 1.971 20.901 2.156 ;
      RECT 20.77 1.976 20.815 2.163 ;
      RECT 20.69 1.981 20.77 2.17 ;
      RECT 20.61 1.987 20.69 2.185 ;
      RECT 20.585 1.991 20.61 2.198 ;
      RECT 20.52 1.994 20.585 2.21 ;
      RECT 20.465 1.999 20.52 2.225 ;
      RECT 20.435 2.002 20.465 2.243 ;
      RECT 20.425 2.004 20.435 2.256 ;
      RECT 20.365 2.019 20.425 2.266 ;
      RECT 20.35 2.036 20.365 2.275 ;
      RECT 20.345 2.045 20.35 2.275 ;
      RECT 20.335 2.055 20.345 2.275 ;
      RECT 20.325 2.072 20.335 2.275 ;
      RECT 20.305 2.082 20.325 2.276 ;
      RECT 20.26 2.092 20.305 2.277 ;
      RECT 20.225 2.101 20.26 2.279 ;
      RECT 20.16 2.106 20.225 2.281 ;
      RECT 20.08 2.107 20.16 2.284 ;
      RECT 20.076 2.105 20.08 2.285 ;
      RECT 19.99 2.102 20.076 2.287 ;
      RECT 19.943 2.099 19.99 2.289 ;
      RECT 19.857 2.095 19.943 2.292 ;
      RECT 19.771 2.091 19.857 2.295 ;
      RECT 19.685 2.087 19.771 2.299 ;
      RECT 23.07 3.71 23.1 3.99 ;
      RECT 22.82 3.6 22.84 3.99 ;
      RECT 22.775 3.6 22.84 3.86 ;
      RECT 22.605 2.225 22.64 2.485 ;
      RECT 22.38 2.225 22.44 2.485 ;
      RECT 23.06 3.69 23.07 3.99 ;
      RECT 23.055 3.65 23.06 3.99 ;
      RECT 23.04 3.605 23.055 3.99 ;
      RECT 23.035 3.57 23.04 3.99 ;
      RECT 23.03 3.55 23.035 3.99 ;
      RECT 23 3.477 23.03 3.99 ;
      RECT 22.98 3.375 23 3.99 ;
      RECT 22.97 3.305 22.98 3.99 ;
      RECT 22.925 3.245 22.97 3.99 ;
      RECT 22.84 3.206 22.925 3.99 ;
      RECT 22.835 3.197 22.84 3.57 ;
      RECT 22.825 3.196 22.835 3.553 ;
      RECT 22.8 3.177 22.825 3.523 ;
      RECT 22.795 3.152 22.8 3.502 ;
      RECT 22.785 3.13 22.795 3.493 ;
      RECT 22.78 3.101 22.785 3.483 ;
      RECT 22.74 3.027 22.78 3.455 ;
      RECT 22.72 2.928 22.74 3.42 ;
      RECT 22.705 2.864 22.72 3.403 ;
      RECT 22.675 2.788 22.705 3.375 ;
      RECT 22.655 2.703 22.675 3.348 ;
      RECT 22.615 2.599 22.655 3.255 ;
      RECT 22.61 2.52 22.615 3.163 ;
      RECT 22.605 2.503 22.61 3.14 ;
      RECT 22.6 2.225 22.605 3.12 ;
      RECT 22.57 2.225 22.6 3.058 ;
      RECT 22.565 2.225 22.57 2.99 ;
      RECT 22.555 2.225 22.565 2.955 ;
      RECT 22.545 2.225 22.555 2.92 ;
      RECT 22.48 2.225 22.545 2.775 ;
      RECT 22.475 2.225 22.48 2.645 ;
      RECT 22.445 2.225 22.475 2.578 ;
      RECT 22.44 2.225 22.445 2.503 ;
      RECT 21.62 3.15 21.9 3.43 ;
      RECT 21.66 3.13 21.92 3.39 ;
      RECT 21.65 3.14 21.92 3.39 ;
      RECT 21.66 3.067 21.875 3.43 ;
      RECT 21.715 2.99 21.87 3.43 ;
      RECT 21.72 2.775 21.87 3.43 ;
      RECT 21.71 2.577 21.86 2.828 ;
      RECT 21.7 2.577 21.86 2.695 ;
      RECT 21.695 2.455 21.855 2.598 ;
      RECT 21.68 2.455 21.855 2.503 ;
      RECT 21.675 2.165 21.85 2.48 ;
      RECT 21.66 2.165 21.85 2.45 ;
      RECT 21.62 2.165 21.88 2.425 ;
      RECT 21.53 3.635 21.61 3.895 ;
      RECT 20.935 2.355 20.94 2.62 ;
      RECT 20.815 2.355 20.94 2.615 ;
      RECT 21.49 3.6 21.53 3.895 ;
      RECT 21.445 3.522 21.49 3.895 ;
      RECT 21.425 3.45 21.445 3.895 ;
      RECT 21.415 3.402 21.425 3.895 ;
      RECT 21.38 3.335 21.415 3.895 ;
      RECT 21.35 3.235 21.38 3.895 ;
      RECT 21.33 3.16 21.35 3.695 ;
      RECT 21.32 3.11 21.33 3.65 ;
      RECT 21.315 3.087 21.32 3.623 ;
      RECT 21.31 3.072 21.315 3.61 ;
      RECT 21.305 3.057 21.31 3.588 ;
      RECT 21.3 3.042 21.305 3.57 ;
      RECT 21.275 2.997 21.3 3.525 ;
      RECT 21.265 2.945 21.275 3.468 ;
      RECT 21.255 2.915 21.265 3.435 ;
      RECT 21.245 2.88 21.255 3.403 ;
      RECT 21.21 2.812 21.245 3.335 ;
      RECT 21.205 2.751 21.21 3.27 ;
      RECT 21.195 2.739 21.205 3.25 ;
      RECT 21.19 2.727 21.195 3.23 ;
      RECT 21.185 2.719 21.19 3.218 ;
      RECT 21.18 2.711 21.185 3.198 ;
      RECT 21.17 2.699 21.18 3.17 ;
      RECT 21.16 2.683 21.17 3.14 ;
      RECT 21.135 2.655 21.16 3.078 ;
      RECT 21.125 2.626 21.135 3.023 ;
      RECT 21.11 2.605 21.125 2.983 ;
      RECT 21.105 2.589 21.11 2.955 ;
      RECT 21.1 2.577 21.105 2.945 ;
      RECT 21.095 2.572 21.1 2.918 ;
      RECT 21.09 2.565 21.095 2.905 ;
      RECT 21.075 2.548 21.09 2.878 ;
      RECT 21.065 2.355 21.075 2.838 ;
      RECT 21.055 2.355 21.065 2.805 ;
      RECT 21.045 2.355 21.055 2.78 ;
      RECT 20.975 2.355 21.045 2.715 ;
      RECT 20.965 2.355 20.975 2.663 ;
      RECT 20.95 2.355 20.965 2.645 ;
      RECT 20.94 2.355 20.95 2.63 ;
      RECT 20.77 3.225 21.03 3.485 ;
      RECT 19.305 3.26 19.31 3.467 ;
      RECT 18.94 3.15 19.015 3.465 ;
      RECT 18.755 3.205 18.91 3.465 ;
      RECT 18.94 3.15 19.045 3.43 ;
      RECT 20.755 3.322 20.77 3.483 ;
      RECT 20.73 3.33 20.755 3.488 ;
      RECT 20.705 3.337 20.73 3.493 ;
      RECT 20.642 3.348 20.705 3.502 ;
      RECT 20.556 3.367 20.642 3.519 ;
      RECT 20.47 3.389 20.556 3.538 ;
      RECT 20.455 3.402 20.47 3.549 ;
      RECT 20.415 3.41 20.455 3.556 ;
      RECT 20.395 3.415 20.415 3.563 ;
      RECT 20.357 3.416 20.395 3.566 ;
      RECT 20.271 3.419 20.357 3.567 ;
      RECT 20.185 3.423 20.271 3.568 ;
      RECT 20.136 3.425 20.185 3.57 ;
      RECT 20.05 3.425 20.136 3.572 ;
      RECT 20.01 3.42 20.05 3.574 ;
      RECT 20 3.414 20.01 3.575 ;
      RECT 19.96 3.409 20 3.572 ;
      RECT 19.95 3.402 19.96 3.568 ;
      RECT 19.935 3.398 19.95 3.566 ;
      RECT 19.918 3.394 19.935 3.564 ;
      RECT 19.832 3.384 19.918 3.556 ;
      RECT 19.746 3.366 19.832 3.542 ;
      RECT 19.66 3.349 19.746 3.528 ;
      RECT 19.635 3.337 19.66 3.519 ;
      RECT 19.565 3.327 19.635 3.512 ;
      RECT 19.52 3.315 19.565 3.503 ;
      RECT 19.46 3.302 19.52 3.495 ;
      RECT 19.455 3.294 19.46 3.49 ;
      RECT 19.42 3.289 19.455 3.488 ;
      RECT 19.365 3.28 19.42 3.481 ;
      RECT 19.325 3.269 19.365 3.473 ;
      RECT 19.31 3.262 19.325 3.469 ;
      RECT 19.29 3.255 19.305 3.466 ;
      RECT 19.275 3.245 19.29 3.464 ;
      RECT 19.26 3.232 19.275 3.461 ;
      RECT 19.235 3.215 19.26 3.457 ;
      RECT 19.22 3.197 19.235 3.454 ;
      RECT 19.195 3.15 19.22 3.452 ;
      RECT 19.171 3.15 19.195 3.449 ;
      RECT 19.085 3.15 19.171 3.441 ;
      RECT 19.045 3.15 19.085 3.433 ;
      RECT 18.91 3.197 18.94 3.465 ;
      RECT 20.59 2.78 20.85 3.04 ;
      RECT 20.55 2.78 20.85 2.918 ;
      RECT 20.515 2.78 20.85 2.903 ;
      RECT 20.46 2.78 20.85 2.883 ;
      RECT 20.38 2.59 20.66 2.87 ;
      RECT 20.38 2.772 20.73 2.87 ;
      RECT 20.38 2.715 20.715 2.87 ;
      RECT 20.38 2.662 20.665 2.87 ;
      RECT 18.21 2.59 18.405 3.375 ;
      RECT 18.29 1.205 18.405 3.375 ;
      RECT 18.145 3.115 18.205 3.375 ;
      RECT 19.515 2.635 19.775 2.895 ;
      RECT 18.2 2.59 18.405 2.87 ;
      RECT 19.51 2.645 19.775 2.83 ;
      RECT 19.225 2.62 19.235 2.77 ;
      RECT 18.46 1.205 18.54 1.55 ;
      RECT 18.195 1.205 18.405 1.55 ;
      RECT 19.5 2.645 19.51 2.829 ;
      RECT 19.49 2.644 19.5 2.826 ;
      RECT 19.481 2.643 19.49 2.824 ;
      RECT 19.395 2.639 19.481 2.814 ;
      RECT 19.321 2.631 19.395 2.796 ;
      RECT 19.235 2.624 19.321 2.779 ;
      RECT 19.175 2.62 19.225 2.769 ;
      RECT 19.14 2.619 19.175 2.766 ;
      RECT 19.085 2.619 19.14 2.768 ;
      RECT 19.05 2.619 19.085 2.772 ;
      RECT 18.964 2.618 19.05 2.779 ;
      RECT 18.878 2.617 18.964 2.789 ;
      RECT 18.792 2.616 18.878 2.8 ;
      RECT 18.706 2.616 18.792 2.81 ;
      RECT 18.62 2.615 18.706 2.82 ;
      RECT 18.585 2.615 18.62 2.86 ;
      RECT 18.58 2.615 18.585 2.903 ;
      RECT 18.555 2.615 18.58 2.92 ;
      RECT 18.48 2.615 18.555 2.935 ;
      RECT 18.46 2.59 18.48 2.948 ;
      RECT 18.455 1.205 18.46 2.958 ;
      RECT 18.43 1.205 18.455 3 ;
      RECT 18.405 1.205 18.43 3.078 ;
      RECT 18.205 2.997 18.21 3.375 ;
      RECT 17.54 2.949 17.555 3.405 ;
      RECT 17.535 3.021 17.641 3.403 ;
      RECT 17.555 2.115 17.69 3.401 ;
      RECT 17.54 2.965 17.695 3.4 ;
      RECT 17.54 3.015 17.7 3.398 ;
      RECT 17.525 3.08 17.7 3.397 ;
      RECT 17.535 3.072 17.705 3.394 ;
      RECT 17.515 3.12 17.705 3.389 ;
      RECT 17.515 3.12 17.72 3.386 ;
      RECT 17.51 3.12 17.72 3.383 ;
      RECT 17.485 3.12 17.745 3.38 ;
      RECT 17.555 2.115 17.715 2.768 ;
      RECT 17.55 2.115 17.715 2.74 ;
      RECT 17.545 2.115 17.715 2.568 ;
      RECT 17.545 2.115 17.735 2.508 ;
      RECT 17.5 2.115 17.76 2.375 ;
      RECT 16.98 2.59 17.26 2.87 ;
      RECT 16.97 2.605 17.26 2.865 ;
      RECT 16.925 2.667 17.26 2.863 ;
      RECT 17 2.582 17.165 2.87 ;
      RECT 17 2.567 17.121 2.87 ;
      RECT 17.035 2.56 17.121 2.87 ;
      RECT 16.5 3.71 16.78 3.99 ;
      RECT 16.46 3.672 16.755 3.783 ;
      RECT 16.445 3.622 16.735 3.678 ;
      RECT 16.39 3.385 16.65 3.645 ;
      RECT 16.39 3.587 16.73 3.645 ;
      RECT 16.39 3.527 16.725 3.645 ;
      RECT 16.39 3.477 16.705 3.645 ;
      RECT 16.39 3.457 16.7 3.645 ;
      RECT 16.39 3.435 16.695 3.645 ;
      RECT 16.39 3.42 16.665 3.645 ;
      RECT 12.12 6.225 12.44 6.545 ;
      RECT 12.15 5.695 12.32 6.545 ;
      RECT 12.15 5.695 12.325 6.045 ;
      RECT 12.15 5.695 13.125 5.87 ;
      RECT 12.95 1.965 13.125 5.87 ;
      RECT 12.895 1.965 13.245 2.315 ;
      RECT 12.92 6.655 13.245 6.98 ;
      RECT 11.805 6.745 13.245 6.915 ;
      RECT 11.805 2.395 11.965 6.915 ;
      RECT 12.12 2.365 12.44 2.685 ;
      RECT 11.805 2.395 12.44 2.565 ;
      RECT 11.065 5.84 11.415 6.19 ;
      RECT 11.14 2.705 11.315 6.19 ;
      RECT 11.075 2.705 11.425 3.055 ;
      RECT 10.475 1.14 10.85 1.51 ;
      RECT 2.395 0.96 2.77 1.33 ;
      RECT 0.96 0.96 1.335 1.33 ;
      RECT 0.96 1.08 10.78 1.25 ;
      RECT 6.905 4.36 10.76 4.53 ;
      RECT 10.59 3.425 10.76 4.53 ;
      RECT 6.905 3.67 7.075 4.53 ;
      RECT 6.855 3.71 7.135 3.99 ;
      RECT 6.875 3.67 7.135 3.99 ;
      RECT 6.515 3.625 6.62 3.885 ;
      RECT 10.5 3.43 10.85 3.78 ;
      RECT 6.37 2.115 6.46 2.375 ;
      RECT 6.91 3.18 6.915 3.22 ;
      RECT 6.905 3.17 6.91 3.305 ;
      RECT 6.9 3.16 6.905 3.398 ;
      RECT 6.89 3.14 6.9 3.454 ;
      RECT 6.81 3.068 6.89 3.534 ;
      RECT 6.845 3.712 6.855 3.937 ;
      RECT 6.84 3.709 6.845 3.932 ;
      RECT 6.825 3.706 6.84 3.925 ;
      RECT 6.79 3.7 6.825 3.907 ;
      RECT 6.805 3.003 6.81 3.608 ;
      RECT 6.785 2.954 6.805 3.623 ;
      RECT 6.775 3.687 6.79 3.89 ;
      RECT 6.78 2.896 6.785 3.638 ;
      RECT 6.775 2.874 6.78 3.648 ;
      RECT 6.74 2.784 6.775 3.885 ;
      RECT 6.725 2.662 6.74 3.885 ;
      RECT 6.72 2.615 6.725 3.885 ;
      RECT 6.695 2.54 6.72 3.885 ;
      RECT 6.68 2.455 6.695 3.885 ;
      RECT 6.675 2.402 6.68 3.885 ;
      RECT 6.67 2.382 6.675 3.885 ;
      RECT 6.665 2.357 6.67 3.119 ;
      RECT 6.65 3.317 6.67 3.885 ;
      RECT 6.66 2.335 6.665 3.096 ;
      RECT 6.65 2.287 6.66 3.061 ;
      RECT 6.645 2.25 6.65 3.027 ;
      RECT 6.645 3.397 6.65 3.885 ;
      RECT 6.63 2.227 6.645 2.982 ;
      RECT 6.625 3.495 6.645 3.885 ;
      RECT 6.575 2.115 6.63 2.824 ;
      RECT 6.62 3.617 6.625 3.885 ;
      RECT 6.56 2.115 6.575 2.663 ;
      RECT 6.555 2.115 6.56 2.615 ;
      RECT 6.55 2.115 6.555 2.603 ;
      RECT 6.505 2.115 6.55 2.54 ;
      RECT 6.48 2.115 6.505 2.458 ;
      RECT 6.465 2.115 6.48 2.41 ;
      RECT 6.46 2.115 6.465 2.38 ;
      RECT 8.85 2.16 9.11 2.42 ;
      RECT 8.845 2.16 9.11 2.368 ;
      RECT 8.84 2.16 9.11 2.338 ;
      RECT 8.815 2.03 9.095 2.31 ;
      RECT -3.325 6.995 -3.035 7.345 ;
      RECT -3.325 7.055 -2.19 7.225 ;
      RECT -2.36 6.685 -2.19 7.225 ;
      RECT 8.365 6.605 8.535 6.96 ;
      RECT 8.315 6.605 8.665 6.955 ;
      RECT -2.36 6.685 8.665 6.855 ;
      RECT 7.855 3.71 8.135 3.99 ;
      RECT 7.895 3.665 8.16 3.925 ;
      RECT 7.885 3.7 8.16 3.925 ;
      RECT 7.89 3.685 8.135 3.99 ;
      RECT 7.895 3.662 8.105 3.99 ;
      RECT 7.895 3.66 8.09 3.99 ;
      RECT 7.935 3.65 8.09 3.99 ;
      RECT 7.905 3.655 8.09 3.99 ;
      RECT 7.935 3.647 8.035 3.99 ;
      RECT 7.96 3.64 8.035 3.99 ;
      RECT 7.94 3.642 8.035 3.99 ;
      RECT 7.27 3.155 7.53 3.415 ;
      RECT 7.32 3.147 7.51 3.415 ;
      RECT 7.325 3.067 7.51 3.415 ;
      RECT 7.445 2.455 7.51 3.415 ;
      RECT 7.35 2.852 7.51 3.415 ;
      RECT 7.425 2.54 7.51 3.415 ;
      RECT 7.46 2.165 7.596 2.893 ;
      RECT 7.405 2.662 7.596 2.893 ;
      RECT 7.42 2.602 7.51 3.415 ;
      RECT 7.46 2.165 7.62 2.558 ;
      RECT 7.46 2.165 7.63 2.455 ;
      RECT 7.45 2.165 7.71 2.425 ;
      RECT 5.785 3.565 5.83 3.825 ;
      RECT 5.69 2.1 5.835 2.36 ;
      RECT 6.195 2.722 6.205 2.813 ;
      RECT 6.18 2.66 6.195 2.869 ;
      RECT 6.175 2.607 6.18 2.915 ;
      RECT 6.125 2.554 6.175 3.041 ;
      RECT 6.12 2.509 6.125 3.188 ;
      RECT 6.11 2.497 6.12 3.23 ;
      RECT 6.075 2.461 6.11 3.335 ;
      RECT 6.07 2.429 6.075 3.441 ;
      RECT 6.055 2.411 6.07 3.486 ;
      RECT 6.05 2.394 6.055 2.72 ;
      RECT 6.045 2.775 6.055 3.543 ;
      RECT 6.04 2.38 6.05 2.693 ;
      RECT 6.035 2.83 6.045 3.825 ;
      RECT 6.03 2.366 6.04 2.678 ;
      RECT 6.03 2.88 6.035 3.825 ;
      RECT 6.015 2.343 6.03 2.658 ;
      RECT 5.995 3.002 6.03 3.825 ;
      RECT 6.01 2.325 6.015 2.64 ;
      RECT 6.005 2.317 6.01 2.63 ;
      RECT 5.975 2.285 6.005 2.594 ;
      RECT 5.985 3.13 5.995 3.825 ;
      RECT 5.98 3.157 5.985 3.825 ;
      RECT 5.975 3.207 5.98 3.825 ;
      RECT 5.965 2.251 5.975 2.559 ;
      RECT 5.925 3.275 5.975 3.825 ;
      RECT 5.95 2.228 5.965 2.535 ;
      RECT 5.925 2.1 5.95 2.498 ;
      RECT 5.92 2.1 5.925 2.47 ;
      RECT 5.89 3.375 5.925 3.825 ;
      RECT 5.915 2.1 5.92 2.463 ;
      RECT 5.91 2.1 5.915 2.453 ;
      RECT 5.895 2.1 5.91 2.438 ;
      RECT 5.88 2.1 5.895 2.41 ;
      RECT 5.845 3.48 5.89 3.825 ;
      RECT 5.865 2.1 5.88 2.383 ;
      RECT 5.835 2.1 5.865 2.368 ;
      RECT 5.83 3.552 5.845 3.825 ;
      RECT 5.755 2.635 5.795 2.895 ;
      RECT 5.53 2.582 5.535 2.84 ;
      RECT 1.485 2.06 1.745 2.32 ;
      RECT 1.485 2.085 1.76 2.3 ;
      RECT 3.875 1.91 3.88 2.055 ;
      RECT 5.745 2.63 5.755 2.895 ;
      RECT 5.725 2.622 5.745 2.895 ;
      RECT 5.707 2.618 5.725 2.895 ;
      RECT 5.621 2.607 5.707 2.895 ;
      RECT 5.535 2.59 5.621 2.895 ;
      RECT 5.48 2.577 5.53 2.825 ;
      RECT 5.446 2.569 5.48 2.8 ;
      RECT 5.36 2.558 5.446 2.765 ;
      RECT 5.325 2.535 5.36 2.73 ;
      RECT 5.315 2.497 5.325 2.716 ;
      RECT 5.31 2.47 5.315 2.712 ;
      RECT 5.305 2.457 5.31 2.709 ;
      RECT 5.295 2.437 5.305 2.705 ;
      RECT 5.29 2.412 5.295 2.701 ;
      RECT 5.265 2.367 5.29 2.695 ;
      RECT 5.255 2.308 5.265 2.687 ;
      RECT 5.245 2.276 5.255 2.678 ;
      RECT 5.225 2.228 5.245 2.658 ;
      RECT 5.22 2.188 5.225 2.628 ;
      RECT 5.205 2.162 5.22 2.602 ;
      RECT 5.2 2.14 5.205 2.578 ;
      RECT 5.185 2.112 5.2 2.554 ;
      RECT 5.17 2.085 5.185 2.518 ;
      RECT 5.155 2.062 5.17 2.48 ;
      RECT 5.15 2.052 5.155 2.455 ;
      RECT 5.14 2.045 5.15 2.438 ;
      RECT 5.125 2.032 5.14 2.408 ;
      RECT 5.12 2.022 5.125 2.383 ;
      RECT 5.115 2.017 5.12 2.37 ;
      RECT 5.105 2.01 5.115 2.35 ;
      RECT 5.1 2.003 5.105 2.335 ;
      RECT 5.075 1.996 5.1 2.293 ;
      RECT 5.06 1.986 5.075 2.243 ;
      RECT 5.05 1.981 5.06 2.213 ;
      RECT 5.04 1.977 5.05 2.188 ;
      RECT 5.025 1.974 5.04 2.178 ;
      RECT 4.975 1.971 5.025 2.163 ;
      RECT 4.955 1.969 4.975 2.148 ;
      RECT 4.906 1.967 4.955 2.143 ;
      RECT 4.82 1.963 4.906 2.138 ;
      RECT 4.781 1.96 4.82 2.134 ;
      RECT 4.695 1.956 4.781 2.129 ;
      RECT 4.645 1.953 4.695 2.123 ;
      RECT 4.596 1.95 4.645 2.118 ;
      RECT 4.51 1.947 4.596 2.113 ;
      RECT 4.506 1.945 4.51 2.11 ;
      RECT 4.42 1.942 4.506 2.105 ;
      RECT 4.371 1.938 4.42 2.098 ;
      RECT 4.285 1.935 4.371 2.093 ;
      RECT 4.261 1.932 4.285 2.089 ;
      RECT 4.175 1.93 4.261 2.084 ;
      RECT 4.11 1.926 4.175 2.077 ;
      RECT 4.107 1.925 4.11 2.074 ;
      RECT 4.021 1.922 4.107 2.071 ;
      RECT 3.935 1.916 4.021 2.064 ;
      RECT 3.905 1.912 3.935 2.06 ;
      RECT 3.88 1.91 3.905 2.058 ;
      RECT 3.825 1.907 3.875 2.055 ;
      RECT 3.745 1.906 3.825 2.055 ;
      RECT 3.69 1.908 3.745 2.058 ;
      RECT 3.675 1.909 3.69 2.062 ;
      RECT 3.62 1.917 3.675 2.072 ;
      RECT 3.59 1.925 3.62 2.085 ;
      RECT 3.571 1.926 3.59 2.091 ;
      RECT 3.485 1.929 3.571 2.096 ;
      RECT 3.415 1.934 3.485 2.105 ;
      RECT 3.396 1.937 3.415 2.111 ;
      RECT 3.31 1.941 3.396 2.116 ;
      RECT 3.27 1.945 3.31 2.123 ;
      RECT 3.261 1.947 3.27 2.126 ;
      RECT 3.175 1.951 3.261 2.131 ;
      RECT 3.172 1.954 3.175 2.135 ;
      RECT 3.086 1.957 3.172 2.139 ;
      RECT 3 1.963 3.086 2.147 ;
      RECT 2.976 1.967 3 2.151 ;
      RECT 2.89 1.971 2.976 2.156 ;
      RECT 2.845 1.976 2.89 2.163 ;
      RECT 2.765 1.981 2.845 2.17 ;
      RECT 2.685 1.987 2.765 2.185 ;
      RECT 2.66 1.991 2.685 2.198 ;
      RECT 2.595 1.994 2.66 2.21 ;
      RECT 2.54 1.999 2.595 2.225 ;
      RECT 2.51 2.002 2.54 2.243 ;
      RECT 2.5 2.004 2.51 2.256 ;
      RECT 2.44 2.019 2.5 2.266 ;
      RECT 2.425 2.036 2.44 2.275 ;
      RECT 2.42 2.045 2.425 2.275 ;
      RECT 2.41 2.055 2.42 2.275 ;
      RECT 2.4 2.072 2.41 2.275 ;
      RECT 2.38 2.082 2.4 2.276 ;
      RECT 2.335 2.092 2.38 2.277 ;
      RECT 2.3 2.101 2.335 2.279 ;
      RECT 2.235 2.106 2.3 2.281 ;
      RECT 2.155 2.107 2.235 2.284 ;
      RECT 2.151 2.105 2.155 2.285 ;
      RECT 2.065 2.102 2.151 2.287 ;
      RECT 2.018 2.099 2.065 2.289 ;
      RECT 1.932 2.095 2.018 2.292 ;
      RECT 1.846 2.091 1.932 2.295 ;
      RECT 1.76 2.087 1.846 2.299 ;
      RECT 5.145 3.71 5.175 3.99 ;
      RECT 4.895 3.6 4.915 3.99 ;
      RECT 4.85 3.6 4.915 3.86 ;
      RECT 4.68 2.225 4.715 2.485 ;
      RECT 4.455 2.225 4.515 2.485 ;
      RECT 5.135 3.69 5.145 3.99 ;
      RECT 5.13 3.65 5.135 3.99 ;
      RECT 5.115 3.605 5.13 3.99 ;
      RECT 5.11 3.57 5.115 3.99 ;
      RECT 5.105 3.55 5.11 3.99 ;
      RECT 5.075 3.477 5.105 3.99 ;
      RECT 5.055 3.375 5.075 3.99 ;
      RECT 5.045 3.305 5.055 3.99 ;
      RECT 5 3.245 5.045 3.99 ;
      RECT 4.915 3.206 5 3.99 ;
      RECT 4.91 3.197 4.915 3.57 ;
      RECT 4.9 3.196 4.91 3.553 ;
      RECT 4.875 3.177 4.9 3.523 ;
      RECT 4.87 3.152 4.875 3.502 ;
      RECT 4.86 3.13 4.87 3.493 ;
      RECT 4.855 3.101 4.86 3.483 ;
      RECT 4.815 3.027 4.855 3.455 ;
      RECT 4.795 2.928 4.815 3.42 ;
      RECT 4.78 2.864 4.795 3.403 ;
      RECT 4.75 2.788 4.78 3.375 ;
      RECT 4.73 2.703 4.75 3.348 ;
      RECT 4.69 2.599 4.73 3.255 ;
      RECT 4.685 2.52 4.69 3.163 ;
      RECT 4.68 2.503 4.685 3.14 ;
      RECT 4.675 2.225 4.68 3.12 ;
      RECT 4.645 2.225 4.675 3.058 ;
      RECT 4.64 2.225 4.645 2.99 ;
      RECT 4.63 2.225 4.64 2.955 ;
      RECT 4.62 2.225 4.63 2.92 ;
      RECT 4.555 2.225 4.62 2.775 ;
      RECT 4.55 2.225 4.555 2.645 ;
      RECT 4.52 2.225 4.55 2.578 ;
      RECT 4.515 2.225 4.52 2.503 ;
      RECT 3.695 3.15 3.975 3.43 ;
      RECT 3.735 3.13 3.995 3.39 ;
      RECT 3.725 3.14 3.995 3.39 ;
      RECT 3.735 3.067 3.95 3.43 ;
      RECT 3.79 2.99 3.945 3.43 ;
      RECT 3.795 2.775 3.945 3.43 ;
      RECT 3.785 2.577 3.935 2.828 ;
      RECT 3.775 2.577 3.935 2.695 ;
      RECT 3.77 2.455 3.93 2.598 ;
      RECT 3.755 2.455 3.93 2.503 ;
      RECT 3.75 2.165 3.925 2.48 ;
      RECT 3.735 2.165 3.925 2.45 ;
      RECT 3.695 2.165 3.955 2.425 ;
      RECT 3.605 3.635 3.685 3.895 ;
      RECT 3.01 2.355 3.015 2.62 ;
      RECT 2.89 2.355 3.015 2.615 ;
      RECT 3.565 3.6 3.605 3.895 ;
      RECT 3.52 3.522 3.565 3.895 ;
      RECT 3.5 3.45 3.52 3.895 ;
      RECT 3.49 3.402 3.5 3.895 ;
      RECT 3.455 3.335 3.49 3.895 ;
      RECT 3.425 3.235 3.455 3.895 ;
      RECT 3.405 3.16 3.425 3.695 ;
      RECT 3.395 3.11 3.405 3.65 ;
      RECT 3.39 3.087 3.395 3.623 ;
      RECT 3.385 3.072 3.39 3.61 ;
      RECT 3.38 3.057 3.385 3.588 ;
      RECT 3.375 3.042 3.38 3.57 ;
      RECT 3.35 2.997 3.375 3.525 ;
      RECT 3.34 2.945 3.35 3.468 ;
      RECT 3.33 2.915 3.34 3.435 ;
      RECT 3.32 2.88 3.33 3.403 ;
      RECT 3.285 2.812 3.32 3.335 ;
      RECT 3.28 2.751 3.285 3.27 ;
      RECT 3.27 2.739 3.28 3.25 ;
      RECT 3.265 2.727 3.27 3.23 ;
      RECT 3.26 2.719 3.265 3.218 ;
      RECT 3.255 2.711 3.26 3.198 ;
      RECT 3.245 2.699 3.255 3.17 ;
      RECT 3.235 2.683 3.245 3.14 ;
      RECT 3.21 2.655 3.235 3.078 ;
      RECT 3.2 2.626 3.21 3.023 ;
      RECT 3.185 2.605 3.2 2.983 ;
      RECT 3.18 2.589 3.185 2.955 ;
      RECT 3.175 2.577 3.18 2.945 ;
      RECT 3.17 2.572 3.175 2.918 ;
      RECT 3.165 2.565 3.17 2.905 ;
      RECT 3.15 2.548 3.165 2.878 ;
      RECT 3.14 2.355 3.15 2.838 ;
      RECT 3.13 2.355 3.14 2.805 ;
      RECT 3.12 2.355 3.13 2.78 ;
      RECT 3.05 2.355 3.12 2.715 ;
      RECT 3.04 2.355 3.05 2.663 ;
      RECT 3.025 2.355 3.04 2.645 ;
      RECT 3.015 2.355 3.025 2.63 ;
      RECT 2.845 3.225 3.105 3.485 ;
      RECT 1.38 3.26 1.385 3.467 ;
      RECT 1.015 3.15 1.09 3.465 ;
      RECT 0.83 3.205 0.985 3.465 ;
      RECT 1.015 3.15 1.12 3.43 ;
      RECT 2.83 3.322 2.845 3.483 ;
      RECT 2.805 3.33 2.83 3.488 ;
      RECT 2.78 3.337 2.805 3.493 ;
      RECT 2.717 3.348 2.78 3.502 ;
      RECT 2.631 3.367 2.717 3.519 ;
      RECT 2.545 3.389 2.631 3.538 ;
      RECT 2.53 3.402 2.545 3.549 ;
      RECT 2.49 3.41 2.53 3.556 ;
      RECT 2.47 3.415 2.49 3.563 ;
      RECT 2.432 3.416 2.47 3.566 ;
      RECT 2.346 3.419 2.432 3.567 ;
      RECT 2.26 3.423 2.346 3.568 ;
      RECT 2.211 3.425 2.26 3.57 ;
      RECT 2.125 3.425 2.211 3.572 ;
      RECT 2.085 3.42 2.125 3.574 ;
      RECT 2.075 3.414 2.085 3.575 ;
      RECT 2.035 3.409 2.075 3.572 ;
      RECT 2.025 3.402 2.035 3.568 ;
      RECT 2.01 3.398 2.025 3.566 ;
      RECT 1.993 3.394 2.01 3.564 ;
      RECT 1.907 3.384 1.993 3.556 ;
      RECT 1.821 3.366 1.907 3.542 ;
      RECT 1.735 3.349 1.821 3.528 ;
      RECT 1.71 3.337 1.735 3.519 ;
      RECT 1.64 3.327 1.71 3.512 ;
      RECT 1.595 3.315 1.64 3.503 ;
      RECT 1.535 3.302 1.595 3.495 ;
      RECT 1.53 3.294 1.535 3.49 ;
      RECT 1.495 3.289 1.53 3.488 ;
      RECT 1.44 3.28 1.495 3.481 ;
      RECT 1.4 3.269 1.44 3.473 ;
      RECT 1.385 3.262 1.4 3.469 ;
      RECT 1.365 3.255 1.38 3.466 ;
      RECT 1.35 3.245 1.365 3.464 ;
      RECT 1.335 3.232 1.35 3.461 ;
      RECT 1.31 3.215 1.335 3.457 ;
      RECT 1.295 3.197 1.31 3.454 ;
      RECT 1.27 3.15 1.295 3.452 ;
      RECT 1.246 3.15 1.27 3.449 ;
      RECT 1.16 3.15 1.246 3.441 ;
      RECT 1.12 3.15 1.16 3.433 ;
      RECT 0.985 3.197 1.015 3.465 ;
      RECT 2.665 2.78 2.925 3.04 ;
      RECT 2.625 2.78 2.925 2.918 ;
      RECT 2.59 2.78 2.925 2.903 ;
      RECT 2.535 2.78 2.925 2.883 ;
      RECT 2.455 2.59 2.735 2.87 ;
      RECT 2.455 2.772 2.805 2.87 ;
      RECT 2.455 2.715 2.79 2.87 ;
      RECT 2.455 2.662 2.74 2.87 ;
      RECT 0.285 2.59 0.48 3.375 ;
      RECT 0.365 1.205 0.48 3.375 ;
      RECT 0.22 3.115 0.28 3.375 ;
      RECT 1.59 2.635 1.85 2.895 ;
      RECT 0.275 2.59 0.48 2.87 ;
      RECT 1.585 2.645 1.85 2.83 ;
      RECT 1.3 2.62 1.31 2.77 ;
      RECT 0.535 1.205 0.615 1.55 ;
      RECT 0.27 1.205 0.48 1.55 ;
      RECT 1.575 2.645 1.585 2.829 ;
      RECT 1.565 2.644 1.575 2.826 ;
      RECT 1.556 2.643 1.565 2.824 ;
      RECT 1.47 2.639 1.556 2.814 ;
      RECT 1.396 2.631 1.47 2.796 ;
      RECT 1.31 2.624 1.396 2.779 ;
      RECT 1.25 2.62 1.3 2.769 ;
      RECT 1.215 2.619 1.25 2.766 ;
      RECT 1.16 2.619 1.215 2.768 ;
      RECT 1.125 2.619 1.16 2.772 ;
      RECT 1.039 2.618 1.125 2.779 ;
      RECT 0.953 2.617 1.039 2.789 ;
      RECT 0.867 2.616 0.953 2.8 ;
      RECT 0.781 2.616 0.867 2.81 ;
      RECT 0.695 2.615 0.781 2.82 ;
      RECT 0.66 2.615 0.695 2.86 ;
      RECT 0.655 2.615 0.66 2.903 ;
      RECT 0.63 2.615 0.655 2.92 ;
      RECT 0.555 2.615 0.63 2.935 ;
      RECT 0.535 2.59 0.555 2.948 ;
      RECT 0.53 1.205 0.535 2.958 ;
      RECT 0.505 1.205 0.53 3 ;
      RECT 0.48 1.205 0.505 3.078 ;
      RECT 0.28 2.997 0.285 3.375 ;
      RECT -0.385 2.949 -0.37 3.405 ;
      RECT -0.39 3.021 -0.284 3.403 ;
      RECT -0.37 2.115 -0.235 3.401 ;
      RECT -0.385 2.965 -0.23 3.4 ;
      RECT -0.385 3.015 -0.225 3.398 ;
      RECT -0.4 3.08 -0.225 3.397 ;
      RECT -0.39 3.072 -0.22 3.394 ;
      RECT -0.41 3.12 -0.22 3.389 ;
      RECT -0.41 3.12 -0.205 3.386 ;
      RECT -0.415 3.12 -0.205 3.383 ;
      RECT -0.44 3.12 -0.18 3.38 ;
      RECT -0.37 2.115 -0.21 2.768 ;
      RECT -0.375 2.115 -0.21 2.74 ;
      RECT -0.38 2.115 -0.21 2.568 ;
      RECT -0.38 2.115 -0.19 2.508 ;
      RECT -0.425 2.115 -0.165 2.375 ;
      RECT -0.945 2.59 -0.665 2.87 ;
      RECT -0.955 2.605 -0.665 2.865 ;
      RECT -1 2.667 -0.665 2.863 ;
      RECT -0.925 2.582 -0.76 2.87 ;
      RECT -0.925 2.567 -0.804 2.87 ;
      RECT -0.89 2.56 -0.804 2.87 ;
      RECT -1.425 3.71 -1.145 3.99 ;
      RECT -1.465 3.672 -1.17 3.783 ;
      RECT -1.48 3.622 -1.19 3.678 ;
      RECT -1.535 3.385 -1.275 3.645 ;
      RECT -1.535 3.587 -1.195 3.645 ;
      RECT -1.535 3.527 -1.2 3.645 ;
      RECT -1.535 3.477 -1.22 3.645 ;
      RECT -1.535 3.457 -1.225 3.645 ;
      RECT -1.535 3.435 -1.23 3.645 ;
      RECT -1.535 3.42 -1.26 3.645 ;
      RECT 79.355 7.055 79.73 7.425 ;
      RECT 70.69 0.93 71.065 1.3 ;
      RECT 61.43 7.055 61.805 7.425 ;
      RECT 52.765 0.93 53.14 1.3 ;
      RECT 43.505 7.055 43.88 7.425 ;
      RECT 34.84 0.93 35.215 1.3 ;
      RECT 25.58 7.055 25.955 7.425 ;
      RECT 16.915 0.93 17.29 1.3 ;
      RECT 7.655 7.055 8.03 7.425 ;
      RECT -1.01 0.93 -0.635 1.3 ;
    LAYER via1 ;
      RECT 87.075 7.375 87.225 7.525 ;
      RECT 84.71 6.74 84.86 6.89 ;
      RECT 84.695 2.065 84.845 2.215 ;
      RECT 83.905 2.45 84.055 2.6 ;
      RECT 83.905 6.325 84.055 6.475 ;
      RECT 82.875 2.805 83.025 2.955 ;
      RECT 82.865 5.94 83.015 6.09 ;
      RECT 82.3 3.53 82.45 3.68 ;
      RECT 82.29 1.25 82.44 1.4 ;
      RECT 80.605 2.215 80.755 2.365 ;
      RECT 80.375 6.71 80.525 6.86 ;
      RECT 79.655 3.72 79.805 3.87 ;
      RECT 79.47 7.165 79.62 7.315 ;
      RECT 79.205 2.22 79.355 2.37 ;
      RECT 79.025 3.21 79.175 3.36 ;
      RECT 78.63 3.725 78.78 3.875 ;
      RECT 78.27 3.68 78.42 3.83 ;
      RECT 78.125 2.17 78.275 2.32 ;
      RECT 77.54 3.62 77.69 3.77 ;
      RECT 77.445 2.155 77.595 2.305 ;
      RECT 77.29 2.69 77.44 2.84 ;
      RECT 76.605 3.655 76.755 3.805 ;
      RECT 76.21 2.28 76.36 2.43 ;
      RECT 75.49 3.185 75.64 3.335 ;
      RECT 75.45 2.22 75.6 2.37 ;
      RECT 75.18 3.69 75.33 3.84 ;
      RECT 74.645 2.41 74.795 2.56 ;
      RECT 74.6 3.28 74.75 3.43 ;
      RECT 74.42 2.835 74.57 2.985 ;
      RECT 73.345 2.69 73.495 2.84 ;
      RECT 73.24 2.115 73.39 2.265 ;
      RECT 72.585 3.26 72.735 3.41 ;
      RECT 72.065 1.3 72.215 1.45 ;
      RECT 71.975 3.17 72.125 3.32 ;
      RECT 71.33 2.17 71.48 2.32 ;
      RECT 71.315 3.175 71.465 3.325 ;
      RECT 70.8 2.66 70.95 2.81 ;
      RECT 70.22 3.44 70.37 3.59 ;
      RECT 69.13 6.755 69.28 6.905 ;
      RECT 66.785 6.74 66.935 6.89 ;
      RECT 66.77 2.065 66.92 2.215 ;
      RECT 65.98 2.45 66.13 2.6 ;
      RECT 65.98 6.325 66.13 6.475 ;
      RECT 64.95 2.805 65.1 2.955 ;
      RECT 64.94 5.94 65.09 6.09 ;
      RECT 64.375 3.53 64.525 3.68 ;
      RECT 64.365 1.25 64.515 1.4 ;
      RECT 62.68 2.215 62.83 2.365 ;
      RECT 62.17 6.71 62.32 6.86 ;
      RECT 61.73 3.72 61.88 3.87 ;
      RECT 61.545 7.165 61.695 7.315 ;
      RECT 61.28 2.22 61.43 2.37 ;
      RECT 61.1 3.21 61.25 3.36 ;
      RECT 60.705 3.725 60.855 3.875 ;
      RECT 60.345 3.68 60.495 3.83 ;
      RECT 60.2 2.17 60.35 2.32 ;
      RECT 59.615 3.62 59.765 3.77 ;
      RECT 59.52 2.155 59.67 2.305 ;
      RECT 59.365 2.69 59.515 2.84 ;
      RECT 58.68 3.655 58.83 3.805 ;
      RECT 58.285 2.28 58.435 2.43 ;
      RECT 57.565 3.185 57.715 3.335 ;
      RECT 57.525 2.22 57.675 2.37 ;
      RECT 57.255 3.69 57.405 3.84 ;
      RECT 56.72 2.41 56.87 2.56 ;
      RECT 56.675 3.28 56.825 3.43 ;
      RECT 56.495 2.835 56.645 2.985 ;
      RECT 55.42 2.69 55.57 2.84 ;
      RECT 55.315 2.115 55.465 2.265 ;
      RECT 54.66 3.26 54.81 3.41 ;
      RECT 54.14 1.3 54.29 1.45 ;
      RECT 54.05 3.17 54.2 3.32 ;
      RECT 53.405 2.17 53.555 2.32 ;
      RECT 53.39 3.175 53.54 3.325 ;
      RECT 52.875 2.66 53.025 2.81 ;
      RECT 52.295 3.44 52.445 3.59 ;
      RECT 51.205 6.755 51.355 6.905 ;
      RECT 48.86 6.74 49.01 6.89 ;
      RECT 48.845 2.065 48.995 2.215 ;
      RECT 48.055 2.45 48.205 2.6 ;
      RECT 48.055 6.325 48.205 6.475 ;
      RECT 47.025 2.805 47.175 2.955 ;
      RECT 47.015 5.94 47.165 6.09 ;
      RECT 46.45 3.53 46.6 3.68 ;
      RECT 46.44 1.25 46.59 1.4 ;
      RECT 44.755 2.215 44.905 2.365 ;
      RECT 44.3 6.715 44.45 6.865 ;
      RECT 43.805 3.72 43.955 3.87 ;
      RECT 43.62 7.165 43.77 7.315 ;
      RECT 43.355 2.22 43.505 2.37 ;
      RECT 43.175 3.21 43.325 3.36 ;
      RECT 42.78 3.725 42.93 3.875 ;
      RECT 42.42 3.68 42.57 3.83 ;
      RECT 42.275 2.17 42.425 2.32 ;
      RECT 41.69 3.62 41.84 3.77 ;
      RECT 41.595 2.155 41.745 2.305 ;
      RECT 41.44 2.69 41.59 2.84 ;
      RECT 40.755 3.655 40.905 3.805 ;
      RECT 40.36 2.28 40.51 2.43 ;
      RECT 39.64 3.185 39.79 3.335 ;
      RECT 39.6 2.22 39.75 2.37 ;
      RECT 39.33 3.69 39.48 3.84 ;
      RECT 38.795 2.41 38.945 2.56 ;
      RECT 38.75 3.28 38.9 3.43 ;
      RECT 38.57 2.835 38.72 2.985 ;
      RECT 37.495 2.69 37.645 2.84 ;
      RECT 37.39 2.115 37.54 2.265 ;
      RECT 36.735 3.26 36.885 3.41 ;
      RECT 36.215 1.3 36.365 1.45 ;
      RECT 36.125 3.17 36.275 3.32 ;
      RECT 35.48 2.17 35.63 2.32 ;
      RECT 35.465 3.175 35.615 3.325 ;
      RECT 34.95 2.66 35.1 2.81 ;
      RECT 34.37 3.44 34.52 3.59 ;
      RECT 33.325 6.76 33.475 6.91 ;
      RECT 30.935 6.74 31.085 6.89 ;
      RECT 30.92 2.065 31.07 2.215 ;
      RECT 30.13 2.45 30.28 2.6 ;
      RECT 30.13 6.325 30.28 6.475 ;
      RECT 29.1 2.805 29.25 2.955 ;
      RECT 29.09 5.94 29.24 6.09 ;
      RECT 28.525 3.53 28.675 3.68 ;
      RECT 28.515 1.25 28.665 1.4 ;
      RECT 26.83 2.215 26.98 2.365 ;
      RECT 26.37 6.71 26.52 6.86 ;
      RECT 25.88 3.72 26.03 3.87 ;
      RECT 25.695 7.165 25.845 7.315 ;
      RECT 25.43 2.22 25.58 2.37 ;
      RECT 25.25 3.21 25.4 3.36 ;
      RECT 24.855 3.725 25.005 3.875 ;
      RECT 24.495 3.68 24.645 3.83 ;
      RECT 24.35 2.17 24.5 2.32 ;
      RECT 23.765 3.62 23.915 3.77 ;
      RECT 23.67 2.155 23.82 2.305 ;
      RECT 23.515 2.69 23.665 2.84 ;
      RECT 22.83 3.655 22.98 3.805 ;
      RECT 22.435 2.28 22.585 2.43 ;
      RECT 21.715 3.185 21.865 3.335 ;
      RECT 21.675 2.22 21.825 2.37 ;
      RECT 21.405 3.69 21.555 3.84 ;
      RECT 20.87 2.41 21.02 2.56 ;
      RECT 20.825 3.28 20.975 3.43 ;
      RECT 20.645 2.835 20.795 2.985 ;
      RECT 19.57 2.69 19.72 2.84 ;
      RECT 19.465 2.115 19.615 2.265 ;
      RECT 18.81 3.26 18.96 3.41 ;
      RECT 18.29 1.3 18.44 1.45 ;
      RECT 18.2 3.17 18.35 3.32 ;
      RECT 17.555 2.17 17.705 2.32 ;
      RECT 17.54 3.175 17.69 3.325 ;
      RECT 17.025 2.66 17.175 2.81 ;
      RECT 16.445 3.44 16.595 3.59 ;
      RECT 15.4 6.755 15.55 6.905 ;
      RECT 13.01 6.74 13.16 6.89 ;
      RECT 12.995 2.065 13.145 2.215 ;
      RECT 12.205 2.45 12.355 2.6 ;
      RECT 12.205 6.325 12.355 6.475 ;
      RECT 11.175 2.805 11.325 2.955 ;
      RECT 11.165 5.94 11.315 6.09 ;
      RECT 10.6 3.53 10.75 3.68 ;
      RECT 10.59 1.25 10.74 1.4 ;
      RECT 8.905 2.215 9.055 2.365 ;
      RECT 8.415 6.705 8.565 6.855 ;
      RECT 7.955 3.72 8.105 3.87 ;
      RECT 7.77 7.165 7.92 7.315 ;
      RECT 7.505 2.22 7.655 2.37 ;
      RECT 7.325 3.21 7.475 3.36 ;
      RECT 6.93 3.725 7.08 3.875 ;
      RECT 6.57 3.68 6.72 3.83 ;
      RECT 6.425 2.17 6.575 2.32 ;
      RECT 5.84 3.62 5.99 3.77 ;
      RECT 5.745 2.155 5.895 2.305 ;
      RECT 5.59 2.69 5.74 2.84 ;
      RECT 4.905 3.655 5.055 3.805 ;
      RECT 4.51 2.28 4.66 2.43 ;
      RECT 3.79 3.185 3.94 3.335 ;
      RECT 3.75 2.22 3.9 2.37 ;
      RECT 3.48 3.69 3.63 3.84 ;
      RECT 2.945 2.41 3.095 2.56 ;
      RECT 2.9 3.28 3.05 3.43 ;
      RECT 2.72 2.835 2.87 2.985 ;
      RECT 1.645 2.69 1.795 2.84 ;
      RECT 1.54 2.115 1.69 2.265 ;
      RECT 0.885 3.26 1.035 3.41 ;
      RECT 0.365 1.3 0.515 1.45 ;
      RECT 0.275 3.17 0.425 3.32 ;
      RECT -0.37 2.17 -0.22 2.32 ;
      RECT -0.385 3.175 -0.235 3.325 ;
      RECT -0.9 2.66 -0.75 2.81 ;
      RECT -1.48 3.44 -1.33 3.59 ;
      RECT -3.255 7.095 -3.105 7.245 ;
      RECT -3.63 6.355 -3.48 6.505 ;
    LAYER met1 ;
      RECT 70 1.285 81.96 1.89 ;
      RECT 74.425 0 81.96 1.89 ;
      RECT 52.075 1.285 64.035 1.89 ;
      RECT 56.5 0 64.035 1.89 ;
      RECT 34.15 1.285 46.11 1.89 ;
      RECT 38.575 0 46.11 1.89 ;
      RECT 16.225 1.285 28.185 1.89 ;
      RECT 20.65 0 28.185 1.89 ;
      RECT -1.7 1.285 10.26 1.89 ;
      RECT 2.725 0 10.26 1.89 ;
      RECT 69.995 0 70.74 1.68 ;
      RECT 52.07 0 52.815 1.68 ;
      RECT 34.145 0 34.89 1.68 ;
      RECT 16.22 0 16.965 1.68 ;
      RECT -1.705 0 -0.96 1.68 ;
      RECT 72.99 0 74.145 1.89 ;
      RECT 69.995 1.255 72.71 1.68 ;
      RECT 71.02 0 72.71 1.89 ;
      RECT 55.065 0 56.22 1.89 ;
      RECT 52.07 1.255 54.785 1.68 ;
      RECT 53.095 0 54.785 1.89 ;
      RECT 37.14 0 38.295 1.89 ;
      RECT 34.145 1.255 36.86 1.68 ;
      RECT 35.17 0 36.86 1.89 ;
      RECT 19.215 0 20.37 1.89 ;
      RECT 16.22 1.255 18.935 1.68 ;
      RECT 17.245 0 18.935 1.89 ;
      RECT 1.29 0 2.445 1.89 ;
      RECT -1.705 1.255 1.01 1.68 ;
      RECT -0.68 0 1.01 1.89 ;
      RECT 71.02 0 81.96 1.005 ;
      RECT 53.095 0 64.035 1.005 ;
      RECT 35.17 0 46.11 1.005 ;
      RECT 17.245 0 28.185 1.005 ;
      RECT -0.68 0 10.26 1.005 ;
      RECT 69.995 0 81.96 0.975 ;
      RECT 52.07 0 64.035 0.975 ;
      RECT 34.145 0 46.11 0.975 ;
      RECT 16.22 0 28.185 0.975 ;
      RECT -1.705 0 10.26 0.975 ;
      RECT -4.865 0 87.55 0.305 ;
      RECT -4.865 4.285 87.55 4.745 ;
      RECT 70 4.135 87.55 4.745 ;
      RECT 52.075 4.135 69.625 4.745 ;
      RECT 34.15 4.135 51.7 4.745 ;
      RECT 16.225 4.135 33.775 4.745 ;
      RECT -1.7 4.135 15.85 4.745 ;
      RECT 70 4.13 81.96 4.745 ;
      RECT 52.075 4.13 64.035 4.745 ;
      RECT 34.15 4.13 46.11 4.745 ;
      RECT 16.225 4.13 28.185 4.745 ;
      RECT -1.7 4.13 10.26 4.745 ;
      RECT -4.885 8.575 87.55 8.88 ;
      RECT 78.695 6.315 78.865 8.88 ;
      RECT 60.77 6.315 60.94 8.88 ;
      RECT 42.845 6.315 43.015 8.88 ;
      RECT 24.92 6.315 25.09 8.88 ;
      RECT 6.995 6.315 7.165 8.88 ;
      RECT 79.03 6.285 79.32 6.515 ;
      RECT 61.105 6.285 61.395 6.515 ;
      RECT 43.18 6.285 43.47 6.515 ;
      RECT 25.255 6.285 25.545 6.515 ;
      RECT 7.33 6.285 7.62 6.515 ;
      RECT 78.695 6.315 79.32 6.485 ;
      RECT 60.77 6.315 61.395 6.485 ;
      RECT 42.845 6.315 43.47 6.485 ;
      RECT 24.92 6.315 25.545 6.485 ;
      RECT 6.995 6.315 7.62 6.485 ;
      RECT 86.95 7.765 87.24 7.995 ;
      RECT 87.01 6.285 87.18 7.995 ;
      RECT 86.975 7.275 87.325 7.625 ;
      RECT 86.95 6.285 87.24 6.515 ;
      RECT 86.95 2.365 87.24 2.595 ;
      RECT 87.01 0.885 87.18 2.595 ;
      RECT 86.95 0.885 87.24 1.115 ;
      RECT 86.54 2.735 86.87 2.965 ;
      RECT 86.54 2.765 87.04 2.935 ;
      RECT 86.54 2.395 86.73 2.965 ;
      RECT 85.96 2.365 86.25 2.595 ;
      RECT 85.96 2.395 86.73 2.565 ;
      RECT 86.02 0.885 86.19 2.595 ;
      RECT 85.96 0.885 86.25 1.115 ;
      RECT 85.96 7.765 86.25 7.995 ;
      RECT 86.02 6.285 86.19 7.995 ;
      RECT 85.96 6.285 86.25 6.515 ;
      RECT 85.96 6.325 86.81 6.485 ;
      RECT 86.64 5.915 86.81 6.485 ;
      RECT 85.96 6.32 86.35 6.485 ;
      RECT 86.58 5.915 86.87 6.145 ;
      RECT 86.58 5.945 87.04 6.115 ;
      RECT 85.59 2.735 85.88 2.965 ;
      RECT 85.59 2.765 86.05 2.935 ;
      RECT 85.65 1.655 85.815 2.965 ;
      RECT 84.165 1.625 84.455 1.855 ;
      RECT 84.165 1.655 85.815 1.825 ;
      RECT 84.225 0.885 84.395 1.855 ;
      RECT 84.165 0.885 84.455 1.115 ;
      RECT 84.165 7.765 84.455 7.995 ;
      RECT 84.225 7.025 84.395 7.995 ;
      RECT 84.225 7.12 85.815 7.29 ;
      RECT 85.645 5.915 85.815 7.29 ;
      RECT 84.165 7.025 84.455 7.255 ;
      RECT 85.59 5.915 85.88 6.145 ;
      RECT 85.59 5.945 86.05 6.115 ;
      RECT 82.2 3.43 82.55 3.78 ;
      RECT 82.29 2.025 82.46 3.78 ;
      RECT 84.595 1.965 84.945 2.315 ;
      RECT 82.29 2.025 83.91 2.2 ;
      RECT 82.29 2.025 84.945 2.195 ;
      RECT 84.62 6.655 84.945 6.98 ;
      RECT 80.275 6.61 80.625 6.96 ;
      RECT 84.595 6.655 84.945 6.885 ;
      RECT 79.835 6.655 80.125 6.885 ;
      RECT 79.665 6.685 84.945 6.855 ;
      RECT 83.82 2.365 84.14 2.685 ;
      RECT 83.79 2.365 84.14 2.595 ;
      RECT 83.62 2.395 84.14 2.565 ;
      RECT 83.82 6.225 84.14 6.545 ;
      RECT 83.79 6.285 84.14 6.515 ;
      RECT 83.62 6.315 84.14 6.485 ;
      RECT 82.775 2.705 83.125 3.055 ;
      RECT 82.775 2.765 83.255 2.935 ;
      RECT 82.765 5.84 83.115 6.19 ;
      RECT 78.035 5.915 78.325 6.145 ;
      RECT 78.035 5.945 83.255 6.115 ;
      RECT 79.6 3.665 79.64 3.925 ;
      RECT 79.64 3.645 79.645 3.655 ;
      RECT 80.97 2.89 80.98 3.111 ;
      RECT 80.9 2.885 80.97 3.236 ;
      RECT 80.89 2.885 80.9 3.363 ;
      RECT 80.865 2.885 80.89 3.41 ;
      RECT 80.84 2.885 80.865 3.488 ;
      RECT 80.82 2.885 80.84 3.558 ;
      RECT 80.795 2.885 80.82 3.598 ;
      RECT 80.785 2.885 80.795 3.618 ;
      RECT 80.775 2.887 80.785 3.626 ;
      RECT 80.77 2.892 80.775 3.083 ;
      RECT 80.77 3.092 80.775 3.627 ;
      RECT 80.765 3.137 80.77 3.628 ;
      RECT 80.755 3.202 80.765 3.629 ;
      RECT 80.745 3.297 80.755 3.631 ;
      RECT 80.74 3.35 80.745 3.633 ;
      RECT 80.735 3.37 80.74 3.634 ;
      RECT 80.68 3.395 80.735 3.64 ;
      RECT 80.64 3.43 80.68 3.649 ;
      RECT 80.63 3.447 80.64 3.654 ;
      RECT 80.621 3.453 80.63 3.656 ;
      RECT 80.535 3.491 80.621 3.667 ;
      RECT 80.53 3.53 80.535 3.677 ;
      RECT 80.455 3.537 80.53 3.687 ;
      RECT 80.435 3.547 80.455 3.698 ;
      RECT 80.405 3.554 80.435 3.706 ;
      RECT 80.38 3.561 80.405 3.713 ;
      RECT 80.356 3.567 80.38 3.718 ;
      RECT 80.27 3.58 80.356 3.73 ;
      RECT 80.192 3.587 80.27 3.748 ;
      RECT 80.106 3.582 80.192 3.766 ;
      RECT 80.02 3.577 80.106 3.786 ;
      RECT 79.94 3.571 80.02 3.803 ;
      RECT 79.875 3.567 79.94 3.832 ;
      RECT 79.87 3.281 79.875 3.305 ;
      RECT 79.86 3.557 79.875 3.86 ;
      RECT 79.865 3.275 79.87 3.345 ;
      RECT 79.86 3.269 79.865 3.415 ;
      RECT 79.855 3.263 79.86 3.493 ;
      RECT 79.855 3.54 79.86 3.925 ;
      RECT 79.847 3.26 79.855 3.925 ;
      RECT 79.761 3.258 79.847 3.925 ;
      RECT 79.675 3.256 79.761 3.925 ;
      RECT 79.665 3.257 79.675 3.925 ;
      RECT 79.66 3.262 79.665 3.925 ;
      RECT 79.65 3.275 79.66 3.925 ;
      RECT 79.645 3.297 79.65 3.925 ;
      RECT 79.64 3.657 79.645 3.925 ;
      RECT 80.27 3.125 80.275 3.345 ;
      RECT 80.775 2.16 80.81 2.42 ;
      RECT 80.76 2.16 80.775 2.428 ;
      RECT 80.731 2.16 80.76 2.45 ;
      RECT 80.645 2.16 80.731 2.51 ;
      RECT 80.625 2.16 80.645 2.575 ;
      RECT 80.565 2.16 80.625 2.74 ;
      RECT 80.56 2.16 80.565 2.888 ;
      RECT 80.555 2.16 80.56 2.9 ;
      RECT 80.55 2.16 80.555 2.926 ;
      RECT 80.52 2.346 80.55 3.006 ;
      RECT 80.515 2.394 80.52 3.095 ;
      RECT 80.51 2.408 80.515 3.11 ;
      RECT 80.505 2.427 80.51 3.14 ;
      RECT 80.5 2.442 80.505 3.156 ;
      RECT 80.495 2.457 80.5 3.178 ;
      RECT 80.49 2.477 80.495 3.2 ;
      RECT 80.48 2.497 80.49 3.233 ;
      RECT 80.465 2.539 80.48 3.295 ;
      RECT 80.46 2.57 80.465 3.335 ;
      RECT 80.455 2.582 80.46 3.34 ;
      RECT 80.45 2.594 80.455 3.345 ;
      RECT 80.445 2.607 80.45 3.345 ;
      RECT 80.44 2.625 80.445 3.345 ;
      RECT 80.435 2.645 80.44 3.345 ;
      RECT 80.43 2.657 80.435 3.345 ;
      RECT 80.425 2.67 80.43 3.345 ;
      RECT 80.405 2.705 80.425 3.345 ;
      RECT 80.355 2.807 80.405 3.345 ;
      RECT 80.35 2.892 80.355 3.345 ;
      RECT 80.345 2.9 80.35 3.345 ;
      RECT 80.34 2.917 80.345 3.345 ;
      RECT 80.335 2.932 80.34 3.345 ;
      RECT 80.3 2.997 80.335 3.345 ;
      RECT 80.285 3.062 80.3 3.345 ;
      RECT 80.28 3.092 80.285 3.345 ;
      RECT 80.275 3.117 80.28 3.345 ;
      RECT 80.26 3.127 80.27 3.345 ;
      RECT 80.245 3.14 80.26 3.338 ;
      RECT 79.99 2.73 80.06 2.94 ;
      RECT 79.78 2.707 79.785 2.9 ;
      RECT 77.235 2.635 77.495 2.895 ;
      RECT 80.07 2.917 80.075 2.92 ;
      RECT 80.06 2.735 80.07 2.935 ;
      RECT 79.961 2.728 79.99 2.94 ;
      RECT 79.875 2.72 79.961 2.94 ;
      RECT 79.86 2.714 79.875 2.938 ;
      RECT 79.84 2.713 79.86 2.925 ;
      RECT 79.835 2.712 79.84 2.908 ;
      RECT 79.785 2.709 79.835 2.903 ;
      RECT 79.755 2.706 79.78 2.898 ;
      RECT 79.735 2.704 79.755 2.893 ;
      RECT 79.72 2.702 79.735 2.89 ;
      RECT 79.69 2.7 79.72 2.888 ;
      RECT 79.625 2.696 79.69 2.88 ;
      RECT 79.595 2.691 79.625 2.875 ;
      RECT 79.575 2.689 79.595 2.873 ;
      RECT 79.545 2.686 79.575 2.868 ;
      RECT 79.485 2.682 79.545 2.86 ;
      RECT 79.48 2.679 79.485 2.855 ;
      RECT 79.41 2.677 79.48 2.85 ;
      RECT 79.381 2.673 79.41 2.843 ;
      RECT 79.295 2.668 79.381 2.835 ;
      RECT 79.261 2.663 79.295 2.827 ;
      RECT 79.175 2.655 79.261 2.819 ;
      RECT 79.136 2.648 79.175 2.811 ;
      RECT 79.05 2.643 79.136 2.803 ;
      RECT 78.985 2.637 79.05 2.793 ;
      RECT 78.965 2.632 78.985 2.788 ;
      RECT 78.956 2.629 78.965 2.787 ;
      RECT 78.87 2.625 78.956 2.781 ;
      RECT 78.83 2.621 78.87 2.773 ;
      RECT 78.81 2.617 78.83 2.771 ;
      RECT 78.75 2.617 78.81 2.768 ;
      RECT 78.73 2.62 78.75 2.766 ;
      RECT 78.709 2.62 78.73 2.766 ;
      RECT 78.623 2.622 78.709 2.77 ;
      RECT 78.537 2.624 78.623 2.776 ;
      RECT 78.451 2.626 78.537 2.783 ;
      RECT 78.365 2.629 78.451 2.789 ;
      RECT 78.331 2.63 78.365 2.794 ;
      RECT 78.245 2.633 78.331 2.799 ;
      RECT 78.216 2.64 78.245 2.804 ;
      RECT 78.13 2.64 78.216 2.809 ;
      RECT 78.097 2.64 78.13 2.814 ;
      RECT 78.011 2.642 78.097 2.819 ;
      RECT 77.925 2.644 78.011 2.826 ;
      RECT 77.861 2.646 77.925 2.832 ;
      RECT 77.775 2.648 77.861 2.838 ;
      RECT 77.772 2.65 77.775 2.841 ;
      RECT 77.686 2.651 77.772 2.845 ;
      RECT 77.6 2.654 77.686 2.852 ;
      RECT 77.581 2.656 77.6 2.856 ;
      RECT 77.495 2.658 77.581 2.861 ;
      RECT 77.225 2.67 77.235 2.865 ;
      RECT 79.405 7.765 79.695 7.995 ;
      RECT 79.465 7.025 79.635 7.995 ;
      RECT 79.355 7.055 79.73 7.425 ;
      RECT 79.405 7.025 79.695 7.425 ;
      RECT 79.46 2.25 79.645 2.46 ;
      RECT 79.455 2.251 79.65 2.458 ;
      RECT 79.45 2.256 79.66 2.453 ;
      RECT 79.445 2.232 79.45 2.45 ;
      RECT 79.415 2.229 79.445 2.443 ;
      RECT 79.41 2.225 79.415 2.434 ;
      RECT 79.375 2.256 79.66 2.429 ;
      RECT 79.15 2.165 79.41 2.425 ;
      RECT 79.45 2.234 79.455 2.453 ;
      RECT 79.455 2.235 79.46 2.458 ;
      RECT 79.15 2.247 79.53 2.425 ;
      RECT 79.15 2.245 79.515 2.425 ;
      RECT 79.15 2.24 79.505 2.425 ;
      RECT 79.105 3.155 79.155 3.44 ;
      RECT 79.05 3.125 79.055 3.44 ;
      RECT 79.02 3.105 79.025 3.44 ;
      RECT 79.17 3.155 79.23 3.415 ;
      RECT 79.165 3.155 79.17 3.423 ;
      RECT 79.155 3.155 79.165 3.435 ;
      RECT 79.07 3.145 79.105 3.44 ;
      RECT 79.065 3.132 79.07 3.44 ;
      RECT 79.055 3.127 79.065 3.44 ;
      RECT 79.035 3.117 79.05 3.44 ;
      RECT 79.025 3.11 79.035 3.44 ;
      RECT 79.015 3.102 79.02 3.44 ;
      RECT 78.985 3.092 79.015 3.44 ;
      RECT 78.97 3.08 78.985 3.44 ;
      RECT 78.955 3.07 78.97 3.435 ;
      RECT 78.935 3.06 78.955 3.41 ;
      RECT 78.925 3.052 78.935 3.387 ;
      RECT 78.895 3.035 78.925 3.377 ;
      RECT 78.89 3.012 78.895 3.368 ;
      RECT 78.885 2.999 78.89 3.366 ;
      RECT 78.87 2.975 78.885 3.36 ;
      RECT 78.865 2.951 78.87 3.354 ;
      RECT 78.855 2.94 78.865 3.349 ;
      RECT 78.85 2.93 78.855 3.345 ;
      RECT 78.845 2.922 78.85 3.342 ;
      RECT 78.835 2.917 78.845 3.338 ;
      RECT 78.83 2.912 78.835 3.334 ;
      RECT 78.745 2.91 78.83 3.309 ;
      RECT 78.715 2.91 78.745 3.275 ;
      RECT 78.7 2.91 78.715 3.258 ;
      RECT 78.645 2.91 78.7 3.203 ;
      RECT 78.64 2.915 78.645 3.152 ;
      RECT 78.63 2.92 78.64 3.142 ;
      RECT 78.625 2.93 78.63 3.128 ;
      RECT 78.575 3.67 78.835 3.93 ;
      RECT 78.495 3.685 78.835 3.906 ;
      RECT 78.475 3.685 78.835 3.901 ;
      RECT 78.451 3.685 78.835 3.899 ;
      RECT 78.365 3.685 78.835 3.894 ;
      RECT 78.215 3.625 78.475 3.89 ;
      RECT 78.17 3.685 78.835 3.885 ;
      RECT 78.165 3.692 78.835 3.88 ;
      RECT 78.18 3.68 78.495 3.89 ;
      RECT 78.07 2.115 78.33 2.375 ;
      RECT 78.07 2.172 78.335 2.368 ;
      RECT 78.07 2.202 78.34 2.3 ;
      RECT 78.13 2.633 78.245 2.635 ;
      RECT 78.216 2.63 78.245 2.635 ;
      RECT 77.24 3.634 77.265 3.874 ;
      RECT 77.225 3.637 77.315 3.868 ;
      RECT 77.22 3.642 77.401 3.863 ;
      RECT 77.215 3.65 77.465 3.861 ;
      RECT 77.215 3.65 77.475 3.86 ;
      RECT 77.21 3.657 77.485 3.853 ;
      RECT 77.21 3.657 77.571 3.842 ;
      RECT 77.205 3.692 77.571 3.838 ;
      RECT 77.205 3.692 77.58 3.827 ;
      RECT 77.485 3.565 77.745 3.825 ;
      RECT 77.195 3.742 77.745 3.823 ;
      RECT 77.465 3.61 77.485 3.858 ;
      RECT 77.401 3.613 77.465 3.862 ;
      RECT 77.315 3.618 77.401 3.867 ;
      RECT 77.245 3.629 77.745 3.825 ;
      RECT 77.265 3.623 77.315 3.872 ;
      RECT 77.39 2.1 77.4 2.362 ;
      RECT 77.38 2.157 77.39 2.365 ;
      RECT 77.355 2.162 77.38 2.371 ;
      RECT 77.33 2.166 77.355 2.383 ;
      RECT 77.32 2.169 77.33 2.393 ;
      RECT 77.315 2.17 77.32 2.398 ;
      RECT 77.31 2.171 77.315 2.403 ;
      RECT 77.305 2.172 77.31 2.405 ;
      RECT 77.28 2.175 77.305 2.408 ;
      RECT 77.25 2.181 77.28 2.411 ;
      RECT 77.185 2.192 77.25 2.414 ;
      RECT 77.14 2.2 77.185 2.418 ;
      RECT 77.125 2.2 77.14 2.426 ;
      RECT 77.12 2.201 77.125 2.433 ;
      RECT 77.115 2.203 77.12 2.436 ;
      RECT 77.11 2.207 77.115 2.439 ;
      RECT 77.1 2.215 77.11 2.443 ;
      RECT 77.095 2.228 77.1 2.448 ;
      RECT 77.09 2.236 77.095 2.45 ;
      RECT 77.085 2.242 77.09 2.45 ;
      RECT 77.08 2.246 77.085 2.453 ;
      RECT 77.075 2.248 77.08 2.456 ;
      RECT 77.07 2.251 77.075 2.459 ;
      RECT 77.06 2.256 77.07 2.463 ;
      RECT 77.055 2.262 77.06 2.468 ;
      RECT 77.045 2.268 77.055 2.472 ;
      RECT 77.03 2.275 77.045 2.478 ;
      RECT 77.001 2.289 77.03 2.488 ;
      RECT 76.915 2.324 77.001 2.52 ;
      RECT 76.895 2.357 76.915 2.549 ;
      RECT 76.875 2.37 76.895 2.56 ;
      RECT 76.855 2.382 76.875 2.571 ;
      RECT 76.805 2.404 76.855 2.591 ;
      RECT 76.79 2.422 76.805 2.608 ;
      RECT 76.785 2.428 76.79 2.611 ;
      RECT 76.78 2.432 76.785 2.614 ;
      RECT 76.775 2.436 76.78 2.618 ;
      RECT 76.77 2.438 76.775 2.621 ;
      RECT 76.76 2.445 76.77 2.624 ;
      RECT 76.755 2.45 76.76 2.628 ;
      RECT 76.75 2.452 76.755 2.631 ;
      RECT 76.745 2.456 76.75 2.634 ;
      RECT 76.74 2.458 76.745 2.638 ;
      RECT 76.725 2.463 76.74 2.643 ;
      RECT 76.72 2.468 76.725 2.646 ;
      RECT 76.715 2.476 76.72 2.649 ;
      RECT 76.71 2.478 76.715 2.652 ;
      RECT 76.705 2.48 76.71 2.655 ;
      RECT 76.695 2.482 76.705 2.661 ;
      RECT 76.66 2.496 76.695 2.673 ;
      RECT 76.65 2.511 76.66 2.683 ;
      RECT 76.575 2.54 76.65 2.707 ;
      RECT 76.57 2.565 76.575 2.73 ;
      RECT 76.555 2.569 76.57 2.736 ;
      RECT 76.545 2.577 76.555 2.741 ;
      RECT 76.515 2.59 76.545 2.745 ;
      RECT 76.505 2.605 76.515 2.75 ;
      RECT 76.495 2.61 76.505 2.753 ;
      RECT 76.49 2.612 76.495 2.755 ;
      RECT 76.475 2.615 76.49 2.758 ;
      RECT 76.47 2.617 76.475 2.761 ;
      RECT 76.45 2.622 76.47 2.765 ;
      RECT 76.42 2.627 76.45 2.773 ;
      RECT 76.395 2.634 76.42 2.781 ;
      RECT 76.39 2.639 76.395 2.786 ;
      RECT 76.36 2.642 76.39 2.79 ;
      RECT 76.32 2.645 76.36 2.8 ;
      RECT 76.285 2.642 76.32 2.812 ;
      RECT 76.275 2.638 76.285 2.819 ;
      RECT 76.25 2.634 76.275 2.825 ;
      RECT 76.245 2.63 76.25 2.83 ;
      RECT 76.205 2.627 76.245 2.83 ;
      RECT 76.19 2.612 76.205 2.831 ;
      RECT 76.167 2.6 76.19 2.831 ;
      RECT 76.081 2.6 76.167 2.832 ;
      RECT 75.995 2.6 76.081 2.834 ;
      RECT 75.975 2.6 75.995 2.831 ;
      RECT 75.97 2.605 75.975 2.826 ;
      RECT 75.965 2.61 75.97 2.824 ;
      RECT 75.955 2.62 75.965 2.822 ;
      RECT 75.95 2.626 75.955 2.815 ;
      RECT 75.945 2.628 75.95 2.8 ;
      RECT 75.94 2.632 75.945 2.79 ;
      RECT 77.4 2.1 77.65 2.36 ;
      RECT 75.125 3.635 75.385 3.895 ;
      RECT 77.42 3.125 77.425 3.335 ;
      RECT 77.425 3.13 77.435 3.33 ;
      RECT 77.375 3.125 77.42 3.35 ;
      RECT 77.365 3.125 77.375 3.37 ;
      RECT 77.346 3.125 77.365 3.375 ;
      RECT 77.26 3.125 77.346 3.372 ;
      RECT 77.23 3.127 77.26 3.37 ;
      RECT 77.175 3.137 77.23 3.368 ;
      RECT 77.11 3.151 77.175 3.366 ;
      RECT 77.105 3.159 77.11 3.365 ;
      RECT 77.09 3.162 77.105 3.363 ;
      RECT 77.025 3.172 77.09 3.359 ;
      RECT 76.977 3.186 77.025 3.36 ;
      RECT 76.891 3.203 76.977 3.374 ;
      RECT 76.805 3.224 76.891 3.391 ;
      RECT 76.785 3.237 76.805 3.401 ;
      RECT 76.74 3.245 76.785 3.408 ;
      RECT 76.705 3.253 76.74 3.416 ;
      RECT 76.671 3.261 76.705 3.424 ;
      RECT 76.585 3.275 76.671 3.436 ;
      RECT 76.55 3.292 76.585 3.448 ;
      RECT 76.541 3.301 76.55 3.452 ;
      RECT 76.455 3.319 76.541 3.469 ;
      RECT 76.396 3.346 76.455 3.496 ;
      RECT 76.31 3.373 76.396 3.524 ;
      RECT 76.29 3.395 76.31 3.544 ;
      RECT 76.23 3.41 76.29 3.56 ;
      RECT 76.22 3.422 76.23 3.573 ;
      RECT 76.215 3.427 76.22 3.576 ;
      RECT 76.205 3.43 76.215 3.579 ;
      RECT 76.2 3.432 76.205 3.582 ;
      RECT 76.17 3.44 76.2 3.589 ;
      RECT 76.155 3.447 76.17 3.597 ;
      RECT 76.145 3.452 76.155 3.601 ;
      RECT 76.14 3.455 76.145 3.604 ;
      RECT 76.13 3.457 76.14 3.607 ;
      RECT 76.095 3.467 76.13 3.616 ;
      RECT 76.02 3.49 76.095 3.638 ;
      RECT 76 3.508 76.02 3.656 ;
      RECT 75.97 3.515 76 3.666 ;
      RECT 75.95 3.523 75.97 3.676 ;
      RECT 75.94 3.529 75.95 3.683 ;
      RECT 75.921 3.534 75.94 3.689 ;
      RECT 75.835 3.554 75.921 3.709 ;
      RECT 75.82 3.574 75.835 3.728 ;
      RECT 75.775 3.586 75.82 3.739 ;
      RECT 75.71 3.607 75.775 3.762 ;
      RECT 75.67 3.627 75.71 3.783 ;
      RECT 75.66 3.637 75.67 3.793 ;
      RECT 75.61 3.649 75.66 3.804 ;
      RECT 75.59 3.665 75.61 3.816 ;
      RECT 75.56 3.675 75.59 3.822 ;
      RECT 75.55 3.68 75.56 3.824 ;
      RECT 75.481 3.681 75.55 3.83 ;
      RECT 75.395 3.683 75.481 3.84 ;
      RECT 75.385 3.684 75.395 3.845 ;
      RECT 76.655 3.71 76.845 3.92 ;
      RECT 76.645 3.715 76.855 3.913 ;
      RECT 76.63 3.715 76.855 3.878 ;
      RECT 76.55 3.6 76.81 3.86 ;
      RECT 75.465 3.13 75.65 3.425 ;
      RECT 75.455 3.13 75.65 3.423 ;
      RECT 75.44 3.13 75.655 3.418 ;
      RECT 75.44 3.13 75.66 3.415 ;
      RECT 75.435 3.13 75.66 3.413 ;
      RECT 75.43 3.385 75.66 3.403 ;
      RECT 75.435 3.13 75.695 3.39 ;
      RECT 75.395 2.165 75.655 2.425 ;
      RECT 75.205 2.09 75.291 2.423 ;
      RECT 75.18 2.094 75.335 2.419 ;
      RECT 75.291 2.086 75.335 2.419 ;
      RECT 75.291 2.087 75.34 2.418 ;
      RECT 75.205 2.092 75.355 2.417 ;
      RECT 75.18 2.1 75.395 2.416 ;
      RECT 75.175 2.095 75.355 2.411 ;
      RECT 75.165 2.11 75.395 2.318 ;
      RECT 75.165 2.162 75.595 2.318 ;
      RECT 75.165 2.155 75.575 2.318 ;
      RECT 75.165 2.142 75.545 2.318 ;
      RECT 75.165 2.13 75.485 2.318 ;
      RECT 75.165 2.115 75.46 2.318 ;
      RECT 74.365 2.745 74.5 3.04 ;
      RECT 74.625 2.768 74.63 2.955 ;
      RECT 75.345 2.665 75.49 2.9 ;
      RECT 75.505 2.665 75.51 2.89 ;
      RECT 75.54 2.676 75.545 2.87 ;
      RECT 75.535 2.668 75.54 2.875 ;
      RECT 75.515 2.665 75.535 2.88 ;
      RECT 75.51 2.665 75.515 2.888 ;
      RECT 75.5 2.665 75.505 2.893 ;
      RECT 75.49 2.665 75.5 2.898 ;
      RECT 75.32 2.667 75.345 2.9 ;
      RECT 75.27 2.674 75.32 2.9 ;
      RECT 75.265 2.679 75.27 2.9 ;
      RECT 75.226 2.684 75.265 2.901 ;
      RECT 75.14 2.696 75.226 2.902 ;
      RECT 75.131 2.706 75.14 2.902 ;
      RECT 75.045 2.715 75.131 2.904 ;
      RECT 75.021 2.725 75.045 2.906 ;
      RECT 74.935 2.736 75.021 2.907 ;
      RECT 74.905 2.747 74.935 2.909 ;
      RECT 74.875 2.752 74.905 2.911 ;
      RECT 74.85 2.758 74.875 2.914 ;
      RECT 74.835 2.763 74.85 2.915 ;
      RECT 74.79 2.769 74.835 2.915 ;
      RECT 74.785 2.774 74.79 2.916 ;
      RECT 74.765 2.774 74.785 2.918 ;
      RECT 74.745 2.772 74.765 2.923 ;
      RECT 74.71 2.771 74.745 2.93 ;
      RECT 74.68 2.77 74.71 2.94 ;
      RECT 74.63 2.769 74.68 2.95 ;
      RECT 74.54 2.766 74.625 3.04 ;
      RECT 74.515 2.76 74.54 3.04 ;
      RECT 74.5 2.75 74.515 3.04 ;
      RECT 74.315 2.745 74.365 2.96 ;
      RECT 74.305 2.75 74.315 2.95 ;
      RECT 74.545 3.225 74.805 3.485 ;
      RECT 74.545 3.225 74.835 3.378 ;
      RECT 74.545 3.225 74.87 3.363 ;
      RECT 74.8 3.145 74.99 3.355 ;
      RECT 74.79 3.15 75 3.348 ;
      RECT 74.755 3.22 75 3.348 ;
      RECT 74.785 3.162 74.805 3.485 ;
      RECT 74.77 3.21 75 3.348 ;
      RECT 74.775 3.182 74.805 3.485 ;
      RECT 73.855 2.25 73.925 3.355 ;
      RECT 74.59 2.355 74.85 2.615 ;
      RECT 74.17 2.401 74.185 2.61 ;
      RECT 74.506 2.414 74.59 2.565 ;
      RECT 74.42 2.411 74.506 2.565 ;
      RECT 74.381 2.409 74.42 2.565 ;
      RECT 74.295 2.407 74.381 2.565 ;
      RECT 74.235 2.405 74.295 2.576 ;
      RECT 74.2 2.403 74.235 2.594 ;
      RECT 74.185 2.401 74.2 2.605 ;
      RECT 74.155 2.401 74.17 2.618 ;
      RECT 74.145 2.401 74.155 2.623 ;
      RECT 74.12 2.4 74.145 2.628 ;
      RECT 74.105 2.395 74.12 2.634 ;
      RECT 74.1 2.388 74.105 2.639 ;
      RECT 74.075 2.379 74.1 2.645 ;
      RECT 74.03 2.358 74.075 2.658 ;
      RECT 74.02 2.342 74.03 2.668 ;
      RECT 74.005 2.335 74.02 2.678 ;
      RECT 73.995 2.328 74.005 2.695 ;
      RECT 73.99 2.325 73.995 2.725 ;
      RECT 73.985 2.323 73.99 2.755 ;
      RECT 73.98 2.321 73.985 2.792 ;
      RECT 73.965 2.317 73.98 2.859 ;
      RECT 73.965 3.15 73.975 3.35 ;
      RECT 73.96 2.313 73.965 2.985 ;
      RECT 73.96 3.137 73.965 3.355 ;
      RECT 73.955 2.311 73.96 3.07 ;
      RECT 73.955 3.127 73.96 3.355 ;
      RECT 73.94 2.282 73.955 3.355 ;
      RECT 73.925 2.255 73.94 3.355 ;
      RECT 73.85 2.25 73.855 2.605 ;
      RECT 73.85 2.66 73.855 3.355 ;
      RECT 73.835 2.25 73.85 2.583 ;
      RECT 73.845 2.682 73.85 3.355 ;
      RECT 73.835 2.722 73.845 3.355 ;
      RECT 73.8 2.25 73.835 2.525 ;
      RECT 73.83 2.757 73.835 3.355 ;
      RECT 73.815 2.812 73.83 3.355 ;
      RECT 73.81 2.877 73.815 3.355 ;
      RECT 73.795 2.925 73.81 3.355 ;
      RECT 73.77 2.25 73.8 2.48 ;
      RECT 73.79 2.98 73.795 3.355 ;
      RECT 73.775 3.04 73.79 3.355 ;
      RECT 73.77 3.088 73.775 3.353 ;
      RECT 73.765 2.25 73.77 2.473 ;
      RECT 73.765 3.12 73.77 3.348 ;
      RECT 73.74 2.25 73.765 2.465 ;
      RECT 73.73 2.255 73.74 2.455 ;
      RECT 73.945 3.53 73.965 3.77 ;
      RECT 73.175 3.46 73.18 3.67 ;
      RECT 74.455 3.533 74.465 3.728 ;
      RECT 74.45 3.523 74.455 3.731 ;
      RECT 74.37 3.52 74.45 3.754 ;
      RECT 74.366 3.52 74.37 3.776 ;
      RECT 74.28 3.52 74.366 3.786 ;
      RECT 74.265 3.52 74.28 3.794 ;
      RECT 74.236 3.521 74.265 3.792 ;
      RECT 74.15 3.526 74.236 3.788 ;
      RECT 74.137 3.53 74.15 3.784 ;
      RECT 74.051 3.53 74.137 3.78 ;
      RECT 73.965 3.53 74.051 3.774 ;
      RECT 73.881 3.53 73.945 3.768 ;
      RECT 73.795 3.53 73.881 3.763 ;
      RECT 73.775 3.53 73.795 3.759 ;
      RECT 73.715 3.525 73.775 3.756 ;
      RECT 73.687 3.519 73.715 3.753 ;
      RECT 73.601 3.514 73.687 3.749 ;
      RECT 73.515 3.508 73.601 3.743 ;
      RECT 73.44 3.49 73.515 3.738 ;
      RECT 73.405 3.467 73.44 3.734 ;
      RECT 73.395 3.457 73.405 3.733 ;
      RECT 73.34 3.455 73.395 3.732 ;
      RECT 73.265 3.455 73.34 3.728 ;
      RECT 73.255 3.455 73.265 3.723 ;
      RECT 73.24 3.455 73.255 3.715 ;
      RECT 73.19 3.457 73.24 3.693 ;
      RECT 73.18 3.46 73.19 3.673 ;
      RECT 73.17 3.465 73.175 3.668 ;
      RECT 73.165 3.47 73.17 3.663 ;
      RECT 73.29 2.635 73.55 2.895 ;
      RECT 73.29 2.65 73.57 2.86 ;
      RECT 73.29 2.655 73.58 2.855 ;
      RECT 71.275 2.115 71.535 2.375 ;
      RECT 71.265 2.145 71.535 2.355 ;
      RECT 73.185 2.06 73.445 2.32 ;
      RECT 73.18 2.135 73.185 2.321 ;
      RECT 73.155 2.14 73.18 2.323 ;
      RECT 73.14 2.147 73.155 2.326 ;
      RECT 73.08 2.165 73.14 2.331 ;
      RECT 73.05 2.185 73.08 2.338 ;
      RECT 73.025 2.193 73.05 2.343 ;
      RECT 73 2.201 73.025 2.345 ;
      RECT 72.982 2.205 73 2.344 ;
      RECT 72.896 2.203 72.982 2.344 ;
      RECT 72.81 2.201 72.896 2.344 ;
      RECT 72.724 2.199 72.81 2.343 ;
      RECT 72.638 2.197 72.724 2.343 ;
      RECT 72.552 2.195 72.638 2.343 ;
      RECT 72.466 2.193 72.552 2.343 ;
      RECT 72.38 2.191 72.466 2.342 ;
      RECT 72.362 2.19 72.38 2.342 ;
      RECT 72.276 2.189 72.362 2.342 ;
      RECT 72.19 2.187 72.276 2.342 ;
      RECT 72.104 2.186 72.19 2.341 ;
      RECT 72.018 2.185 72.104 2.341 ;
      RECT 71.932 2.183 72.018 2.341 ;
      RECT 71.846 2.182 71.932 2.341 ;
      RECT 71.76 2.18 71.846 2.34 ;
      RECT 71.736 2.178 71.76 2.34 ;
      RECT 71.65 2.171 71.736 2.34 ;
      RECT 71.621 2.163 71.65 2.34 ;
      RECT 71.535 2.155 71.621 2.34 ;
      RECT 71.255 2.152 71.265 2.35 ;
      RECT 72.76 3.115 72.765 3.465 ;
      RECT 72.53 3.205 72.67 3.465 ;
      RECT 73.005 2.89 73.05 3.1 ;
      RECT 73.06 2.901 73.07 3.095 ;
      RECT 73.05 2.893 73.06 3.1 ;
      RECT 72.985 2.89 73.005 3.105 ;
      RECT 72.955 2.89 72.985 3.128 ;
      RECT 72.945 2.89 72.955 3.153 ;
      RECT 72.94 2.89 72.945 3.163 ;
      RECT 72.885 2.89 72.94 3.203 ;
      RECT 72.88 2.89 72.885 3.243 ;
      RECT 72.875 2.892 72.88 3.248 ;
      RECT 72.86 2.902 72.875 3.259 ;
      RECT 72.815 2.96 72.86 3.295 ;
      RECT 72.805 3.015 72.815 3.329 ;
      RECT 72.79 3.042 72.805 3.345 ;
      RECT 72.78 3.069 72.79 3.465 ;
      RECT 72.765 3.092 72.78 3.465 ;
      RECT 72.755 3.132 72.76 3.465 ;
      RECT 72.75 3.142 72.755 3.465 ;
      RECT 72.745 3.157 72.75 3.465 ;
      RECT 72.735 3.162 72.745 3.465 ;
      RECT 72.67 3.185 72.735 3.465 ;
      RECT 72.17 2.68 72.36 2.89 ;
      RECT 70.745 2.605 71.005 2.865 ;
      RECT 71.095 2.6 71.19 2.81 ;
      RECT 71.07 2.615 71.08 2.81 ;
      RECT 72.36 2.687 72.37 2.885 ;
      RECT 72.16 2.687 72.17 2.885 ;
      RECT 72.145 2.702 72.16 2.875 ;
      RECT 72.14 2.71 72.145 2.868 ;
      RECT 72.13 2.713 72.14 2.865 ;
      RECT 72.095 2.712 72.13 2.863 ;
      RECT 72.066 2.708 72.095 2.86 ;
      RECT 71.98 2.703 72.066 2.857 ;
      RECT 71.92 2.697 71.98 2.853 ;
      RECT 71.891 2.693 71.92 2.85 ;
      RECT 71.805 2.685 71.891 2.847 ;
      RECT 71.796 2.679 71.805 2.845 ;
      RECT 71.71 2.674 71.796 2.843 ;
      RECT 71.687 2.669 71.71 2.84 ;
      RECT 71.601 2.663 71.687 2.837 ;
      RECT 71.515 2.654 71.601 2.832 ;
      RECT 71.505 2.649 71.515 2.83 ;
      RECT 71.486 2.648 71.505 2.829 ;
      RECT 71.4 2.643 71.486 2.825 ;
      RECT 71.38 2.638 71.4 2.821 ;
      RECT 71.32 2.633 71.38 2.818 ;
      RECT 71.295 2.623 71.32 2.816 ;
      RECT 71.29 2.616 71.295 2.815 ;
      RECT 71.28 2.607 71.29 2.814 ;
      RECT 71.276 2.6 71.28 2.814 ;
      RECT 71.19 2.6 71.276 2.812 ;
      RECT 71.08 2.607 71.095 2.81 ;
      RECT 71.065 2.617 71.07 2.81 ;
      RECT 71.045 2.62 71.065 2.807 ;
      RECT 71.015 2.62 71.045 2.803 ;
      RECT 71.005 2.62 71.015 2.803 ;
      RECT 71.92 3.115 72.18 3.375 ;
      RECT 71.85 3.125 72.18 3.335 ;
      RECT 71.84 3.132 72.18 3.33 ;
      RECT 71.26 3.12 71.52 3.38 ;
      RECT 71.26 3.16 71.625 3.37 ;
      RECT 71.26 3.162 71.63 3.369 ;
      RECT 71.26 3.17 71.635 3.366 ;
      RECT 70.185 2.245 70.285 3.77 ;
      RECT 70.375 3.385 70.425 3.645 ;
      RECT 70.37 2.258 70.375 2.445 ;
      RECT 70.365 3.366 70.375 3.645 ;
      RECT 70.365 2.255 70.37 2.453 ;
      RECT 70.35 2.249 70.365 2.46 ;
      RECT 70.36 3.354 70.365 3.728 ;
      RECT 70.35 3.342 70.36 3.765 ;
      RECT 70.34 2.245 70.35 2.467 ;
      RECT 70.34 3.327 70.35 3.77 ;
      RECT 70.335 2.245 70.34 2.475 ;
      RECT 70.315 3.297 70.34 3.77 ;
      RECT 70.295 2.245 70.335 2.523 ;
      RECT 70.305 3.257 70.315 3.77 ;
      RECT 70.295 3.212 70.305 3.77 ;
      RECT 70.29 2.245 70.295 2.593 ;
      RECT 70.29 3.17 70.295 3.77 ;
      RECT 70.285 2.245 70.29 3.07 ;
      RECT 70.285 3.152 70.29 3.77 ;
      RECT 70.175 2.248 70.185 3.77 ;
      RECT 70.16 2.255 70.175 3.766 ;
      RECT 70.155 2.265 70.16 3.761 ;
      RECT 70.15 2.465 70.155 3.653 ;
      RECT 70.145 2.55 70.15 3.205 ;
      RECT 69.025 7.765 69.315 7.995 ;
      RECT 69.085 6.285 69.255 7.995 ;
      RECT 69.03 6.655 69.38 7.005 ;
      RECT 69.025 6.285 69.315 6.515 ;
      RECT 69.025 2.365 69.315 2.595 ;
      RECT 69.085 0.885 69.255 2.595 ;
      RECT 69.025 0.885 69.315 1.115 ;
      RECT 68.615 2.735 68.945 2.965 ;
      RECT 68.615 2.765 69.115 2.935 ;
      RECT 68.615 2.395 68.805 2.965 ;
      RECT 68.035 2.365 68.325 2.595 ;
      RECT 68.035 2.395 68.805 2.565 ;
      RECT 68.095 0.885 68.265 2.595 ;
      RECT 68.035 0.885 68.325 1.115 ;
      RECT 68.035 7.765 68.325 7.995 ;
      RECT 68.095 6.285 68.265 7.995 ;
      RECT 68.035 6.285 68.325 6.515 ;
      RECT 68.035 6.325 68.885 6.485 ;
      RECT 68.715 5.915 68.885 6.485 ;
      RECT 68.035 6.32 68.425 6.485 ;
      RECT 68.655 5.915 68.945 6.145 ;
      RECT 68.655 5.945 69.115 6.115 ;
      RECT 67.665 2.735 67.955 2.965 ;
      RECT 67.665 2.765 68.125 2.935 ;
      RECT 67.725 1.655 67.89 2.965 ;
      RECT 66.24 1.625 66.53 1.855 ;
      RECT 66.24 1.655 67.89 1.825 ;
      RECT 66.3 0.885 66.47 1.855 ;
      RECT 66.24 0.885 66.53 1.115 ;
      RECT 66.24 7.765 66.53 7.995 ;
      RECT 66.3 7.025 66.47 7.995 ;
      RECT 66.3 7.12 67.89 7.29 ;
      RECT 67.72 5.915 67.89 7.29 ;
      RECT 66.24 7.025 66.53 7.255 ;
      RECT 67.665 5.915 67.955 6.145 ;
      RECT 67.665 5.945 68.125 6.115 ;
      RECT 64.275 3.43 64.625 3.78 ;
      RECT 64.365 2.025 64.535 3.78 ;
      RECT 66.67 1.965 67.02 2.315 ;
      RECT 64.365 2.025 65.985 2.2 ;
      RECT 64.365 2.025 67.02 2.195 ;
      RECT 66.695 6.655 67.02 6.98 ;
      RECT 62.07 6.61 62.42 6.96 ;
      RECT 66.67 6.655 67.02 6.885 ;
      RECT 61.91 6.655 62.42 6.885 ;
      RECT 61.74 6.685 67.02 6.855 ;
      RECT 65.895 2.365 66.215 2.685 ;
      RECT 65.865 2.365 66.215 2.595 ;
      RECT 65.695 2.395 66.215 2.565 ;
      RECT 65.895 6.225 66.215 6.545 ;
      RECT 65.865 6.285 66.215 6.515 ;
      RECT 65.695 6.315 66.215 6.485 ;
      RECT 64.85 2.705 65.2 3.055 ;
      RECT 64.85 2.765 65.33 2.935 ;
      RECT 64.84 5.84 65.19 6.19 ;
      RECT 60.11 5.915 60.4 6.145 ;
      RECT 60.11 5.945 65.33 6.115 ;
      RECT 61.675 3.665 61.715 3.925 ;
      RECT 61.715 3.645 61.72 3.655 ;
      RECT 63.045 2.89 63.055 3.111 ;
      RECT 62.975 2.885 63.045 3.236 ;
      RECT 62.965 2.885 62.975 3.363 ;
      RECT 62.94 2.885 62.965 3.41 ;
      RECT 62.915 2.885 62.94 3.488 ;
      RECT 62.895 2.885 62.915 3.558 ;
      RECT 62.87 2.885 62.895 3.598 ;
      RECT 62.86 2.885 62.87 3.618 ;
      RECT 62.85 2.887 62.86 3.626 ;
      RECT 62.845 2.892 62.85 3.083 ;
      RECT 62.845 3.092 62.85 3.627 ;
      RECT 62.84 3.137 62.845 3.628 ;
      RECT 62.83 3.202 62.84 3.629 ;
      RECT 62.82 3.297 62.83 3.631 ;
      RECT 62.815 3.35 62.82 3.633 ;
      RECT 62.81 3.37 62.815 3.634 ;
      RECT 62.755 3.395 62.81 3.64 ;
      RECT 62.715 3.43 62.755 3.649 ;
      RECT 62.705 3.447 62.715 3.654 ;
      RECT 62.696 3.453 62.705 3.656 ;
      RECT 62.61 3.491 62.696 3.667 ;
      RECT 62.605 3.53 62.61 3.677 ;
      RECT 62.53 3.537 62.605 3.687 ;
      RECT 62.51 3.547 62.53 3.698 ;
      RECT 62.48 3.554 62.51 3.706 ;
      RECT 62.455 3.561 62.48 3.713 ;
      RECT 62.431 3.567 62.455 3.718 ;
      RECT 62.345 3.58 62.431 3.73 ;
      RECT 62.267 3.587 62.345 3.748 ;
      RECT 62.181 3.582 62.267 3.766 ;
      RECT 62.095 3.577 62.181 3.786 ;
      RECT 62.015 3.571 62.095 3.803 ;
      RECT 61.95 3.567 62.015 3.832 ;
      RECT 61.945 3.281 61.95 3.305 ;
      RECT 61.935 3.557 61.95 3.86 ;
      RECT 61.94 3.275 61.945 3.345 ;
      RECT 61.935 3.269 61.94 3.415 ;
      RECT 61.93 3.263 61.935 3.493 ;
      RECT 61.93 3.54 61.935 3.925 ;
      RECT 61.922 3.26 61.93 3.925 ;
      RECT 61.836 3.258 61.922 3.925 ;
      RECT 61.75 3.256 61.836 3.925 ;
      RECT 61.74 3.257 61.75 3.925 ;
      RECT 61.735 3.262 61.74 3.925 ;
      RECT 61.725 3.275 61.735 3.925 ;
      RECT 61.72 3.297 61.725 3.925 ;
      RECT 61.715 3.657 61.72 3.925 ;
      RECT 62.345 3.125 62.35 3.345 ;
      RECT 62.85 2.16 62.885 2.42 ;
      RECT 62.835 2.16 62.85 2.428 ;
      RECT 62.806 2.16 62.835 2.45 ;
      RECT 62.72 2.16 62.806 2.51 ;
      RECT 62.7 2.16 62.72 2.575 ;
      RECT 62.64 2.16 62.7 2.74 ;
      RECT 62.635 2.16 62.64 2.888 ;
      RECT 62.63 2.16 62.635 2.9 ;
      RECT 62.625 2.16 62.63 2.926 ;
      RECT 62.595 2.346 62.625 3.006 ;
      RECT 62.59 2.394 62.595 3.095 ;
      RECT 62.585 2.408 62.59 3.11 ;
      RECT 62.58 2.427 62.585 3.14 ;
      RECT 62.575 2.442 62.58 3.156 ;
      RECT 62.57 2.457 62.575 3.178 ;
      RECT 62.565 2.477 62.57 3.2 ;
      RECT 62.555 2.497 62.565 3.233 ;
      RECT 62.54 2.539 62.555 3.295 ;
      RECT 62.535 2.57 62.54 3.335 ;
      RECT 62.53 2.582 62.535 3.34 ;
      RECT 62.525 2.594 62.53 3.345 ;
      RECT 62.52 2.607 62.525 3.345 ;
      RECT 62.515 2.625 62.52 3.345 ;
      RECT 62.51 2.645 62.515 3.345 ;
      RECT 62.505 2.657 62.51 3.345 ;
      RECT 62.5 2.67 62.505 3.345 ;
      RECT 62.48 2.705 62.5 3.345 ;
      RECT 62.43 2.807 62.48 3.345 ;
      RECT 62.425 2.892 62.43 3.345 ;
      RECT 62.42 2.9 62.425 3.345 ;
      RECT 62.415 2.917 62.42 3.345 ;
      RECT 62.41 2.932 62.415 3.345 ;
      RECT 62.375 2.997 62.41 3.345 ;
      RECT 62.36 3.062 62.375 3.345 ;
      RECT 62.355 3.092 62.36 3.345 ;
      RECT 62.35 3.117 62.355 3.345 ;
      RECT 62.335 3.127 62.345 3.345 ;
      RECT 62.32 3.14 62.335 3.338 ;
      RECT 62.065 2.73 62.135 2.94 ;
      RECT 61.855 2.707 61.86 2.9 ;
      RECT 59.31 2.635 59.57 2.895 ;
      RECT 62.145 2.917 62.15 2.92 ;
      RECT 62.135 2.735 62.145 2.935 ;
      RECT 62.036 2.728 62.065 2.94 ;
      RECT 61.95 2.72 62.036 2.94 ;
      RECT 61.935 2.714 61.95 2.938 ;
      RECT 61.915 2.713 61.935 2.925 ;
      RECT 61.91 2.712 61.915 2.908 ;
      RECT 61.86 2.709 61.91 2.903 ;
      RECT 61.83 2.706 61.855 2.898 ;
      RECT 61.81 2.704 61.83 2.893 ;
      RECT 61.795 2.702 61.81 2.89 ;
      RECT 61.765 2.7 61.795 2.888 ;
      RECT 61.7 2.696 61.765 2.88 ;
      RECT 61.67 2.691 61.7 2.875 ;
      RECT 61.65 2.689 61.67 2.873 ;
      RECT 61.62 2.686 61.65 2.868 ;
      RECT 61.56 2.682 61.62 2.86 ;
      RECT 61.555 2.679 61.56 2.855 ;
      RECT 61.485 2.677 61.555 2.85 ;
      RECT 61.456 2.673 61.485 2.843 ;
      RECT 61.37 2.668 61.456 2.835 ;
      RECT 61.336 2.663 61.37 2.827 ;
      RECT 61.25 2.655 61.336 2.819 ;
      RECT 61.211 2.648 61.25 2.811 ;
      RECT 61.125 2.643 61.211 2.803 ;
      RECT 61.06 2.637 61.125 2.793 ;
      RECT 61.04 2.632 61.06 2.788 ;
      RECT 61.031 2.629 61.04 2.787 ;
      RECT 60.945 2.625 61.031 2.781 ;
      RECT 60.905 2.621 60.945 2.773 ;
      RECT 60.885 2.617 60.905 2.771 ;
      RECT 60.825 2.617 60.885 2.768 ;
      RECT 60.805 2.62 60.825 2.766 ;
      RECT 60.784 2.62 60.805 2.766 ;
      RECT 60.698 2.622 60.784 2.77 ;
      RECT 60.612 2.624 60.698 2.776 ;
      RECT 60.526 2.626 60.612 2.783 ;
      RECT 60.44 2.629 60.526 2.789 ;
      RECT 60.406 2.63 60.44 2.794 ;
      RECT 60.32 2.633 60.406 2.799 ;
      RECT 60.291 2.64 60.32 2.804 ;
      RECT 60.205 2.64 60.291 2.809 ;
      RECT 60.172 2.64 60.205 2.814 ;
      RECT 60.086 2.642 60.172 2.819 ;
      RECT 60 2.644 60.086 2.826 ;
      RECT 59.936 2.646 60 2.832 ;
      RECT 59.85 2.648 59.936 2.838 ;
      RECT 59.847 2.65 59.85 2.841 ;
      RECT 59.761 2.651 59.847 2.845 ;
      RECT 59.675 2.654 59.761 2.852 ;
      RECT 59.656 2.656 59.675 2.856 ;
      RECT 59.57 2.658 59.656 2.861 ;
      RECT 59.3 2.67 59.31 2.865 ;
      RECT 61.48 7.765 61.77 7.995 ;
      RECT 61.54 7.025 61.71 7.995 ;
      RECT 61.43 7.055 61.805 7.425 ;
      RECT 61.48 7.025 61.77 7.425 ;
      RECT 61.535 2.25 61.72 2.46 ;
      RECT 61.53 2.251 61.725 2.458 ;
      RECT 61.525 2.256 61.735 2.453 ;
      RECT 61.52 2.232 61.525 2.45 ;
      RECT 61.49 2.229 61.52 2.443 ;
      RECT 61.485 2.225 61.49 2.434 ;
      RECT 61.45 2.256 61.735 2.429 ;
      RECT 61.225 2.165 61.485 2.425 ;
      RECT 61.525 2.234 61.53 2.453 ;
      RECT 61.53 2.235 61.535 2.458 ;
      RECT 61.225 2.247 61.605 2.425 ;
      RECT 61.225 2.245 61.59 2.425 ;
      RECT 61.225 2.24 61.58 2.425 ;
      RECT 61.18 3.155 61.23 3.44 ;
      RECT 61.125 3.125 61.13 3.44 ;
      RECT 61.095 3.105 61.1 3.44 ;
      RECT 61.245 3.155 61.305 3.415 ;
      RECT 61.24 3.155 61.245 3.423 ;
      RECT 61.23 3.155 61.24 3.435 ;
      RECT 61.145 3.145 61.18 3.44 ;
      RECT 61.14 3.132 61.145 3.44 ;
      RECT 61.13 3.127 61.14 3.44 ;
      RECT 61.11 3.117 61.125 3.44 ;
      RECT 61.1 3.11 61.11 3.44 ;
      RECT 61.09 3.102 61.095 3.44 ;
      RECT 61.06 3.092 61.09 3.44 ;
      RECT 61.045 3.08 61.06 3.44 ;
      RECT 61.03 3.07 61.045 3.435 ;
      RECT 61.01 3.06 61.03 3.41 ;
      RECT 61 3.052 61.01 3.387 ;
      RECT 60.97 3.035 61 3.377 ;
      RECT 60.965 3.012 60.97 3.368 ;
      RECT 60.96 2.999 60.965 3.366 ;
      RECT 60.945 2.975 60.96 3.36 ;
      RECT 60.94 2.951 60.945 3.354 ;
      RECT 60.93 2.94 60.94 3.349 ;
      RECT 60.925 2.93 60.93 3.345 ;
      RECT 60.92 2.922 60.925 3.342 ;
      RECT 60.91 2.917 60.92 3.338 ;
      RECT 60.905 2.912 60.91 3.334 ;
      RECT 60.82 2.91 60.905 3.309 ;
      RECT 60.79 2.91 60.82 3.275 ;
      RECT 60.775 2.91 60.79 3.258 ;
      RECT 60.72 2.91 60.775 3.203 ;
      RECT 60.715 2.915 60.72 3.152 ;
      RECT 60.705 2.92 60.715 3.142 ;
      RECT 60.7 2.93 60.705 3.128 ;
      RECT 60.65 3.67 60.91 3.93 ;
      RECT 60.57 3.685 60.91 3.906 ;
      RECT 60.55 3.685 60.91 3.901 ;
      RECT 60.526 3.685 60.91 3.899 ;
      RECT 60.44 3.685 60.91 3.894 ;
      RECT 60.29 3.625 60.55 3.89 ;
      RECT 60.245 3.685 60.91 3.885 ;
      RECT 60.24 3.692 60.91 3.88 ;
      RECT 60.255 3.68 60.57 3.89 ;
      RECT 60.145 2.115 60.405 2.375 ;
      RECT 60.145 2.172 60.41 2.368 ;
      RECT 60.145 2.202 60.415 2.3 ;
      RECT 60.205 2.633 60.32 2.635 ;
      RECT 60.291 2.63 60.32 2.635 ;
      RECT 59.315 3.634 59.34 3.874 ;
      RECT 59.3 3.637 59.39 3.868 ;
      RECT 59.295 3.642 59.476 3.863 ;
      RECT 59.29 3.65 59.54 3.861 ;
      RECT 59.29 3.65 59.55 3.86 ;
      RECT 59.285 3.657 59.56 3.853 ;
      RECT 59.285 3.657 59.646 3.842 ;
      RECT 59.28 3.692 59.646 3.838 ;
      RECT 59.28 3.692 59.655 3.827 ;
      RECT 59.56 3.565 59.82 3.825 ;
      RECT 59.27 3.742 59.82 3.823 ;
      RECT 59.54 3.61 59.56 3.858 ;
      RECT 59.476 3.613 59.54 3.862 ;
      RECT 59.39 3.618 59.476 3.867 ;
      RECT 59.32 3.629 59.82 3.825 ;
      RECT 59.34 3.623 59.39 3.872 ;
      RECT 59.465 2.1 59.475 2.362 ;
      RECT 59.455 2.157 59.465 2.365 ;
      RECT 59.43 2.162 59.455 2.371 ;
      RECT 59.405 2.166 59.43 2.383 ;
      RECT 59.395 2.169 59.405 2.393 ;
      RECT 59.39 2.17 59.395 2.398 ;
      RECT 59.385 2.171 59.39 2.403 ;
      RECT 59.38 2.172 59.385 2.405 ;
      RECT 59.355 2.175 59.38 2.408 ;
      RECT 59.325 2.181 59.355 2.411 ;
      RECT 59.26 2.192 59.325 2.414 ;
      RECT 59.215 2.2 59.26 2.418 ;
      RECT 59.2 2.2 59.215 2.426 ;
      RECT 59.195 2.201 59.2 2.433 ;
      RECT 59.19 2.203 59.195 2.436 ;
      RECT 59.185 2.207 59.19 2.439 ;
      RECT 59.175 2.215 59.185 2.443 ;
      RECT 59.17 2.228 59.175 2.448 ;
      RECT 59.165 2.236 59.17 2.45 ;
      RECT 59.16 2.242 59.165 2.45 ;
      RECT 59.155 2.246 59.16 2.453 ;
      RECT 59.15 2.248 59.155 2.456 ;
      RECT 59.145 2.251 59.15 2.459 ;
      RECT 59.135 2.256 59.145 2.463 ;
      RECT 59.13 2.262 59.135 2.468 ;
      RECT 59.12 2.268 59.13 2.472 ;
      RECT 59.105 2.275 59.12 2.478 ;
      RECT 59.076 2.289 59.105 2.488 ;
      RECT 58.99 2.324 59.076 2.52 ;
      RECT 58.97 2.357 58.99 2.549 ;
      RECT 58.95 2.37 58.97 2.56 ;
      RECT 58.93 2.382 58.95 2.571 ;
      RECT 58.88 2.404 58.93 2.591 ;
      RECT 58.865 2.422 58.88 2.608 ;
      RECT 58.86 2.428 58.865 2.611 ;
      RECT 58.855 2.432 58.86 2.614 ;
      RECT 58.85 2.436 58.855 2.618 ;
      RECT 58.845 2.438 58.85 2.621 ;
      RECT 58.835 2.445 58.845 2.624 ;
      RECT 58.83 2.45 58.835 2.628 ;
      RECT 58.825 2.452 58.83 2.631 ;
      RECT 58.82 2.456 58.825 2.634 ;
      RECT 58.815 2.458 58.82 2.638 ;
      RECT 58.8 2.463 58.815 2.643 ;
      RECT 58.795 2.468 58.8 2.646 ;
      RECT 58.79 2.476 58.795 2.649 ;
      RECT 58.785 2.478 58.79 2.652 ;
      RECT 58.78 2.48 58.785 2.655 ;
      RECT 58.77 2.482 58.78 2.661 ;
      RECT 58.735 2.496 58.77 2.673 ;
      RECT 58.725 2.511 58.735 2.683 ;
      RECT 58.65 2.54 58.725 2.707 ;
      RECT 58.645 2.565 58.65 2.73 ;
      RECT 58.63 2.569 58.645 2.736 ;
      RECT 58.62 2.577 58.63 2.741 ;
      RECT 58.59 2.59 58.62 2.745 ;
      RECT 58.58 2.605 58.59 2.75 ;
      RECT 58.57 2.61 58.58 2.753 ;
      RECT 58.565 2.612 58.57 2.755 ;
      RECT 58.55 2.615 58.565 2.758 ;
      RECT 58.545 2.617 58.55 2.761 ;
      RECT 58.525 2.622 58.545 2.765 ;
      RECT 58.495 2.627 58.525 2.773 ;
      RECT 58.47 2.634 58.495 2.781 ;
      RECT 58.465 2.639 58.47 2.786 ;
      RECT 58.435 2.642 58.465 2.79 ;
      RECT 58.395 2.645 58.435 2.8 ;
      RECT 58.36 2.642 58.395 2.812 ;
      RECT 58.35 2.638 58.36 2.819 ;
      RECT 58.325 2.634 58.35 2.825 ;
      RECT 58.32 2.63 58.325 2.83 ;
      RECT 58.28 2.627 58.32 2.83 ;
      RECT 58.265 2.612 58.28 2.831 ;
      RECT 58.242 2.6 58.265 2.831 ;
      RECT 58.156 2.6 58.242 2.832 ;
      RECT 58.07 2.6 58.156 2.834 ;
      RECT 58.05 2.6 58.07 2.831 ;
      RECT 58.045 2.605 58.05 2.826 ;
      RECT 58.04 2.61 58.045 2.824 ;
      RECT 58.03 2.62 58.04 2.822 ;
      RECT 58.025 2.626 58.03 2.815 ;
      RECT 58.02 2.628 58.025 2.8 ;
      RECT 58.015 2.632 58.02 2.79 ;
      RECT 59.475 2.1 59.725 2.36 ;
      RECT 57.2 3.635 57.46 3.895 ;
      RECT 59.495 3.125 59.5 3.335 ;
      RECT 59.5 3.13 59.51 3.33 ;
      RECT 59.45 3.125 59.495 3.35 ;
      RECT 59.44 3.125 59.45 3.37 ;
      RECT 59.421 3.125 59.44 3.375 ;
      RECT 59.335 3.125 59.421 3.372 ;
      RECT 59.305 3.127 59.335 3.37 ;
      RECT 59.25 3.137 59.305 3.368 ;
      RECT 59.185 3.151 59.25 3.366 ;
      RECT 59.18 3.159 59.185 3.365 ;
      RECT 59.165 3.162 59.18 3.363 ;
      RECT 59.1 3.172 59.165 3.359 ;
      RECT 59.052 3.186 59.1 3.36 ;
      RECT 58.966 3.203 59.052 3.374 ;
      RECT 58.88 3.224 58.966 3.391 ;
      RECT 58.86 3.237 58.88 3.401 ;
      RECT 58.815 3.245 58.86 3.408 ;
      RECT 58.78 3.253 58.815 3.416 ;
      RECT 58.746 3.261 58.78 3.424 ;
      RECT 58.66 3.275 58.746 3.436 ;
      RECT 58.625 3.292 58.66 3.448 ;
      RECT 58.616 3.301 58.625 3.452 ;
      RECT 58.53 3.319 58.616 3.469 ;
      RECT 58.471 3.346 58.53 3.496 ;
      RECT 58.385 3.373 58.471 3.524 ;
      RECT 58.365 3.395 58.385 3.544 ;
      RECT 58.305 3.41 58.365 3.56 ;
      RECT 58.295 3.422 58.305 3.573 ;
      RECT 58.29 3.427 58.295 3.576 ;
      RECT 58.28 3.43 58.29 3.579 ;
      RECT 58.275 3.432 58.28 3.582 ;
      RECT 58.245 3.44 58.275 3.589 ;
      RECT 58.23 3.447 58.245 3.597 ;
      RECT 58.22 3.452 58.23 3.601 ;
      RECT 58.215 3.455 58.22 3.604 ;
      RECT 58.205 3.457 58.215 3.607 ;
      RECT 58.17 3.467 58.205 3.616 ;
      RECT 58.095 3.49 58.17 3.638 ;
      RECT 58.075 3.508 58.095 3.656 ;
      RECT 58.045 3.515 58.075 3.666 ;
      RECT 58.025 3.523 58.045 3.676 ;
      RECT 58.015 3.529 58.025 3.683 ;
      RECT 57.996 3.534 58.015 3.689 ;
      RECT 57.91 3.554 57.996 3.709 ;
      RECT 57.895 3.574 57.91 3.728 ;
      RECT 57.85 3.586 57.895 3.739 ;
      RECT 57.785 3.607 57.85 3.762 ;
      RECT 57.745 3.627 57.785 3.783 ;
      RECT 57.735 3.637 57.745 3.793 ;
      RECT 57.685 3.649 57.735 3.804 ;
      RECT 57.665 3.665 57.685 3.816 ;
      RECT 57.635 3.675 57.665 3.822 ;
      RECT 57.625 3.68 57.635 3.824 ;
      RECT 57.556 3.681 57.625 3.83 ;
      RECT 57.47 3.683 57.556 3.84 ;
      RECT 57.46 3.684 57.47 3.845 ;
      RECT 58.73 3.71 58.92 3.92 ;
      RECT 58.72 3.715 58.93 3.913 ;
      RECT 58.705 3.715 58.93 3.878 ;
      RECT 58.625 3.6 58.885 3.86 ;
      RECT 57.54 3.13 57.725 3.425 ;
      RECT 57.53 3.13 57.725 3.423 ;
      RECT 57.515 3.13 57.73 3.418 ;
      RECT 57.515 3.13 57.735 3.415 ;
      RECT 57.51 3.13 57.735 3.413 ;
      RECT 57.505 3.385 57.735 3.403 ;
      RECT 57.51 3.13 57.77 3.39 ;
      RECT 57.47 2.165 57.73 2.425 ;
      RECT 57.28 2.09 57.366 2.423 ;
      RECT 57.255 2.094 57.41 2.419 ;
      RECT 57.366 2.086 57.41 2.419 ;
      RECT 57.366 2.087 57.415 2.418 ;
      RECT 57.28 2.092 57.43 2.417 ;
      RECT 57.255 2.1 57.47 2.416 ;
      RECT 57.25 2.095 57.43 2.411 ;
      RECT 57.24 2.11 57.47 2.318 ;
      RECT 57.24 2.162 57.67 2.318 ;
      RECT 57.24 2.155 57.65 2.318 ;
      RECT 57.24 2.142 57.62 2.318 ;
      RECT 57.24 2.13 57.56 2.318 ;
      RECT 57.24 2.115 57.535 2.318 ;
      RECT 56.44 2.745 56.575 3.04 ;
      RECT 56.7 2.768 56.705 2.955 ;
      RECT 57.42 2.665 57.565 2.9 ;
      RECT 57.58 2.665 57.585 2.89 ;
      RECT 57.615 2.676 57.62 2.87 ;
      RECT 57.61 2.668 57.615 2.875 ;
      RECT 57.59 2.665 57.61 2.88 ;
      RECT 57.585 2.665 57.59 2.888 ;
      RECT 57.575 2.665 57.58 2.893 ;
      RECT 57.565 2.665 57.575 2.898 ;
      RECT 57.395 2.667 57.42 2.9 ;
      RECT 57.345 2.674 57.395 2.9 ;
      RECT 57.34 2.679 57.345 2.9 ;
      RECT 57.301 2.684 57.34 2.901 ;
      RECT 57.215 2.696 57.301 2.902 ;
      RECT 57.206 2.706 57.215 2.902 ;
      RECT 57.12 2.715 57.206 2.904 ;
      RECT 57.096 2.725 57.12 2.906 ;
      RECT 57.01 2.736 57.096 2.907 ;
      RECT 56.98 2.747 57.01 2.909 ;
      RECT 56.95 2.752 56.98 2.911 ;
      RECT 56.925 2.758 56.95 2.914 ;
      RECT 56.91 2.763 56.925 2.915 ;
      RECT 56.865 2.769 56.91 2.915 ;
      RECT 56.86 2.774 56.865 2.916 ;
      RECT 56.84 2.774 56.86 2.918 ;
      RECT 56.82 2.772 56.84 2.923 ;
      RECT 56.785 2.771 56.82 2.93 ;
      RECT 56.755 2.77 56.785 2.94 ;
      RECT 56.705 2.769 56.755 2.95 ;
      RECT 56.615 2.766 56.7 3.04 ;
      RECT 56.59 2.76 56.615 3.04 ;
      RECT 56.575 2.75 56.59 3.04 ;
      RECT 56.39 2.745 56.44 2.96 ;
      RECT 56.38 2.75 56.39 2.95 ;
      RECT 56.62 3.225 56.88 3.485 ;
      RECT 56.62 3.225 56.91 3.378 ;
      RECT 56.62 3.225 56.945 3.363 ;
      RECT 56.875 3.145 57.065 3.355 ;
      RECT 56.865 3.15 57.075 3.348 ;
      RECT 56.83 3.22 57.075 3.348 ;
      RECT 56.86 3.162 56.88 3.485 ;
      RECT 56.845 3.21 57.075 3.348 ;
      RECT 56.85 3.182 56.88 3.485 ;
      RECT 55.93 2.25 56 3.355 ;
      RECT 56.665 2.355 56.925 2.615 ;
      RECT 56.245 2.401 56.26 2.61 ;
      RECT 56.581 2.414 56.665 2.565 ;
      RECT 56.495 2.411 56.581 2.565 ;
      RECT 56.456 2.409 56.495 2.565 ;
      RECT 56.37 2.407 56.456 2.565 ;
      RECT 56.31 2.405 56.37 2.576 ;
      RECT 56.275 2.403 56.31 2.594 ;
      RECT 56.26 2.401 56.275 2.605 ;
      RECT 56.23 2.401 56.245 2.618 ;
      RECT 56.22 2.401 56.23 2.623 ;
      RECT 56.195 2.4 56.22 2.628 ;
      RECT 56.18 2.395 56.195 2.634 ;
      RECT 56.175 2.388 56.18 2.639 ;
      RECT 56.15 2.379 56.175 2.645 ;
      RECT 56.105 2.358 56.15 2.658 ;
      RECT 56.095 2.342 56.105 2.668 ;
      RECT 56.08 2.335 56.095 2.678 ;
      RECT 56.07 2.328 56.08 2.695 ;
      RECT 56.065 2.325 56.07 2.725 ;
      RECT 56.06 2.323 56.065 2.755 ;
      RECT 56.055 2.321 56.06 2.792 ;
      RECT 56.04 2.317 56.055 2.859 ;
      RECT 56.04 3.15 56.05 3.35 ;
      RECT 56.035 2.313 56.04 2.985 ;
      RECT 56.035 3.137 56.04 3.355 ;
      RECT 56.03 2.311 56.035 3.07 ;
      RECT 56.03 3.127 56.035 3.355 ;
      RECT 56.015 2.282 56.03 3.355 ;
      RECT 56 2.255 56.015 3.355 ;
      RECT 55.925 2.25 55.93 2.605 ;
      RECT 55.925 2.66 55.93 3.355 ;
      RECT 55.91 2.25 55.925 2.583 ;
      RECT 55.92 2.682 55.925 3.355 ;
      RECT 55.91 2.722 55.92 3.355 ;
      RECT 55.875 2.25 55.91 2.525 ;
      RECT 55.905 2.757 55.91 3.355 ;
      RECT 55.89 2.812 55.905 3.355 ;
      RECT 55.885 2.877 55.89 3.355 ;
      RECT 55.87 2.925 55.885 3.355 ;
      RECT 55.845 2.25 55.875 2.48 ;
      RECT 55.865 2.98 55.87 3.355 ;
      RECT 55.85 3.04 55.865 3.355 ;
      RECT 55.845 3.088 55.85 3.353 ;
      RECT 55.84 2.25 55.845 2.473 ;
      RECT 55.84 3.12 55.845 3.348 ;
      RECT 55.815 2.25 55.84 2.465 ;
      RECT 55.805 2.255 55.815 2.455 ;
      RECT 56.02 3.53 56.04 3.77 ;
      RECT 55.25 3.46 55.255 3.67 ;
      RECT 56.53 3.533 56.54 3.728 ;
      RECT 56.525 3.523 56.53 3.731 ;
      RECT 56.445 3.52 56.525 3.754 ;
      RECT 56.441 3.52 56.445 3.776 ;
      RECT 56.355 3.52 56.441 3.786 ;
      RECT 56.34 3.52 56.355 3.794 ;
      RECT 56.311 3.521 56.34 3.792 ;
      RECT 56.225 3.526 56.311 3.788 ;
      RECT 56.212 3.53 56.225 3.784 ;
      RECT 56.126 3.53 56.212 3.78 ;
      RECT 56.04 3.53 56.126 3.774 ;
      RECT 55.956 3.53 56.02 3.768 ;
      RECT 55.87 3.53 55.956 3.763 ;
      RECT 55.85 3.53 55.87 3.759 ;
      RECT 55.79 3.525 55.85 3.756 ;
      RECT 55.762 3.519 55.79 3.753 ;
      RECT 55.676 3.514 55.762 3.749 ;
      RECT 55.59 3.508 55.676 3.743 ;
      RECT 55.515 3.49 55.59 3.738 ;
      RECT 55.48 3.467 55.515 3.734 ;
      RECT 55.47 3.457 55.48 3.733 ;
      RECT 55.415 3.455 55.47 3.732 ;
      RECT 55.34 3.455 55.415 3.728 ;
      RECT 55.33 3.455 55.34 3.723 ;
      RECT 55.315 3.455 55.33 3.715 ;
      RECT 55.265 3.457 55.315 3.693 ;
      RECT 55.255 3.46 55.265 3.673 ;
      RECT 55.245 3.465 55.25 3.668 ;
      RECT 55.24 3.47 55.245 3.663 ;
      RECT 55.365 2.635 55.625 2.895 ;
      RECT 55.365 2.65 55.645 2.86 ;
      RECT 55.365 2.655 55.655 2.855 ;
      RECT 53.35 2.115 53.61 2.375 ;
      RECT 53.34 2.145 53.61 2.355 ;
      RECT 55.26 2.06 55.52 2.32 ;
      RECT 55.255 2.135 55.26 2.321 ;
      RECT 55.23 2.14 55.255 2.323 ;
      RECT 55.215 2.147 55.23 2.326 ;
      RECT 55.155 2.165 55.215 2.331 ;
      RECT 55.125 2.185 55.155 2.338 ;
      RECT 55.1 2.193 55.125 2.343 ;
      RECT 55.075 2.201 55.1 2.345 ;
      RECT 55.057 2.205 55.075 2.344 ;
      RECT 54.971 2.203 55.057 2.344 ;
      RECT 54.885 2.201 54.971 2.344 ;
      RECT 54.799 2.199 54.885 2.343 ;
      RECT 54.713 2.197 54.799 2.343 ;
      RECT 54.627 2.195 54.713 2.343 ;
      RECT 54.541 2.193 54.627 2.343 ;
      RECT 54.455 2.191 54.541 2.342 ;
      RECT 54.437 2.19 54.455 2.342 ;
      RECT 54.351 2.189 54.437 2.342 ;
      RECT 54.265 2.187 54.351 2.342 ;
      RECT 54.179 2.186 54.265 2.341 ;
      RECT 54.093 2.185 54.179 2.341 ;
      RECT 54.007 2.183 54.093 2.341 ;
      RECT 53.921 2.182 54.007 2.341 ;
      RECT 53.835 2.18 53.921 2.34 ;
      RECT 53.811 2.178 53.835 2.34 ;
      RECT 53.725 2.171 53.811 2.34 ;
      RECT 53.696 2.163 53.725 2.34 ;
      RECT 53.61 2.155 53.696 2.34 ;
      RECT 53.33 2.152 53.34 2.35 ;
      RECT 54.835 3.115 54.84 3.465 ;
      RECT 54.605 3.205 54.745 3.465 ;
      RECT 55.08 2.89 55.125 3.1 ;
      RECT 55.135 2.901 55.145 3.095 ;
      RECT 55.125 2.893 55.135 3.1 ;
      RECT 55.06 2.89 55.08 3.105 ;
      RECT 55.03 2.89 55.06 3.128 ;
      RECT 55.02 2.89 55.03 3.153 ;
      RECT 55.015 2.89 55.02 3.163 ;
      RECT 54.96 2.89 55.015 3.203 ;
      RECT 54.955 2.89 54.96 3.243 ;
      RECT 54.95 2.892 54.955 3.248 ;
      RECT 54.935 2.902 54.95 3.259 ;
      RECT 54.89 2.96 54.935 3.295 ;
      RECT 54.88 3.015 54.89 3.329 ;
      RECT 54.865 3.042 54.88 3.345 ;
      RECT 54.855 3.069 54.865 3.465 ;
      RECT 54.84 3.092 54.855 3.465 ;
      RECT 54.83 3.132 54.835 3.465 ;
      RECT 54.825 3.142 54.83 3.465 ;
      RECT 54.82 3.157 54.825 3.465 ;
      RECT 54.81 3.162 54.82 3.465 ;
      RECT 54.745 3.185 54.81 3.465 ;
      RECT 54.245 2.68 54.435 2.89 ;
      RECT 52.82 2.605 53.08 2.865 ;
      RECT 53.17 2.6 53.265 2.81 ;
      RECT 53.145 2.615 53.155 2.81 ;
      RECT 54.435 2.687 54.445 2.885 ;
      RECT 54.235 2.687 54.245 2.885 ;
      RECT 54.22 2.702 54.235 2.875 ;
      RECT 54.215 2.71 54.22 2.868 ;
      RECT 54.205 2.713 54.215 2.865 ;
      RECT 54.17 2.712 54.205 2.863 ;
      RECT 54.141 2.708 54.17 2.86 ;
      RECT 54.055 2.703 54.141 2.857 ;
      RECT 53.995 2.697 54.055 2.853 ;
      RECT 53.966 2.693 53.995 2.85 ;
      RECT 53.88 2.685 53.966 2.847 ;
      RECT 53.871 2.679 53.88 2.845 ;
      RECT 53.785 2.674 53.871 2.843 ;
      RECT 53.762 2.669 53.785 2.84 ;
      RECT 53.676 2.663 53.762 2.837 ;
      RECT 53.59 2.654 53.676 2.832 ;
      RECT 53.58 2.649 53.59 2.83 ;
      RECT 53.561 2.648 53.58 2.829 ;
      RECT 53.475 2.643 53.561 2.825 ;
      RECT 53.455 2.638 53.475 2.821 ;
      RECT 53.395 2.633 53.455 2.818 ;
      RECT 53.37 2.623 53.395 2.816 ;
      RECT 53.365 2.616 53.37 2.815 ;
      RECT 53.355 2.607 53.365 2.814 ;
      RECT 53.351 2.6 53.355 2.814 ;
      RECT 53.265 2.6 53.351 2.812 ;
      RECT 53.155 2.607 53.17 2.81 ;
      RECT 53.14 2.617 53.145 2.81 ;
      RECT 53.12 2.62 53.14 2.807 ;
      RECT 53.09 2.62 53.12 2.803 ;
      RECT 53.08 2.62 53.09 2.803 ;
      RECT 53.995 3.115 54.255 3.375 ;
      RECT 53.925 3.125 54.255 3.335 ;
      RECT 53.915 3.132 54.255 3.33 ;
      RECT 53.335 3.12 53.595 3.38 ;
      RECT 53.335 3.16 53.7 3.37 ;
      RECT 53.335 3.162 53.705 3.369 ;
      RECT 53.335 3.17 53.71 3.366 ;
      RECT 52.26 2.245 52.36 3.77 ;
      RECT 52.45 3.385 52.5 3.645 ;
      RECT 52.445 2.258 52.45 2.445 ;
      RECT 52.44 3.366 52.45 3.645 ;
      RECT 52.44 2.255 52.445 2.453 ;
      RECT 52.425 2.249 52.44 2.46 ;
      RECT 52.435 3.354 52.44 3.728 ;
      RECT 52.425 3.342 52.435 3.765 ;
      RECT 52.415 2.245 52.425 2.467 ;
      RECT 52.415 3.327 52.425 3.77 ;
      RECT 52.41 2.245 52.415 2.475 ;
      RECT 52.39 3.297 52.415 3.77 ;
      RECT 52.37 2.245 52.41 2.523 ;
      RECT 52.38 3.257 52.39 3.77 ;
      RECT 52.37 3.212 52.38 3.77 ;
      RECT 52.365 2.245 52.37 2.593 ;
      RECT 52.365 3.17 52.37 3.77 ;
      RECT 52.36 2.245 52.365 3.07 ;
      RECT 52.36 3.152 52.365 3.77 ;
      RECT 52.25 2.248 52.26 3.77 ;
      RECT 52.235 2.255 52.25 3.766 ;
      RECT 52.23 2.265 52.235 3.761 ;
      RECT 52.225 2.465 52.23 3.653 ;
      RECT 52.22 2.55 52.225 3.205 ;
      RECT 51.1 7.765 51.39 7.995 ;
      RECT 51.16 6.285 51.33 7.995 ;
      RECT 51.105 6.655 51.455 7.005 ;
      RECT 51.1 6.285 51.39 6.515 ;
      RECT 51.1 2.365 51.39 2.595 ;
      RECT 51.16 0.885 51.33 2.595 ;
      RECT 51.1 0.885 51.39 1.115 ;
      RECT 50.69 2.735 51.02 2.965 ;
      RECT 50.69 2.765 51.19 2.935 ;
      RECT 50.69 2.395 50.88 2.965 ;
      RECT 50.11 2.365 50.4 2.595 ;
      RECT 50.11 2.395 50.88 2.565 ;
      RECT 50.17 0.885 50.34 2.595 ;
      RECT 50.11 0.885 50.4 1.115 ;
      RECT 50.11 7.765 50.4 7.995 ;
      RECT 50.17 6.285 50.34 7.995 ;
      RECT 50.11 6.285 50.4 6.515 ;
      RECT 50.11 6.325 50.96 6.485 ;
      RECT 50.79 5.915 50.96 6.485 ;
      RECT 50.11 6.32 50.5 6.485 ;
      RECT 50.73 5.915 51.02 6.145 ;
      RECT 50.73 5.945 51.19 6.115 ;
      RECT 49.74 2.735 50.03 2.965 ;
      RECT 49.74 2.765 50.2 2.935 ;
      RECT 49.8 1.655 49.965 2.965 ;
      RECT 48.315 1.625 48.605 1.855 ;
      RECT 48.315 1.655 49.965 1.825 ;
      RECT 48.375 0.885 48.545 1.855 ;
      RECT 48.315 0.885 48.605 1.115 ;
      RECT 48.315 7.765 48.605 7.995 ;
      RECT 48.375 7.025 48.545 7.995 ;
      RECT 48.375 7.12 49.965 7.29 ;
      RECT 49.795 5.915 49.965 7.29 ;
      RECT 48.315 7.025 48.605 7.255 ;
      RECT 49.74 5.915 50.03 6.145 ;
      RECT 49.74 5.945 50.2 6.115 ;
      RECT 46.35 3.43 46.7 3.78 ;
      RECT 46.44 2.025 46.61 3.78 ;
      RECT 48.745 1.965 49.095 2.315 ;
      RECT 46.44 2.025 48.06 2.2 ;
      RECT 46.44 2.025 49.095 2.195 ;
      RECT 48.77 6.655 49.095 6.98 ;
      RECT 44.2 6.615 44.55 6.965 ;
      RECT 48.745 6.655 49.095 6.885 ;
      RECT 43.985 6.655 44.55 6.885 ;
      RECT 43.815 6.685 49.095 6.855 ;
      RECT 47.97 2.365 48.29 2.685 ;
      RECT 47.94 2.365 48.29 2.595 ;
      RECT 47.77 2.395 48.29 2.565 ;
      RECT 47.97 6.225 48.29 6.545 ;
      RECT 47.94 6.285 48.29 6.515 ;
      RECT 47.77 6.315 48.29 6.485 ;
      RECT 46.925 2.705 47.275 3.055 ;
      RECT 46.925 2.765 47.405 2.935 ;
      RECT 46.915 5.84 47.265 6.19 ;
      RECT 42.185 5.915 42.475 6.145 ;
      RECT 42.185 5.945 47.405 6.115 ;
      RECT 43.75 3.665 43.79 3.925 ;
      RECT 43.79 3.645 43.795 3.655 ;
      RECT 45.12 2.89 45.13 3.111 ;
      RECT 45.05 2.885 45.12 3.236 ;
      RECT 45.04 2.885 45.05 3.363 ;
      RECT 45.015 2.885 45.04 3.41 ;
      RECT 44.99 2.885 45.015 3.488 ;
      RECT 44.97 2.885 44.99 3.558 ;
      RECT 44.945 2.885 44.97 3.598 ;
      RECT 44.935 2.885 44.945 3.618 ;
      RECT 44.925 2.887 44.935 3.626 ;
      RECT 44.92 2.892 44.925 3.083 ;
      RECT 44.92 3.092 44.925 3.627 ;
      RECT 44.915 3.137 44.92 3.628 ;
      RECT 44.905 3.202 44.915 3.629 ;
      RECT 44.895 3.297 44.905 3.631 ;
      RECT 44.89 3.35 44.895 3.633 ;
      RECT 44.885 3.37 44.89 3.634 ;
      RECT 44.83 3.395 44.885 3.64 ;
      RECT 44.79 3.43 44.83 3.649 ;
      RECT 44.78 3.447 44.79 3.654 ;
      RECT 44.771 3.453 44.78 3.656 ;
      RECT 44.685 3.491 44.771 3.667 ;
      RECT 44.68 3.53 44.685 3.677 ;
      RECT 44.605 3.537 44.68 3.687 ;
      RECT 44.585 3.547 44.605 3.698 ;
      RECT 44.555 3.554 44.585 3.706 ;
      RECT 44.53 3.561 44.555 3.713 ;
      RECT 44.506 3.567 44.53 3.718 ;
      RECT 44.42 3.58 44.506 3.73 ;
      RECT 44.342 3.587 44.42 3.748 ;
      RECT 44.256 3.582 44.342 3.766 ;
      RECT 44.17 3.577 44.256 3.786 ;
      RECT 44.09 3.571 44.17 3.803 ;
      RECT 44.025 3.567 44.09 3.832 ;
      RECT 44.02 3.281 44.025 3.305 ;
      RECT 44.01 3.557 44.025 3.86 ;
      RECT 44.015 3.275 44.02 3.345 ;
      RECT 44.01 3.269 44.015 3.415 ;
      RECT 44.005 3.263 44.01 3.493 ;
      RECT 44.005 3.54 44.01 3.925 ;
      RECT 43.997 3.26 44.005 3.925 ;
      RECT 43.911 3.258 43.997 3.925 ;
      RECT 43.825 3.256 43.911 3.925 ;
      RECT 43.815 3.257 43.825 3.925 ;
      RECT 43.81 3.262 43.815 3.925 ;
      RECT 43.8 3.275 43.81 3.925 ;
      RECT 43.795 3.297 43.8 3.925 ;
      RECT 43.79 3.657 43.795 3.925 ;
      RECT 44.42 3.125 44.425 3.345 ;
      RECT 44.925 2.16 44.96 2.42 ;
      RECT 44.91 2.16 44.925 2.428 ;
      RECT 44.881 2.16 44.91 2.45 ;
      RECT 44.795 2.16 44.881 2.51 ;
      RECT 44.775 2.16 44.795 2.575 ;
      RECT 44.715 2.16 44.775 2.74 ;
      RECT 44.71 2.16 44.715 2.888 ;
      RECT 44.705 2.16 44.71 2.9 ;
      RECT 44.7 2.16 44.705 2.926 ;
      RECT 44.67 2.346 44.7 3.006 ;
      RECT 44.665 2.394 44.67 3.095 ;
      RECT 44.66 2.408 44.665 3.11 ;
      RECT 44.655 2.427 44.66 3.14 ;
      RECT 44.65 2.442 44.655 3.156 ;
      RECT 44.645 2.457 44.65 3.178 ;
      RECT 44.64 2.477 44.645 3.2 ;
      RECT 44.63 2.497 44.64 3.233 ;
      RECT 44.615 2.539 44.63 3.295 ;
      RECT 44.61 2.57 44.615 3.335 ;
      RECT 44.605 2.582 44.61 3.34 ;
      RECT 44.6 2.594 44.605 3.345 ;
      RECT 44.595 2.607 44.6 3.345 ;
      RECT 44.59 2.625 44.595 3.345 ;
      RECT 44.585 2.645 44.59 3.345 ;
      RECT 44.58 2.657 44.585 3.345 ;
      RECT 44.575 2.67 44.58 3.345 ;
      RECT 44.555 2.705 44.575 3.345 ;
      RECT 44.505 2.807 44.555 3.345 ;
      RECT 44.5 2.892 44.505 3.345 ;
      RECT 44.495 2.9 44.5 3.345 ;
      RECT 44.49 2.917 44.495 3.345 ;
      RECT 44.485 2.932 44.49 3.345 ;
      RECT 44.45 2.997 44.485 3.345 ;
      RECT 44.435 3.062 44.45 3.345 ;
      RECT 44.43 3.092 44.435 3.345 ;
      RECT 44.425 3.117 44.43 3.345 ;
      RECT 44.41 3.127 44.42 3.345 ;
      RECT 44.395 3.14 44.41 3.338 ;
      RECT 44.14 2.73 44.21 2.94 ;
      RECT 43.93 2.707 43.935 2.9 ;
      RECT 41.385 2.635 41.645 2.895 ;
      RECT 44.22 2.917 44.225 2.92 ;
      RECT 44.21 2.735 44.22 2.935 ;
      RECT 44.111 2.728 44.14 2.94 ;
      RECT 44.025 2.72 44.111 2.94 ;
      RECT 44.01 2.714 44.025 2.938 ;
      RECT 43.99 2.713 44.01 2.925 ;
      RECT 43.985 2.712 43.99 2.908 ;
      RECT 43.935 2.709 43.985 2.903 ;
      RECT 43.905 2.706 43.93 2.898 ;
      RECT 43.885 2.704 43.905 2.893 ;
      RECT 43.87 2.702 43.885 2.89 ;
      RECT 43.84 2.7 43.87 2.888 ;
      RECT 43.775 2.696 43.84 2.88 ;
      RECT 43.745 2.691 43.775 2.875 ;
      RECT 43.725 2.689 43.745 2.873 ;
      RECT 43.695 2.686 43.725 2.868 ;
      RECT 43.635 2.682 43.695 2.86 ;
      RECT 43.63 2.679 43.635 2.855 ;
      RECT 43.56 2.677 43.63 2.85 ;
      RECT 43.531 2.673 43.56 2.843 ;
      RECT 43.445 2.668 43.531 2.835 ;
      RECT 43.411 2.663 43.445 2.827 ;
      RECT 43.325 2.655 43.411 2.819 ;
      RECT 43.286 2.648 43.325 2.811 ;
      RECT 43.2 2.643 43.286 2.803 ;
      RECT 43.135 2.637 43.2 2.793 ;
      RECT 43.115 2.632 43.135 2.788 ;
      RECT 43.106 2.629 43.115 2.787 ;
      RECT 43.02 2.625 43.106 2.781 ;
      RECT 42.98 2.621 43.02 2.773 ;
      RECT 42.96 2.617 42.98 2.771 ;
      RECT 42.9 2.617 42.96 2.768 ;
      RECT 42.88 2.62 42.9 2.766 ;
      RECT 42.859 2.62 42.88 2.766 ;
      RECT 42.773 2.622 42.859 2.77 ;
      RECT 42.687 2.624 42.773 2.776 ;
      RECT 42.601 2.626 42.687 2.783 ;
      RECT 42.515 2.629 42.601 2.789 ;
      RECT 42.481 2.63 42.515 2.794 ;
      RECT 42.395 2.633 42.481 2.799 ;
      RECT 42.366 2.64 42.395 2.804 ;
      RECT 42.28 2.64 42.366 2.809 ;
      RECT 42.247 2.64 42.28 2.814 ;
      RECT 42.161 2.642 42.247 2.819 ;
      RECT 42.075 2.644 42.161 2.826 ;
      RECT 42.011 2.646 42.075 2.832 ;
      RECT 41.925 2.648 42.011 2.838 ;
      RECT 41.922 2.65 41.925 2.841 ;
      RECT 41.836 2.651 41.922 2.845 ;
      RECT 41.75 2.654 41.836 2.852 ;
      RECT 41.731 2.656 41.75 2.856 ;
      RECT 41.645 2.658 41.731 2.861 ;
      RECT 41.375 2.67 41.385 2.865 ;
      RECT 43.555 7.765 43.845 7.995 ;
      RECT 43.615 7.025 43.785 7.995 ;
      RECT 43.505 7.055 43.88 7.425 ;
      RECT 43.555 7.025 43.845 7.425 ;
      RECT 43.61 2.25 43.795 2.46 ;
      RECT 43.605 2.251 43.8 2.458 ;
      RECT 43.6 2.256 43.81 2.453 ;
      RECT 43.595 2.232 43.6 2.45 ;
      RECT 43.565 2.229 43.595 2.443 ;
      RECT 43.56 2.225 43.565 2.434 ;
      RECT 43.525 2.256 43.81 2.429 ;
      RECT 43.3 2.165 43.56 2.425 ;
      RECT 43.6 2.234 43.605 2.453 ;
      RECT 43.605 2.235 43.61 2.458 ;
      RECT 43.3 2.247 43.68 2.425 ;
      RECT 43.3 2.245 43.665 2.425 ;
      RECT 43.3 2.24 43.655 2.425 ;
      RECT 43.255 3.155 43.305 3.44 ;
      RECT 43.2 3.125 43.205 3.44 ;
      RECT 43.17 3.105 43.175 3.44 ;
      RECT 43.32 3.155 43.38 3.415 ;
      RECT 43.315 3.155 43.32 3.423 ;
      RECT 43.305 3.155 43.315 3.435 ;
      RECT 43.22 3.145 43.255 3.44 ;
      RECT 43.215 3.132 43.22 3.44 ;
      RECT 43.205 3.127 43.215 3.44 ;
      RECT 43.185 3.117 43.2 3.44 ;
      RECT 43.175 3.11 43.185 3.44 ;
      RECT 43.165 3.102 43.17 3.44 ;
      RECT 43.135 3.092 43.165 3.44 ;
      RECT 43.12 3.08 43.135 3.44 ;
      RECT 43.105 3.07 43.12 3.435 ;
      RECT 43.085 3.06 43.105 3.41 ;
      RECT 43.075 3.052 43.085 3.387 ;
      RECT 43.045 3.035 43.075 3.377 ;
      RECT 43.04 3.012 43.045 3.368 ;
      RECT 43.035 2.999 43.04 3.366 ;
      RECT 43.02 2.975 43.035 3.36 ;
      RECT 43.015 2.951 43.02 3.354 ;
      RECT 43.005 2.94 43.015 3.349 ;
      RECT 43 2.93 43.005 3.345 ;
      RECT 42.995 2.922 43 3.342 ;
      RECT 42.985 2.917 42.995 3.338 ;
      RECT 42.98 2.912 42.985 3.334 ;
      RECT 42.895 2.91 42.98 3.309 ;
      RECT 42.865 2.91 42.895 3.275 ;
      RECT 42.85 2.91 42.865 3.258 ;
      RECT 42.795 2.91 42.85 3.203 ;
      RECT 42.79 2.915 42.795 3.152 ;
      RECT 42.78 2.92 42.79 3.142 ;
      RECT 42.775 2.93 42.78 3.128 ;
      RECT 42.725 3.67 42.985 3.93 ;
      RECT 42.645 3.685 42.985 3.906 ;
      RECT 42.625 3.685 42.985 3.901 ;
      RECT 42.601 3.685 42.985 3.899 ;
      RECT 42.515 3.685 42.985 3.894 ;
      RECT 42.365 3.625 42.625 3.89 ;
      RECT 42.32 3.685 42.985 3.885 ;
      RECT 42.315 3.692 42.985 3.88 ;
      RECT 42.33 3.68 42.645 3.89 ;
      RECT 42.22 2.115 42.48 2.375 ;
      RECT 42.22 2.172 42.485 2.368 ;
      RECT 42.22 2.202 42.49 2.3 ;
      RECT 42.28 2.633 42.395 2.635 ;
      RECT 42.366 2.63 42.395 2.635 ;
      RECT 41.39 3.634 41.415 3.874 ;
      RECT 41.375 3.637 41.465 3.868 ;
      RECT 41.37 3.642 41.551 3.863 ;
      RECT 41.365 3.65 41.615 3.861 ;
      RECT 41.365 3.65 41.625 3.86 ;
      RECT 41.36 3.657 41.635 3.853 ;
      RECT 41.36 3.657 41.721 3.842 ;
      RECT 41.355 3.692 41.721 3.838 ;
      RECT 41.355 3.692 41.73 3.827 ;
      RECT 41.635 3.565 41.895 3.825 ;
      RECT 41.345 3.742 41.895 3.823 ;
      RECT 41.615 3.61 41.635 3.858 ;
      RECT 41.551 3.613 41.615 3.862 ;
      RECT 41.465 3.618 41.551 3.867 ;
      RECT 41.395 3.629 41.895 3.825 ;
      RECT 41.415 3.623 41.465 3.872 ;
      RECT 41.54 2.1 41.55 2.362 ;
      RECT 41.53 2.157 41.54 2.365 ;
      RECT 41.505 2.162 41.53 2.371 ;
      RECT 41.48 2.166 41.505 2.383 ;
      RECT 41.47 2.169 41.48 2.393 ;
      RECT 41.465 2.17 41.47 2.398 ;
      RECT 41.46 2.171 41.465 2.403 ;
      RECT 41.455 2.172 41.46 2.405 ;
      RECT 41.43 2.175 41.455 2.408 ;
      RECT 41.4 2.181 41.43 2.411 ;
      RECT 41.335 2.192 41.4 2.414 ;
      RECT 41.29 2.2 41.335 2.418 ;
      RECT 41.275 2.2 41.29 2.426 ;
      RECT 41.27 2.201 41.275 2.433 ;
      RECT 41.265 2.203 41.27 2.436 ;
      RECT 41.26 2.207 41.265 2.439 ;
      RECT 41.25 2.215 41.26 2.443 ;
      RECT 41.245 2.228 41.25 2.448 ;
      RECT 41.24 2.236 41.245 2.45 ;
      RECT 41.235 2.242 41.24 2.45 ;
      RECT 41.23 2.246 41.235 2.453 ;
      RECT 41.225 2.248 41.23 2.456 ;
      RECT 41.22 2.251 41.225 2.459 ;
      RECT 41.21 2.256 41.22 2.463 ;
      RECT 41.205 2.262 41.21 2.468 ;
      RECT 41.195 2.268 41.205 2.472 ;
      RECT 41.18 2.275 41.195 2.478 ;
      RECT 41.151 2.289 41.18 2.488 ;
      RECT 41.065 2.324 41.151 2.52 ;
      RECT 41.045 2.357 41.065 2.549 ;
      RECT 41.025 2.37 41.045 2.56 ;
      RECT 41.005 2.382 41.025 2.571 ;
      RECT 40.955 2.404 41.005 2.591 ;
      RECT 40.94 2.422 40.955 2.608 ;
      RECT 40.935 2.428 40.94 2.611 ;
      RECT 40.93 2.432 40.935 2.614 ;
      RECT 40.925 2.436 40.93 2.618 ;
      RECT 40.92 2.438 40.925 2.621 ;
      RECT 40.91 2.445 40.92 2.624 ;
      RECT 40.905 2.45 40.91 2.628 ;
      RECT 40.9 2.452 40.905 2.631 ;
      RECT 40.895 2.456 40.9 2.634 ;
      RECT 40.89 2.458 40.895 2.638 ;
      RECT 40.875 2.463 40.89 2.643 ;
      RECT 40.87 2.468 40.875 2.646 ;
      RECT 40.865 2.476 40.87 2.649 ;
      RECT 40.86 2.478 40.865 2.652 ;
      RECT 40.855 2.48 40.86 2.655 ;
      RECT 40.845 2.482 40.855 2.661 ;
      RECT 40.81 2.496 40.845 2.673 ;
      RECT 40.8 2.511 40.81 2.683 ;
      RECT 40.725 2.54 40.8 2.707 ;
      RECT 40.72 2.565 40.725 2.73 ;
      RECT 40.705 2.569 40.72 2.736 ;
      RECT 40.695 2.577 40.705 2.741 ;
      RECT 40.665 2.59 40.695 2.745 ;
      RECT 40.655 2.605 40.665 2.75 ;
      RECT 40.645 2.61 40.655 2.753 ;
      RECT 40.64 2.612 40.645 2.755 ;
      RECT 40.625 2.615 40.64 2.758 ;
      RECT 40.62 2.617 40.625 2.761 ;
      RECT 40.6 2.622 40.62 2.765 ;
      RECT 40.57 2.627 40.6 2.773 ;
      RECT 40.545 2.634 40.57 2.781 ;
      RECT 40.54 2.639 40.545 2.786 ;
      RECT 40.51 2.642 40.54 2.79 ;
      RECT 40.47 2.645 40.51 2.8 ;
      RECT 40.435 2.642 40.47 2.812 ;
      RECT 40.425 2.638 40.435 2.819 ;
      RECT 40.4 2.634 40.425 2.825 ;
      RECT 40.395 2.63 40.4 2.83 ;
      RECT 40.355 2.627 40.395 2.83 ;
      RECT 40.34 2.612 40.355 2.831 ;
      RECT 40.317 2.6 40.34 2.831 ;
      RECT 40.231 2.6 40.317 2.832 ;
      RECT 40.145 2.6 40.231 2.834 ;
      RECT 40.125 2.6 40.145 2.831 ;
      RECT 40.12 2.605 40.125 2.826 ;
      RECT 40.115 2.61 40.12 2.824 ;
      RECT 40.105 2.62 40.115 2.822 ;
      RECT 40.1 2.626 40.105 2.815 ;
      RECT 40.095 2.628 40.1 2.8 ;
      RECT 40.09 2.632 40.095 2.79 ;
      RECT 41.55 2.1 41.8 2.36 ;
      RECT 39.275 3.635 39.535 3.895 ;
      RECT 41.57 3.125 41.575 3.335 ;
      RECT 41.575 3.13 41.585 3.33 ;
      RECT 41.525 3.125 41.57 3.35 ;
      RECT 41.515 3.125 41.525 3.37 ;
      RECT 41.496 3.125 41.515 3.375 ;
      RECT 41.41 3.125 41.496 3.372 ;
      RECT 41.38 3.127 41.41 3.37 ;
      RECT 41.325 3.137 41.38 3.368 ;
      RECT 41.26 3.151 41.325 3.366 ;
      RECT 41.255 3.159 41.26 3.365 ;
      RECT 41.24 3.162 41.255 3.363 ;
      RECT 41.175 3.172 41.24 3.359 ;
      RECT 41.127 3.186 41.175 3.36 ;
      RECT 41.041 3.203 41.127 3.374 ;
      RECT 40.955 3.224 41.041 3.391 ;
      RECT 40.935 3.237 40.955 3.401 ;
      RECT 40.89 3.245 40.935 3.408 ;
      RECT 40.855 3.253 40.89 3.416 ;
      RECT 40.821 3.261 40.855 3.424 ;
      RECT 40.735 3.275 40.821 3.436 ;
      RECT 40.7 3.292 40.735 3.448 ;
      RECT 40.691 3.301 40.7 3.452 ;
      RECT 40.605 3.319 40.691 3.469 ;
      RECT 40.546 3.346 40.605 3.496 ;
      RECT 40.46 3.373 40.546 3.524 ;
      RECT 40.44 3.395 40.46 3.544 ;
      RECT 40.38 3.41 40.44 3.56 ;
      RECT 40.37 3.422 40.38 3.573 ;
      RECT 40.365 3.427 40.37 3.576 ;
      RECT 40.355 3.43 40.365 3.579 ;
      RECT 40.35 3.432 40.355 3.582 ;
      RECT 40.32 3.44 40.35 3.589 ;
      RECT 40.305 3.447 40.32 3.597 ;
      RECT 40.295 3.452 40.305 3.601 ;
      RECT 40.29 3.455 40.295 3.604 ;
      RECT 40.28 3.457 40.29 3.607 ;
      RECT 40.245 3.467 40.28 3.616 ;
      RECT 40.17 3.49 40.245 3.638 ;
      RECT 40.15 3.508 40.17 3.656 ;
      RECT 40.12 3.515 40.15 3.666 ;
      RECT 40.1 3.523 40.12 3.676 ;
      RECT 40.09 3.529 40.1 3.683 ;
      RECT 40.071 3.534 40.09 3.689 ;
      RECT 39.985 3.554 40.071 3.709 ;
      RECT 39.97 3.574 39.985 3.728 ;
      RECT 39.925 3.586 39.97 3.739 ;
      RECT 39.86 3.607 39.925 3.762 ;
      RECT 39.82 3.627 39.86 3.783 ;
      RECT 39.81 3.637 39.82 3.793 ;
      RECT 39.76 3.649 39.81 3.804 ;
      RECT 39.74 3.665 39.76 3.816 ;
      RECT 39.71 3.675 39.74 3.822 ;
      RECT 39.7 3.68 39.71 3.824 ;
      RECT 39.631 3.681 39.7 3.83 ;
      RECT 39.545 3.683 39.631 3.84 ;
      RECT 39.535 3.684 39.545 3.845 ;
      RECT 40.805 3.71 40.995 3.92 ;
      RECT 40.795 3.715 41.005 3.913 ;
      RECT 40.78 3.715 41.005 3.878 ;
      RECT 40.7 3.6 40.96 3.86 ;
      RECT 39.615 3.13 39.8 3.425 ;
      RECT 39.605 3.13 39.8 3.423 ;
      RECT 39.59 3.13 39.805 3.418 ;
      RECT 39.59 3.13 39.81 3.415 ;
      RECT 39.585 3.13 39.81 3.413 ;
      RECT 39.58 3.385 39.81 3.403 ;
      RECT 39.585 3.13 39.845 3.39 ;
      RECT 39.545 2.165 39.805 2.425 ;
      RECT 39.355 2.09 39.441 2.423 ;
      RECT 39.33 2.094 39.485 2.419 ;
      RECT 39.441 2.086 39.485 2.419 ;
      RECT 39.441 2.087 39.49 2.418 ;
      RECT 39.355 2.092 39.505 2.417 ;
      RECT 39.33 2.1 39.545 2.416 ;
      RECT 39.325 2.095 39.505 2.411 ;
      RECT 39.315 2.11 39.545 2.318 ;
      RECT 39.315 2.162 39.745 2.318 ;
      RECT 39.315 2.155 39.725 2.318 ;
      RECT 39.315 2.142 39.695 2.318 ;
      RECT 39.315 2.13 39.635 2.318 ;
      RECT 39.315 2.115 39.61 2.318 ;
      RECT 38.515 2.745 38.65 3.04 ;
      RECT 38.775 2.768 38.78 2.955 ;
      RECT 39.495 2.665 39.64 2.9 ;
      RECT 39.655 2.665 39.66 2.89 ;
      RECT 39.69 2.676 39.695 2.87 ;
      RECT 39.685 2.668 39.69 2.875 ;
      RECT 39.665 2.665 39.685 2.88 ;
      RECT 39.66 2.665 39.665 2.888 ;
      RECT 39.65 2.665 39.655 2.893 ;
      RECT 39.64 2.665 39.65 2.898 ;
      RECT 39.47 2.667 39.495 2.9 ;
      RECT 39.42 2.674 39.47 2.9 ;
      RECT 39.415 2.679 39.42 2.9 ;
      RECT 39.376 2.684 39.415 2.901 ;
      RECT 39.29 2.696 39.376 2.902 ;
      RECT 39.281 2.706 39.29 2.902 ;
      RECT 39.195 2.715 39.281 2.904 ;
      RECT 39.171 2.725 39.195 2.906 ;
      RECT 39.085 2.736 39.171 2.907 ;
      RECT 39.055 2.747 39.085 2.909 ;
      RECT 39.025 2.752 39.055 2.911 ;
      RECT 39 2.758 39.025 2.914 ;
      RECT 38.985 2.763 39 2.915 ;
      RECT 38.94 2.769 38.985 2.915 ;
      RECT 38.935 2.774 38.94 2.916 ;
      RECT 38.915 2.774 38.935 2.918 ;
      RECT 38.895 2.772 38.915 2.923 ;
      RECT 38.86 2.771 38.895 2.93 ;
      RECT 38.83 2.77 38.86 2.94 ;
      RECT 38.78 2.769 38.83 2.95 ;
      RECT 38.69 2.766 38.775 3.04 ;
      RECT 38.665 2.76 38.69 3.04 ;
      RECT 38.65 2.75 38.665 3.04 ;
      RECT 38.465 2.745 38.515 2.96 ;
      RECT 38.455 2.75 38.465 2.95 ;
      RECT 38.695 3.225 38.955 3.485 ;
      RECT 38.695 3.225 38.985 3.378 ;
      RECT 38.695 3.225 39.02 3.363 ;
      RECT 38.95 3.145 39.14 3.355 ;
      RECT 38.94 3.15 39.15 3.348 ;
      RECT 38.905 3.22 39.15 3.348 ;
      RECT 38.935 3.162 38.955 3.485 ;
      RECT 38.92 3.21 39.15 3.348 ;
      RECT 38.925 3.182 38.955 3.485 ;
      RECT 38.005 2.25 38.075 3.355 ;
      RECT 38.74 2.355 39 2.615 ;
      RECT 38.32 2.401 38.335 2.61 ;
      RECT 38.656 2.414 38.74 2.565 ;
      RECT 38.57 2.411 38.656 2.565 ;
      RECT 38.531 2.409 38.57 2.565 ;
      RECT 38.445 2.407 38.531 2.565 ;
      RECT 38.385 2.405 38.445 2.576 ;
      RECT 38.35 2.403 38.385 2.594 ;
      RECT 38.335 2.401 38.35 2.605 ;
      RECT 38.305 2.401 38.32 2.618 ;
      RECT 38.295 2.401 38.305 2.623 ;
      RECT 38.27 2.4 38.295 2.628 ;
      RECT 38.255 2.395 38.27 2.634 ;
      RECT 38.25 2.388 38.255 2.639 ;
      RECT 38.225 2.379 38.25 2.645 ;
      RECT 38.18 2.358 38.225 2.658 ;
      RECT 38.17 2.342 38.18 2.668 ;
      RECT 38.155 2.335 38.17 2.678 ;
      RECT 38.145 2.328 38.155 2.695 ;
      RECT 38.14 2.325 38.145 2.725 ;
      RECT 38.135 2.323 38.14 2.755 ;
      RECT 38.13 2.321 38.135 2.792 ;
      RECT 38.115 2.317 38.13 2.859 ;
      RECT 38.115 3.15 38.125 3.35 ;
      RECT 38.11 2.313 38.115 2.985 ;
      RECT 38.11 3.137 38.115 3.355 ;
      RECT 38.105 2.311 38.11 3.07 ;
      RECT 38.105 3.127 38.11 3.355 ;
      RECT 38.09 2.282 38.105 3.355 ;
      RECT 38.075 2.255 38.09 3.355 ;
      RECT 38 2.25 38.005 2.605 ;
      RECT 38 2.66 38.005 3.355 ;
      RECT 37.985 2.25 38 2.583 ;
      RECT 37.995 2.682 38 3.355 ;
      RECT 37.985 2.722 37.995 3.355 ;
      RECT 37.95 2.25 37.985 2.525 ;
      RECT 37.98 2.757 37.985 3.355 ;
      RECT 37.965 2.812 37.98 3.355 ;
      RECT 37.96 2.877 37.965 3.355 ;
      RECT 37.945 2.925 37.96 3.355 ;
      RECT 37.92 2.25 37.95 2.48 ;
      RECT 37.94 2.98 37.945 3.355 ;
      RECT 37.925 3.04 37.94 3.355 ;
      RECT 37.92 3.088 37.925 3.353 ;
      RECT 37.915 2.25 37.92 2.473 ;
      RECT 37.915 3.12 37.92 3.348 ;
      RECT 37.89 2.25 37.915 2.465 ;
      RECT 37.88 2.255 37.89 2.455 ;
      RECT 38.095 3.53 38.115 3.77 ;
      RECT 37.325 3.46 37.33 3.67 ;
      RECT 38.605 3.533 38.615 3.728 ;
      RECT 38.6 3.523 38.605 3.731 ;
      RECT 38.52 3.52 38.6 3.754 ;
      RECT 38.516 3.52 38.52 3.776 ;
      RECT 38.43 3.52 38.516 3.786 ;
      RECT 38.415 3.52 38.43 3.794 ;
      RECT 38.386 3.521 38.415 3.792 ;
      RECT 38.3 3.526 38.386 3.788 ;
      RECT 38.287 3.53 38.3 3.784 ;
      RECT 38.201 3.53 38.287 3.78 ;
      RECT 38.115 3.53 38.201 3.774 ;
      RECT 38.031 3.53 38.095 3.768 ;
      RECT 37.945 3.53 38.031 3.763 ;
      RECT 37.925 3.53 37.945 3.759 ;
      RECT 37.865 3.525 37.925 3.756 ;
      RECT 37.837 3.519 37.865 3.753 ;
      RECT 37.751 3.514 37.837 3.749 ;
      RECT 37.665 3.508 37.751 3.743 ;
      RECT 37.59 3.49 37.665 3.738 ;
      RECT 37.555 3.467 37.59 3.734 ;
      RECT 37.545 3.457 37.555 3.733 ;
      RECT 37.49 3.455 37.545 3.732 ;
      RECT 37.415 3.455 37.49 3.728 ;
      RECT 37.405 3.455 37.415 3.723 ;
      RECT 37.39 3.455 37.405 3.715 ;
      RECT 37.34 3.457 37.39 3.693 ;
      RECT 37.33 3.46 37.34 3.673 ;
      RECT 37.32 3.465 37.325 3.668 ;
      RECT 37.315 3.47 37.32 3.663 ;
      RECT 37.44 2.635 37.7 2.895 ;
      RECT 37.44 2.65 37.72 2.86 ;
      RECT 37.44 2.655 37.73 2.855 ;
      RECT 35.425 2.115 35.685 2.375 ;
      RECT 35.415 2.145 35.685 2.355 ;
      RECT 37.335 2.06 37.595 2.32 ;
      RECT 37.33 2.135 37.335 2.321 ;
      RECT 37.305 2.14 37.33 2.323 ;
      RECT 37.29 2.147 37.305 2.326 ;
      RECT 37.23 2.165 37.29 2.331 ;
      RECT 37.2 2.185 37.23 2.338 ;
      RECT 37.175 2.193 37.2 2.343 ;
      RECT 37.15 2.201 37.175 2.345 ;
      RECT 37.132 2.205 37.15 2.344 ;
      RECT 37.046 2.203 37.132 2.344 ;
      RECT 36.96 2.201 37.046 2.344 ;
      RECT 36.874 2.199 36.96 2.343 ;
      RECT 36.788 2.197 36.874 2.343 ;
      RECT 36.702 2.195 36.788 2.343 ;
      RECT 36.616 2.193 36.702 2.343 ;
      RECT 36.53 2.191 36.616 2.342 ;
      RECT 36.512 2.19 36.53 2.342 ;
      RECT 36.426 2.189 36.512 2.342 ;
      RECT 36.34 2.187 36.426 2.342 ;
      RECT 36.254 2.186 36.34 2.341 ;
      RECT 36.168 2.185 36.254 2.341 ;
      RECT 36.082 2.183 36.168 2.341 ;
      RECT 35.996 2.182 36.082 2.341 ;
      RECT 35.91 2.18 35.996 2.34 ;
      RECT 35.886 2.178 35.91 2.34 ;
      RECT 35.8 2.171 35.886 2.34 ;
      RECT 35.771 2.163 35.8 2.34 ;
      RECT 35.685 2.155 35.771 2.34 ;
      RECT 35.405 2.152 35.415 2.35 ;
      RECT 36.91 3.115 36.915 3.465 ;
      RECT 36.68 3.205 36.82 3.465 ;
      RECT 37.155 2.89 37.2 3.1 ;
      RECT 37.21 2.901 37.22 3.095 ;
      RECT 37.2 2.893 37.21 3.1 ;
      RECT 37.135 2.89 37.155 3.105 ;
      RECT 37.105 2.89 37.135 3.128 ;
      RECT 37.095 2.89 37.105 3.153 ;
      RECT 37.09 2.89 37.095 3.163 ;
      RECT 37.035 2.89 37.09 3.203 ;
      RECT 37.03 2.89 37.035 3.243 ;
      RECT 37.025 2.892 37.03 3.248 ;
      RECT 37.01 2.902 37.025 3.259 ;
      RECT 36.965 2.96 37.01 3.295 ;
      RECT 36.955 3.015 36.965 3.329 ;
      RECT 36.94 3.042 36.955 3.345 ;
      RECT 36.93 3.069 36.94 3.465 ;
      RECT 36.915 3.092 36.93 3.465 ;
      RECT 36.905 3.132 36.91 3.465 ;
      RECT 36.9 3.142 36.905 3.465 ;
      RECT 36.895 3.157 36.9 3.465 ;
      RECT 36.885 3.162 36.895 3.465 ;
      RECT 36.82 3.185 36.885 3.465 ;
      RECT 36.32 2.68 36.51 2.89 ;
      RECT 34.895 2.605 35.155 2.865 ;
      RECT 35.245 2.6 35.34 2.81 ;
      RECT 35.22 2.615 35.23 2.81 ;
      RECT 36.51 2.687 36.52 2.885 ;
      RECT 36.31 2.687 36.32 2.885 ;
      RECT 36.295 2.702 36.31 2.875 ;
      RECT 36.29 2.71 36.295 2.868 ;
      RECT 36.28 2.713 36.29 2.865 ;
      RECT 36.245 2.712 36.28 2.863 ;
      RECT 36.216 2.708 36.245 2.86 ;
      RECT 36.13 2.703 36.216 2.857 ;
      RECT 36.07 2.697 36.13 2.853 ;
      RECT 36.041 2.693 36.07 2.85 ;
      RECT 35.955 2.685 36.041 2.847 ;
      RECT 35.946 2.679 35.955 2.845 ;
      RECT 35.86 2.674 35.946 2.843 ;
      RECT 35.837 2.669 35.86 2.84 ;
      RECT 35.751 2.663 35.837 2.837 ;
      RECT 35.665 2.654 35.751 2.832 ;
      RECT 35.655 2.649 35.665 2.83 ;
      RECT 35.636 2.648 35.655 2.829 ;
      RECT 35.55 2.643 35.636 2.825 ;
      RECT 35.53 2.638 35.55 2.821 ;
      RECT 35.47 2.633 35.53 2.818 ;
      RECT 35.445 2.623 35.47 2.816 ;
      RECT 35.44 2.616 35.445 2.815 ;
      RECT 35.43 2.607 35.44 2.814 ;
      RECT 35.426 2.6 35.43 2.814 ;
      RECT 35.34 2.6 35.426 2.812 ;
      RECT 35.23 2.607 35.245 2.81 ;
      RECT 35.215 2.617 35.22 2.81 ;
      RECT 35.195 2.62 35.215 2.807 ;
      RECT 35.165 2.62 35.195 2.803 ;
      RECT 35.155 2.62 35.165 2.803 ;
      RECT 36.07 3.115 36.33 3.375 ;
      RECT 36 3.125 36.33 3.335 ;
      RECT 35.99 3.132 36.33 3.33 ;
      RECT 35.41 3.12 35.67 3.38 ;
      RECT 35.41 3.16 35.775 3.37 ;
      RECT 35.41 3.162 35.78 3.369 ;
      RECT 35.41 3.17 35.785 3.366 ;
      RECT 34.335 2.245 34.435 3.77 ;
      RECT 34.525 3.385 34.575 3.645 ;
      RECT 34.52 2.258 34.525 2.445 ;
      RECT 34.515 3.366 34.525 3.645 ;
      RECT 34.515 2.255 34.52 2.453 ;
      RECT 34.5 2.249 34.515 2.46 ;
      RECT 34.51 3.354 34.515 3.728 ;
      RECT 34.5 3.342 34.51 3.765 ;
      RECT 34.49 2.245 34.5 2.467 ;
      RECT 34.49 3.327 34.5 3.77 ;
      RECT 34.485 2.245 34.49 2.475 ;
      RECT 34.465 3.297 34.49 3.77 ;
      RECT 34.445 2.245 34.485 2.523 ;
      RECT 34.455 3.257 34.465 3.77 ;
      RECT 34.445 3.212 34.455 3.77 ;
      RECT 34.44 2.245 34.445 2.593 ;
      RECT 34.44 3.17 34.445 3.77 ;
      RECT 34.435 2.245 34.44 3.07 ;
      RECT 34.435 3.152 34.44 3.77 ;
      RECT 34.325 2.248 34.335 3.77 ;
      RECT 34.31 2.255 34.325 3.766 ;
      RECT 34.305 2.265 34.31 3.761 ;
      RECT 34.3 2.465 34.305 3.653 ;
      RECT 34.295 2.55 34.3 3.205 ;
      RECT 33.175 7.765 33.465 7.995 ;
      RECT 33.235 6.285 33.405 7.995 ;
      RECT 33.22 6.66 33.575 7.015 ;
      RECT 33.175 6.285 33.465 6.515 ;
      RECT 33.175 2.365 33.465 2.595 ;
      RECT 33.235 0.885 33.405 2.595 ;
      RECT 33.175 0.885 33.465 1.115 ;
      RECT 32.765 2.735 33.095 2.965 ;
      RECT 32.765 2.765 33.265 2.935 ;
      RECT 32.765 2.395 32.955 2.965 ;
      RECT 32.185 2.365 32.475 2.595 ;
      RECT 32.185 2.395 32.955 2.565 ;
      RECT 32.245 0.885 32.415 2.595 ;
      RECT 32.185 0.885 32.475 1.115 ;
      RECT 32.185 7.765 32.475 7.995 ;
      RECT 32.245 6.285 32.415 7.995 ;
      RECT 32.185 6.285 32.475 6.515 ;
      RECT 32.185 6.325 33.035 6.485 ;
      RECT 32.865 5.915 33.035 6.485 ;
      RECT 32.185 6.32 32.575 6.485 ;
      RECT 32.805 5.915 33.095 6.145 ;
      RECT 32.805 5.945 33.265 6.115 ;
      RECT 31.815 2.735 32.105 2.965 ;
      RECT 31.815 2.765 32.275 2.935 ;
      RECT 31.875 1.655 32.04 2.965 ;
      RECT 30.39 1.625 30.68 1.855 ;
      RECT 30.39 1.655 32.04 1.825 ;
      RECT 30.45 0.885 30.62 1.855 ;
      RECT 30.39 0.885 30.68 1.115 ;
      RECT 30.39 7.765 30.68 7.995 ;
      RECT 30.45 7.025 30.62 7.995 ;
      RECT 30.45 7.12 32.04 7.29 ;
      RECT 31.87 5.915 32.04 7.29 ;
      RECT 30.39 7.025 30.68 7.255 ;
      RECT 31.815 5.915 32.105 6.145 ;
      RECT 31.815 5.945 32.275 6.115 ;
      RECT 28.425 3.43 28.775 3.78 ;
      RECT 28.515 2.025 28.685 3.78 ;
      RECT 30.82 1.965 31.17 2.315 ;
      RECT 28.515 2.025 30.135 2.2 ;
      RECT 28.515 2.025 31.17 2.195 ;
      RECT 30.845 6.655 31.17 6.98 ;
      RECT 26.27 6.61 26.62 6.96 ;
      RECT 30.82 6.655 31.17 6.885 ;
      RECT 26.06 6.655 26.62 6.885 ;
      RECT 25.89 6.685 31.17 6.855 ;
      RECT 30.045 2.365 30.365 2.685 ;
      RECT 30.015 2.365 30.365 2.595 ;
      RECT 29.845 2.395 30.365 2.565 ;
      RECT 30.045 6.225 30.365 6.545 ;
      RECT 30.015 6.285 30.365 6.515 ;
      RECT 29.845 6.315 30.365 6.485 ;
      RECT 29 2.705 29.35 3.055 ;
      RECT 29 2.765 29.48 2.935 ;
      RECT 28.99 5.84 29.34 6.19 ;
      RECT 24.26 5.915 24.55 6.145 ;
      RECT 24.26 5.945 29.48 6.115 ;
      RECT 25.825 3.665 25.865 3.925 ;
      RECT 25.865 3.645 25.87 3.655 ;
      RECT 27.195 2.89 27.205 3.111 ;
      RECT 27.125 2.885 27.195 3.236 ;
      RECT 27.115 2.885 27.125 3.363 ;
      RECT 27.09 2.885 27.115 3.41 ;
      RECT 27.065 2.885 27.09 3.488 ;
      RECT 27.045 2.885 27.065 3.558 ;
      RECT 27.02 2.885 27.045 3.598 ;
      RECT 27.01 2.885 27.02 3.618 ;
      RECT 27 2.887 27.01 3.626 ;
      RECT 26.995 2.892 27 3.083 ;
      RECT 26.995 3.092 27 3.627 ;
      RECT 26.99 3.137 26.995 3.628 ;
      RECT 26.98 3.202 26.99 3.629 ;
      RECT 26.97 3.297 26.98 3.631 ;
      RECT 26.965 3.35 26.97 3.633 ;
      RECT 26.96 3.37 26.965 3.634 ;
      RECT 26.905 3.395 26.96 3.64 ;
      RECT 26.865 3.43 26.905 3.649 ;
      RECT 26.855 3.447 26.865 3.654 ;
      RECT 26.846 3.453 26.855 3.656 ;
      RECT 26.76 3.491 26.846 3.667 ;
      RECT 26.755 3.53 26.76 3.677 ;
      RECT 26.68 3.537 26.755 3.687 ;
      RECT 26.66 3.547 26.68 3.698 ;
      RECT 26.63 3.554 26.66 3.706 ;
      RECT 26.605 3.561 26.63 3.713 ;
      RECT 26.581 3.567 26.605 3.718 ;
      RECT 26.495 3.58 26.581 3.73 ;
      RECT 26.417 3.587 26.495 3.748 ;
      RECT 26.331 3.582 26.417 3.766 ;
      RECT 26.245 3.577 26.331 3.786 ;
      RECT 26.165 3.571 26.245 3.803 ;
      RECT 26.1 3.567 26.165 3.832 ;
      RECT 26.095 3.281 26.1 3.305 ;
      RECT 26.085 3.557 26.1 3.86 ;
      RECT 26.09 3.275 26.095 3.345 ;
      RECT 26.085 3.269 26.09 3.415 ;
      RECT 26.08 3.263 26.085 3.493 ;
      RECT 26.08 3.54 26.085 3.925 ;
      RECT 26.072 3.26 26.08 3.925 ;
      RECT 25.986 3.258 26.072 3.925 ;
      RECT 25.9 3.256 25.986 3.925 ;
      RECT 25.89 3.257 25.9 3.925 ;
      RECT 25.885 3.262 25.89 3.925 ;
      RECT 25.875 3.275 25.885 3.925 ;
      RECT 25.87 3.297 25.875 3.925 ;
      RECT 25.865 3.657 25.87 3.925 ;
      RECT 26.495 3.125 26.5 3.345 ;
      RECT 27 2.16 27.035 2.42 ;
      RECT 26.985 2.16 27 2.428 ;
      RECT 26.956 2.16 26.985 2.45 ;
      RECT 26.87 2.16 26.956 2.51 ;
      RECT 26.85 2.16 26.87 2.575 ;
      RECT 26.79 2.16 26.85 2.74 ;
      RECT 26.785 2.16 26.79 2.888 ;
      RECT 26.78 2.16 26.785 2.9 ;
      RECT 26.775 2.16 26.78 2.926 ;
      RECT 26.745 2.346 26.775 3.006 ;
      RECT 26.74 2.394 26.745 3.095 ;
      RECT 26.735 2.408 26.74 3.11 ;
      RECT 26.73 2.427 26.735 3.14 ;
      RECT 26.725 2.442 26.73 3.156 ;
      RECT 26.72 2.457 26.725 3.178 ;
      RECT 26.715 2.477 26.72 3.2 ;
      RECT 26.705 2.497 26.715 3.233 ;
      RECT 26.69 2.539 26.705 3.295 ;
      RECT 26.685 2.57 26.69 3.335 ;
      RECT 26.68 2.582 26.685 3.34 ;
      RECT 26.675 2.594 26.68 3.345 ;
      RECT 26.67 2.607 26.675 3.345 ;
      RECT 26.665 2.625 26.67 3.345 ;
      RECT 26.66 2.645 26.665 3.345 ;
      RECT 26.655 2.657 26.66 3.345 ;
      RECT 26.65 2.67 26.655 3.345 ;
      RECT 26.63 2.705 26.65 3.345 ;
      RECT 26.58 2.807 26.63 3.345 ;
      RECT 26.575 2.892 26.58 3.345 ;
      RECT 26.57 2.9 26.575 3.345 ;
      RECT 26.565 2.917 26.57 3.345 ;
      RECT 26.56 2.932 26.565 3.345 ;
      RECT 26.525 2.997 26.56 3.345 ;
      RECT 26.51 3.062 26.525 3.345 ;
      RECT 26.505 3.092 26.51 3.345 ;
      RECT 26.5 3.117 26.505 3.345 ;
      RECT 26.485 3.127 26.495 3.345 ;
      RECT 26.47 3.14 26.485 3.338 ;
      RECT 26.215 2.73 26.285 2.94 ;
      RECT 26.005 2.707 26.01 2.9 ;
      RECT 23.46 2.635 23.72 2.895 ;
      RECT 26.295 2.917 26.3 2.92 ;
      RECT 26.285 2.735 26.295 2.935 ;
      RECT 26.186 2.728 26.215 2.94 ;
      RECT 26.1 2.72 26.186 2.94 ;
      RECT 26.085 2.714 26.1 2.938 ;
      RECT 26.065 2.713 26.085 2.925 ;
      RECT 26.06 2.712 26.065 2.908 ;
      RECT 26.01 2.709 26.06 2.903 ;
      RECT 25.98 2.706 26.005 2.898 ;
      RECT 25.96 2.704 25.98 2.893 ;
      RECT 25.945 2.702 25.96 2.89 ;
      RECT 25.915 2.7 25.945 2.888 ;
      RECT 25.85 2.696 25.915 2.88 ;
      RECT 25.82 2.691 25.85 2.875 ;
      RECT 25.8 2.689 25.82 2.873 ;
      RECT 25.77 2.686 25.8 2.868 ;
      RECT 25.71 2.682 25.77 2.86 ;
      RECT 25.705 2.679 25.71 2.855 ;
      RECT 25.635 2.677 25.705 2.85 ;
      RECT 25.606 2.673 25.635 2.843 ;
      RECT 25.52 2.668 25.606 2.835 ;
      RECT 25.486 2.663 25.52 2.827 ;
      RECT 25.4 2.655 25.486 2.819 ;
      RECT 25.361 2.648 25.4 2.811 ;
      RECT 25.275 2.643 25.361 2.803 ;
      RECT 25.21 2.637 25.275 2.793 ;
      RECT 25.19 2.632 25.21 2.788 ;
      RECT 25.181 2.629 25.19 2.787 ;
      RECT 25.095 2.625 25.181 2.781 ;
      RECT 25.055 2.621 25.095 2.773 ;
      RECT 25.035 2.617 25.055 2.771 ;
      RECT 24.975 2.617 25.035 2.768 ;
      RECT 24.955 2.62 24.975 2.766 ;
      RECT 24.934 2.62 24.955 2.766 ;
      RECT 24.848 2.622 24.934 2.77 ;
      RECT 24.762 2.624 24.848 2.776 ;
      RECT 24.676 2.626 24.762 2.783 ;
      RECT 24.59 2.629 24.676 2.789 ;
      RECT 24.556 2.63 24.59 2.794 ;
      RECT 24.47 2.633 24.556 2.799 ;
      RECT 24.441 2.64 24.47 2.804 ;
      RECT 24.355 2.64 24.441 2.809 ;
      RECT 24.322 2.64 24.355 2.814 ;
      RECT 24.236 2.642 24.322 2.819 ;
      RECT 24.15 2.644 24.236 2.826 ;
      RECT 24.086 2.646 24.15 2.832 ;
      RECT 24 2.648 24.086 2.838 ;
      RECT 23.997 2.65 24 2.841 ;
      RECT 23.911 2.651 23.997 2.845 ;
      RECT 23.825 2.654 23.911 2.852 ;
      RECT 23.806 2.656 23.825 2.856 ;
      RECT 23.72 2.658 23.806 2.861 ;
      RECT 23.45 2.67 23.46 2.865 ;
      RECT 25.63 7.765 25.92 7.995 ;
      RECT 25.69 7.025 25.86 7.995 ;
      RECT 25.58 7.055 25.955 7.425 ;
      RECT 25.63 7.025 25.92 7.425 ;
      RECT 25.685 2.25 25.87 2.46 ;
      RECT 25.68 2.251 25.875 2.458 ;
      RECT 25.675 2.256 25.885 2.453 ;
      RECT 25.67 2.232 25.675 2.45 ;
      RECT 25.64 2.229 25.67 2.443 ;
      RECT 25.635 2.225 25.64 2.434 ;
      RECT 25.6 2.256 25.885 2.429 ;
      RECT 25.375 2.165 25.635 2.425 ;
      RECT 25.675 2.234 25.68 2.453 ;
      RECT 25.68 2.235 25.685 2.458 ;
      RECT 25.375 2.247 25.755 2.425 ;
      RECT 25.375 2.245 25.74 2.425 ;
      RECT 25.375 2.24 25.73 2.425 ;
      RECT 25.33 3.155 25.38 3.44 ;
      RECT 25.275 3.125 25.28 3.44 ;
      RECT 25.245 3.105 25.25 3.44 ;
      RECT 25.395 3.155 25.455 3.415 ;
      RECT 25.39 3.155 25.395 3.423 ;
      RECT 25.38 3.155 25.39 3.435 ;
      RECT 25.295 3.145 25.33 3.44 ;
      RECT 25.29 3.132 25.295 3.44 ;
      RECT 25.28 3.127 25.29 3.44 ;
      RECT 25.26 3.117 25.275 3.44 ;
      RECT 25.25 3.11 25.26 3.44 ;
      RECT 25.24 3.102 25.245 3.44 ;
      RECT 25.21 3.092 25.24 3.44 ;
      RECT 25.195 3.08 25.21 3.44 ;
      RECT 25.18 3.07 25.195 3.435 ;
      RECT 25.16 3.06 25.18 3.41 ;
      RECT 25.15 3.052 25.16 3.387 ;
      RECT 25.12 3.035 25.15 3.377 ;
      RECT 25.115 3.012 25.12 3.368 ;
      RECT 25.11 2.999 25.115 3.366 ;
      RECT 25.095 2.975 25.11 3.36 ;
      RECT 25.09 2.951 25.095 3.354 ;
      RECT 25.08 2.94 25.09 3.349 ;
      RECT 25.075 2.93 25.08 3.345 ;
      RECT 25.07 2.922 25.075 3.342 ;
      RECT 25.06 2.917 25.07 3.338 ;
      RECT 25.055 2.912 25.06 3.334 ;
      RECT 24.97 2.91 25.055 3.309 ;
      RECT 24.94 2.91 24.97 3.275 ;
      RECT 24.925 2.91 24.94 3.258 ;
      RECT 24.87 2.91 24.925 3.203 ;
      RECT 24.865 2.915 24.87 3.152 ;
      RECT 24.855 2.92 24.865 3.142 ;
      RECT 24.85 2.93 24.855 3.128 ;
      RECT 24.8 3.67 25.06 3.93 ;
      RECT 24.72 3.685 25.06 3.906 ;
      RECT 24.7 3.685 25.06 3.901 ;
      RECT 24.676 3.685 25.06 3.899 ;
      RECT 24.59 3.685 25.06 3.894 ;
      RECT 24.44 3.625 24.7 3.89 ;
      RECT 24.395 3.685 25.06 3.885 ;
      RECT 24.39 3.692 25.06 3.88 ;
      RECT 24.405 3.68 24.72 3.89 ;
      RECT 24.295 2.115 24.555 2.375 ;
      RECT 24.295 2.172 24.56 2.368 ;
      RECT 24.295 2.202 24.565 2.3 ;
      RECT 24.355 2.633 24.47 2.635 ;
      RECT 24.441 2.63 24.47 2.635 ;
      RECT 23.465 3.634 23.49 3.874 ;
      RECT 23.45 3.637 23.54 3.868 ;
      RECT 23.445 3.642 23.626 3.863 ;
      RECT 23.44 3.65 23.69 3.861 ;
      RECT 23.44 3.65 23.7 3.86 ;
      RECT 23.435 3.657 23.71 3.853 ;
      RECT 23.435 3.657 23.796 3.842 ;
      RECT 23.43 3.692 23.796 3.838 ;
      RECT 23.43 3.692 23.805 3.827 ;
      RECT 23.71 3.565 23.97 3.825 ;
      RECT 23.42 3.742 23.97 3.823 ;
      RECT 23.69 3.61 23.71 3.858 ;
      RECT 23.626 3.613 23.69 3.862 ;
      RECT 23.54 3.618 23.626 3.867 ;
      RECT 23.47 3.629 23.97 3.825 ;
      RECT 23.49 3.623 23.54 3.872 ;
      RECT 23.615 2.1 23.625 2.362 ;
      RECT 23.605 2.157 23.615 2.365 ;
      RECT 23.58 2.162 23.605 2.371 ;
      RECT 23.555 2.166 23.58 2.383 ;
      RECT 23.545 2.169 23.555 2.393 ;
      RECT 23.54 2.17 23.545 2.398 ;
      RECT 23.535 2.171 23.54 2.403 ;
      RECT 23.53 2.172 23.535 2.405 ;
      RECT 23.505 2.175 23.53 2.408 ;
      RECT 23.475 2.181 23.505 2.411 ;
      RECT 23.41 2.192 23.475 2.414 ;
      RECT 23.365 2.2 23.41 2.418 ;
      RECT 23.35 2.2 23.365 2.426 ;
      RECT 23.345 2.201 23.35 2.433 ;
      RECT 23.34 2.203 23.345 2.436 ;
      RECT 23.335 2.207 23.34 2.439 ;
      RECT 23.325 2.215 23.335 2.443 ;
      RECT 23.32 2.228 23.325 2.448 ;
      RECT 23.315 2.236 23.32 2.45 ;
      RECT 23.31 2.242 23.315 2.45 ;
      RECT 23.305 2.246 23.31 2.453 ;
      RECT 23.3 2.248 23.305 2.456 ;
      RECT 23.295 2.251 23.3 2.459 ;
      RECT 23.285 2.256 23.295 2.463 ;
      RECT 23.28 2.262 23.285 2.468 ;
      RECT 23.27 2.268 23.28 2.472 ;
      RECT 23.255 2.275 23.27 2.478 ;
      RECT 23.226 2.289 23.255 2.488 ;
      RECT 23.14 2.324 23.226 2.52 ;
      RECT 23.12 2.357 23.14 2.549 ;
      RECT 23.1 2.37 23.12 2.56 ;
      RECT 23.08 2.382 23.1 2.571 ;
      RECT 23.03 2.404 23.08 2.591 ;
      RECT 23.015 2.422 23.03 2.608 ;
      RECT 23.01 2.428 23.015 2.611 ;
      RECT 23.005 2.432 23.01 2.614 ;
      RECT 23 2.436 23.005 2.618 ;
      RECT 22.995 2.438 23 2.621 ;
      RECT 22.985 2.445 22.995 2.624 ;
      RECT 22.98 2.45 22.985 2.628 ;
      RECT 22.975 2.452 22.98 2.631 ;
      RECT 22.97 2.456 22.975 2.634 ;
      RECT 22.965 2.458 22.97 2.638 ;
      RECT 22.95 2.463 22.965 2.643 ;
      RECT 22.945 2.468 22.95 2.646 ;
      RECT 22.94 2.476 22.945 2.649 ;
      RECT 22.935 2.478 22.94 2.652 ;
      RECT 22.93 2.48 22.935 2.655 ;
      RECT 22.92 2.482 22.93 2.661 ;
      RECT 22.885 2.496 22.92 2.673 ;
      RECT 22.875 2.511 22.885 2.683 ;
      RECT 22.8 2.54 22.875 2.707 ;
      RECT 22.795 2.565 22.8 2.73 ;
      RECT 22.78 2.569 22.795 2.736 ;
      RECT 22.77 2.577 22.78 2.741 ;
      RECT 22.74 2.59 22.77 2.745 ;
      RECT 22.73 2.605 22.74 2.75 ;
      RECT 22.72 2.61 22.73 2.753 ;
      RECT 22.715 2.612 22.72 2.755 ;
      RECT 22.7 2.615 22.715 2.758 ;
      RECT 22.695 2.617 22.7 2.761 ;
      RECT 22.675 2.622 22.695 2.765 ;
      RECT 22.645 2.627 22.675 2.773 ;
      RECT 22.62 2.634 22.645 2.781 ;
      RECT 22.615 2.639 22.62 2.786 ;
      RECT 22.585 2.642 22.615 2.79 ;
      RECT 22.545 2.645 22.585 2.8 ;
      RECT 22.51 2.642 22.545 2.812 ;
      RECT 22.5 2.638 22.51 2.819 ;
      RECT 22.475 2.634 22.5 2.825 ;
      RECT 22.47 2.63 22.475 2.83 ;
      RECT 22.43 2.627 22.47 2.83 ;
      RECT 22.415 2.612 22.43 2.831 ;
      RECT 22.392 2.6 22.415 2.831 ;
      RECT 22.306 2.6 22.392 2.832 ;
      RECT 22.22 2.6 22.306 2.834 ;
      RECT 22.2 2.6 22.22 2.831 ;
      RECT 22.195 2.605 22.2 2.826 ;
      RECT 22.19 2.61 22.195 2.824 ;
      RECT 22.18 2.62 22.19 2.822 ;
      RECT 22.175 2.626 22.18 2.815 ;
      RECT 22.17 2.628 22.175 2.8 ;
      RECT 22.165 2.632 22.17 2.79 ;
      RECT 23.625 2.1 23.875 2.36 ;
      RECT 21.35 3.635 21.61 3.895 ;
      RECT 23.645 3.125 23.65 3.335 ;
      RECT 23.65 3.13 23.66 3.33 ;
      RECT 23.6 3.125 23.645 3.35 ;
      RECT 23.59 3.125 23.6 3.37 ;
      RECT 23.571 3.125 23.59 3.375 ;
      RECT 23.485 3.125 23.571 3.372 ;
      RECT 23.455 3.127 23.485 3.37 ;
      RECT 23.4 3.137 23.455 3.368 ;
      RECT 23.335 3.151 23.4 3.366 ;
      RECT 23.33 3.159 23.335 3.365 ;
      RECT 23.315 3.162 23.33 3.363 ;
      RECT 23.25 3.172 23.315 3.359 ;
      RECT 23.202 3.186 23.25 3.36 ;
      RECT 23.116 3.203 23.202 3.374 ;
      RECT 23.03 3.224 23.116 3.391 ;
      RECT 23.01 3.237 23.03 3.401 ;
      RECT 22.965 3.245 23.01 3.408 ;
      RECT 22.93 3.253 22.965 3.416 ;
      RECT 22.896 3.261 22.93 3.424 ;
      RECT 22.81 3.275 22.896 3.436 ;
      RECT 22.775 3.292 22.81 3.448 ;
      RECT 22.766 3.301 22.775 3.452 ;
      RECT 22.68 3.319 22.766 3.469 ;
      RECT 22.621 3.346 22.68 3.496 ;
      RECT 22.535 3.373 22.621 3.524 ;
      RECT 22.515 3.395 22.535 3.544 ;
      RECT 22.455 3.41 22.515 3.56 ;
      RECT 22.445 3.422 22.455 3.573 ;
      RECT 22.44 3.427 22.445 3.576 ;
      RECT 22.43 3.43 22.44 3.579 ;
      RECT 22.425 3.432 22.43 3.582 ;
      RECT 22.395 3.44 22.425 3.589 ;
      RECT 22.38 3.447 22.395 3.597 ;
      RECT 22.37 3.452 22.38 3.601 ;
      RECT 22.365 3.455 22.37 3.604 ;
      RECT 22.355 3.457 22.365 3.607 ;
      RECT 22.32 3.467 22.355 3.616 ;
      RECT 22.245 3.49 22.32 3.638 ;
      RECT 22.225 3.508 22.245 3.656 ;
      RECT 22.195 3.515 22.225 3.666 ;
      RECT 22.175 3.523 22.195 3.676 ;
      RECT 22.165 3.529 22.175 3.683 ;
      RECT 22.146 3.534 22.165 3.689 ;
      RECT 22.06 3.554 22.146 3.709 ;
      RECT 22.045 3.574 22.06 3.728 ;
      RECT 22 3.586 22.045 3.739 ;
      RECT 21.935 3.607 22 3.762 ;
      RECT 21.895 3.627 21.935 3.783 ;
      RECT 21.885 3.637 21.895 3.793 ;
      RECT 21.835 3.649 21.885 3.804 ;
      RECT 21.815 3.665 21.835 3.816 ;
      RECT 21.785 3.675 21.815 3.822 ;
      RECT 21.775 3.68 21.785 3.824 ;
      RECT 21.706 3.681 21.775 3.83 ;
      RECT 21.62 3.683 21.706 3.84 ;
      RECT 21.61 3.684 21.62 3.845 ;
      RECT 22.88 3.71 23.07 3.92 ;
      RECT 22.87 3.715 23.08 3.913 ;
      RECT 22.855 3.715 23.08 3.878 ;
      RECT 22.775 3.6 23.035 3.86 ;
      RECT 21.69 3.13 21.875 3.425 ;
      RECT 21.68 3.13 21.875 3.423 ;
      RECT 21.665 3.13 21.88 3.418 ;
      RECT 21.665 3.13 21.885 3.415 ;
      RECT 21.66 3.13 21.885 3.413 ;
      RECT 21.655 3.385 21.885 3.403 ;
      RECT 21.66 3.13 21.92 3.39 ;
      RECT 21.62 2.165 21.88 2.425 ;
      RECT 21.43 2.09 21.516 2.423 ;
      RECT 21.405 2.094 21.56 2.419 ;
      RECT 21.516 2.086 21.56 2.419 ;
      RECT 21.516 2.087 21.565 2.418 ;
      RECT 21.43 2.092 21.58 2.417 ;
      RECT 21.405 2.1 21.62 2.416 ;
      RECT 21.4 2.095 21.58 2.411 ;
      RECT 21.39 2.11 21.62 2.318 ;
      RECT 21.39 2.162 21.82 2.318 ;
      RECT 21.39 2.155 21.8 2.318 ;
      RECT 21.39 2.142 21.77 2.318 ;
      RECT 21.39 2.13 21.71 2.318 ;
      RECT 21.39 2.115 21.685 2.318 ;
      RECT 20.59 2.745 20.725 3.04 ;
      RECT 20.85 2.768 20.855 2.955 ;
      RECT 21.57 2.665 21.715 2.9 ;
      RECT 21.73 2.665 21.735 2.89 ;
      RECT 21.765 2.676 21.77 2.87 ;
      RECT 21.76 2.668 21.765 2.875 ;
      RECT 21.74 2.665 21.76 2.88 ;
      RECT 21.735 2.665 21.74 2.888 ;
      RECT 21.725 2.665 21.73 2.893 ;
      RECT 21.715 2.665 21.725 2.898 ;
      RECT 21.545 2.667 21.57 2.9 ;
      RECT 21.495 2.674 21.545 2.9 ;
      RECT 21.49 2.679 21.495 2.9 ;
      RECT 21.451 2.684 21.49 2.901 ;
      RECT 21.365 2.696 21.451 2.902 ;
      RECT 21.356 2.706 21.365 2.902 ;
      RECT 21.27 2.715 21.356 2.904 ;
      RECT 21.246 2.725 21.27 2.906 ;
      RECT 21.16 2.736 21.246 2.907 ;
      RECT 21.13 2.747 21.16 2.909 ;
      RECT 21.1 2.752 21.13 2.911 ;
      RECT 21.075 2.758 21.1 2.914 ;
      RECT 21.06 2.763 21.075 2.915 ;
      RECT 21.015 2.769 21.06 2.915 ;
      RECT 21.01 2.774 21.015 2.916 ;
      RECT 20.99 2.774 21.01 2.918 ;
      RECT 20.97 2.772 20.99 2.923 ;
      RECT 20.935 2.771 20.97 2.93 ;
      RECT 20.905 2.77 20.935 2.94 ;
      RECT 20.855 2.769 20.905 2.95 ;
      RECT 20.765 2.766 20.85 3.04 ;
      RECT 20.74 2.76 20.765 3.04 ;
      RECT 20.725 2.75 20.74 3.04 ;
      RECT 20.54 2.745 20.59 2.96 ;
      RECT 20.53 2.75 20.54 2.95 ;
      RECT 20.77 3.225 21.03 3.485 ;
      RECT 20.77 3.225 21.06 3.378 ;
      RECT 20.77 3.225 21.095 3.363 ;
      RECT 21.025 3.145 21.215 3.355 ;
      RECT 21.015 3.15 21.225 3.348 ;
      RECT 20.98 3.22 21.225 3.348 ;
      RECT 21.01 3.162 21.03 3.485 ;
      RECT 20.995 3.21 21.225 3.348 ;
      RECT 21 3.182 21.03 3.485 ;
      RECT 20.08 2.25 20.15 3.355 ;
      RECT 20.815 2.355 21.075 2.615 ;
      RECT 20.395 2.401 20.41 2.61 ;
      RECT 20.731 2.414 20.815 2.565 ;
      RECT 20.645 2.411 20.731 2.565 ;
      RECT 20.606 2.409 20.645 2.565 ;
      RECT 20.52 2.407 20.606 2.565 ;
      RECT 20.46 2.405 20.52 2.576 ;
      RECT 20.425 2.403 20.46 2.594 ;
      RECT 20.41 2.401 20.425 2.605 ;
      RECT 20.38 2.401 20.395 2.618 ;
      RECT 20.37 2.401 20.38 2.623 ;
      RECT 20.345 2.4 20.37 2.628 ;
      RECT 20.33 2.395 20.345 2.634 ;
      RECT 20.325 2.388 20.33 2.639 ;
      RECT 20.3 2.379 20.325 2.645 ;
      RECT 20.255 2.358 20.3 2.658 ;
      RECT 20.245 2.342 20.255 2.668 ;
      RECT 20.23 2.335 20.245 2.678 ;
      RECT 20.22 2.328 20.23 2.695 ;
      RECT 20.215 2.325 20.22 2.725 ;
      RECT 20.21 2.323 20.215 2.755 ;
      RECT 20.205 2.321 20.21 2.792 ;
      RECT 20.19 2.317 20.205 2.859 ;
      RECT 20.19 3.15 20.2 3.35 ;
      RECT 20.185 2.313 20.19 2.985 ;
      RECT 20.185 3.137 20.19 3.355 ;
      RECT 20.18 2.311 20.185 3.07 ;
      RECT 20.18 3.127 20.185 3.355 ;
      RECT 20.165 2.282 20.18 3.355 ;
      RECT 20.15 2.255 20.165 3.355 ;
      RECT 20.075 2.25 20.08 2.605 ;
      RECT 20.075 2.66 20.08 3.355 ;
      RECT 20.06 2.25 20.075 2.583 ;
      RECT 20.07 2.682 20.075 3.355 ;
      RECT 20.06 2.722 20.07 3.355 ;
      RECT 20.025 2.25 20.06 2.525 ;
      RECT 20.055 2.757 20.06 3.355 ;
      RECT 20.04 2.812 20.055 3.355 ;
      RECT 20.035 2.877 20.04 3.355 ;
      RECT 20.02 2.925 20.035 3.355 ;
      RECT 19.995 2.25 20.025 2.48 ;
      RECT 20.015 2.98 20.02 3.355 ;
      RECT 20 3.04 20.015 3.355 ;
      RECT 19.995 3.088 20 3.353 ;
      RECT 19.99 2.25 19.995 2.473 ;
      RECT 19.99 3.12 19.995 3.348 ;
      RECT 19.965 2.25 19.99 2.465 ;
      RECT 19.955 2.255 19.965 2.455 ;
      RECT 20.17 3.53 20.19 3.77 ;
      RECT 19.4 3.46 19.405 3.67 ;
      RECT 20.68 3.533 20.69 3.728 ;
      RECT 20.675 3.523 20.68 3.731 ;
      RECT 20.595 3.52 20.675 3.754 ;
      RECT 20.591 3.52 20.595 3.776 ;
      RECT 20.505 3.52 20.591 3.786 ;
      RECT 20.49 3.52 20.505 3.794 ;
      RECT 20.461 3.521 20.49 3.792 ;
      RECT 20.375 3.526 20.461 3.788 ;
      RECT 20.362 3.53 20.375 3.784 ;
      RECT 20.276 3.53 20.362 3.78 ;
      RECT 20.19 3.53 20.276 3.774 ;
      RECT 20.106 3.53 20.17 3.768 ;
      RECT 20.02 3.53 20.106 3.763 ;
      RECT 20 3.53 20.02 3.759 ;
      RECT 19.94 3.525 20 3.756 ;
      RECT 19.912 3.519 19.94 3.753 ;
      RECT 19.826 3.514 19.912 3.749 ;
      RECT 19.74 3.508 19.826 3.743 ;
      RECT 19.665 3.49 19.74 3.738 ;
      RECT 19.63 3.467 19.665 3.734 ;
      RECT 19.62 3.457 19.63 3.733 ;
      RECT 19.565 3.455 19.62 3.732 ;
      RECT 19.49 3.455 19.565 3.728 ;
      RECT 19.48 3.455 19.49 3.723 ;
      RECT 19.465 3.455 19.48 3.715 ;
      RECT 19.415 3.457 19.465 3.693 ;
      RECT 19.405 3.46 19.415 3.673 ;
      RECT 19.395 3.465 19.4 3.668 ;
      RECT 19.39 3.47 19.395 3.663 ;
      RECT 19.515 2.635 19.775 2.895 ;
      RECT 19.515 2.65 19.795 2.86 ;
      RECT 19.515 2.655 19.805 2.855 ;
      RECT 17.5 2.115 17.76 2.375 ;
      RECT 17.49 2.145 17.76 2.355 ;
      RECT 19.41 2.06 19.67 2.32 ;
      RECT 19.405 2.135 19.41 2.321 ;
      RECT 19.38 2.14 19.405 2.323 ;
      RECT 19.365 2.147 19.38 2.326 ;
      RECT 19.305 2.165 19.365 2.331 ;
      RECT 19.275 2.185 19.305 2.338 ;
      RECT 19.25 2.193 19.275 2.343 ;
      RECT 19.225 2.201 19.25 2.345 ;
      RECT 19.207 2.205 19.225 2.344 ;
      RECT 19.121 2.203 19.207 2.344 ;
      RECT 19.035 2.201 19.121 2.344 ;
      RECT 18.949 2.199 19.035 2.343 ;
      RECT 18.863 2.197 18.949 2.343 ;
      RECT 18.777 2.195 18.863 2.343 ;
      RECT 18.691 2.193 18.777 2.343 ;
      RECT 18.605 2.191 18.691 2.342 ;
      RECT 18.587 2.19 18.605 2.342 ;
      RECT 18.501 2.189 18.587 2.342 ;
      RECT 18.415 2.187 18.501 2.342 ;
      RECT 18.329 2.186 18.415 2.341 ;
      RECT 18.243 2.185 18.329 2.341 ;
      RECT 18.157 2.183 18.243 2.341 ;
      RECT 18.071 2.182 18.157 2.341 ;
      RECT 17.985 2.18 18.071 2.34 ;
      RECT 17.961 2.178 17.985 2.34 ;
      RECT 17.875 2.171 17.961 2.34 ;
      RECT 17.846 2.163 17.875 2.34 ;
      RECT 17.76 2.155 17.846 2.34 ;
      RECT 17.48 2.152 17.49 2.35 ;
      RECT 18.985 3.115 18.99 3.465 ;
      RECT 18.755 3.205 18.895 3.465 ;
      RECT 19.23 2.89 19.275 3.1 ;
      RECT 19.285 2.901 19.295 3.095 ;
      RECT 19.275 2.893 19.285 3.1 ;
      RECT 19.21 2.89 19.23 3.105 ;
      RECT 19.18 2.89 19.21 3.128 ;
      RECT 19.17 2.89 19.18 3.153 ;
      RECT 19.165 2.89 19.17 3.163 ;
      RECT 19.11 2.89 19.165 3.203 ;
      RECT 19.105 2.89 19.11 3.243 ;
      RECT 19.1 2.892 19.105 3.248 ;
      RECT 19.085 2.902 19.1 3.259 ;
      RECT 19.04 2.96 19.085 3.295 ;
      RECT 19.03 3.015 19.04 3.329 ;
      RECT 19.015 3.042 19.03 3.345 ;
      RECT 19.005 3.069 19.015 3.465 ;
      RECT 18.99 3.092 19.005 3.465 ;
      RECT 18.98 3.132 18.985 3.465 ;
      RECT 18.975 3.142 18.98 3.465 ;
      RECT 18.97 3.157 18.975 3.465 ;
      RECT 18.96 3.162 18.97 3.465 ;
      RECT 18.895 3.185 18.96 3.465 ;
      RECT 18.395 2.68 18.585 2.89 ;
      RECT 16.97 2.605 17.23 2.865 ;
      RECT 17.32 2.6 17.415 2.81 ;
      RECT 17.295 2.615 17.305 2.81 ;
      RECT 18.585 2.687 18.595 2.885 ;
      RECT 18.385 2.687 18.395 2.885 ;
      RECT 18.37 2.702 18.385 2.875 ;
      RECT 18.365 2.71 18.37 2.868 ;
      RECT 18.355 2.713 18.365 2.865 ;
      RECT 18.32 2.712 18.355 2.863 ;
      RECT 18.291 2.708 18.32 2.86 ;
      RECT 18.205 2.703 18.291 2.857 ;
      RECT 18.145 2.697 18.205 2.853 ;
      RECT 18.116 2.693 18.145 2.85 ;
      RECT 18.03 2.685 18.116 2.847 ;
      RECT 18.021 2.679 18.03 2.845 ;
      RECT 17.935 2.674 18.021 2.843 ;
      RECT 17.912 2.669 17.935 2.84 ;
      RECT 17.826 2.663 17.912 2.837 ;
      RECT 17.74 2.654 17.826 2.832 ;
      RECT 17.73 2.649 17.74 2.83 ;
      RECT 17.711 2.648 17.73 2.829 ;
      RECT 17.625 2.643 17.711 2.825 ;
      RECT 17.605 2.638 17.625 2.821 ;
      RECT 17.545 2.633 17.605 2.818 ;
      RECT 17.52 2.623 17.545 2.816 ;
      RECT 17.515 2.616 17.52 2.815 ;
      RECT 17.505 2.607 17.515 2.814 ;
      RECT 17.501 2.6 17.505 2.814 ;
      RECT 17.415 2.6 17.501 2.812 ;
      RECT 17.305 2.607 17.32 2.81 ;
      RECT 17.29 2.617 17.295 2.81 ;
      RECT 17.27 2.62 17.29 2.807 ;
      RECT 17.24 2.62 17.27 2.803 ;
      RECT 17.23 2.62 17.24 2.803 ;
      RECT 18.145 3.115 18.405 3.375 ;
      RECT 18.075 3.125 18.405 3.335 ;
      RECT 18.065 3.132 18.405 3.33 ;
      RECT 17.485 3.12 17.745 3.38 ;
      RECT 17.485 3.16 17.85 3.37 ;
      RECT 17.485 3.162 17.855 3.369 ;
      RECT 17.485 3.17 17.86 3.366 ;
      RECT 16.41 2.245 16.51 3.77 ;
      RECT 16.6 3.385 16.65 3.645 ;
      RECT 16.595 2.258 16.6 2.445 ;
      RECT 16.59 3.366 16.6 3.645 ;
      RECT 16.59 2.255 16.595 2.453 ;
      RECT 16.575 2.249 16.59 2.46 ;
      RECT 16.585 3.354 16.59 3.728 ;
      RECT 16.575 3.342 16.585 3.765 ;
      RECT 16.565 2.245 16.575 2.467 ;
      RECT 16.565 3.327 16.575 3.77 ;
      RECT 16.56 2.245 16.565 2.475 ;
      RECT 16.54 3.297 16.565 3.77 ;
      RECT 16.52 2.245 16.56 2.523 ;
      RECT 16.53 3.257 16.54 3.77 ;
      RECT 16.52 3.212 16.53 3.77 ;
      RECT 16.515 2.245 16.52 2.593 ;
      RECT 16.515 3.17 16.52 3.77 ;
      RECT 16.51 2.245 16.515 3.07 ;
      RECT 16.51 3.152 16.515 3.77 ;
      RECT 16.4 2.248 16.41 3.77 ;
      RECT 16.385 2.255 16.4 3.766 ;
      RECT 16.38 2.265 16.385 3.761 ;
      RECT 16.375 2.465 16.38 3.653 ;
      RECT 16.37 2.55 16.375 3.205 ;
      RECT 15.25 7.765 15.54 7.995 ;
      RECT 15.31 6.285 15.48 7.995 ;
      RECT 15.3 6.655 15.65 7.005 ;
      RECT 15.25 6.285 15.54 6.515 ;
      RECT 15.25 2.365 15.54 2.595 ;
      RECT 15.31 0.885 15.48 2.595 ;
      RECT 15.25 0.885 15.54 1.115 ;
      RECT 14.84 2.735 15.17 2.965 ;
      RECT 14.84 2.765 15.34 2.935 ;
      RECT 14.84 2.395 15.03 2.965 ;
      RECT 14.26 2.365 14.55 2.595 ;
      RECT 14.26 2.395 15.03 2.565 ;
      RECT 14.32 0.885 14.49 2.595 ;
      RECT 14.26 0.885 14.55 1.115 ;
      RECT 14.26 7.765 14.55 7.995 ;
      RECT 14.32 6.285 14.49 7.995 ;
      RECT 14.26 6.285 14.55 6.515 ;
      RECT 14.26 6.325 15.11 6.485 ;
      RECT 14.94 5.915 15.11 6.485 ;
      RECT 14.26 6.32 14.65 6.485 ;
      RECT 14.88 5.915 15.17 6.145 ;
      RECT 14.88 5.945 15.34 6.115 ;
      RECT 13.89 2.735 14.18 2.965 ;
      RECT 13.89 2.765 14.35 2.935 ;
      RECT 13.95 1.655 14.115 2.965 ;
      RECT 12.465 1.625 12.755 1.855 ;
      RECT 12.465 1.655 14.115 1.825 ;
      RECT 12.525 0.885 12.695 1.855 ;
      RECT 12.465 0.885 12.755 1.115 ;
      RECT 12.465 7.765 12.755 7.995 ;
      RECT 12.525 7.025 12.695 7.995 ;
      RECT 12.525 7.12 14.115 7.29 ;
      RECT 13.945 5.915 14.115 7.29 ;
      RECT 12.465 7.025 12.755 7.255 ;
      RECT 13.89 5.915 14.18 6.145 ;
      RECT 13.89 5.945 14.35 6.115 ;
      RECT 10.5 3.43 10.85 3.78 ;
      RECT 10.59 2.025 10.76 3.78 ;
      RECT 12.895 1.965 13.245 2.315 ;
      RECT 10.59 2.025 12.21 2.2 ;
      RECT 10.59 2.025 13.245 2.195 ;
      RECT 12.92 6.655 13.245 6.98 ;
      RECT 8.315 6.605 8.665 6.955 ;
      RECT 12.895 6.655 13.245 6.885 ;
      RECT 8.135 6.655 8.665 6.885 ;
      RECT 7.965 6.685 13.245 6.855 ;
      RECT 12.12 2.365 12.44 2.685 ;
      RECT 12.09 2.365 12.44 2.595 ;
      RECT 11.92 2.395 12.44 2.565 ;
      RECT 12.12 6.225 12.44 6.545 ;
      RECT 12.09 6.285 12.44 6.515 ;
      RECT 11.92 6.315 12.44 6.485 ;
      RECT 11.075 2.705 11.425 3.055 ;
      RECT 11.075 2.765 11.555 2.935 ;
      RECT 11.065 5.84 11.415 6.19 ;
      RECT 6.335 5.915 6.625 6.145 ;
      RECT 6.335 5.945 11.555 6.115 ;
      RECT 7.9 3.665 7.94 3.925 ;
      RECT 7.94 3.645 7.945 3.655 ;
      RECT 9.27 2.89 9.28 3.111 ;
      RECT 9.2 2.885 9.27 3.236 ;
      RECT 9.19 2.885 9.2 3.363 ;
      RECT 9.165 2.885 9.19 3.41 ;
      RECT 9.14 2.885 9.165 3.488 ;
      RECT 9.12 2.885 9.14 3.558 ;
      RECT 9.095 2.885 9.12 3.598 ;
      RECT 9.085 2.885 9.095 3.618 ;
      RECT 9.075 2.887 9.085 3.626 ;
      RECT 9.07 2.892 9.075 3.083 ;
      RECT 9.07 3.092 9.075 3.627 ;
      RECT 9.065 3.137 9.07 3.628 ;
      RECT 9.055 3.202 9.065 3.629 ;
      RECT 9.045 3.297 9.055 3.631 ;
      RECT 9.04 3.35 9.045 3.633 ;
      RECT 9.035 3.37 9.04 3.634 ;
      RECT 8.98 3.395 9.035 3.64 ;
      RECT 8.94 3.43 8.98 3.649 ;
      RECT 8.93 3.447 8.94 3.654 ;
      RECT 8.921 3.453 8.93 3.656 ;
      RECT 8.835 3.491 8.921 3.667 ;
      RECT 8.83 3.53 8.835 3.677 ;
      RECT 8.755 3.537 8.83 3.687 ;
      RECT 8.735 3.547 8.755 3.698 ;
      RECT 8.705 3.554 8.735 3.706 ;
      RECT 8.68 3.561 8.705 3.713 ;
      RECT 8.656 3.567 8.68 3.718 ;
      RECT 8.57 3.58 8.656 3.73 ;
      RECT 8.492 3.587 8.57 3.748 ;
      RECT 8.406 3.582 8.492 3.766 ;
      RECT 8.32 3.577 8.406 3.786 ;
      RECT 8.24 3.571 8.32 3.803 ;
      RECT 8.175 3.567 8.24 3.832 ;
      RECT 8.17 3.281 8.175 3.305 ;
      RECT 8.16 3.557 8.175 3.86 ;
      RECT 8.165 3.275 8.17 3.345 ;
      RECT 8.16 3.269 8.165 3.415 ;
      RECT 8.155 3.263 8.16 3.493 ;
      RECT 8.155 3.54 8.16 3.925 ;
      RECT 8.147 3.26 8.155 3.925 ;
      RECT 8.061 3.258 8.147 3.925 ;
      RECT 7.975 3.256 8.061 3.925 ;
      RECT 7.965 3.257 7.975 3.925 ;
      RECT 7.96 3.262 7.965 3.925 ;
      RECT 7.95 3.275 7.96 3.925 ;
      RECT 7.945 3.297 7.95 3.925 ;
      RECT 7.94 3.657 7.945 3.925 ;
      RECT 8.57 3.125 8.575 3.345 ;
      RECT 9.075 2.16 9.11 2.42 ;
      RECT 9.06 2.16 9.075 2.428 ;
      RECT 9.031 2.16 9.06 2.45 ;
      RECT 8.945 2.16 9.031 2.51 ;
      RECT 8.925 2.16 8.945 2.575 ;
      RECT 8.865 2.16 8.925 2.74 ;
      RECT 8.86 2.16 8.865 2.888 ;
      RECT 8.855 2.16 8.86 2.9 ;
      RECT 8.85 2.16 8.855 2.926 ;
      RECT 8.82 2.346 8.85 3.006 ;
      RECT 8.815 2.394 8.82 3.095 ;
      RECT 8.81 2.408 8.815 3.11 ;
      RECT 8.805 2.427 8.81 3.14 ;
      RECT 8.8 2.442 8.805 3.156 ;
      RECT 8.795 2.457 8.8 3.178 ;
      RECT 8.79 2.477 8.795 3.2 ;
      RECT 8.78 2.497 8.79 3.233 ;
      RECT 8.765 2.539 8.78 3.295 ;
      RECT 8.76 2.57 8.765 3.335 ;
      RECT 8.755 2.582 8.76 3.34 ;
      RECT 8.75 2.594 8.755 3.345 ;
      RECT 8.745 2.607 8.75 3.345 ;
      RECT 8.74 2.625 8.745 3.345 ;
      RECT 8.735 2.645 8.74 3.345 ;
      RECT 8.73 2.657 8.735 3.345 ;
      RECT 8.725 2.67 8.73 3.345 ;
      RECT 8.705 2.705 8.725 3.345 ;
      RECT 8.655 2.807 8.705 3.345 ;
      RECT 8.65 2.892 8.655 3.345 ;
      RECT 8.645 2.9 8.65 3.345 ;
      RECT 8.64 2.917 8.645 3.345 ;
      RECT 8.635 2.932 8.64 3.345 ;
      RECT 8.6 2.997 8.635 3.345 ;
      RECT 8.585 3.062 8.6 3.345 ;
      RECT 8.58 3.092 8.585 3.345 ;
      RECT 8.575 3.117 8.58 3.345 ;
      RECT 8.56 3.127 8.57 3.345 ;
      RECT 8.545 3.14 8.56 3.338 ;
      RECT 8.29 2.73 8.36 2.94 ;
      RECT 8.08 2.707 8.085 2.9 ;
      RECT 5.535 2.635 5.795 2.895 ;
      RECT 8.37 2.917 8.375 2.92 ;
      RECT 8.36 2.735 8.37 2.935 ;
      RECT 8.261 2.728 8.29 2.94 ;
      RECT 8.175 2.72 8.261 2.94 ;
      RECT 8.16 2.714 8.175 2.938 ;
      RECT 8.14 2.713 8.16 2.925 ;
      RECT 8.135 2.712 8.14 2.908 ;
      RECT 8.085 2.709 8.135 2.903 ;
      RECT 8.055 2.706 8.08 2.898 ;
      RECT 8.035 2.704 8.055 2.893 ;
      RECT 8.02 2.702 8.035 2.89 ;
      RECT 7.99 2.7 8.02 2.888 ;
      RECT 7.925 2.696 7.99 2.88 ;
      RECT 7.895 2.691 7.925 2.875 ;
      RECT 7.875 2.689 7.895 2.873 ;
      RECT 7.845 2.686 7.875 2.868 ;
      RECT 7.785 2.682 7.845 2.86 ;
      RECT 7.78 2.679 7.785 2.855 ;
      RECT 7.71 2.677 7.78 2.85 ;
      RECT 7.681 2.673 7.71 2.843 ;
      RECT 7.595 2.668 7.681 2.835 ;
      RECT 7.561 2.663 7.595 2.827 ;
      RECT 7.475 2.655 7.561 2.819 ;
      RECT 7.436 2.648 7.475 2.811 ;
      RECT 7.35 2.643 7.436 2.803 ;
      RECT 7.285 2.637 7.35 2.793 ;
      RECT 7.265 2.632 7.285 2.788 ;
      RECT 7.256 2.629 7.265 2.787 ;
      RECT 7.17 2.625 7.256 2.781 ;
      RECT 7.13 2.621 7.17 2.773 ;
      RECT 7.11 2.617 7.13 2.771 ;
      RECT 7.05 2.617 7.11 2.768 ;
      RECT 7.03 2.62 7.05 2.766 ;
      RECT 7.009 2.62 7.03 2.766 ;
      RECT 6.923 2.622 7.009 2.77 ;
      RECT 6.837 2.624 6.923 2.776 ;
      RECT 6.751 2.626 6.837 2.783 ;
      RECT 6.665 2.629 6.751 2.789 ;
      RECT 6.631 2.63 6.665 2.794 ;
      RECT 6.545 2.633 6.631 2.799 ;
      RECT 6.516 2.64 6.545 2.804 ;
      RECT 6.43 2.64 6.516 2.809 ;
      RECT 6.397 2.64 6.43 2.814 ;
      RECT 6.311 2.642 6.397 2.819 ;
      RECT 6.225 2.644 6.311 2.826 ;
      RECT 6.161 2.646 6.225 2.832 ;
      RECT 6.075 2.648 6.161 2.838 ;
      RECT 6.072 2.65 6.075 2.841 ;
      RECT 5.986 2.651 6.072 2.845 ;
      RECT 5.9 2.654 5.986 2.852 ;
      RECT 5.881 2.656 5.9 2.856 ;
      RECT 5.795 2.658 5.881 2.861 ;
      RECT 5.525 2.67 5.535 2.865 ;
      RECT 7.705 7.765 7.995 7.995 ;
      RECT 7.765 7.025 7.935 7.995 ;
      RECT 7.655 7.055 8.03 7.425 ;
      RECT 7.705 7.025 7.995 7.425 ;
      RECT 7.76 2.25 7.945 2.46 ;
      RECT 7.755 2.251 7.95 2.458 ;
      RECT 7.75 2.256 7.96 2.453 ;
      RECT 7.745 2.232 7.75 2.45 ;
      RECT 7.715 2.229 7.745 2.443 ;
      RECT 7.71 2.225 7.715 2.434 ;
      RECT 7.675 2.256 7.96 2.429 ;
      RECT 7.45 2.165 7.71 2.425 ;
      RECT 7.75 2.234 7.755 2.453 ;
      RECT 7.755 2.235 7.76 2.458 ;
      RECT 7.45 2.247 7.83 2.425 ;
      RECT 7.45 2.245 7.815 2.425 ;
      RECT 7.45 2.24 7.805 2.425 ;
      RECT 7.405 3.155 7.455 3.44 ;
      RECT 7.35 3.125 7.355 3.44 ;
      RECT 7.32 3.105 7.325 3.44 ;
      RECT 7.47 3.155 7.53 3.415 ;
      RECT 7.465 3.155 7.47 3.423 ;
      RECT 7.455 3.155 7.465 3.435 ;
      RECT 7.37 3.145 7.405 3.44 ;
      RECT 7.365 3.132 7.37 3.44 ;
      RECT 7.355 3.127 7.365 3.44 ;
      RECT 7.335 3.117 7.35 3.44 ;
      RECT 7.325 3.11 7.335 3.44 ;
      RECT 7.315 3.102 7.32 3.44 ;
      RECT 7.285 3.092 7.315 3.44 ;
      RECT 7.27 3.08 7.285 3.44 ;
      RECT 7.255 3.07 7.27 3.435 ;
      RECT 7.235 3.06 7.255 3.41 ;
      RECT 7.225 3.052 7.235 3.387 ;
      RECT 7.195 3.035 7.225 3.377 ;
      RECT 7.19 3.012 7.195 3.368 ;
      RECT 7.185 2.999 7.19 3.366 ;
      RECT 7.17 2.975 7.185 3.36 ;
      RECT 7.165 2.951 7.17 3.354 ;
      RECT 7.155 2.94 7.165 3.349 ;
      RECT 7.15 2.93 7.155 3.345 ;
      RECT 7.145 2.922 7.15 3.342 ;
      RECT 7.135 2.917 7.145 3.338 ;
      RECT 7.13 2.912 7.135 3.334 ;
      RECT 7.045 2.91 7.13 3.309 ;
      RECT 7.015 2.91 7.045 3.275 ;
      RECT 7 2.91 7.015 3.258 ;
      RECT 6.945 2.91 7 3.203 ;
      RECT 6.94 2.915 6.945 3.152 ;
      RECT 6.93 2.92 6.94 3.142 ;
      RECT 6.925 2.93 6.93 3.128 ;
      RECT 6.875 3.67 7.135 3.93 ;
      RECT 6.795 3.685 7.135 3.906 ;
      RECT 6.775 3.685 7.135 3.901 ;
      RECT 6.751 3.685 7.135 3.899 ;
      RECT 6.665 3.685 7.135 3.894 ;
      RECT 6.515 3.625 6.775 3.89 ;
      RECT 6.47 3.685 7.135 3.885 ;
      RECT 6.465 3.692 7.135 3.88 ;
      RECT 6.48 3.68 6.795 3.89 ;
      RECT 6.37 2.115 6.63 2.375 ;
      RECT 6.37 2.172 6.635 2.368 ;
      RECT 6.37 2.202 6.64 2.3 ;
      RECT 6.43 2.633 6.545 2.635 ;
      RECT 6.516 2.63 6.545 2.635 ;
      RECT 5.54 3.634 5.565 3.874 ;
      RECT 5.525 3.637 5.615 3.868 ;
      RECT 5.52 3.642 5.701 3.863 ;
      RECT 5.515 3.65 5.765 3.861 ;
      RECT 5.515 3.65 5.775 3.86 ;
      RECT 5.51 3.657 5.785 3.853 ;
      RECT 5.51 3.657 5.871 3.842 ;
      RECT 5.505 3.692 5.871 3.838 ;
      RECT 5.505 3.692 5.88 3.827 ;
      RECT 5.785 3.565 6.045 3.825 ;
      RECT 5.495 3.742 6.045 3.823 ;
      RECT 5.765 3.61 5.785 3.858 ;
      RECT 5.701 3.613 5.765 3.862 ;
      RECT 5.615 3.618 5.701 3.867 ;
      RECT 5.545 3.629 6.045 3.825 ;
      RECT 5.565 3.623 5.615 3.872 ;
      RECT 5.69 2.1 5.7 2.362 ;
      RECT 5.68 2.157 5.69 2.365 ;
      RECT 5.655 2.162 5.68 2.371 ;
      RECT 5.63 2.166 5.655 2.383 ;
      RECT 5.62 2.169 5.63 2.393 ;
      RECT 5.615 2.17 5.62 2.398 ;
      RECT 5.61 2.171 5.615 2.403 ;
      RECT 5.605 2.172 5.61 2.405 ;
      RECT 5.58 2.175 5.605 2.408 ;
      RECT 5.55 2.181 5.58 2.411 ;
      RECT 5.485 2.192 5.55 2.414 ;
      RECT 5.44 2.2 5.485 2.418 ;
      RECT 5.425 2.2 5.44 2.426 ;
      RECT 5.42 2.201 5.425 2.433 ;
      RECT 5.415 2.203 5.42 2.436 ;
      RECT 5.41 2.207 5.415 2.439 ;
      RECT 5.4 2.215 5.41 2.443 ;
      RECT 5.395 2.228 5.4 2.448 ;
      RECT 5.39 2.236 5.395 2.45 ;
      RECT 5.385 2.242 5.39 2.45 ;
      RECT 5.38 2.246 5.385 2.453 ;
      RECT 5.375 2.248 5.38 2.456 ;
      RECT 5.37 2.251 5.375 2.459 ;
      RECT 5.36 2.256 5.37 2.463 ;
      RECT 5.355 2.262 5.36 2.468 ;
      RECT 5.345 2.268 5.355 2.472 ;
      RECT 5.33 2.275 5.345 2.478 ;
      RECT 5.301 2.289 5.33 2.488 ;
      RECT 5.215 2.324 5.301 2.52 ;
      RECT 5.195 2.357 5.215 2.549 ;
      RECT 5.175 2.37 5.195 2.56 ;
      RECT 5.155 2.382 5.175 2.571 ;
      RECT 5.105 2.404 5.155 2.591 ;
      RECT 5.09 2.422 5.105 2.608 ;
      RECT 5.085 2.428 5.09 2.611 ;
      RECT 5.08 2.432 5.085 2.614 ;
      RECT 5.075 2.436 5.08 2.618 ;
      RECT 5.07 2.438 5.075 2.621 ;
      RECT 5.06 2.445 5.07 2.624 ;
      RECT 5.055 2.45 5.06 2.628 ;
      RECT 5.05 2.452 5.055 2.631 ;
      RECT 5.045 2.456 5.05 2.634 ;
      RECT 5.04 2.458 5.045 2.638 ;
      RECT 5.025 2.463 5.04 2.643 ;
      RECT 5.02 2.468 5.025 2.646 ;
      RECT 5.015 2.476 5.02 2.649 ;
      RECT 5.01 2.478 5.015 2.652 ;
      RECT 5.005 2.48 5.01 2.655 ;
      RECT 4.995 2.482 5.005 2.661 ;
      RECT 4.96 2.496 4.995 2.673 ;
      RECT 4.95 2.511 4.96 2.683 ;
      RECT 4.875 2.54 4.95 2.707 ;
      RECT 4.87 2.565 4.875 2.73 ;
      RECT 4.855 2.569 4.87 2.736 ;
      RECT 4.845 2.577 4.855 2.741 ;
      RECT 4.815 2.59 4.845 2.745 ;
      RECT 4.805 2.605 4.815 2.75 ;
      RECT 4.795 2.61 4.805 2.753 ;
      RECT 4.79 2.612 4.795 2.755 ;
      RECT 4.775 2.615 4.79 2.758 ;
      RECT 4.77 2.617 4.775 2.761 ;
      RECT 4.75 2.622 4.77 2.765 ;
      RECT 4.72 2.627 4.75 2.773 ;
      RECT 4.695 2.634 4.72 2.781 ;
      RECT 4.69 2.639 4.695 2.786 ;
      RECT 4.66 2.642 4.69 2.79 ;
      RECT 4.62 2.645 4.66 2.8 ;
      RECT 4.585 2.642 4.62 2.812 ;
      RECT 4.575 2.638 4.585 2.819 ;
      RECT 4.55 2.634 4.575 2.825 ;
      RECT 4.545 2.63 4.55 2.83 ;
      RECT 4.505 2.627 4.545 2.83 ;
      RECT 4.49 2.612 4.505 2.831 ;
      RECT 4.467 2.6 4.49 2.831 ;
      RECT 4.381 2.6 4.467 2.832 ;
      RECT 4.295 2.6 4.381 2.834 ;
      RECT 4.275 2.6 4.295 2.831 ;
      RECT 4.27 2.605 4.275 2.826 ;
      RECT 4.265 2.61 4.27 2.824 ;
      RECT 4.255 2.62 4.265 2.822 ;
      RECT 4.25 2.626 4.255 2.815 ;
      RECT 4.245 2.628 4.25 2.8 ;
      RECT 4.24 2.632 4.245 2.79 ;
      RECT 5.7 2.1 5.95 2.36 ;
      RECT 3.425 3.635 3.685 3.895 ;
      RECT 5.72 3.125 5.725 3.335 ;
      RECT 5.725 3.13 5.735 3.33 ;
      RECT 5.675 3.125 5.72 3.35 ;
      RECT 5.665 3.125 5.675 3.37 ;
      RECT 5.646 3.125 5.665 3.375 ;
      RECT 5.56 3.125 5.646 3.372 ;
      RECT 5.53 3.127 5.56 3.37 ;
      RECT 5.475 3.137 5.53 3.368 ;
      RECT 5.41 3.151 5.475 3.366 ;
      RECT 5.405 3.159 5.41 3.365 ;
      RECT 5.39 3.162 5.405 3.363 ;
      RECT 5.325 3.172 5.39 3.359 ;
      RECT 5.277 3.186 5.325 3.36 ;
      RECT 5.191 3.203 5.277 3.374 ;
      RECT 5.105 3.224 5.191 3.391 ;
      RECT 5.085 3.237 5.105 3.401 ;
      RECT 5.04 3.245 5.085 3.408 ;
      RECT 5.005 3.253 5.04 3.416 ;
      RECT 4.971 3.261 5.005 3.424 ;
      RECT 4.885 3.275 4.971 3.436 ;
      RECT 4.85 3.292 4.885 3.448 ;
      RECT 4.841 3.301 4.85 3.452 ;
      RECT 4.755 3.319 4.841 3.469 ;
      RECT 4.696 3.346 4.755 3.496 ;
      RECT 4.61 3.373 4.696 3.524 ;
      RECT 4.59 3.395 4.61 3.544 ;
      RECT 4.53 3.41 4.59 3.56 ;
      RECT 4.52 3.422 4.53 3.573 ;
      RECT 4.515 3.427 4.52 3.576 ;
      RECT 4.505 3.43 4.515 3.579 ;
      RECT 4.5 3.432 4.505 3.582 ;
      RECT 4.47 3.44 4.5 3.589 ;
      RECT 4.455 3.447 4.47 3.597 ;
      RECT 4.445 3.452 4.455 3.601 ;
      RECT 4.44 3.455 4.445 3.604 ;
      RECT 4.43 3.457 4.44 3.607 ;
      RECT 4.395 3.467 4.43 3.616 ;
      RECT 4.32 3.49 4.395 3.638 ;
      RECT 4.3 3.508 4.32 3.656 ;
      RECT 4.27 3.515 4.3 3.666 ;
      RECT 4.25 3.523 4.27 3.676 ;
      RECT 4.24 3.529 4.25 3.683 ;
      RECT 4.221 3.534 4.24 3.689 ;
      RECT 4.135 3.554 4.221 3.709 ;
      RECT 4.12 3.574 4.135 3.728 ;
      RECT 4.075 3.586 4.12 3.739 ;
      RECT 4.01 3.607 4.075 3.762 ;
      RECT 3.97 3.627 4.01 3.783 ;
      RECT 3.96 3.637 3.97 3.793 ;
      RECT 3.91 3.649 3.96 3.804 ;
      RECT 3.89 3.665 3.91 3.816 ;
      RECT 3.86 3.675 3.89 3.822 ;
      RECT 3.85 3.68 3.86 3.824 ;
      RECT 3.781 3.681 3.85 3.83 ;
      RECT 3.695 3.683 3.781 3.84 ;
      RECT 3.685 3.684 3.695 3.845 ;
      RECT 4.955 3.71 5.145 3.92 ;
      RECT 4.945 3.715 5.155 3.913 ;
      RECT 4.93 3.715 5.155 3.878 ;
      RECT 4.85 3.6 5.11 3.86 ;
      RECT 3.765 3.13 3.95 3.425 ;
      RECT 3.755 3.13 3.95 3.423 ;
      RECT 3.74 3.13 3.955 3.418 ;
      RECT 3.74 3.13 3.96 3.415 ;
      RECT 3.735 3.13 3.96 3.413 ;
      RECT 3.73 3.385 3.96 3.403 ;
      RECT 3.735 3.13 3.995 3.39 ;
      RECT 3.695 2.165 3.955 2.425 ;
      RECT 3.505 2.09 3.591 2.423 ;
      RECT 3.48 2.094 3.635 2.419 ;
      RECT 3.591 2.086 3.635 2.419 ;
      RECT 3.591 2.087 3.64 2.418 ;
      RECT 3.505 2.092 3.655 2.417 ;
      RECT 3.48 2.1 3.695 2.416 ;
      RECT 3.475 2.095 3.655 2.411 ;
      RECT 3.465 2.11 3.695 2.318 ;
      RECT 3.465 2.162 3.895 2.318 ;
      RECT 3.465 2.155 3.875 2.318 ;
      RECT 3.465 2.142 3.845 2.318 ;
      RECT 3.465 2.13 3.785 2.318 ;
      RECT 3.465 2.115 3.76 2.318 ;
      RECT 2.665 2.745 2.8 3.04 ;
      RECT 2.925 2.768 2.93 2.955 ;
      RECT 3.645 2.665 3.79 2.9 ;
      RECT 3.805 2.665 3.81 2.89 ;
      RECT 3.84 2.676 3.845 2.87 ;
      RECT 3.835 2.668 3.84 2.875 ;
      RECT 3.815 2.665 3.835 2.88 ;
      RECT 3.81 2.665 3.815 2.888 ;
      RECT 3.8 2.665 3.805 2.893 ;
      RECT 3.79 2.665 3.8 2.898 ;
      RECT 3.62 2.667 3.645 2.9 ;
      RECT 3.57 2.674 3.62 2.9 ;
      RECT 3.565 2.679 3.57 2.9 ;
      RECT 3.526 2.684 3.565 2.901 ;
      RECT 3.44 2.696 3.526 2.902 ;
      RECT 3.431 2.706 3.44 2.902 ;
      RECT 3.345 2.715 3.431 2.904 ;
      RECT 3.321 2.725 3.345 2.906 ;
      RECT 3.235 2.736 3.321 2.907 ;
      RECT 3.205 2.747 3.235 2.909 ;
      RECT 3.175 2.752 3.205 2.911 ;
      RECT 3.15 2.758 3.175 2.914 ;
      RECT 3.135 2.763 3.15 2.915 ;
      RECT 3.09 2.769 3.135 2.915 ;
      RECT 3.085 2.774 3.09 2.916 ;
      RECT 3.065 2.774 3.085 2.918 ;
      RECT 3.045 2.772 3.065 2.923 ;
      RECT 3.01 2.771 3.045 2.93 ;
      RECT 2.98 2.77 3.01 2.94 ;
      RECT 2.93 2.769 2.98 2.95 ;
      RECT 2.84 2.766 2.925 3.04 ;
      RECT 2.815 2.76 2.84 3.04 ;
      RECT 2.8 2.75 2.815 3.04 ;
      RECT 2.615 2.745 2.665 2.96 ;
      RECT 2.605 2.75 2.615 2.95 ;
      RECT 2.845 3.225 3.105 3.485 ;
      RECT 2.845 3.225 3.135 3.378 ;
      RECT 2.845 3.225 3.17 3.363 ;
      RECT 3.1 3.145 3.29 3.355 ;
      RECT 3.09 3.15 3.3 3.348 ;
      RECT 3.055 3.22 3.3 3.348 ;
      RECT 3.085 3.162 3.105 3.485 ;
      RECT 3.07 3.21 3.3 3.348 ;
      RECT 3.075 3.182 3.105 3.485 ;
      RECT 2.155 2.25 2.225 3.355 ;
      RECT 2.89 2.355 3.15 2.615 ;
      RECT 2.47 2.401 2.485 2.61 ;
      RECT 2.806 2.414 2.89 2.565 ;
      RECT 2.72 2.411 2.806 2.565 ;
      RECT 2.681 2.409 2.72 2.565 ;
      RECT 2.595 2.407 2.681 2.565 ;
      RECT 2.535 2.405 2.595 2.576 ;
      RECT 2.5 2.403 2.535 2.594 ;
      RECT 2.485 2.401 2.5 2.605 ;
      RECT 2.455 2.401 2.47 2.618 ;
      RECT 2.445 2.401 2.455 2.623 ;
      RECT 2.42 2.4 2.445 2.628 ;
      RECT 2.405 2.395 2.42 2.634 ;
      RECT 2.4 2.388 2.405 2.639 ;
      RECT 2.375 2.379 2.4 2.645 ;
      RECT 2.33 2.358 2.375 2.658 ;
      RECT 2.32 2.342 2.33 2.668 ;
      RECT 2.305 2.335 2.32 2.678 ;
      RECT 2.295 2.328 2.305 2.695 ;
      RECT 2.29 2.325 2.295 2.725 ;
      RECT 2.285 2.323 2.29 2.755 ;
      RECT 2.28 2.321 2.285 2.792 ;
      RECT 2.265 2.317 2.28 2.859 ;
      RECT 2.265 3.15 2.275 3.35 ;
      RECT 2.26 2.313 2.265 2.985 ;
      RECT 2.26 3.137 2.265 3.355 ;
      RECT 2.255 2.311 2.26 3.07 ;
      RECT 2.255 3.127 2.26 3.355 ;
      RECT 2.24 2.282 2.255 3.355 ;
      RECT 2.225 2.255 2.24 3.355 ;
      RECT 2.15 2.25 2.155 2.605 ;
      RECT 2.15 2.66 2.155 3.355 ;
      RECT 2.135 2.25 2.15 2.583 ;
      RECT 2.145 2.682 2.15 3.355 ;
      RECT 2.135 2.722 2.145 3.355 ;
      RECT 2.1 2.25 2.135 2.525 ;
      RECT 2.13 2.757 2.135 3.355 ;
      RECT 2.115 2.812 2.13 3.355 ;
      RECT 2.11 2.877 2.115 3.355 ;
      RECT 2.095 2.925 2.11 3.355 ;
      RECT 2.07 2.25 2.1 2.48 ;
      RECT 2.09 2.98 2.095 3.355 ;
      RECT 2.075 3.04 2.09 3.355 ;
      RECT 2.07 3.088 2.075 3.353 ;
      RECT 2.065 2.25 2.07 2.473 ;
      RECT 2.065 3.12 2.07 3.348 ;
      RECT 2.04 2.25 2.065 2.465 ;
      RECT 2.03 2.255 2.04 2.455 ;
      RECT 2.245 3.53 2.265 3.77 ;
      RECT 1.475 3.46 1.48 3.67 ;
      RECT 2.755 3.533 2.765 3.728 ;
      RECT 2.75 3.523 2.755 3.731 ;
      RECT 2.67 3.52 2.75 3.754 ;
      RECT 2.666 3.52 2.67 3.776 ;
      RECT 2.58 3.52 2.666 3.786 ;
      RECT 2.565 3.52 2.58 3.794 ;
      RECT 2.536 3.521 2.565 3.792 ;
      RECT 2.45 3.526 2.536 3.788 ;
      RECT 2.437 3.53 2.45 3.784 ;
      RECT 2.351 3.53 2.437 3.78 ;
      RECT 2.265 3.53 2.351 3.774 ;
      RECT 2.181 3.53 2.245 3.768 ;
      RECT 2.095 3.53 2.181 3.763 ;
      RECT 2.075 3.53 2.095 3.759 ;
      RECT 2.015 3.525 2.075 3.756 ;
      RECT 1.987 3.519 2.015 3.753 ;
      RECT 1.901 3.514 1.987 3.749 ;
      RECT 1.815 3.508 1.901 3.743 ;
      RECT 1.74 3.49 1.815 3.738 ;
      RECT 1.705 3.467 1.74 3.734 ;
      RECT 1.695 3.457 1.705 3.733 ;
      RECT 1.64 3.455 1.695 3.732 ;
      RECT 1.565 3.455 1.64 3.728 ;
      RECT 1.555 3.455 1.565 3.723 ;
      RECT 1.54 3.455 1.555 3.715 ;
      RECT 1.49 3.457 1.54 3.693 ;
      RECT 1.48 3.46 1.49 3.673 ;
      RECT 1.47 3.465 1.475 3.668 ;
      RECT 1.465 3.47 1.47 3.663 ;
      RECT 1.59 2.635 1.85 2.895 ;
      RECT 1.59 2.65 1.87 2.86 ;
      RECT 1.59 2.655 1.88 2.855 ;
      RECT -0.425 2.115 -0.165 2.375 ;
      RECT -0.435 2.145 -0.165 2.355 ;
      RECT 1.485 2.06 1.745 2.32 ;
      RECT 1.48 2.135 1.485 2.321 ;
      RECT 1.455 2.14 1.48 2.323 ;
      RECT 1.44 2.147 1.455 2.326 ;
      RECT 1.38 2.165 1.44 2.331 ;
      RECT 1.35 2.185 1.38 2.338 ;
      RECT 1.325 2.193 1.35 2.343 ;
      RECT 1.3 2.201 1.325 2.345 ;
      RECT 1.282 2.205 1.3 2.344 ;
      RECT 1.196 2.203 1.282 2.344 ;
      RECT 1.11 2.201 1.196 2.344 ;
      RECT 1.024 2.199 1.11 2.343 ;
      RECT 0.938 2.197 1.024 2.343 ;
      RECT 0.852 2.195 0.938 2.343 ;
      RECT 0.766 2.193 0.852 2.343 ;
      RECT 0.68 2.191 0.766 2.342 ;
      RECT 0.662 2.19 0.68 2.342 ;
      RECT 0.576 2.189 0.662 2.342 ;
      RECT 0.49 2.187 0.576 2.342 ;
      RECT 0.404 2.186 0.49 2.341 ;
      RECT 0.318 2.185 0.404 2.341 ;
      RECT 0.232 2.183 0.318 2.341 ;
      RECT 0.146 2.182 0.232 2.341 ;
      RECT 0.06 2.18 0.146 2.34 ;
      RECT 0.036 2.178 0.06 2.34 ;
      RECT -0.05 2.171 0.036 2.34 ;
      RECT -0.079 2.163 -0.05 2.34 ;
      RECT -0.165 2.155 -0.079 2.34 ;
      RECT -0.445 2.152 -0.435 2.35 ;
      RECT 1.06 3.115 1.065 3.465 ;
      RECT 0.83 3.205 0.97 3.465 ;
      RECT 1.305 2.89 1.35 3.1 ;
      RECT 1.36 2.901 1.37 3.095 ;
      RECT 1.35 2.893 1.36 3.1 ;
      RECT 1.285 2.89 1.305 3.105 ;
      RECT 1.255 2.89 1.285 3.128 ;
      RECT 1.245 2.89 1.255 3.153 ;
      RECT 1.24 2.89 1.245 3.163 ;
      RECT 1.185 2.89 1.24 3.203 ;
      RECT 1.18 2.89 1.185 3.243 ;
      RECT 1.175 2.892 1.18 3.248 ;
      RECT 1.16 2.902 1.175 3.259 ;
      RECT 1.115 2.96 1.16 3.295 ;
      RECT 1.105 3.015 1.115 3.329 ;
      RECT 1.09 3.042 1.105 3.345 ;
      RECT 1.08 3.069 1.09 3.465 ;
      RECT 1.065 3.092 1.08 3.465 ;
      RECT 1.055 3.132 1.06 3.465 ;
      RECT 1.05 3.142 1.055 3.465 ;
      RECT 1.045 3.157 1.05 3.465 ;
      RECT 1.035 3.162 1.045 3.465 ;
      RECT 0.97 3.185 1.035 3.465 ;
      RECT 0.47 2.68 0.66 2.89 ;
      RECT -0.955 2.605 -0.695 2.865 ;
      RECT -0.605 2.6 -0.51 2.81 ;
      RECT -0.63 2.615 -0.62 2.81 ;
      RECT 0.66 2.687 0.67 2.885 ;
      RECT 0.46 2.687 0.47 2.885 ;
      RECT 0.445 2.702 0.46 2.875 ;
      RECT 0.44 2.71 0.445 2.868 ;
      RECT 0.43 2.713 0.44 2.865 ;
      RECT 0.395 2.712 0.43 2.863 ;
      RECT 0.366 2.708 0.395 2.86 ;
      RECT 0.28 2.703 0.366 2.857 ;
      RECT 0.22 2.697 0.28 2.853 ;
      RECT 0.191 2.693 0.22 2.85 ;
      RECT 0.105 2.685 0.191 2.847 ;
      RECT 0.096 2.679 0.105 2.845 ;
      RECT 0.01 2.674 0.096 2.843 ;
      RECT -0.013 2.669 0.01 2.84 ;
      RECT -0.099 2.663 -0.013 2.837 ;
      RECT -0.185 2.654 -0.099 2.832 ;
      RECT -0.195 2.649 -0.185 2.83 ;
      RECT -0.214 2.648 -0.195 2.829 ;
      RECT -0.3 2.643 -0.214 2.825 ;
      RECT -0.32 2.638 -0.3 2.821 ;
      RECT -0.38 2.633 -0.32 2.818 ;
      RECT -0.405 2.623 -0.38 2.816 ;
      RECT -0.41 2.616 -0.405 2.815 ;
      RECT -0.42 2.607 -0.41 2.814 ;
      RECT -0.424 2.6 -0.42 2.814 ;
      RECT -0.51 2.6 -0.424 2.812 ;
      RECT -0.62 2.607 -0.605 2.81 ;
      RECT -0.635 2.617 -0.63 2.81 ;
      RECT -0.655 2.62 -0.635 2.807 ;
      RECT -0.685 2.62 -0.655 2.803 ;
      RECT -0.695 2.62 -0.685 2.803 ;
      RECT 0.22 3.115 0.48 3.375 ;
      RECT 0.15 3.125 0.48 3.335 ;
      RECT 0.14 3.132 0.48 3.33 ;
      RECT -0.44 3.12 -0.18 3.38 ;
      RECT -0.44 3.16 -0.075 3.37 ;
      RECT -0.44 3.162 -0.07 3.369 ;
      RECT -0.44 3.17 -0.065 3.366 ;
      RECT -1.515 2.245 -1.415 3.77 ;
      RECT -1.325 3.385 -1.275 3.645 ;
      RECT -1.33 2.258 -1.325 2.445 ;
      RECT -1.335 3.366 -1.325 3.645 ;
      RECT -1.335 2.255 -1.33 2.453 ;
      RECT -1.35 2.249 -1.335 2.46 ;
      RECT -1.34 3.354 -1.335 3.728 ;
      RECT -1.35 3.342 -1.34 3.765 ;
      RECT -1.36 2.245 -1.35 2.467 ;
      RECT -1.36 3.327 -1.35 3.77 ;
      RECT -1.365 2.245 -1.36 2.475 ;
      RECT -1.385 3.297 -1.36 3.77 ;
      RECT -1.405 2.245 -1.365 2.523 ;
      RECT -1.395 3.257 -1.385 3.77 ;
      RECT -1.405 3.212 -1.395 3.77 ;
      RECT -1.41 2.245 -1.405 2.593 ;
      RECT -1.41 3.17 -1.405 3.77 ;
      RECT -1.415 2.245 -1.41 3.07 ;
      RECT -1.415 3.152 -1.41 3.77 ;
      RECT -1.525 2.248 -1.515 3.77 ;
      RECT -1.54 2.255 -1.525 3.766 ;
      RECT -1.545 2.265 -1.54 3.761 ;
      RECT -1.55 2.465 -1.545 3.653 ;
      RECT -1.555 2.55 -1.55 3.205 ;
      RECT -2.895 6.655 -2.605 6.885 ;
      RECT -3.065 6.685 -2.605 6.855 ;
      RECT -3.325 7.765 -3.035 7.995 ;
      RECT -3.265 7.025 -3.095 7.995 ;
      RECT -3.355 7.025 -3.005 7.315 ;
      RECT -3.73 6.285 -3.38 6.575 ;
      RECT -3.87 6.315 -3.38 6.485 ;
      RECT -4.695 5.915 -4.405 6.145 ;
      RECT -4.695 5.945 -4.235 6.115 ;
      RECT 82.175 1.14 82.55 1.51 ;
      RECT 76.155 2.225 76.415 2.485 ;
      RECT 64.25 1.14 64.625 1.51 ;
      RECT 58.23 2.225 58.49 2.485 ;
      RECT 46.325 1.14 46.7 1.51 ;
      RECT 40.305 2.225 40.565 2.485 ;
      RECT 28.4 1.14 28.775 1.51 ;
      RECT 22.38 2.225 22.64 2.485 ;
      RECT 10.475 1.14 10.85 1.51 ;
      RECT 4.455 2.225 4.715 2.485 ;
    LAYER mcon ;
      RECT 87.01 0.915 87.18 1.085 ;
      RECT 87.01 2.395 87.18 2.565 ;
      RECT 87.01 6.315 87.18 6.485 ;
      RECT 87.01 7.795 87.18 7.965 ;
      RECT 86.66 0.105 86.83 0.275 ;
      RECT 86.66 4.165 86.83 4.335 ;
      RECT 86.66 4.545 86.83 4.715 ;
      RECT 86.66 8.605 86.83 8.775 ;
      RECT 86.64 2.765 86.81 2.935 ;
      RECT 86.64 5.945 86.81 6.115 ;
      RECT 86.02 0.915 86.19 1.085 ;
      RECT 86.02 2.395 86.19 2.565 ;
      RECT 86.02 6.315 86.19 6.485 ;
      RECT 86.02 7.795 86.19 7.965 ;
      RECT 85.67 0.105 85.84 0.275 ;
      RECT 85.67 4.165 85.84 4.335 ;
      RECT 85.67 4.545 85.84 4.715 ;
      RECT 85.67 8.605 85.84 8.775 ;
      RECT 85.65 2.765 85.82 2.935 ;
      RECT 85.65 5.945 85.82 6.115 ;
      RECT 84.965 0.105 85.135 0.275 ;
      RECT 84.965 4.165 85.135 4.335 ;
      RECT 84.965 4.545 85.135 4.715 ;
      RECT 84.965 8.605 85.135 8.775 ;
      RECT 84.655 2.025 84.825 2.195 ;
      RECT 84.655 6.685 84.825 6.855 ;
      RECT 84.285 0.105 84.455 0.275 ;
      RECT 84.285 8.605 84.455 8.775 ;
      RECT 84.225 0.915 84.395 1.085 ;
      RECT 84.225 1.655 84.395 1.825 ;
      RECT 84.225 7.055 84.395 7.225 ;
      RECT 84.225 7.795 84.395 7.965 ;
      RECT 83.85 2.395 84.02 2.565 ;
      RECT 83.85 6.315 84.02 6.485 ;
      RECT 83.605 0.105 83.775 0.275 ;
      RECT 83.605 8.605 83.775 8.775 ;
      RECT 82.925 0.105 83.095 0.275 ;
      RECT 82.925 8.605 83.095 8.775 ;
      RECT 82.855 2.765 83.025 2.935 ;
      RECT 82.855 5.945 83.025 6.115 ;
      RECT 81.645 1.565 81.815 1.735 ;
      RECT 81.645 4.285 81.815 4.455 ;
      RECT 81.185 1.565 81.355 1.735 ;
      RECT 81.185 4.285 81.355 4.455 ;
      RECT 80.79 2.905 80.96 3.075 ;
      RECT 80.725 1.565 80.895 1.735 ;
      RECT 80.725 4.285 80.895 4.455 ;
      RECT 80.58 2.245 80.75 2.415 ;
      RECT 80.265 1.565 80.435 1.735 ;
      RECT 80.265 3.155 80.435 3.325 ;
      RECT 80.265 4.285 80.435 4.455 ;
      RECT 80.205 4.545 80.375 4.715 ;
      RECT 80.205 8.605 80.375 8.775 ;
      RECT 79.895 6.685 80.065 6.855 ;
      RECT 79.88 2.75 80.05 2.92 ;
      RECT 79.805 1.565 79.975 1.735 ;
      RECT 79.805 4.285 79.975 4.455 ;
      RECT 79.665 3.315 79.835 3.485 ;
      RECT 79.645 3.715 79.815 3.885 ;
      RECT 79.525 8.605 79.695 8.775 ;
      RECT 79.47 2.27 79.64 2.44 ;
      RECT 79.465 7.055 79.635 7.225 ;
      RECT 79.465 7.795 79.635 7.965 ;
      RECT 79.345 1.565 79.515 1.735 ;
      RECT 79.345 4.285 79.515 4.455 ;
      RECT 79.09 6.315 79.26 6.485 ;
      RECT 78.975 3.25 79.145 3.42 ;
      RECT 78.885 1.565 79.055 1.735 ;
      RECT 78.885 4.285 79.055 4.455 ;
      RECT 78.845 8.605 79.015 8.775 ;
      RECT 78.65 2.935 78.82 3.105 ;
      RECT 78.585 3.715 78.755 3.885 ;
      RECT 78.425 1.565 78.595 1.735 ;
      RECT 78.425 4.285 78.595 4.455 ;
      RECT 78.185 3.7 78.355 3.87 ;
      RECT 78.165 8.605 78.335 8.775 ;
      RECT 78.145 2.185 78.315 2.355 ;
      RECT 78.095 5.945 78.265 6.115 ;
      RECT 77.965 1.565 78.135 1.735 ;
      RECT 77.965 4.285 78.135 4.455 ;
      RECT 77.505 1.565 77.675 1.735 ;
      RECT 77.505 4.285 77.675 4.455 ;
      RECT 77.245 2.685 77.415 2.855 ;
      RECT 77.245 3.145 77.415 3.315 ;
      RECT 77.245 3.66 77.415 3.83 ;
      RECT 77.13 2.22 77.3 2.39 ;
      RECT 77.045 1.565 77.215 1.735 ;
      RECT 77.045 4.285 77.215 4.455 ;
      RECT 76.665 3.73 76.835 3.9 ;
      RECT 76.585 1.565 76.755 1.735 ;
      RECT 76.585 4.285 76.755 4.455 ;
      RECT 76.185 2.26 76.355 2.43 ;
      RECT 76.125 1.565 76.295 1.735 ;
      RECT 76.125 4.285 76.295 4.455 ;
      RECT 75.97 2.635 76.14 2.805 ;
      RECT 75.665 1.565 75.835 1.735 ;
      RECT 75.665 4.285 75.835 4.455 ;
      RECT 75.47 3.235 75.64 3.405 ;
      RECT 75.355 2.685 75.525 2.855 ;
      RECT 75.205 1.565 75.375 1.735 ;
      RECT 75.205 4.285 75.375 4.455 ;
      RECT 75.185 2.135 75.355 2.305 ;
      RECT 74.81 3.165 74.98 3.335 ;
      RECT 74.745 1.565 74.915 1.735 ;
      RECT 74.745 4.285 74.915 4.455 ;
      RECT 74.325 2.765 74.495 2.935 ;
      RECT 74.285 1.565 74.455 1.735 ;
      RECT 74.285 4.285 74.455 4.455 ;
      RECT 74.275 3.54 74.445 3.71 ;
      RECT 73.825 1.565 73.995 1.735 ;
      RECT 73.825 4.285 73.995 4.455 ;
      RECT 73.785 3.165 73.955 3.335 ;
      RECT 73.75 2.27 73.92 2.44 ;
      RECT 73.39 2.67 73.56 2.84 ;
      RECT 73.365 1.565 73.535 1.735 ;
      RECT 73.365 4.285 73.535 4.455 ;
      RECT 73.185 3.48 73.355 3.65 ;
      RECT 72.905 1.565 73.075 1.735 ;
      RECT 72.905 4.285 73.075 4.455 ;
      RECT 72.88 2.91 73.05 3.08 ;
      RECT 72.445 1.565 72.615 1.735 ;
      RECT 72.445 4.285 72.615 4.455 ;
      RECT 72.18 2.7 72.35 2.87 ;
      RECT 71.985 1.565 72.155 1.735 ;
      RECT 71.985 4.285 72.155 4.455 ;
      RECT 71.86 3.145 72.03 3.315 ;
      RECT 71.525 1.565 71.695 1.735 ;
      RECT 71.525 4.285 71.695 4.455 ;
      RECT 71.445 3.18 71.615 3.35 ;
      RECT 71.275 2.165 71.445 2.335 ;
      RECT 71.1 2.62 71.27 2.79 ;
      RECT 71.065 1.565 71.235 1.735 ;
      RECT 71.065 4.285 71.235 4.455 ;
      RECT 70.605 1.565 70.775 1.735 ;
      RECT 70.605 4.285 70.775 4.455 ;
      RECT 70.18 2.27 70.35 2.44 ;
      RECT 70.175 3.585 70.345 3.755 ;
      RECT 70.145 1.565 70.315 1.735 ;
      RECT 70.145 4.285 70.315 4.455 ;
      RECT 69.085 0.915 69.255 1.085 ;
      RECT 69.085 2.395 69.255 2.565 ;
      RECT 69.085 6.315 69.255 6.485 ;
      RECT 69.085 7.795 69.255 7.965 ;
      RECT 68.735 0.105 68.905 0.275 ;
      RECT 68.735 4.165 68.905 4.335 ;
      RECT 68.735 4.545 68.905 4.715 ;
      RECT 68.735 8.605 68.905 8.775 ;
      RECT 68.715 2.765 68.885 2.935 ;
      RECT 68.715 5.945 68.885 6.115 ;
      RECT 68.095 0.915 68.265 1.085 ;
      RECT 68.095 2.395 68.265 2.565 ;
      RECT 68.095 6.315 68.265 6.485 ;
      RECT 68.095 7.795 68.265 7.965 ;
      RECT 67.745 0.105 67.915 0.275 ;
      RECT 67.745 4.165 67.915 4.335 ;
      RECT 67.745 4.545 67.915 4.715 ;
      RECT 67.745 8.605 67.915 8.775 ;
      RECT 67.725 2.765 67.895 2.935 ;
      RECT 67.725 5.945 67.895 6.115 ;
      RECT 67.04 0.105 67.21 0.275 ;
      RECT 67.04 4.165 67.21 4.335 ;
      RECT 67.04 4.545 67.21 4.715 ;
      RECT 67.04 8.605 67.21 8.775 ;
      RECT 66.73 2.025 66.9 2.195 ;
      RECT 66.73 6.685 66.9 6.855 ;
      RECT 66.36 0.105 66.53 0.275 ;
      RECT 66.36 8.605 66.53 8.775 ;
      RECT 66.3 0.915 66.47 1.085 ;
      RECT 66.3 1.655 66.47 1.825 ;
      RECT 66.3 7.055 66.47 7.225 ;
      RECT 66.3 7.795 66.47 7.965 ;
      RECT 65.925 2.395 66.095 2.565 ;
      RECT 65.925 6.315 66.095 6.485 ;
      RECT 65.68 0.105 65.85 0.275 ;
      RECT 65.68 8.605 65.85 8.775 ;
      RECT 65 0.105 65.17 0.275 ;
      RECT 65 8.605 65.17 8.775 ;
      RECT 64.93 2.765 65.1 2.935 ;
      RECT 64.93 5.945 65.1 6.115 ;
      RECT 63.72 1.565 63.89 1.735 ;
      RECT 63.72 4.285 63.89 4.455 ;
      RECT 63.26 1.565 63.43 1.735 ;
      RECT 63.26 4.285 63.43 4.455 ;
      RECT 62.865 2.905 63.035 3.075 ;
      RECT 62.8 1.565 62.97 1.735 ;
      RECT 62.8 4.285 62.97 4.455 ;
      RECT 62.655 2.245 62.825 2.415 ;
      RECT 62.34 1.565 62.51 1.735 ;
      RECT 62.34 3.155 62.51 3.325 ;
      RECT 62.34 4.285 62.51 4.455 ;
      RECT 62.28 4.545 62.45 4.715 ;
      RECT 62.28 8.605 62.45 8.775 ;
      RECT 61.97 6.685 62.14 6.855 ;
      RECT 61.955 2.75 62.125 2.92 ;
      RECT 61.88 1.565 62.05 1.735 ;
      RECT 61.88 4.285 62.05 4.455 ;
      RECT 61.74 3.315 61.91 3.485 ;
      RECT 61.72 3.715 61.89 3.885 ;
      RECT 61.6 8.605 61.77 8.775 ;
      RECT 61.545 2.27 61.715 2.44 ;
      RECT 61.54 7.055 61.71 7.225 ;
      RECT 61.54 7.795 61.71 7.965 ;
      RECT 61.42 1.565 61.59 1.735 ;
      RECT 61.42 4.285 61.59 4.455 ;
      RECT 61.165 6.315 61.335 6.485 ;
      RECT 61.05 3.25 61.22 3.42 ;
      RECT 60.96 1.565 61.13 1.735 ;
      RECT 60.96 4.285 61.13 4.455 ;
      RECT 60.92 8.605 61.09 8.775 ;
      RECT 60.725 2.935 60.895 3.105 ;
      RECT 60.66 3.715 60.83 3.885 ;
      RECT 60.5 1.565 60.67 1.735 ;
      RECT 60.5 4.285 60.67 4.455 ;
      RECT 60.26 3.7 60.43 3.87 ;
      RECT 60.24 8.605 60.41 8.775 ;
      RECT 60.22 2.185 60.39 2.355 ;
      RECT 60.17 5.945 60.34 6.115 ;
      RECT 60.04 1.565 60.21 1.735 ;
      RECT 60.04 4.285 60.21 4.455 ;
      RECT 59.58 1.565 59.75 1.735 ;
      RECT 59.58 4.285 59.75 4.455 ;
      RECT 59.32 2.685 59.49 2.855 ;
      RECT 59.32 3.145 59.49 3.315 ;
      RECT 59.32 3.66 59.49 3.83 ;
      RECT 59.205 2.22 59.375 2.39 ;
      RECT 59.12 1.565 59.29 1.735 ;
      RECT 59.12 4.285 59.29 4.455 ;
      RECT 58.74 3.73 58.91 3.9 ;
      RECT 58.66 1.565 58.83 1.735 ;
      RECT 58.66 4.285 58.83 4.455 ;
      RECT 58.26 2.26 58.43 2.43 ;
      RECT 58.2 1.565 58.37 1.735 ;
      RECT 58.2 4.285 58.37 4.455 ;
      RECT 58.045 2.635 58.215 2.805 ;
      RECT 57.74 1.565 57.91 1.735 ;
      RECT 57.74 4.285 57.91 4.455 ;
      RECT 57.545 3.235 57.715 3.405 ;
      RECT 57.43 2.685 57.6 2.855 ;
      RECT 57.28 1.565 57.45 1.735 ;
      RECT 57.28 4.285 57.45 4.455 ;
      RECT 57.26 2.135 57.43 2.305 ;
      RECT 56.885 3.165 57.055 3.335 ;
      RECT 56.82 1.565 56.99 1.735 ;
      RECT 56.82 4.285 56.99 4.455 ;
      RECT 56.4 2.765 56.57 2.935 ;
      RECT 56.36 1.565 56.53 1.735 ;
      RECT 56.36 4.285 56.53 4.455 ;
      RECT 56.35 3.54 56.52 3.71 ;
      RECT 55.9 1.565 56.07 1.735 ;
      RECT 55.9 4.285 56.07 4.455 ;
      RECT 55.86 3.165 56.03 3.335 ;
      RECT 55.825 2.27 55.995 2.44 ;
      RECT 55.465 2.67 55.635 2.84 ;
      RECT 55.44 1.565 55.61 1.735 ;
      RECT 55.44 4.285 55.61 4.455 ;
      RECT 55.26 3.48 55.43 3.65 ;
      RECT 54.98 1.565 55.15 1.735 ;
      RECT 54.98 4.285 55.15 4.455 ;
      RECT 54.955 2.91 55.125 3.08 ;
      RECT 54.52 1.565 54.69 1.735 ;
      RECT 54.52 4.285 54.69 4.455 ;
      RECT 54.255 2.7 54.425 2.87 ;
      RECT 54.06 1.565 54.23 1.735 ;
      RECT 54.06 4.285 54.23 4.455 ;
      RECT 53.935 3.145 54.105 3.315 ;
      RECT 53.6 1.565 53.77 1.735 ;
      RECT 53.6 4.285 53.77 4.455 ;
      RECT 53.52 3.18 53.69 3.35 ;
      RECT 53.35 2.165 53.52 2.335 ;
      RECT 53.175 2.62 53.345 2.79 ;
      RECT 53.14 1.565 53.31 1.735 ;
      RECT 53.14 4.285 53.31 4.455 ;
      RECT 52.68 1.565 52.85 1.735 ;
      RECT 52.68 4.285 52.85 4.455 ;
      RECT 52.255 2.27 52.425 2.44 ;
      RECT 52.25 3.585 52.42 3.755 ;
      RECT 52.22 1.565 52.39 1.735 ;
      RECT 52.22 4.285 52.39 4.455 ;
      RECT 51.16 0.915 51.33 1.085 ;
      RECT 51.16 2.395 51.33 2.565 ;
      RECT 51.16 6.315 51.33 6.485 ;
      RECT 51.16 7.795 51.33 7.965 ;
      RECT 50.81 0.105 50.98 0.275 ;
      RECT 50.81 4.165 50.98 4.335 ;
      RECT 50.81 4.545 50.98 4.715 ;
      RECT 50.81 8.605 50.98 8.775 ;
      RECT 50.79 2.765 50.96 2.935 ;
      RECT 50.79 5.945 50.96 6.115 ;
      RECT 50.17 0.915 50.34 1.085 ;
      RECT 50.17 2.395 50.34 2.565 ;
      RECT 50.17 6.315 50.34 6.485 ;
      RECT 50.17 7.795 50.34 7.965 ;
      RECT 49.82 0.105 49.99 0.275 ;
      RECT 49.82 4.165 49.99 4.335 ;
      RECT 49.82 4.545 49.99 4.715 ;
      RECT 49.82 8.605 49.99 8.775 ;
      RECT 49.8 2.765 49.97 2.935 ;
      RECT 49.8 5.945 49.97 6.115 ;
      RECT 49.115 0.105 49.285 0.275 ;
      RECT 49.115 4.165 49.285 4.335 ;
      RECT 49.115 4.545 49.285 4.715 ;
      RECT 49.115 8.605 49.285 8.775 ;
      RECT 48.805 2.025 48.975 2.195 ;
      RECT 48.805 6.685 48.975 6.855 ;
      RECT 48.435 0.105 48.605 0.275 ;
      RECT 48.435 8.605 48.605 8.775 ;
      RECT 48.375 0.915 48.545 1.085 ;
      RECT 48.375 1.655 48.545 1.825 ;
      RECT 48.375 7.055 48.545 7.225 ;
      RECT 48.375 7.795 48.545 7.965 ;
      RECT 48 2.395 48.17 2.565 ;
      RECT 48 6.315 48.17 6.485 ;
      RECT 47.755 0.105 47.925 0.275 ;
      RECT 47.755 8.605 47.925 8.775 ;
      RECT 47.075 0.105 47.245 0.275 ;
      RECT 47.075 8.605 47.245 8.775 ;
      RECT 47.005 2.765 47.175 2.935 ;
      RECT 47.005 5.945 47.175 6.115 ;
      RECT 45.795 1.565 45.965 1.735 ;
      RECT 45.795 4.285 45.965 4.455 ;
      RECT 45.335 1.565 45.505 1.735 ;
      RECT 45.335 4.285 45.505 4.455 ;
      RECT 44.94 2.905 45.11 3.075 ;
      RECT 44.875 1.565 45.045 1.735 ;
      RECT 44.875 4.285 45.045 4.455 ;
      RECT 44.73 2.245 44.9 2.415 ;
      RECT 44.415 1.565 44.585 1.735 ;
      RECT 44.415 3.155 44.585 3.325 ;
      RECT 44.415 4.285 44.585 4.455 ;
      RECT 44.355 4.545 44.525 4.715 ;
      RECT 44.355 8.605 44.525 8.775 ;
      RECT 44.045 6.685 44.215 6.855 ;
      RECT 44.03 2.75 44.2 2.92 ;
      RECT 43.955 1.565 44.125 1.735 ;
      RECT 43.955 4.285 44.125 4.455 ;
      RECT 43.815 3.315 43.985 3.485 ;
      RECT 43.795 3.715 43.965 3.885 ;
      RECT 43.675 8.605 43.845 8.775 ;
      RECT 43.62 2.27 43.79 2.44 ;
      RECT 43.615 7.055 43.785 7.225 ;
      RECT 43.615 7.795 43.785 7.965 ;
      RECT 43.495 1.565 43.665 1.735 ;
      RECT 43.495 4.285 43.665 4.455 ;
      RECT 43.24 6.315 43.41 6.485 ;
      RECT 43.125 3.25 43.295 3.42 ;
      RECT 43.035 1.565 43.205 1.735 ;
      RECT 43.035 4.285 43.205 4.455 ;
      RECT 42.995 8.605 43.165 8.775 ;
      RECT 42.8 2.935 42.97 3.105 ;
      RECT 42.735 3.715 42.905 3.885 ;
      RECT 42.575 1.565 42.745 1.735 ;
      RECT 42.575 4.285 42.745 4.455 ;
      RECT 42.335 3.7 42.505 3.87 ;
      RECT 42.315 8.605 42.485 8.775 ;
      RECT 42.295 2.185 42.465 2.355 ;
      RECT 42.245 5.945 42.415 6.115 ;
      RECT 42.115 1.565 42.285 1.735 ;
      RECT 42.115 4.285 42.285 4.455 ;
      RECT 41.655 1.565 41.825 1.735 ;
      RECT 41.655 4.285 41.825 4.455 ;
      RECT 41.395 2.685 41.565 2.855 ;
      RECT 41.395 3.145 41.565 3.315 ;
      RECT 41.395 3.66 41.565 3.83 ;
      RECT 41.28 2.22 41.45 2.39 ;
      RECT 41.195 1.565 41.365 1.735 ;
      RECT 41.195 4.285 41.365 4.455 ;
      RECT 40.815 3.73 40.985 3.9 ;
      RECT 40.735 1.565 40.905 1.735 ;
      RECT 40.735 4.285 40.905 4.455 ;
      RECT 40.335 2.26 40.505 2.43 ;
      RECT 40.275 1.565 40.445 1.735 ;
      RECT 40.275 4.285 40.445 4.455 ;
      RECT 40.12 2.635 40.29 2.805 ;
      RECT 39.815 1.565 39.985 1.735 ;
      RECT 39.815 4.285 39.985 4.455 ;
      RECT 39.62 3.235 39.79 3.405 ;
      RECT 39.505 2.685 39.675 2.855 ;
      RECT 39.355 1.565 39.525 1.735 ;
      RECT 39.355 4.285 39.525 4.455 ;
      RECT 39.335 2.135 39.505 2.305 ;
      RECT 38.96 3.165 39.13 3.335 ;
      RECT 38.895 1.565 39.065 1.735 ;
      RECT 38.895 4.285 39.065 4.455 ;
      RECT 38.475 2.765 38.645 2.935 ;
      RECT 38.435 1.565 38.605 1.735 ;
      RECT 38.435 4.285 38.605 4.455 ;
      RECT 38.425 3.54 38.595 3.71 ;
      RECT 37.975 1.565 38.145 1.735 ;
      RECT 37.975 4.285 38.145 4.455 ;
      RECT 37.935 3.165 38.105 3.335 ;
      RECT 37.9 2.27 38.07 2.44 ;
      RECT 37.54 2.67 37.71 2.84 ;
      RECT 37.515 1.565 37.685 1.735 ;
      RECT 37.515 4.285 37.685 4.455 ;
      RECT 37.335 3.48 37.505 3.65 ;
      RECT 37.055 1.565 37.225 1.735 ;
      RECT 37.055 4.285 37.225 4.455 ;
      RECT 37.03 2.91 37.2 3.08 ;
      RECT 36.595 1.565 36.765 1.735 ;
      RECT 36.595 4.285 36.765 4.455 ;
      RECT 36.33 2.7 36.5 2.87 ;
      RECT 36.135 1.565 36.305 1.735 ;
      RECT 36.135 4.285 36.305 4.455 ;
      RECT 36.01 3.145 36.18 3.315 ;
      RECT 35.675 1.565 35.845 1.735 ;
      RECT 35.675 4.285 35.845 4.455 ;
      RECT 35.595 3.18 35.765 3.35 ;
      RECT 35.425 2.165 35.595 2.335 ;
      RECT 35.25 2.62 35.42 2.79 ;
      RECT 35.215 1.565 35.385 1.735 ;
      RECT 35.215 4.285 35.385 4.455 ;
      RECT 34.755 1.565 34.925 1.735 ;
      RECT 34.755 4.285 34.925 4.455 ;
      RECT 34.33 2.27 34.5 2.44 ;
      RECT 34.325 3.585 34.495 3.755 ;
      RECT 34.295 1.565 34.465 1.735 ;
      RECT 34.295 4.285 34.465 4.455 ;
      RECT 33.235 0.915 33.405 1.085 ;
      RECT 33.235 2.395 33.405 2.565 ;
      RECT 33.235 6.315 33.405 6.485 ;
      RECT 33.235 7.795 33.405 7.965 ;
      RECT 32.885 0.105 33.055 0.275 ;
      RECT 32.885 4.165 33.055 4.335 ;
      RECT 32.885 4.545 33.055 4.715 ;
      RECT 32.885 8.605 33.055 8.775 ;
      RECT 32.865 2.765 33.035 2.935 ;
      RECT 32.865 5.945 33.035 6.115 ;
      RECT 32.245 0.915 32.415 1.085 ;
      RECT 32.245 2.395 32.415 2.565 ;
      RECT 32.245 6.315 32.415 6.485 ;
      RECT 32.245 7.795 32.415 7.965 ;
      RECT 31.895 0.105 32.065 0.275 ;
      RECT 31.895 4.165 32.065 4.335 ;
      RECT 31.895 4.545 32.065 4.715 ;
      RECT 31.895 8.605 32.065 8.775 ;
      RECT 31.875 2.765 32.045 2.935 ;
      RECT 31.875 5.945 32.045 6.115 ;
      RECT 31.19 0.105 31.36 0.275 ;
      RECT 31.19 4.165 31.36 4.335 ;
      RECT 31.19 4.545 31.36 4.715 ;
      RECT 31.19 8.605 31.36 8.775 ;
      RECT 30.88 2.025 31.05 2.195 ;
      RECT 30.88 6.685 31.05 6.855 ;
      RECT 30.51 0.105 30.68 0.275 ;
      RECT 30.51 8.605 30.68 8.775 ;
      RECT 30.45 0.915 30.62 1.085 ;
      RECT 30.45 1.655 30.62 1.825 ;
      RECT 30.45 7.055 30.62 7.225 ;
      RECT 30.45 7.795 30.62 7.965 ;
      RECT 30.075 2.395 30.245 2.565 ;
      RECT 30.075 6.315 30.245 6.485 ;
      RECT 29.83 0.105 30 0.275 ;
      RECT 29.83 8.605 30 8.775 ;
      RECT 29.15 0.105 29.32 0.275 ;
      RECT 29.15 8.605 29.32 8.775 ;
      RECT 29.08 2.765 29.25 2.935 ;
      RECT 29.08 5.945 29.25 6.115 ;
      RECT 27.87 1.565 28.04 1.735 ;
      RECT 27.87 4.285 28.04 4.455 ;
      RECT 27.41 1.565 27.58 1.735 ;
      RECT 27.41 4.285 27.58 4.455 ;
      RECT 27.015 2.905 27.185 3.075 ;
      RECT 26.95 1.565 27.12 1.735 ;
      RECT 26.95 4.285 27.12 4.455 ;
      RECT 26.805 2.245 26.975 2.415 ;
      RECT 26.49 1.565 26.66 1.735 ;
      RECT 26.49 3.155 26.66 3.325 ;
      RECT 26.49 4.285 26.66 4.455 ;
      RECT 26.43 4.545 26.6 4.715 ;
      RECT 26.43 8.605 26.6 8.775 ;
      RECT 26.12 6.685 26.29 6.855 ;
      RECT 26.105 2.75 26.275 2.92 ;
      RECT 26.03 1.565 26.2 1.735 ;
      RECT 26.03 4.285 26.2 4.455 ;
      RECT 25.89 3.315 26.06 3.485 ;
      RECT 25.87 3.715 26.04 3.885 ;
      RECT 25.75 8.605 25.92 8.775 ;
      RECT 25.695 2.27 25.865 2.44 ;
      RECT 25.69 7.055 25.86 7.225 ;
      RECT 25.69 7.795 25.86 7.965 ;
      RECT 25.57 1.565 25.74 1.735 ;
      RECT 25.57 4.285 25.74 4.455 ;
      RECT 25.315 6.315 25.485 6.485 ;
      RECT 25.2 3.25 25.37 3.42 ;
      RECT 25.11 1.565 25.28 1.735 ;
      RECT 25.11 4.285 25.28 4.455 ;
      RECT 25.07 8.605 25.24 8.775 ;
      RECT 24.875 2.935 25.045 3.105 ;
      RECT 24.81 3.715 24.98 3.885 ;
      RECT 24.65 1.565 24.82 1.735 ;
      RECT 24.65 4.285 24.82 4.455 ;
      RECT 24.41 3.7 24.58 3.87 ;
      RECT 24.39 8.605 24.56 8.775 ;
      RECT 24.37 2.185 24.54 2.355 ;
      RECT 24.32 5.945 24.49 6.115 ;
      RECT 24.19 1.565 24.36 1.735 ;
      RECT 24.19 4.285 24.36 4.455 ;
      RECT 23.73 1.565 23.9 1.735 ;
      RECT 23.73 4.285 23.9 4.455 ;
      RECT 23.47 2.685 23.64 2.855 ;
      RECT 23.47 3.145 23.64 3.315 ;
      RECT 23.47 3.66 23.64 3.83 ;
      RECT 23.355 2.22 23.525 2.39 ;
      RECT 23.27 1.565 23.44 1.735 ;
      RECT 23.27 4.285 23.44 4.455 ;
      RECT 22.89 3.73 23.06 3.9 ;
      RECT 22.81 1.565 22.98 1.735 ;
      RECT 22.81 4.285 22.98 4.455 ;
      RECT 22.41 2.26 22.58 2.43 ;
      RECT 22.35 1.565 22.52 1.735 ;
      RECT 22.35 4.285 22.52 4.455 ;
      RECT 22.195 2.635 22.365 2.805 ;
      RECT 21.89 1.565 22.06 1.735 ;
      RECT 21.89 4.285 22.06 4.455 ;
      RECT 21.695 3.235 21.865 3.405 ;
      RECT 21.58 2.685 21.75 2.855 ;
      RECT 21.43 1.565 21.6 1.735 ;
      RECT 21.43 4.285 21.6 4.455 ;
      RECT 21.41 2.135 21.58 2.305 ;
      RECT 21.035 3.165 21.205 3.335 ;
      RECT 20.97 1.565 21.14 1.735 ;
      RECT 20.97 4.285 21.14 4.455 ;
      RECT 20.55 2.765 20.72 2.935 ;
      RECT 20.51 1.565 20.68 1.735 ;
      RECT 20.51 4.285 20.68 4.455 ;
      RECT 20.5 3.54 20.67 3.71 ;
      RECT 20.05 1.565 20.22 1.735 ;
      RECT 20.05 4.285 20.22 4.455 ;
      RECT 20.01 3.165 20.18 3.335 ;
      RECT 19.975 2.27 20.145 2.44 ;
      RECT 19.615 2.67 19.785 2.84 ;
      RECT 19.59 1.565 19.76 1.735 ;
      RECT 19.59 4.285 19.76 4.455 ;
      RECT 19.41 3.48 19.58 3.65 ;
      RECT 19.13 1.565 19.3 1.735 ;
      RECT 19.13 4.285 19.3 4.455 ;
      RECT 19.105 2.91 19.275 3.08 ;
      RECT 18.67 1.565 18.84 1.735 ;
      RECT 18.67 4.285 18.84 4.455 ;
      RECT 18.405 2.7 18.575 2.87 ;
      RECT 18.21 1.565 18.38 1.735 ;
      RECT 18.21 4.285 18.38 4.455 ;
      RECT 18.085 3.145 18.255 3.315 ;
      RECT 17.75 1.565 17.92 1.735 ;
      RECT 17.75 4.285 17.92 4.455 ;
      RECT 17.67 3.18 17.84 3.35 ;
      RECT 17.5 2.165 17.67 2.335 ;
      RECT 17.325 2.62 17.495 2.79 ;
      RECT 17.29 1.565 17.46 1.735 ;
      RECT 17.29 4.285 17.46 4.455 ;
      RECT 16.83 1.565 17 1.735 ;
      RECT 16.83 4.285 17 4.455 ;
      RECT 16.405 2.27 16.575 2.44 ;
      RECT 16.4 3.585 16.57 3.755 ;
      RECT 16.37 1.565 16.54 1.735 ;
      RECT 16.37 4.285 16.54 4.455 ;
      RECT 15.31 0.915 15.48 1.085 ;
      RECT 15.31 2.395 15.48 2.565 ;
      RECT 15.31 6.315 15.48 6.485 ;
      RECT 15.31 7.795 15.48 7.965 ;
      RECT 14.96 0.105 15.13 0.275 ;
      RECT 14.96 4.165 15.13 4.335 ;
      RECT 14.96 4.545 15.13 4.715 ;
      RECT 14.96 8.605 15.13 8.775 ;
      RECT 14.94 2.765 15.11 2.935 ;
      RECT 14.94 5.945 15.11 6.115 ;
      RECT 14.32 0.915 14.49 1.085 ;
      RECT 14.32 2.395 14.49 2.565 ;
      RECT 14.32 6.315 14.49 6.485 ;
      RECT 14.32 7.795 14.49 7.965 ;
      RECT 13.97 0.105 14.14 0.275 ;
      RECT 13.97 4.165 14.14 4.335 ;
      RECT 13.97 4.545 14.14 4.715 ;
      RECT 13.97 8.605 14.14 8.775 ;
      RECT 13.95 2.765 14.12 2.935 ;
      RECT 13.95 5.945 14.12 6.115 ;
      RECT 13.265 0.105 13.435 0.275 ;
      RECT 13.265 4.165 13.435 4.335 ;
      RECT 13.265 4.545 13.435 4.715 ;
      RECT 13.265 8.605 13.435 8.775 ;
      RECT 12.955 2.025 13.125 2.195 ;
      RECT 12.955 6.685 13.125 6.855 ;
      RECT 12.585 0.105 12.755 0.275 ;
      RECT 12.585 8.605 12.755 8.775 ;
      RECT 12.525 0.915 12.695 1.085 ;
      RECT 12.525 1.655 12.695 1.825 ;
      RECT 12.525 7.055 12.695 7.225 ;
      RECT 12.525 7.795 12.695 7.965 ;
      RECT 12.15 2.395 12.32 2.565 ;
      RECT 12.15 6.315 12.32 6.485 ;
      RECT 11.905 0.105 12.075 0.275 ;
      RECT 11.905 8.605 12.075 8.775 ;
      RECT 11.225 0.105 11.395 0.275 ;
      RECT 11.225 8.605 11.395 8.775 ;
      RECT 11.155 2.765 11.325 2.935 ;
      RECT 11.155 5.945 11.325 6.115 ;
      RECT 9.945 1.565 10.115 1.735 ;
      RECT 9.945 4.285 10.115 4.455 ;
      RECT 9.485 1.565 9.655 1.735 ;
      RECT 9.485 4.285 9.655 4.455 ;
      RECT 9.09 2.905 9.26 3.075 ;
      RECT 9.025 1.565 9.195 1.735 ;
      RECT 9.025 4.285 9.195 4.455 ;
      RECT 8.88 2.245 9.05 2.415 ;
      RECT 8.565 1.565 8.735 1.735 ;
      RECT 8.565 3.155 8.735 3.325 ;
      RECT 8.565 4.285 8.735 4.455 ;
      RECT 8.505 4.545 8.675 4.715 ;
      RECT 8.505 8.605 8.675 8.775 ;
      RECT 8.195 6.685 8.365 6.855 ;
      RECT 8.18 2.75 8.35 2.92 ;
      RECT 8.105 1.565 8.275 1.735 ;
      RECT 8.105 4.285 8.275 4.455 ;
      RECT 7.965 3.315 8.135 3.485 ;
      RECT 7.945 3.715 8.115 3.885 ;
      RECT 7.825 8.605 7.995 8.775 ;
      RECT 7.77 2.27 7.94 2.44 ;
      RECT 7.765 7.055 7.935 7.225 ;
      RECT 7.765 7.795 7.935 7.965 ;
      RECT 7.645 1.565 7.815 1.735 ;
      RECT 7.645 4.285 7.815 4.455 ;
      RECT 7.39 6.315 7.56 6.485 ;
      RECT 7.275 3.25 7.445 3.42 ;
      RECT 7.185 1.565 7.355 1.735 ;
      RECT 7.185 4.285 7.355 4.455 ;
      RECT 7.145 8.605 7.315 8.775 ;
      RECT 6.95 2.935 7.12 3.105 ;
      RECT 6.885 3.715 7.055 3.885 ;
      RECT 6.725 1.565 6.895 1.735 ;
      RECT 6.725 4.285 6.895 4.455 ;
      RECT 6.485 3.7 6.655 3.87 ;
      RECT 6.465 8.605 6.635 8.775 ;
      RECT 6.445 2.185 6.615 2.355 ;
      RECT 6.395 5.945 6.565 6.115 ;
      RECT 6.265 1.565 6.435 1.735 ;
      RECT 6.265 4.285 6.435 4.455 ;
      RECT 5.805 1.565 5.975 1.735 ;
      RECT 5.805 4.285 5.975 4.455 ;
      RECT 5.545 2.685 5.715 2.855 ;
      RECT 5.545 3.145 5.715 3.315 ;
      RECT 5.545 3.66 5.715 3.83 ;
      RECT 5.43 2.22 5.6 2.39 ;
      RECT 5.345 1.565 5.515 1.735 ;
      RECT 5.345 4.285 5.515 4.455 ;
      RECT 4.965 3.73 5.135 3.9 ;
      RECT 4.885 1.565 5.055 1.735 ;
      RECT 4.885 4.285 5.055 4.455 ;
      RECT 4.485 2.26 4.655 2.43 ;
      RECT 4.425 1.565 4.595 1.735 ;
      RECT 4.425 4.285 4.595 4.455 ;
      RECT 4.27 2.635 4.44 2.805 ;
      RECT 3.965 1.565 4.135 1.735 ;
      RECT 3.965 4.285 4.135 4.455 ;
      RECT 3.77 3.235 3.94 3.405 ;
      RECT 3.655 2.685 3.825 2.855 ;
      RECT 3.505 1.565 3.675 1.735 ;
      RECT 3.505 4.285 3.675 4.455 ;
      RECT 3.485 2.135 3.655 2.305 ;
      RECT 3.11 3.165 3.28 3.335 ;
      RECT 3.045 1.565 3.215 1.735 ;
      RECT 3.045 4.285 3.215 4.455 ;
      RECT 2.625 2.765 2.795 2.935 ;
      RECT 2.585 1.565 2.755 1.735 ;
      RECT 2.585 4.285 2.755 4.455 ;
      RECT 2.575 3.54 2.745 3.71 ;
      RECT 2.125 1.565 2.295 1.735 ;
      RECT 2.125 4.285 2.295 4.455 ;
      RECT 2.085 3.165 2.255 3.335 ;
      RECT 2.05 2.27 2.22 2.44 ;
      RECT 1.69 2.67 1.86 2.84 ;
      RECT 1.665 1.565 1.835 1.735 ;
      RECT 1.665 4.285 1.835 4.455 ;
      RECT 1.485 3.48 1.655 3.65 ;
      RECT 1.205 1.565 1.375 1.735 ;
      RECT 1.205 4.285 1.375 4.455 ;
      RECT 1.18 2.91 1.35 3.08 ;
      RECT 0.745 1.565 0.915 1.735 ;
      RECT 0.745 4.285 0.915 4.455 ;
      RECT 0.48 2.7 0.65 2.87 ;
      RECT 0.285 1.565 0.455 1.735 ;
      RECT 0.285 4.285 0.455 4.455 ;
      RECT 0.16 3.145 0.33 3.315 ;
      RECT -0.175 1.565 -0.005 1.735 ;
      RECT -0.175 4.285 -0.005 4.455 ;
      RECT -0.255 3.18 -0.085 3.35 ;
      RECT -0.425 2.165 -0.255 2.335 ;
      RECT -0.6 2.62 -0.43 2.79 ;
      RECT -0.635 1.565 -0.465 1.735 ;
      RECT -0.635 4.285 -0.465 4.455 ;
      RECT -1.095 1.565 -0.925 1.735 ;
      RECT -1.095 4.285 -0.925 4.455 ;
      RECT -1.52 2.27 -1.35 2.44 ;
      RECT -1.525 3.585 -1.355 3.755 ;
      RECT -1.555 1.565 -1.385 1.735 ;
      RECT -1.555 4.285 -1.385 4.455 ;
      RECT -2.525 4.545 -2.355 4.715 ;
      RECT -2.525 8.605 -2.355 8.775 ;
      RECT -2.835 6.685 -2.665 6.855 ;
      RECT -3.205 8.605 -3.035 8.775 ;
      RECT -3.265 7.055 -3.095 7.225 ;
      RECT -3.265 7.795 -3.095 7.965 ;
      RECT -3.64 6.315 -3.47 6.485 ;
      RECT -3.885 8.605 -3.715 8.775 ;
      RECT -4.565 8.605 -4.395 8.775 ;
      RECT -4.635 5.945 -4.465 6.115 ;
    LAYER li ;
      RECT 81.05 0 81.22 2.235 ;
      RECT 80.09 0 80.26 2.235 ;
      RECT 79.13 0 79.3 2.235 ;
      RECT 78.61 0 78.78 2.235 ;
      RECT 77.65 0 77.82 2.235 ;
      RECT 76.65 0 76.82 2.235 ;
      RECT 75.69 0 75.86 2.235 ;
      RECT 74.21 0 74.38 2.235 ;
      RECT 72.29 0 72.46 2.235 ;
      RECT 70.81 0 70.98 2.235 ;
      RECT 63.125 0 63.295 2.235 ;
      RECT 62.165 0 62.335 2.235 ;
      RECT 61.205 0 61.375 2.235 ;
      RECT 60.685 0 60.855 2.235 ;
      RECT 59.725 0 59.895 2.235 ;
      RECT 58.725 0 58.895 2.235 ;
      RECT 57.765 0 57.935 2.235 ;
      RECT 56.285 0 56.455 2.235 ;
      RECT 54.365 0 54.535 2.235 ;
      RECT 52.885 0 53.055 2.235 ;
      RECT 45.2 0 45.37 2.235 ;
      RECT 44.24 0 44.41 2.235 ;
      RECT 43.28 0 43.45 2.235 ;
      RECT 42.76 0 42.93 2.235 ;
      RECT 41.8 0 41.97 2.235 ;
      RECT 40.8 0 40.97 2.235 ;
      RECT 39.84 0 40.01 2.235 ;
      RECT 38.36 0 38.53 2.235 ;
      RECT 36.44 0 36.61 2.235 ;
      RECT 34.96 0 35.13 2.235 ;
      RECT 27.275 0 27.445 2.235 ;
      RECT 26.315 0 26.485 2.235 ;
      RECT 25.355 0 25.525 2.235 ;
      RECT 24.835 0 25.005 2.235 ;
      RECT 23.875 0 24.045 2.235 ;
      RECT 22.875 0 23.045 2.235 ;
      RECT 21.915 0 22.085 2.235 ;
      RECT 20.435 0 20.605 2.235 ;
      RECT 18.515 0 18.685 2.235 ;
      RECT 17.035 0 17.205 2.235 ;
      RECT 9.35 0 9.52 2.235 ;
      RECT 8.39 0 8.56 2.235 ;
      RECT 7.43 0 7.6 2.235 ;
      RECT 6.91 0 7.08 2.235 ;
      RECT 5.95 0 6.12 2.235 ;
      RECT 4.95 0 5.12 2.235 ;
      RECT 3.99 0 4.16 2.235 ;
      RECT 2.51 0 2.68 2.235 ;
      RECT 0.59 0 0.76 2.235 ;
      RECT -0.89 0 -0.72 2.235 ;
      RECT 70 0 81.96 1.735 ;
      RECT 52.075 0 64.035 1.735 ;
      RECT 34.15 0 46.11 1.735 ;
      RECT 16.225 0 28.185 1.735 ;
      RECT -1.7 0 10.26 1.735 ;
      RECT 69.995 0 81.96 1.68 ;
      RECT 52.07 0 64.035 1.68 ;
      RECT 34.145 0 46.11 1.68 ;
      RECT 16.22 0 28.185 1.68 ;
      RECT -1.705 0 10.26 1.68 ;
      RECT 86.58 0 86.75 0.935 ;
      RECT 85.59 0 85.76 0.935 ;
      RECT 82.845 0 83.015 0.935 ;
      RECT 68.655 0 68.825 0.935 ;
      RECT 67.665 0 67.835 0.935 ;
      RECT 64.92 0 65.09 0.935 ;
      RECT 50.73 0 50.9 0.935 ;
      RECT 49.74 0 49.91 0.935 ;
      RECT 46.995 0 47.165 0.935 ;
      RECT 32.805 0 32.975 0.935 ;
      RECT 31.815 0 31.985 0.935 ;
      RECT 29.07 0 29.24 0.935 ;
      RECT 14.88 0 15.05 0.935 ;
      RECT 13.89 0 14.06 0.935 ;
      RECT 11.145 0 11.315 0.935 ;
      RECT -4.865 0 87.55 0.305 ;
      RECT -2.835 4.285 -2.665 8.305 ;
      RECT 86.58 3.405 86.75 5.475 ;
      RECT 85.59 3.405 85.76 5.475 ;
      RECT 82.845 3.405 83.015 5.475 ;
      RECT 78.085 4.285 78.255 5.475 ;
      RECT 68.655 3.405 68.825 5.475 ;
      RECT 67.665 3.405 67.835 5.475 ;
      RECT 64.92 3.405 65.09 5.475 ;
      RECT 60.16 4.285 60.33 5.475 ;
      RECT 50.73 3.405 50.9 5.475 ;
      RECT 49.74 3.405 49.91 5.475 ;
      RECT 46.995 3.405 47.165 5.475 ;
      RECT 42.235 4.285 42.405 5.475 ;
      RECT 32.805 3.405 32.975 5.475 ;
      RECT 31.815 3.405 31.985 5.475 ;
      RECT 29.07 3.405 29.24 5.475 ;
      RECT 24.31 4.285 24.48 5.475 ;
      RECT 14.88 3.405 15.05 5.475 ;
      RECT 13.89 3.405 14.06 5.475 ;
      RECT 11.145 3.405 11.315 5.475 ;
      RECT 6.385 4.285 6.555 5.475 ;
      RECT -4.645 4.285 -4.475 5.475 ;
      RECT -4.865 4.285 87.55 4.745 ;
      RECT 81.59 4.135 87.55 4.745 ;
      RECT 80.09 3.785 80.26 4.745 ;
      RECT 77.65 3.785 77.82 4.745 ;
      RECT 75.69 3.785 75.86 4.745 ;
      RECT 74.73 3.785 74.9 4.745 ;
      RECT 72.77 3.785 72.94 4.745 ;
      RECT 71.77 3.785 71.94 4.745 ;
      RECT 70.81 3.785 70.98 4.745 ;
      RECT 63.665 4.135 69.625 4.745 ;
      RECT 62.165 3.785 62.335 4.745 ;
      RECT 59.725 3.785 59.895 4.745 ;
      RECT 57.765 3.785 57.935 4.745 ;
      RECT 56.805 3.785 56.975 4.745 ;
      RECT 54.845 3.785 55.015 4.745 ;
      RECT 53.845 3.785 54.015 4.745 ;
      RECT 52.885 3.785 53.055 4.745 ;
      RECT 45.74 4.135 51.7 4.745 ;
      RECT 44.24 3.785 44.41 4.745 ;
      RECT 41.8 3.785 41.97 4.745 ;
      RECT 39.84 3.785 40.01 4.745 ;
      RECT 38.88 3.785 39.05 4.745 ;
      RECT 36.92 3.785 37.09 4.745 ;
      RECT 35.92 3.785 36.09 4.745 ;
      RECT 34.96 3.785 35.13 4.745 ;
      RECT 27.815 4.135 33.775 4.745 ;
      RECT 26.315 3.785 26.485 4.745 ;
      RECT 23.875 3.785 24.045 4.745 ;
      RECT 21.915 3.785 22.085 4.745 ;
      RECT 20.955 3.785 21.125 4.745 ;
      RECT 18.995 3.785 19.165 4.745 ;
      RECT 17.995 3.785 18.165 4.745 ;
      RECT 17.035 3.785 17.205 4.745 ;
      RECT 9.89 4.135 15.85 4.745 ;
      RECT 8.39 3.785 8.56 4.745 ;
      RECT 5.95 3.785 6.12 4.745 ;
      RECT 3.99 3.785 4.16 4.745 ;
      RECT 3.03 3.785 3.2 4.745 ;
      RECT 1.07 3.785 1.24 4.745 ;
      RECT 0.07 3.785 0.24 4.745 ;
      RECT -0.89 3.785 -0.72 4.745 ;
      RECT -4.885 8.575 87.55 8.88 ;
      RECT 86.58 7.945 86.75 8.88 ;
      RECT 85.59 7.945 85.76 8.88 ;
      RECT 82.845 7.945 83.015 8.88 ;
      RECT 78.085 7.945 78.255 8.88 ;
      RECT 68.655 7.945 68.825 8.88 ;
      RECT 67.665 7.945 67.835 8.88 ;
      RECT 64.92 7.945 65.09 8.88 ;
      RECT 60.16 7.945 60.33 8.88 ;
      RECT 50.73 7.945 50.9 8.88 ;
      RECT 49.74 7.945 49.91 8.88 ;
      RECT 46.995 7.945 47.165 8.88 ;
      RECT 42.235 7.945 42.405 8.88 ;
      RECT 32.805 7.945 32.975 8.88 ;
      RECT 31.815 7.945 31.985 8.88 ;
      RECT 29.07 7.945 29.24 8.88 ;
      RECT 24.31 7.945 24.48 8.88 ;
      RECT 14.88 7.945 15.05 8.88 ;
      RECT 13.89 7.945 14.06 8.88 ;
      RECT 11.145 7.945 11.315 8.88 ;
      RECT 6.385 7.945 6.555 8.88 ;
      RECT -4.645 7.945 -4.475 8.88 ;
      RECT 86.64 1.74 86.81 2.935 ;
      RECT 86.64 1.74 87.105 1.91 ;
      RECT 86.64 6.97 87.105 7.14 ;
      RECT 86.64 5.945 86.81 7.14 ;
      RECT 85.65 1.74 85.82 2.935 ;
      RECT 85.65 1.74 86.115 1.91 ;
      RECT 85.65 6.97 86.115 7.14 ;
      RECT 85.65 5.945 85.82 7.14 ;
      RECT 83.795 2.635 83.965 3.865 ;
      RECT 83.85 0.855 84.02 2.805 ;
      RECT 83.795 0.575 83.965 1.025 ;
      RECT 83.795 7.855 83.965 8.305 ;
      RECT 83.85 6.075 84.02 8.025 ;
      RECT 83.795 5.015 83.965 6.245 ;
      RECT 83.275 0.575 83.445 3.865 ;
      RECT 83.275 2.075 83.68 2.405 ;
      RECT 83.275 1.235 83.68 1.565 ;
      RECT 83.275 5.015 83.445 8.305 ;
      RECT 83.275 7.315 83.68 7.645 ;
      RECT 83.275 6.475 83.68 6.805 ;
      RECT 81.375 3.392 81.39 3.443 ;
      RECT 81.37 3.372 81.375 3.49 ;
      RECT 81.355 3.362 81.37 3.558 ;
      RECT 81.33 3.342 81.355 3.613 ;
      RECT 81.29 3.327 81.33 3.633 ;
      RECT 81.245 3.321 81.29 3.661 ;
      RECT 81.175 3.311 81.245 3.678 ;
      RECT 81.155 3.303 81.175 3.678 ;
      RECT 81.095 3.297 81.155 3.67 ;
      RECT 81.036 3.288 81.095 3.658 ;
      RECT 80.95 3.277 81.036 3.641 ;
      RECT 80.928 3.268 80.95 3.629 ;
      RECT 80.842 3.261 80.928 3.616 ;
      RECT 80.756 3.248 80.842 3.597 ;
      RECT 80.67 3.236 80.756 3.577 ;
      RECT 80.64 3.225 80.67 3.564 ;
      RECT 80.59 3.211 80.64 3.556 ;
      RECT 80.57 3.2 80.59 3.548 ;
      RECT 80.521 3.189 80.57 3.54 ;
      RECT 80.435 3.168 80.521 3.525 ;
      RECT 80.39 3.155 80.435 3.51 ;
      RECT 80.345 3.155 80.39 3.49 ;
      RECT 80.29 3.155 80.345 3.425 ;
      RECT 80.265 3.155 80.29 3.348 ;
      RECT 80.79 2.892 80.96 3.075 ;
      RECT 80.79 2.892 80.975 3.033 ;
      RECT 80.79 2.892 80.98 2.975 ;
      RECT 80.85 2.66 80.985 2.951 ;
      RECT 80.85 2.664 80.99 2.934 ;
      RECT 80.795 2.827 80.99 2.934 ;
      RECT 80.82 2.672 80.96 3.075 ;
      RECT 80.82 2.676 81 2.875 ;
      RECT 80.805 2.762 81 2.875 ;
      RECT 80.815 2.692 80.96 3.075 ;
      RECT 80.815 2.695 81.01 2.788 ;
      RECT 80.81 2.712 81.01 2.788 ;
      RECT 80.58 1.932 80.75 2.415 ;
      RECT 80.575 1.927 80.725 2.405 ;
      RECT 80.575 1.934 80.755 2.399 ;
      RECT 80.565 1.928 80.725 2.378 ;
      RECT 80.565 1.944 80.77 2.337 ;
      RECT 80.535 1.929 80.725 2.3 ;
      RECT 80.535 1.959 80.78 2.24 ;
      RECT 80.53 1.931 80.725 2.238 ;
      RECT 80.51 1.94 80.755 2.195 ;
      RECT 80.485 1.956 80.77 2.107 ;
      RECT 80.485 1.975 80.795 2.098 ;
      RECT 80.48 2.012 80.795 2.05 ;
      RECT 80.485 1.992 80.8 2.018 ;
      RECT 80.58 1.926 80.69 2.415 ;
      RECT 80.666 1.925 80.69 2.415 ;
      RECT 79.9 2.71 79.905 2.921 ;
      RECT 80.5 2.71 80.505 2.895 ;
      RECT 80.565 2.75 80.57 2.863 ;
      RECT 80.56 2.742 80.565 2.869 ;
      RECT 80.555 2.732 80.56 2.877 ;
      RECT 80.55 2.722 80.555 2.886 ;
      RECT 80.545 2.712 80.55 2.89 ;
      RECT 80.505 2.71 80.545 2.893 ;
      RECT 80.477 2.709 80.5 2.897 ;
      RECT 80.391 2.706 80.477 2.904 ;
      RECT 80.305 2.702 80.391 2.915 ;
      RECT 80.285 2.7 80.305 2.921 ;
      RECT 80.267 2.699 80.285 2.924 ;
      RECT 80.181 2.697 80.267 2.931 ;
      RECT 80.095 2.692 80.181 2.944 ;
      RECT 80.076 2.689 80.095 2.949 ;
      RECT 79.99 2.687 80.076 2.94 ;
      RECT 79.98 2.687 79.99 2.933 ;
      RECT 79.905 2.7 79.98 2.927 ;
      RECT 79.89 2.711 79.9 2.921 ;
      RECT 79.88 2.713 79.89 2.92 ;
      RECT 79.87 2.717 79.88 2.916 ;
      RECT 79.865 2.72 79.87 2.91 ;
      RECT 79.855 2.722 79.865 2.904 ;
      RECT 79.85 2.725 79.855 2.898 ;
      RECT 79.83 3.311 79.835 3.515 ;
      RECT 79.815 3.298 79.83 3.608 ;
      RECT 79.8 3.279 79.815 3.885 ;
      RECT 79.765 3.245 79.8 3.885 ;
      RECT 79.761 3.215 79.765 3.885 ;
      RECT 79.675 3.097 79.761 3.885 ;
      RECT 79.665 2.972 79.675 3.885 ;
      RECT 79.65 2.94 79.665 3.885 ;
      RECT 79.645 2.915 79.65 3.885 ;
      RECT 79.64 2.905 79.645 3.841 ;
      RECT 79.625 2.877 79.64 3.746 ;
      RECT 79.61 2.843 79.625 3.645 ;
      RECT 79.605 2.821 79.61 3.598 ;
      RECT 79.6 2.81 79.605 3.568 ;
      RECT 79.595 2.8 79.6 3.534 ;
      RECT 79.585 2.787 79.595 3.502 ;
      RECT 79.56 2.763 79.585 3.428 ;
      RECT 79.555 2.743 79.56 3.353 ;
      RECT 79.55 2.737 79.555 3.328 ;
      RECT 79.545 2.732 79.55 3.293 ;
      RECT 79.54 2.727 79.545 3.268 ;
      RECT 79.535 2.725 79.54 3.248 ;
      RECT 79.53 2.725 79.535 3.233 ;
      RECT 79.525 2.725 79.53 3.193 ;
      RECT 79.515 2.725 79.525 3.165 ;
      RECT 79.505 2.725 79.515 3.11 ;
      RECT 79.49 2.725 79.505 3.048 ;
      RECT 79.485 2.724 79.49 2.993 ;
      RECT 79.47 2.723 79.485 2.973 ;
      RECT 79.41 2.721 79.47 2.947 ;
      RECT 79.375 2.722 79.41 2.927 ;
      RECT 79.37 2.724 79.375 2.917 ;
      RECT 79.36 2.743 79.37 2.907 ;
      RECT 79.355 2.77 79.36 2.838 ;
      RECT 79.47 2.195 79.64 2.44 ;
      RECT 79.505 1.966 79.64 2.44 ;
      RECT 79.505 1.968 79.65 2.435 ;
      RECT 79.505 1.97 79.675 2.423 ;
      RECT 79.505 1.973 79.7 2.405 ;
      RECT 79.505 1.978 79.75 2.378 ;
      RECT 79.505 1.983 79.77 2.343 ;
      RECT 79.485 1.985 79.78 2.318 ;
      RECT 79.475 2.08 79.78 2.318 ;
      RECT 79.505 1.965 79.615 2.44 ;
      RECT 79.515 1.962 79.61 2.44 ;
      RECT 79.035 3.227 79.225 3.585 ;
      RECT 79.035 3.239 79.26 3.584 ;
      RECT 79.035 3.267 79.28 3.582 ;
      RECT 79.035 3.292 79.285 3.581 ;
      RECT 79.035 3.35 79.3 3.58 ;
      RECT 79.02 3.223 79.18 3.565 ;
      RECT 79 3.232 79.225 3.518 ;
      RECT 78.975 3.243 79.26 3.455 ;
      RECT 78.975 3.327 79.295 3.455 ;
      RECT 78.975 3.302 79.29 3.455 ;
      RECT 79.035 3.218 79.18 3.585 ;
      RECT 79.121 3.217 79.18 3.585 ;
      RECT 79.121 3.216 79.165 3.585 ;
      RECT 79.035 7.855 79.205 8.305 ;
      RECT 79.09 6.075 79.26 8.025 ;
      RECT 79.035 5.015 79.205 6.245 ;
      RECT 78.515 5.015 78.685 8.305 ;
      RECT 78.515 7.315 78.92 7.645 ;
      RECT 78.515 6.475 78.92 6.805 ;
      RECT 78.82 2.732 78.825 3.11 ;
      RECT 78.815 2.7 78.82 3.11 ;
      RECT 78.81 2.672 78.815 3.11 ;
      RECT 78.805 2.652 78.81 3.11 ;
      RECT 78.75 2.635 78.805 3.11 ;
      RECT 78.71 2.62 78.75 3.11 ;
      RECT 78.655 2.607 78.71 3.11 ;
      RECT 78.62 2.598 78.655 3.11 ;
      RECT 78.616 2.596 78.62 3.109 ;
      RECT 78.53 2.592 78.616 3.092 ;
      RECT 78.445 2.584 78.53 3.055 ;
      RECT 78.435 2.58 78.445 3.028 ;
      RECT 78.425 2.58 78.435 3.01 ;
      RECT 78.415 2.582 78.425 2.993 ;
      RECT 78.41 2.587 78.415 2.979 ;
      RECT 78.405 2.591 78.41 2.966 ;
      RECT 78.395 2.596 78.405 2.95 ;
      RECT 78.38 2.61 78.395 2.925 ;
      RECT 78.375 2.616 78.38 2.905 ;
      RECT 78.37 2.618 78.375 2.898 ;
      RECT 78.365 2.622 78.37 2.773 ;
      RECT 78.545 3.422 78.79 3.885 ;
      RECT 78.465 3.395 78.785 3.881 ;
      RECT 78.395 3.43 78.79 3.874 ;
      RECT 78.185 3.685 78.79 3.87 ;
      RECT 78.365 3.453 78.79 3.87 ;
      RECT 78.205 3.645 78.79 3.87 ;
      RECT 78.355 3.465 78.79 3.87 ;
      RECT 78.24 3.582 78.79 3.87 ;
      RECT 78.295 3.507 78.79 3.87 ;
      RECT 78.545 3.372 78.785 3.885 ;
      RECT 78.575 3.365 78.785 3.885 ;
      RECT 78.565 3.367 78.785 3.885 ;
      RECT 78.575 3.362 78.705 3.885 ;
      RECT 78.13 1.925 78.216 2.364 ;
      RECT 78.125 1.925 78.216 2.362 ;
      RECT 78.125 1.925 78.285 2.361 ;
      RECT 78.125 1.925 78.315 2.358 ;
      RECT 78.11 1.932 78.315 2.349 ;
      RECT 78.11 1.932 78.32 2.345 ;
      RECT 78.105 1.942 78.32 2.338 ;
      RECT 78.1 1.947 78.32 2.313 ;
      RECT 78.1 1.947 78.335 2.295 ;
      RECT 78.125 1.925 78.355 2.21 ;
      RECT 78.095 1.952 78.355 2.208 ;
      RECT 78.105 1.945 78.36 2.146 ;
      RECT 78.095 2.067 78.365 2.129 ;
      RECT 78.08 1.962 78.36 2.08 ;
      RECT 78.075 1.972 78.36 1.98 ;
      RECT 78.155 2.743 78.16 2.82 ;
      RECT 78.145 2.737 78.155 3.01 ;
      RECT 78.135 2.729 78.145 3.031 ;
      RECT 78.125 2.72 78.135 3.053 ;
      RECT 78.12 2.715 78.125 3.07 ;
      RECT 78.08 2.715 78.12 3.11 ;
      RECT 78.06 2.715 78.08 3.165 ;
      RECT 78.055 2.715 78.06 3.193 ;
      RECT 78.045 2.715 78.055 3.208 ;
      RECT 78.01 2.715 78.045 3.25 ;
      RECT 78.005 2.715 78.01 3.293 ;
      RECT 77.995 2.715 78.005 3.308 ;
      RECT 77.98 2.715 77.995 3.328 ;
      RECT 77.965 2.715 77.98 3.355 ;
      RECT 77.96 2.716 77.965 3.373 ;
      RECT 77.94 2.717 77.96 3.38 ;
      RECT 77.885 2.718 77.94 3.4 ;
      RECT 77.875 2.719 77.885 3.414 ;
      RECT 77.87 2.722 77.875 3.413 ;
      RECT 77.83 2.795 77.87 3.411 ;
      RECT 77.815 2.875 77.83 3.409 ;
      RECT 77.79 2.93 77.815 3.407 ;
      RECT 77.775 2.995 77.79 3.406 ;
      RECT 77.73 3.027 77.775 3.403 ;
      RECT 77.645 3.05 77.73 3.398 ;
      RECT 77.62 3.07 77.645 3.393 ;
      RECT 77.55 3.075 77.62 3.389 ;
      RECT 77.53 3.077 77.55 3.386 ;
      RECT 77.445 3.088 77.53 3.38 ;
      RECT 77.44 3.099 77.445 3.375 ;
      RECT 77.43 3.101 77.44 3.375 ;
      RECT 77.395 3.105 77.43 3.373 ;
      RECT 77.345 3.115 77.395 3.36 ;
      RECT 77.325 3.123 77.345 3.345 ;
      RECT 77.245 3.135 77.325 3.328 ;
      RECT 77.41 2.685 77.58 2.895 ;
      RECT 77.526 2.681 77.58 2.895 ;
      RECT 77.331 2.685 77.58 2.886 ;
      RECT 77.331 2.685 77.585 2.875 ;
      RECT 77.245 2.685 77.585 2.866 ;
      RECT 77.245 2.693 77.595 2.81 ;
      RECT 77.245 2.705 77.6 2.723 ;
      RECT 77.245 2.712 77.605 2.715 ;
      RECT 77.44 2.683 77.58 2.895 ;
      RECT 77.195 3.628 77.44 3.96 ;
      RECT 77.19 3.62 77.195 3.957 ;
      RECT 77.16 3.64 77.44 3.938 ;
      RECT 77.14 3.672 77.44 3.911 ;
      RECT 77.19 3.625 77.367 3.957 ;
      RECT 77.19 3.622 77.281 3.957 ;
      RECT 77.13 1.97 77.3 2.39 ;
      RECT 77.125 1.97 77.3 2.388 ;
      RECT 77.125 1.97 77.325 2.378 ;
      RECT 77.125 1.97 77.345 2.353 ;
      RECT 77.12 1.97 77.345 2.348 ;
      RECT 77.12 1.97 77.355 2.338 ;
      RECT 77.12 1.97 77.36 2.333 ;
      RECT 77.12 1.975 77.365 2.328 ;
      RECT 77.12 2.007 77.38 2.318 ;
      RECT 77.12 2.077 77.405 2.301 ;
      RECT 77.1 2.077 77.405 2.293 ;
      RECT 77.1 2.137 77.415 2.27 ;
      RECT 77.1 2.177 77.425 2.215 ;
      RECT 77.085 1.97 77.36 2.195 ;
      RECT 77.075 1.985 77.365 2.093 ;
      RECT 76.665 3.375 76.835 3.9 ;
      RECT 76.66 3.375 76.835 3.893 ;
      RECT 76.65 3.375 76.84 3.858 ;
      RECT 76.645 3.385 76.84 3.83 ;
      RECT 76.64 3.405 76.84 3.813 ;
      RECT 76.65 3.38 76.845 3.803 ;
      RECT 76.635 3.425 76.845 3.795 ;
      RECT 76.63 3.445 76.845 3.78 ;
      RECT 76.625 3.475 76.845 3.77 ;
      RECT 76.615 3.52 76.845 3.745 ;
      RECT 76.645 3.39 76.85 3.728 ;
      RECT 76.61 3.572 76.85 3.723 ;
      RECT 76.645 3.4 76.855 3.693 ;
      RECT 76.605 3.605 76.855 3.69 ;
      RECT 76.6 3.63 76.855 3.67 ;
      RECT 76.64 3.417 76.865 3.61 ;
      RECT 76.635 3.439 76.875 3.503 ;
      RECT 76.585 2.686 76.6 2.955 ;
      RECT 76.54 2.67 76.585 3 ;
      RECT 76.535 2.658 76.54 3.05 ;
      RECT 76.525 2.654 76.535 3.083 ;
      RECT 76.52 2.651 76.525 3.111 ;
      RECT 76.505 2.653 76.52 3.153 ;
      RECT 76.5 2.657 76.505 3.193 ;
      RECT 76.48 2.662 76.5 3.245 ;
      RECT 76.476 2.667 76.48 3.302 ;
      RECT 76.39 2.686 76.476 3.339 ;
      RECT 76.38 2.707 76.39 3.375 ;
      RECT 76.375 2.715 76.38 3.376 ;
      RECT 76.37 2.757 76.375 3.377 ;
      RECT 76.355 2.845 76.37 3.378 ;
      RECT 76.345 2.995 76.355 3.38 ;
      RECT 76.34 3.04 76.345 3.382 ;
      RECT 76.305 3.082 76.34 3.385 ;
      RECT 76.3 3.1 76.305 3.388 ;
      RECT 76.223 3.106 76.3 3.394 ;
      RECT 76.137 3.12 76.223 3.407 ;
      RECT 76.051 3.134 76.137 3.421 ;
      RECT 75.965 3.148 76.051 3.434 ;
      RECT 75.905 3.16 75.965 3.446 ;
      RECT 75.88 3.167 75.905 3.453 ;
      RECT 75.866 3.17 75.88 3.458 ;
      RECT 75.78 3.178 75.866 3.474 ;
      RECT 75.775 3.185 75.78 3.489 ;
      RECT 75.751 3.185 75.775 3.496 ;
      RECT 75.665 3.188 75.751 3.524 ;
      RECT 75.58 3.192 75.665 3.568 ;
      RECT 75.515 3.196 75.58 3.605 ;
      RECT 75.49 3.199 75.515 3.621 ;
      RECT 75.415 3.212 75.49 3.625 ;
      RECT 75.39 3.23 75.415 3.629 ;
      RECT 75.38 3.237 75.39 3.631 ;
      RECT 75.365 3.24 75.38 3.632 ;
      RECT 75.305 3.252 75.365 3.636 ;
      RECT 75.295 3.266 75.305 3.64 ;
      RECT 75.24 3.276 75.295 3.628 ;
      RECT 75.215 3.297 75.24 3.611 ;
      RECT 75.195 3.317 75.215 3.602 ;
      RECT 75.19 3.33 75.195 3.597 ;
      RECT 75.175 3.342 75.19 3.593 ;
      RECT 76.41 1.997 76.415 2.02 ;
      RECT 76.405 1.988 76.41 2.06 ;
      RECT 76.4 1.986 76.405 2.103 ;
      RECT 76.395 1.977 76.4 2.138 ;
      RECT 76.39 1.967 76.395 2.21 ;
      RECT 76.385 1.957 76.39 2.275 ;
      RECT 76.38 1.954 76.385 2.315 ;
      RECT 76.355 1.948 76.38 2.405 ;
      RECT 76.32 1.936 76.355 2.43 ;
      RECT 76.31 1.927 76.32 2.43 ;
      RECT 76.175 1.925 76.185 2.413 ;
      RECT 76.165 1.925 76.175 2.38 ;
      RECT 76.16 1.925 76.165 2.355 ;
      RECT 76.155 1.925 76.16 2.343 ;
      RECT 76.15 1.925 76.155 2.325 ;
      RECT 76.14 1.925 76.15 2.29 ;
      RECT 76.135 1.927 76.14 2.268 ;
      RECT 76.13 1.933 76.135 2.253 ;
      RECT 76.125 1.939 76.13 2.238 ;
      RECT 76.11 1.951 76.125 2.211 ;
      RECT 76.105 1.962 76.11 2.179 ;
      RECT 76.1 1.972 76.105 2.163 ;
      RECT 76.09 1.98 76.1 2.132 ;
      RECT 76.085 1.99 76.09 2.106 ;
      RECT 76.08 2.047 76.085 2.089 ;
      RECT 76.185 1.925 76.31 2.43 ;
      RECT 75.9 2.612 76.16 2.91 ;
      RECT 75.895 2.619 76.16 2.908 ;
      RECT 75.9 2.614 76.175 2.903 ;
      RECT 75.89 2.627 76.175 2.9 ;
      RECT 75.89 2.632 76.18 2.893 ;
      RECT 75.885 2.64 76.18 2.89 ;
      RECT 75.885 2.657 76.185 2.688 ;
      RECT 75.9 2.609 76.131 2.91 ;
      RECT 75.955 2.608 76.131 2.91 ;
      RECT 75.955 2.605 76.045 2.91 ;
      RECT 75.955 2.602 76.041 2.91 ;
      RECT 75.645 2.875 75.65 2.888 ;
      RECT 75.64 2.842 75.645 2.893 ;
      RECT 75.635 2.797 75.64 2.9 ;
      RECT 75.63 2.752 75.635 2.908 ;
      RECT 75.625 2.72 75.63 2.916 ;
      RECT 75.62 2.68 75.625 2.917 ;
      RECT 75.605 2.66 75.62 2.919 ;
      RECT 75.53 2.642 75.605 2.931 ;
      RECT 75.52 2.635 75.53 2.942 ;
      RECT 75.515 2.635 75.52 2.944 ;
      RECT 75.485 2.641 75.515 2.948 ;
      RECT 75.445 2.654 75.485 2.948 ;
      RECT 75.42 2.665 75.445 2.934 ;
      RECT 75.405 2.671 75.42 2.917 ;
      RECT 75.395 2.673 75.405 2.908 ;
      RECT 75.39 2.674 75.395 2.903 ;
      RECT 75.385 2.675 75.39 2.898 ;
      RECT 75.38 2.676 75.385 2.895 ;
      RECT 75.355 2.681 75.38 2.885 ;
      RECT 75.345 2.697 75.355 2.872 ;
      RECT 75.34 2.717 75.345 2.867 ;
      RECT 75.35 2.11 75.355 2.306 ;
      RECT 75.335 2.074 75.35 2.308 ;
      RECT 75.325 2.056 75.335 2.313 ;
      RECT 75.315 2.042 75.325 2.317 ;
      RECT 75.27 2.026 75.315 2.327 ;
      RECT 75.265 2.016 75.27 2.336 ;
      RECT 75.22 2.005 75.265 2.342 ;
      RECT 75.215 1.993 75.22 2.349 ;
      RECT 75.2 1.988 75.215 2.353 ;
      RECT 75.185 1.98 75.2 2.358 ;
      RECT 75.175 1.973 75.185 2.363 ;
      RECT 75.165 1.97 75.175 2.368 ;
      RECT 75.155 1.97 75.165 2.369 ;
      RECT 75.15 1.967 75.155 2.368 ;
      RECT 75.115 1.962 75.14 2.367 ;
      RECT 75.091 1.958 75.115 2.366 ;
      RECT 75.005 1.949 75.091 2.363 ;
      RECT 74.99 1.941 75.005 2.36 ;
      RECT 74.968 1.94 74.99 2.359 ;
      RECT 74.882 1.94 74.968 2.357 ;
      RECT 74.796 1.94 74.882 2.355 ;
      RECT 74.71 1.94 74.796 2.352 ;
      RECT 74.7 1.94 74.71 2.343 ;
      RECT 74.67 1.94 74.7 2.303 ;
      RECT 74.66 1.95 74.67 2.258 ;
      RECT 74.655 1.99 74.66 2.243 ;
      RECT 74.65 2.005 74.655 2.23 ;
      RECT 74.62 2.085 74.65 2.192 ;
      RECT 75.14 1.965 75.15 2.368 ;
      RECT 74.965 2.73 74.98 3.335 ;
      RECT 74.97 2.725 74.98 3.335 ;
      RECT 75.135 2.725 75.14 2.908 ;
      RECT 75.125 2.725 75.135 2.938 ;
      RECT 75.11 2.725 75.125 2.998 ;
      RECT 75.105 2.725 75.11 3.043 ;
      RECT 75.1 2.725 75.105 3.073 ;
      RECT 75.095 2.725 75.1 3.093 ;
      RECT 75.085 2.725 75.095 3.128 ;
      RECT 75.07 2.725 75.085 3.16 ;
      RECT 75.025 2.725 75.07 3.188 ;
      RECT 75.02 2.725 75.025 3.218 ;
      RECT 75.015 2.725 75.02 3.23 ;
      RECT 75.01 2.725 75.015 3.238 ;
      RECT 75 2.725 75.01 3.253 ;
      RECT 74.995 2.725 75 3.275 ;
      RECT 74.985 2.725 74.995 3.298 ;
      RECT 74.98 2.725 74.985 3.318 ;
      RECT 74.945 2.74 74.965 3.335 ;
      RECT 74.92 2.757 74.945 3.335 ;
      RECT 74.915 2.767 74.92 3.335 ;
      RECT 74.885 2.782 74.915 3.335 ;
      RECT 74.81 2.824 74.885 3.335 ;
      RECT 74.805 2.855 74.81 3.318 ;
      RECT 74.8 2.859 74.805 3.3 ;
      RECT 74.795 2.863 74.8 3.263 ;
      RECT 74.79 3.047 74.795 3.23 ;
      RECT 74.275 3.236 74.361 3.801 ;
      RECT 74.23 3.238 74.395 3.795 ;
      RECT 74.361 3.235 74.395 3.795 ;
      RECT 74.275 3.237 74.48 3.789 ;
      RECT 74.23 3.247 74.49 3.785 ;
      RECT 74.205 3.239 74.48 3.781 ;
      RECT 74.2 3.242 74.48 3.776 ;
      RECT 74.175 3.257 74.49 3.77 ;
      RECT 74.175 3.282 74.53 3.765 ;
      RECT 74.135 3.29 74.53 3.74 ;
      RECT 74.135 3.317 74.545 3.738 ;
      RECT 74.135 3.347 74.555 3.725 ;
      RECT 74.13 3.492 74.555 3.713 ;
      RECT 74.135 3.421 74.575 3.71 ;
      RECT 74.135 3.478 74.58 3.518 ;
      RECT 74.325 2.757 74.495 2.935 ;
      RECT 74.275 2.696 74.325 2.92 ;
      RECT 74.01 2.676 74.275 2.905 ;
      RECT 73.97 2.74 74.445 2.905 ;
      RECT 73.97 2.73 74.4 2.905 ;
      RECT 73.97 2.727 74.39 2.905 ;
      RECT 73.97 2.715 74.38 2.905 ;
      RECT 73.97 2.7 74.325 2.905 ;
      RECT 74.01 2.672 74.211 2.905 ;
      RECT 74.02 2.65 74.211 2.905 ;
      RECT 74.045 2.635 74.125 2.905 ;
      RECT 73.8 3.165 73.92 3.61 ;
      RECT 73.785 3.165 73.92 3.609 ;
      RECT 73.74 3.187 73.92 3.604 ;
      RECT 73.7 3.236 73.92 3.598 ;
      RECT 73.7 3.236 73.925 3.573 ;
      RECT 73.7 3.236 73.945 3.463 ;
      RECT 73.695 3.266 73.945 3.46 ;
      RECT 73.785 3.165 73.955 3.355 ;
      RECT 73.445 1.95 73.45 2.395 ;
      RECT 73.255 1.95 73.275 2.36 ;
      RECT 73.225 1.95 73.23 2.335 ;
      RECT 73.905 2.257 73.92 2.445 ;
      RECT 73.9 2.242 73.905 2.451 ;
      RECT 73.88 2.215 73.9 2.454 ;
      RECT 73.83 2.182 73.88 2.463 ;
      RECT 73.8 2.162 73.83 2.467 ;
      RECT 73.781 2.15 73.8 2.463 ;
      RECT 73.695 2.122 73.781 2.453 ;
      RECT 73.685 2.097 73.695 2.443 ;
      RECT 73.615 2.065 73.685 2.435 ;
      RECT 73.59 2.025 73.615 2.427 ;
      RECT 73.57 2.007 73.59 2.421 ;
      RECT 73.56 1.997 73.57 2.418 ;
      RECT 73.55 1.99 73.56 2.416 ;
      RECT 73.53 1.977 73.55 2.413 ;
      RECT 73.52 1.967 73.53 2.41 ;
      RECT 73.51 1.96 73.52 2.408 ;
      RECT 73.46 1.952 73.51 2.402 ;
      RECT 73.45 1.95 73.46 2.396 ;
      RECT 73.42 1.95 73.445 2.393 ;
      RECT 73.391 1.95 73.42 2.388 ;
      RECT 73.305 1.95 73.391 2.378 ;
      RECT 73.275 1.95 73.305 2.365 ;
      RECT 73.23 1.95 73.255 2.348 ;
      RECT 73.215 1.95 73.225 2.33 ;
      RECT 73.195 1.957 73.215 2.315 ;
      RECT 73.19 1.972 73.195 2.303 ;
      RECT 73.185 1.977 73.19 2.243 ;
      RECT 73.18 1.982 73.185 2.085 ;
      RECT 73.175 1.985 73.18 2.003 ;
      RECT 73.44 2.67 73.526 2.991 ;
      RECT 73.44 2.67 73.56 2.984 ;
      RECT 73.39 2.67 73.56 2.98 ;
      RECT 73.39 2.672 73.646 2.978 ;
      RECT 73.39 2.674 73.67 2.972 ;
      RECT 73.39 2.681 73.68 2.971 ;
      RECT 73.39 2.69 73.685 2.968 ;
      RECT 73.39 2.696 73.69 2.963 ;
      RECT 73.39 2.74 73.695 2.96 ;
      RECT 73.39 2.832 73.7 2.957 ;
      RECT 72.915 3.275 72.95 3.595 ;
      RECT 73.5 3.46 73.505 3.642 ;
      RECT 73.455 3.342 73.5 3.661 ;
      RECT 73.44 3.319 73.455 3.684 ;
      RECT 73.43 3.309 73.44 3.694 ;
      RECT 73.41 3.304 73.43 3.707 ;
      RECT 73.385 3.302 73.41 3.728 ;
      RECT 73.366 3.301 73.385 3.74 ;
      RECT 73.28 3.298 73.366 3.74 ;
      RECT 73.21 3.293 73.28 3.728 ;
      RECT 73.135 3.289 73.21 3.703 ;
      RECT 73.07 3.285 73.135 3.67 ;
      RECT 73 3.282 73.07 3.63 ;
      RECT 72.97 3.278 73 3.605 ;
      RECT 72.95 3.276 72.97 3.598 ;
      RECT 72.866 3.274 72.915 3.596 ;
      RECT 72.78 3.271 72.866 3.597 ;
      RECT 72.705 3.27 72.78 3.599 ;
      RECT 72.62 3.27 72.705 3.625 ;
      RECT 72.543 3.271 72.62 3.65 ;
      RECT 72.457 3.272 72.543 3.65 ;
      RECT 72.371 3.272 72.457 3.65 ;
      RECT 72.285 3.273 72.371 3.65 ;
      RECT 72.265 3.274 72.285 3.642 ;
      RECT 72.25 3.28 72.265 3.627 ;
      RECT 72.215 3.3 72.25 3.607 ;
      RECT 72.205 3.32 72.215 3.589 ;
      RECT 73.175 2.625 73.18 2.895 ;
      RECT 73.17 2.616 73.175 2.9 ;
      RECT 73.16 2.606 73.17 2.912 ;
      RECT 73.155 2.595 73.16 2.923 ;
      RECT 73.135 2.589 73.155 2.941 ;
      RECT 73.09 2.586 73.135 2.99 ;
      RECT 73.075 2.585 73.09 3.035 ;
      RECT 73.07 2.585 73.075 3.048 ;
      RECT 73.06 2.585 73.07 3.06 ;
      RECT 73.055 2.586 73.06 3.075 ;
      RECT 73.035 2.594 73.055 3.08 ;
      RECT 73.005 2.61 73.035 3.08 ;
      RECT 72.995 2.622 73 3.08 ;
      RECT 72.96 2.637 72.995 3.08 ;
      RECT 72.93 2.657 72.96 3.08 ;
      RECT 72.92 2.682 72.93 3.08 ;
      RECT 72.915 2.71 72.92 3.08 ;
      RECT 72.91 2.74 72.915 3.08 ;
      RECT 72.905 2.757 72.91 3.08 ;
      RECT 72.895 2.785 72.905 3.08 ;
      RECT 72.885 2.82 72.895 3.08 ;
      RECT 72.88 2.855 72.885 3.08 ;
      RECT 73 2.62 73.005 3.08 ;
      RECT 72.515 2.722 72.7 2.895 ;
      RECT 72.475 2.64 72.66 2.893 ;
      RECT 72.436 2.645 72.66 2.889 ;
      RECT 72.35 2.654 72.66 2.884 ;
      RECT 72.266 2.67 72.665 2.879 ;
      RECT 72.18 2.69 72.69 2.873 ;
      RECT 72.18 2.71 72.695 2.873 ;
      RECT 72.266 2.68 72.69 2.879 ;
      RECT 72.35 2.655 72.665 2.884 ;
      RECT 72.515 2.637 72.66 2.895 ;
      RECT 72.515 2.632 72.615 2.895 ;
      RECT 72.601 2.626 72.615 2.895 ;
      RECT 71.99 1.95 71.995 2.349 ;
      RECT 71.735 1.95 71.77 2.347 ;
      RECT 71.33 1.985 71.335 2.341 ;
      RECT 72.075 1.988 72.08 2.243 ;
      RECT 72.07 1.986 72.075 2.249 ;
      RECT 72.065 1.985 72.07 2.256 ;
      RECT 72.04 1.978 72.065 2.28 ;
      RECT 72.035 1.971 72.04 2.304 ;
      RECT 72.03 1.967 72.035 2.313 ;
      RECT 72.02 1.962 72.03 2.326 ;
      RECT 72.015 1.959 72.02 2.335 ;
      RECT 72.01 1.957 72.015 2.34 ;
      RECT 71.995 1.953 72.01 2.35 ;
      RECT 71.98 1.947 71.99 2.349 ;
      RECT 71.942 1.945 71.98 2.349 ;
      RECT 71.856 1.947 71.942 2.349 ;
      RECT 71.77 1.949 71.856 2.348 ;
      RECT 71.699 1.95 71.735 2.347 ;
      RECT 71.613 1.952 71.699 2.347 ;
      RECT 71.527 1.954 71.613 2.346 ;
      RECT 71.441 1.956 71.527 2.346 ;
      RECT 71.355 1.959 71.441 2.345 ;
      RECT 71.345 1.965 71.355 2.344 ;
      RECT 71.335 1.977 71.345 2.342 ;
      RECT 71.275 2.012 71.33 2.338 ;
      RECT 71.27 2.042 71.275 2.1 ;
      RECT 72.015 3.122 72.03 3.315 ;
      RECT 72.01 3.09 72.015 3.315 ;
      RECT 72 3.065 72.01 3.315 ;
      RECT 71.995 3.037 72 3.315 ;
      RECT 71.965 2.96 71.995 3.315 ;
      RECT 71.94 2.842 71.965 3.315 ;
      RECT 71.935 2.78 71.94 3.315 ;
      RECT 71.925 2.767 71.935 3.315 ;
      RECT 71.905 2.757 71.925 3.315 ;
      RECT 71.89 2.74 71.905 3.315 ;
      RECT 71.86 2.728 71.89 3.315 ;
      RECT 71.855 2.727 71.86 3.26 ;
      RECT 71.85 2.727 71.855 3.218 ;
      RECT 71.835 2.726 71.85 3.17 ;
      RECT 71.82 2.726 71.835 3.108 ;
      RECT 71.8 2.726 71.82 3.068 ;
      RECT 71.795 2.726 71.8 3.053 ;
      RECT 71.77 2.725 71.795 3.048 ;
      RECT 71.7 2.724 71.77 3.035 ;
      RECT 71.685 2.723 71.7 3.02 ;
      RECT 71.655 2.722 71.685 3.003 ;
      RECT 71.65 2.722 71.655 2.988 ;
      RECT 71.6 2.721 71.65 2.968 ;
      RECT 71.535 2.72 71.6 2.923 ;
      RECT 71.53 2.72 71.535 2.895 ;
      RECT 71.615 3.257 71.62 3.514 ;
      RECT 71.595 3.176 71.615 3.531 ;
      RECT 71.575 3.17 71.595 3.56 ;
      RECT 71.515 3.157 71.575 3.58 ;
      RECT 71.47 3.141 71.515 3.581 ;
      RECT 71.386 3.129 71.47 3.569 ;
      RECT 71.3 3.116 71.386 3.553 ;
      RECT 71.29 3.109 71.3 3.545 ;
      RECT 71.245 3.106 71.29 3.485 ;
      RECT 71.225 3.102 71.245 3.4 ;
      RECT 71.21 3.1 71.225 3.353 ;
      RECT 71.18 3.097 71.21 3.323 ;
      RECT 71.145 3.093 71.18 3.3 ;
      RECT 71.102 3.088 71.145 3.288 ;
      RECT 71.016 3.079 71.102 3.297 ;
      RECT 70.93 3.068 71.016 3.309 ;
      RECT 70.865 3.059 70.93 3.318 ;
      RECT 70.845 3.05 70.865 3.323 ;
      RECT 70.84 3.043 70.845 3.325 ;
      RECT 70.8 3.028 70.84 3.322 ;
      RECT 70.78 3.007 70.8 3.317 ;
      RECT 70.765 2.995 70.78 3.31 ;
      RECT 70.76 2.987 70.765 3.303 ;
      RECT 70.745 2.967 70.76 3.296 ;
      RECT 70.74 2.83 70.745 3.29 ;
      RECT 70.66 2.719 70.74 3.262 ;
      RECT 70.651 2.712 70.66 3.228 ;
      RECT 70.565 2.706 70.651 3.153 ;
      RECT 70.54 2.697 70.565 3.065 ;
      RECT 70.51 2.692 70.54 3.04 ;
      RECT 70.445 2.701 70.51 3.025 ;
      RECT 70.425 2.717 70.445 3 ;
      RECT 70.415 2.723 70.425 2.948 ;
      RECT 70.395 2.745 70.415 2.83 ;
      RECT 71.05 2.71 71.22 2.895 ;
      RECT 71.05 2.71 71.255 2.893 ;
      RECT 71.1 2.62 71.27 2.884 ;
      RECT 71.05 2.777 71.275 2.877 ;
      RECT 71.065 2.655 71.27 2.884 ;
      RECT 70.265 3.388 70.33 3.831 ;
      RECT 70.205 3.413 70.33 3.829 ;
      RECT 70.205 3.413 70.385 3.823 ;
      RECT 70.19 3.438 70.385 3.822 ;
      RECT 70.33 3.375 70.405 3.819 ;
      RECT 70.265 3.4 70.485 3.813 ;
      RECT 70.19 3.439 70.53 3.807 ;
      RECT 70.175 3.466 70.53 3.798 ;
      RECT 70.19 3.459 70.55 3.79 ;
      RECT 70.175 3.468 70.555 3.773 ;
      RECT 70.17 3.485 70.555 3.6 ;
      RECT 70.175 2.207 70.21 2.445 ;
      RECT 70.175 2.207 70.24 2.444 ;
      RECT 70.175 2.207 70.355 2.44 ;
      RECT 70.175 2.207 70.41 2.418 ;
      RECT 70.185 2.15 70.465 2.318 ;
      RECT 70.29 1.99 70.32 2.441 ;
      RECT 70.32 1.985 70.5 2.198 ;
      RECT 70.19 2.126 70.5 2.198 ;
      RECT 70.24 2.022 70.29 2.442 ;
      RECT 70.21 2.078 70.5 2.198 ;
      RECT 68.715 1.74 68.885 2.935 ;
      RECT 68.715 1.74 69.18 1.91 ;
      RECT 68.715 6.97 69.18 7.14 ;
      RECT 68.715 5.945 68.885 7.14 ;
      RECT 67.725 1.74 67.895 2.935 ;
      RECT 67.725 1.74 68.19 1.91 ;
      RECT 67.725 6.97 68.19 7.14 ;
      RECT 67.725 5.945 67.895 7.14 ;
      RECT 65.87 2.635 66.04 3.865 ;
      RECT 65.925 0.855 66.095 2.805 ;
      RECT 65.87 0.575 66.04 1.025 ;
      RECT 65.87 7.855 66.04 8.305 ;
      RECT 65.925 6.075 66.095 8.025 ;
      RECT 65.87 5.015 66.04 6.245 ;
      RECT 65.35 0.575 65.52 3.865 ;
      RECT 65.35 2.075 65.755 2.405 ;
      RECT 65.35 1.235 65.755 1.565 ;
      RECT 65.35 5.015 65.52 8.305 ;
      RECT 65.35 7.315 65.755 7.645 ;
      RECT 65.35 6.475 65.755 6.805 ;
      RECT 63.45 3.392 63.465 3.443 ;
      RECT 63.445 3.372 63.45 3.49 ;
      RECT 63.43 3.362 63.445 3.558 ;
      RECT 63.405 3.342 63.43 3.613 ;
      RECT 63.365 3.327 63.405 3.633 ;
      RECT 63.32 3.321 63.365 3.661 ;
      RECT 63.25 3.311 63.32 3.678 ;
      RECT 63.23 3.303 63.25 3.678 ;
      RECT 63.17 3.297 63.23 3.67 ;
      RECT 63.111 3.288 63.17 3.658 ;
      RECT 63.025 3.277 63.111 3.641 ;
      RECT 63.003 3.268 63.025 3.629 ;
      RECT 62.917 3.261 63.003 3.616 ;
      RECT 62.831 3.248 62.917 3.597 ;
      RECT 62.745 3.236 62.831 3.577 ;
      RECT 62.715 3.225 62.745 3.564 ;
      RECT 62.665 3.211 62.715 3.556 ;
      RECT 62.645 3.2 62.665 3.548 ;
      RECT 62.596 3.189 62.645 3.54 ;
      RECT 62.51 3.168 62.596 3.525 ;
      RECT 62.465 3.155 62.51 3.51 ;
      RECT 62.42 3.155 62.465 3.49 ;
      RECT 62.365 3.155 62.42 3.425 ;
      RECT 62.34 3.155 62.365 3.348 ;
      RECT 62.865 2.892 63.035 3.075 ;
      RECT 62.865 2.892 63.05 3.033 ;
      RECT 62.865 2.892 63.055 2.975 ;
      RECT 62.925 2.66 63.06 2.951 ;
      RECT 62.925 2.664 63.065 2.934 ;
      RECT 62.87 2.827 63.065 2.934 ;
      RECT 62.895 2.672 63.035 3.075 ;
      RECT 62.895 2.676 63.075 2.875 ;
      RECT 62.88 2.762 63.075 2.875 ;
      RECT 62.89 2.692 63.035 3.075 ;
      RECT 62.89 2.695 63.085 2.788 ;
      RECT 62.885 2.712 63.085 2.788 ;
      RECT 62.655 1.932 62.825 2.415 ;
      RECT 62.65 1.927 62.8 2.405 ;
      RECT 62.65 1.934 62.83 2.399 ;
      RECT 62.64 1.928 62.8 2.378 ;
      RECT 62.64 1.944 62.845 2.337 ;
      RECT 62.61 1.929 62.8 2.3 ;
      RECT 62.61 1.959 62.855 2.24 ;
      RECT 62.605 1.931 62.8 2.238 ;
      RECT 62.585 1.94 62.83 2.195 ;
      RECT 62.56 1.956 62.845 2.107 ;
      RECT 62.56 1.975 62.87 2.098 ;
      RECT 62.555 2.012 62.87 2.05 ;
      RECT 62.56 1.992 62.875 2.018 ;
      RECT 62.655 1.926 62.765 2.415 ;
      RECT 62.741 1.925 62.765 2.415 ;
      RECT 61.975 2.71 61.98 2.921 ;
      RECT 62.575 2.71 62.58 2.895 ;
      RECT 62.64 2.75 62.645 2.863 ;
      RECT 62.635 2.742 62.64 2.869 ;
      RECT 62.63 2.732 62.635 2.877 ;
      RECT 62.625 2.722 62.63 2.886 ;
      RECT 62.62 2.712 62.625 2.89 ;
      RECT 62.58 2.71 62.62 2.893 ;
      RECT 62.552 2.709 62.575 2.897 ;
      RECT 62.466 2.706 62.552 2.904 ;
      RECT 62.38 2.702 62.466 2.915 ;
      RECT 62.36 2.7 62.38 2.921 ;
      RECT 62.342 2.699 62.36 2.924 ;
      RECT 62.256 2.697 62.342 2.931 ;
      RECT 62.17 2.692 62.256 2.944 ;
      RECT 62.151 2.689 62.17 2.949 ;
      RECT 62.065 2.687 62.151 2.94 ;
      RECT 62.055 2.687 62.065 2.933 ;
      RECT 61.98 2.7 62.055 2.927 ;
      RECT 61.965 2.711 61.975 2.921 ;
      RECT 61.955 2.713 61.965 2.92 ;
      RECT 61.945 2.717 61.955 2.916 ;
      RECT 61.94 2.72 61.945 2.91 ;
      RECT 61.93 2.722 61.94 2.904 ;
      RECT 61.925 2.725 61.93 2.898 ;
      RECT 61.905 3.311 61.91 3.515 ;
      RECT 61.89 3.298 61.905 3.608 ;
      RECT 61.875 3.279 61.89 3.885 ;
      RECT 61.84 3.245 61.875 3.885 ;
      RECT 61.836 3.215 61.84 3.885 ;
      RECT 61.75 3.097 61.836 3.885 ;
      RECT 61.74 2.972 61.75 3.885 ;
      RECT 61.725 2.94 61.74 3.885 ;
      RECT 61.72 2.915 61.725 3.885 ;
      RECT 61.715 2.905 61.72 3.841 ;
      RECT 61.7 2.877 61.715 3.746 ;
      RECT 61.685 2.843 61.7 3.645 ;
      RECT 61.68 2.821 61.685 3.598 ;
      RECT 61.675 2.81 61.68 3.568 ;
      RECT 61.67 2.8 61.675 3.534 ;
      RECT 61.66 2.787 61.67 3.502 ;
      RECT 61.635 2.763 61.66 3.428 ;
      RECT 61.63 2.743 61.635 3.353 ;
      RECT 61.625 2.737 61.63 3.328 ;
      RECT 61.62 2.732 61.625 3.293 ;
      RECT 61.615 2.727 61.62 3.268 ;
      RECT 61.61 2.725 61.615 3.248 ;
      RECT 61.605 2.725 61.61 3.233 ;
      RECT 61.6 2.725 61.605 3.193 ;
      RECT 61.59 2.725 61.6 3.165 ;
      RECT 61.58 2.725 61.59 3.11 ;
      RECT 61.565 2.725 61.58 3.048 ;
      RECT 61.56 2.724 61.565 2.993 ;
      RECT 61.545 2.723 61.56 2.973 ;
      RECT 61.485 2.721 61.545 2.947 ;
      RECT 61.45 2.722 61.485 2.927 ;
      RECT 61.445 2.724 61.45 2.917 ;
      RECT 61.435 2.743 61.445 2.907 ;
      RECT 61.43 2.77 61.435 2.838 ;
      RECT 61.545 2.195 61.715 2.44 ;
      RECT 61.58 1.966 61.715 2.44 ;
      RECT 61.58 1.968 61.725 2.435 ;
      RECT 61.58 1.97 61.75 2.423 ;
      RECT 61.58 1.973 61.775 2.405 ;
      RECT 61.58 1.978 61.825 2.378 ;
      RECT 61.58 1.983 61.845 2.343 ;
      RECT 61.56 1.985 61.855 2.318 ;
      RECT 61.55 2.08 61.855 2.318 ;
      RECT 61.58 1.965 61.69 2.44 ;
      RECT 61.59 1.962 61.685 2.44 ;
      RECT 61.11 3.227 61.3 3.585 ;
      RECT 61.11 3.239 61.335 3.584 ;
      RECT 61.11 3.267 61.355 3.582 ;
      RECT 61.11 3.292 61.36 3.581 ;
      RECT 61.11 3.35 61.375 3.58 ;
      RECT 61.095 3.223 61.255 3.565 ;
      RECT 61.075 3.232 61.3 3.518 ;
      RECT 61.05 3.243 61.335 3.455 ;
      RECT 61.05 3.327 61.37 3.455 ;
      RECT 61.05 3.302 61.365 3.455 ;
      RECT 61.11 3.218 61.255 3.585 ;
      RECT 61.196 3.217 61.255 3.585 ;
      RECT 61.196 3.216 61.24 3.585 ;
      RECT 61.11 7.855 61.28 8.305 ;
      RECT 61.165 6.075 61.335 8.025 ;
      RECT 61.11 5.015 61.28 6.245 ;
      RECT 60.59 5.015 60.76 8.305 ;
      RECT 60.59 7.315 60.995 7.645 ;
      RECT 60.59 6.475 60.995 6.805 ;
      RECT 60.895 2.732 60.9 3.11 ;
      RECT 60.89 2.7 60.895 3.11 ;
      RECT 60.885 2.672 60.89 3.11 ;
      RECT 60.88 2.652 60.885 3.11 ;
      RECT 60.825 2.635 60.88 3.11 ;
      RECT 60.785 2.62 60.825 3.11 ;
      RECT 60.73 2.607 60.785 3.11 ;
      RECT 60.695 2.598 60.73 3.11 ;
      RECT 60.691 2.596 60.695 3.109 ;
      RECT 60.605 2.592 60.691 3.092 ;
      RECT 60.52 2.584 60.605 3.055 ;
      RECT 60.51 2.58 60.52 3.028 ;
      RECT 60.5 2.58 60.51 3.01 ;
      RECT 60.49 2.582 60.5 2.993 ;
      RECT 60.485 2.587 60.49 2.979 ;
      RECT 60.48 2.591 60.485 2.966 ;
      RECT 60.47 2.596 60.48 2.95 ;
      RECT 60.455 2.61 60.47 2.925 ;
      RECT 60.45 2.616 60.455 2.905 ;
      RECT 60.445 2.618 60.45 2.898 ;
      RECT 60.44 2.622 60.445 2.773 ;
      RECT 60.62 3.422 60.865 3.885 ;
      RECT 60.54 3.395 60.86 3.881 ;
      RECT 60.47 3.43 60.865 3.874 ;
      RECT 60.26 3.685 60.865 3.87 ;
      RECT 60.44 3.453 60.865 3.87 ;
      RECT 60.28 3.645 60.865 3.87 ;
      RECT 60.43 3.465 60.865 3.87 ;
      RECT 60.315 3.582 60.865 3.87 ;
      RECT 60.37 3.507 60.865 3.87 ;
      RECT 60.62 3.372 60.86 3.885 ;
      RECT 60.65 3.365 60.86 3.885 ;
      RECT 60.64 3.367 60.86 3.885 ;
      RECT 60.65 3.362 60.78 3.885 ;
      RECT 60.205 1.925 60.291 2.364 ;
      RECT 60.2 1.925 60.291 2.362 ;
      RECT 60.2 1.925 60.36 2.361 ;
      RECT 60.2 1.925 60.39 2.358 ;
      RECT 60.185 1.932 60.39 2.349 ;
      RECT 60.185 1.932 60.395 2.345 ;
      RECT 60.18 1.942 60.395 2.338 ;
      RECT 60.175 1.947 60.395 2.313 ;
      RECT 60.175 1.947 60.41 2.295 ;
      RECT 60.2 1.925 60.43 2.21 ;
      RECT 60.17 1.952 60.43 2.208 ;
      RECT 60.18 1.945 60.435 2.146 ;
      RECT 60.17 2.067 60.44 2.129 ;
      RECT 60.155 1.962 60.435 2.08 ;
      RECT 60.15 1.972 60.435 1.98 ;
      RECT 60.23 2.743 60.235 2.82 ;
      RECT 60.22 2.737 60.23 3.01 ;
      RECT 60.21 2.729 60.22 3.031 ;
      RECT 60.2 2.72 60.21 3.053 ;
      RECT 60.195 2.715 60.2 3.07 ;
      RECT 60.155 2.715 60.195 3.11 ;
      RECT 60.135 2.715 60.155 3.165 ;
      RECT 60.13 2.715 60.135 3.193 ;
      RECT 60.12 2.715 60.13 3.208 ;
      RECT 60.085 2.715 60.12 3.25 ;
      RECT 60.08 2.715 60.085 3.293 ;
      RECT 60.07 2.715 60.08 3.308 ;
      RECT 60.055 2.715 60.07 3.328 ;
      RECT 60.04 2.715 60.055 3.355 ;
      RECT 60.035 2.716 60.04 3.373 ;
      RECT 60.015 2.717 60.035 3.38 ;
      RECT 59.96 2.718 60.015 3.4 ;
      RECT 59.95 2.719 59.96 3.414 ;
      RECT 59.945 2.722 59.95 3.413 ;
      RECT 59.905 2.795 59.945 3.411 ;
      RECT 59.89 2.875 59.905 3.409 ;
      RECT 59.865 2.93 59.89 3.407 ;
      RECT 59.85 2.995 59.865 3.406 ;
      RECT 59.805 3.027 59.85 3.403 ;
      RECT 59.72 3.05 59.805 3.398 ;
      RECT 59.695 3.07 59.72 3.393 ;
      RECT 59.625 3.075 59.695 3.389 ;
      RECT 59.605 3.077 59.625 3.386 ;
      RECT 59.52 3.088 59.605 3.38 ;
      RECT 59.515 3.099 59.52 3.375 ;
      RECT 59.505 3.101 59.515 3.375 ;
      RECT 59.47 3.105 59.505 3.373 ;
      RECT 59.42 3.115 59.47 3.36 ;
      RECT 59.4 3.123 59.42 3.345 ;
      RECT 59.32 3.135 59.4 3.328 ;
      RECT 59.485 2.685 59.655 2.895 ;
      RECT 59.601 2.681 59.655 2.895 ;
      RECT 59.406 2.685 59.655 2.886 ;
      RECT 59.406 2.685 59.66 2.875 ;
      RECT 59.32 2.685 59.66 2.866 ;
      RECT 59.32 2.693 59.67 2.81 ;
      RECT 59.32 2.705 59.675 2.723 ;
      RECT 59.32 2.712 59.68 2.715 ;
      RECT 59.515 2.683 59.655 2.895 ;
      RECT 59.27 3.628 59.515 3.96 ;
      RECT 59.265 3.62 59.27 3.957 ;
      RECT 59.235 3.64 59.515 3.938 ;
      RECT 59.215 3.672 59.515 3.911 ;
      RECT 59.265 3.625 59.442 3.957 ;
      RECT 59.265 3.622 59.356 3.957 ;
      RECT 59.205 1.97 59.375 2.39 ;
      RECT 59.2 1.97 59.375 2.388 ;
      RECT 59.2 1.97 59.4 2.378 ;
      RECT 59.2 1.97 59.42 2.353 ;
      RECT 59.195 1.97 59.42 2.348 ;
      RECT 59.195 1.97 59.43 2.338 ;
      RECT 59.195 1.97 59.435 2.333 ;
      RECT 59.195 1.975 59.44 2.328 ;
      RECT 59.195 2.007 59.455 2.318 ;
      RECT 59.195 2.077 59.48 2.301 ;
      RECT 59.175 2.077 59.48 2.293 ;
      RECT 59.175 2.137 59.49 2.27 ;
      RECT 59.175 2.177 59.5 2.215 ;
      RECT 59.16 1.97 59.435 2.195 ;
      RECT 59.15 1.985 59.44 2.093 ;
      RECT 58.74 3.375 58.91 3.9 ;
      RECT 58.735 3.375 58.91 3.893 ;
      RECT 58.725 3.375 58.915 3.858 ;
      RECT 58.72 3.385 58.915 3.83 ;
      RECT 58.715 3.405 58.915 3.813 ;
      RECT 58.725 3.38 58.92 3.803 ;
      RECT 58.71 3.425 58.92 3.795 ;
      RECT 58.705 3.445 58.92 3.78 ;
      RECT 58.7 3.475 58.92 3.77 ;
      RECT 58.69 3.52 58.92 3.745 ;
      RECT 58.72 3.39 58.925 3.728 ;
      RECT 58.685 3.572 58.925 3.723 ;
      RECT 58.72 3.4 58.93 3.693 ;
      RECT 58.68 3.605 58.93 3.69 ;
      RECT 58.675 3.63 58.93 3.67 ;
      RECT 58.715 3.417 58.94 3.61 ;
      RECT 58.71 3.439 58.95 3.503 ;
      RECT 58.66 2.686 58.675 2.955 ;
      RECT 58.615 2.67 58.66 3 ;
      RECT 58.61 2.658 58.615 3.05 ;
      RECT 58.6 2.654 58.61 3.083 ;
      RECT 58.595 2.651 58.6 3.111 ;
      RECT 58.58 2.653 58.595 3.153 ;
      RECT 58.575 2.657 58.58 3.193 ;
      RECT 58.555 2.662 58.575 3.245 ;
      RECT 58.551 2.667 58.555 3.302 ;
      RECT 58.465 2.686 58.551 3.339 ;
      RECT 58.455 2.707 58.465 3.375 ;
      RECT 58.45 2.715 58.455 3.376 ;
      RECT 58.445 2.757 58.45 3.377 ;
      RECT 58.43 2.845 58.445 3.378 ;
      RECT 58.42 2.995 58.43 3.38 ;
      RECT 58.415 3.04 58.42 3.382 ;
      RECT 58.38 3.082 58.415 3.385 ;
      RECT 58.375 3.1 58.38 3.388 ;
      RECT 58.298 3.106 58.375 3.394 ;
      RECT 58.212 3.12 58.298 3.407 ;
      RECT 58.126 3.134 58.212 3.421 ;
      RECT 58.04 3.148 58.126 3.434 ;
      RECT 57.98 3.16 58.04 3.446 ;
      RECT 57.955 3.167 57.98 3.453 ;
      RECT 57.941 3.17 57.955 3.458 ;
      RECT 57.855 3.178 57.941 3.474 ;
      RECT 57.85 3.185 57.855 3.489 ;
      RECT 57.826 3.185 57.85 3.496 ;
      RECT 57.74 3.188 57.826 3.524 ;
      RECT 57.655 3.192 57.74 3.568 ;
      RECT 57.59 3.196 57.655 3.605 ;
      RECT 57.565 3.199 57.59 3.621 ;
      RECT 57.49 3.212 57.565 3.625 ;
      RECT 57.465 3.23 57.49 3.629 ;
      RECT 57.455 3.237 57.465 3.631 ;
      RECT 57.44 3.24 57.455 3.632 ;
      RECT 57.38 3.252 57.44 3.636 ;
      RECT 57.37 3.266 57.38 3.64 ;
      RECT 57.315 3.276 57.37 3.628 ;
      RECT 57.29 3.297 57.315 3.611 ;
      RECT 57.27 3.317 57.29 3.602 ;
      RECT 57.265 3.33 57.27 3.597 ;
      RECT 57.25 3.342 57.265 3.593 ;
      RECT 58.485 1.997 58.49 2.02 ;
      RECT 58.48 1.988 58.485 2.06 ;
      RECT 58.475 1.986 58.48 2.103 ;
      RECT 58.47 1.977 58.475 2.138 ;
      RECT 58.465 1.967 58.47 2.21 ;
      RECT 58.46 1.957 58.465 2.275 ;
      RECT 58.455 1.954 58.46 2.315 ;
      RECT 58.43 1.948 58.455 2.405 ;
      RECT 58.395 1.936 58.43 2.43 ;
      RECT 58.385 1.927 58.395 2.43 ;
      RECT 58.25 1.925 58.26 2.413 ;
      RECT 58.24 1.925 58.25 2.38 ;
      RECT 58.235 1.925 58.24 2.355 ;
      RECT 58.23 1.925 58.235 2.343 ;
      RECT 58.225 1.925 58.23 2.325 ;
      RECT 58.215 1.925 58.225 2.29 ;
      RECT 58.21 1.927 58.215 2.268 ;
      RECT 58.205 1.933 58.21 2.253 ;
      RECT 58.2 1.939 58.205 2.238 ;
      RECT 58.185 1.951 58.2 2.211 ;
      RECT 58.18 1.962 58.185 2.179 ;
      RECT 58.175 1.972 58.18 2.163 ;
      RECT 58.165 1.98 58.175 2.132 ;
      RECT 58.16 1.99 58.165 2.106 ;
      RECT 58.155 2.047 58.16 2.089 ;
      RECT 58.26 1.925 58.385 2.43 ;
      RECT 57.975 2.612 58.235 2.91 ;
      RECT 57.97 2.619 58.235 2.908 ;
      RECT 57.975 2.614 58.25 2.903 ;
      RECT 57.965 2.627 58.25 2.9 ;
      RECT 57.965 2.632 58.255 2.893 ;
      RECT 57.96 2.64 58.255 2.89 ;
      RECT 57.96 2.657 58.26 2.688 ;
      RECT 57.975 2.609 58.206 2.91 ;
      RECT 58.03 2.608 58.206 2.91 ;
      RECT 58.03 2.605 58.12 2.91 ;
      RECT 58.03 2.602 58.116 2.91 ;
      RECT 57.72 2.875 57.725 2.888 ;
      RECT 57.715 2.842 57.72 2.893 ;
      RECT 57.71 2.797 57.715 2.9 ;
      RECT 57.705 2.752 57.71 2.908 ;
      RECT 57.7 2.72 57.705 2.916 ;
      RECT 57.695 2.68 57.7 2.917 ;
      RECT 57.68 2.66 57.695 2.919 ;
      RECT 57.605 2.642 57.68 2.931 ;
      RECT 57.595 2.635 57.605 2.942 ;
      RECT 57.59 2.635 57.595 2.944 ;
      RECT 57.56 2.641 57.59 2.948 ;
      RECT 57.52 2.654 57.56 2.948 ;
      RECT 57.495 2.665 57.52 2.934 ;
      RECT 57.48 2.671 57.495 2.917 ;
      RECT 57.47 2.673 57.48 2.908 ;
      RECT 57.465 2.674 57.47 2.903 ;
      RECT 57.46 2.675 57.465 2.898 ;
      RECT 57.455 2.676 57.46 2.895 ;
      RECT 57.43 2.681 57.455 2.885 ;
      RECT 57.42 2.697 57.43 2.872 ;
      RECT 57.415 2.717 57.42 2.867 ;
      RECT 57.425 2.11 57.43 2.306 ;
      RECT 57.41 2.074 57.425 2.308 ;
      RECT 57.4 2.056 57.41 2.313 ;
      RECT 57.39 2.042 57.4 2.317 ;
      RECT 57.345 2.026 57.39 2.327 ;
      RECT 57.34 2.016 57.345 2.336 ;
      RECT 57.295 2.005 57.34 2.342 ;
      RECT 57.29 1.993 57.295 2.349 ;
      RECT 57.275 1.988 57.29 2.353 ;
      RECT 57.26 1.98 57.275 2.358 ;
      RECT 57.25 1.973 57.26 2.363 ;
      RECT 57.24 1.97 57.25 2.368 ;
      RECT 57.23 1.97 57.24 2.369 ;
      RECT 57.225 1.967 57.23 2.368 ;
      RECT 57.19 1.962 57.215 2.367 ;
      RECT 57.166 1.958 57.19 2.366 ;
      RECT 57.08 1.949 57.166 2.363 ;
      RECT 57.065 1.941 57.08 2.36 ;
      RECT 57.043 1.94 57.065 2.359 ;
      RECT 56.957 1.94 57.043 2.357 ;
      RECT 56.871 1.94 56.957 2.355 ;
      RECT 56.785 1.94 56.871 2.352 ;
      RECT 56.775 1.94 56.785 2.343 ;
      RECT 56.745 1.94 56.775 2.303 ;
      RECT 56.735 1.95 56.745 2.258 ;
      RECT 56.73 1.99 56.735 2.243 ;
      RECT 56.725 2.005 56.73 2.23 ;
      RECT 56.695 2.085 56.725 2.192 ;
      RECT 57.215 1.965 57.225 2.368 ;
      RECT 57.04 2.73 57.055 3.335 ;
      RECT 57.045 2.725 57.055 3.335 ;
      RECT 57.21 2.725 57.215 2.908 ;
      RECT 57.2 2.725 57.21 2.938 ;
      RECT 57.185 2.725 57.2 2.998 ;
      RECT 57.18 2.725 57.185 3.043 ;
      RECT 57.175 2.725 57.18 3.073 ;
      RECT 57.17 2.725 57.175 3.093 ;
      RECT 57.16 2.725 57.17 3.128 ;
      RECT 57.145 2.725 57.16 3.16 ;
      RECT 57.1 2.725 57.145 3.188 ;
      RECT 57.095 2.725 57.1 3.218 ;
      RECT 57.09 2.725 57.095 3.23 ;
      RECT 57.085 2.725 57.09 3.238 ;
      RECT 57.075 2.725 57.085 3.253 ;
      RECT 57.07 2.725 57.075 3.275 ;
      RECT 57.06 2.725 57.07 3.298 ;
      RECT 57.055 2.725 57.06 3.318 ;
      RECT 57.02 2.74 57.04 3.335 ;
      RECT 56.995 2.757 57.02 3.335 ;
      RECT 56.99 2.767 56.995 3.335 ;
      RECT 56.96 2.782 56.99 3.335 ;
      RECT 56.885 2.824 56.96 3.335 ;
      RECT 56.88 2.855 56.885 3.318 ;
      RECT 56.875 2.859 56.88 3.3 ;
      RECT 56.87 2.863 56.875 3.263 ;
      RECT 56.865 3.047 56.87 3.23 ;
      RECT 56.35 3.236 56.436 3.801 ;
      RECT 56.305 3.238 56.47 3.795 ;
      RECT 56.436 3.235 56.47 3.795 ;
      RECT 56.35 3.237 56.555 3.789 ;
      RECT 56.305 3.247 56.565 3.785 ;
      RECT 56.28 3.239 56.555 3.781 ;
      RECT 56.275 3.242 56.555 3.776 ;
      RECT 56.25 3.257 56.565 3.77 ;
      RECT 56.25 3.282 56.605 3.765 ;
      RECT 56.21 3.29 56.605 3.74 ;
      RECT 56.21 3.317 56.62 3.738 ;
      RECT 56.21 3.347 56.63 3.725 ;
      RECT 56.205 3.492 56.63 3.713 ;
      RECT 56.21 3.421 56.65 3.71 ;
      RECT 56.21 3.478 56.655 3.518 ;
      RECT 56.4 2.757 56.57 2.935 ;
      RECT 56.35 2.696 56.4 2.92 ;
      RECT 56.085 2.676 56.35 2.905 ;
      RECT 56.045 2.74 56.52 2.905 ;
      RECT 56.045 2.73 56.475 2.905 ;
      RECT 56.045 2.727 56.465 2.905 ;
      RECT 56.045 2.715 56.455 2.905 ;
      RECT 56.045 2.7 56.4 2.905 ;
      RECT 56.085 2.672 56.286 2.905 ;
      RECT 56.095 2.65 56.286 2.905 ;
      RECT 56.12 2.635 56.2 2.905 ;
      RECT 55.875 3.165 55.995 3.61 ;
      RECT 55.86 3.165 55.995 3.609 ;
      RECT 55.815 3.187 55.995 3.604 ;
      RECT 55.775 3.236 55.995 3.598 ;
      RECT 55.775 3.236 56 3.573 ;
      RECT 55.775 3.236 56.02 3.463 ;
      RECT 55.77 3.266 56.02 3.46 ;
      RECT 55.86 3.165 56.03 3.355 ;
      RECT 55.52 1.95 55.525 2.395 ;
      RECT 55.33 1.95 55.35 2.36 ;
      RECT 55.3 1.95 55.305 2.335 ;
      RECT 55.98 2.257 55.995 2.445 ;
      RECT 55.975 2.242 55.98 2.451 ;
      RECT 55.955 2.215 55.975 2.454 ;
      RECT 55.905 2.182 55.955 2.463 ;
      RECT 55.875 2.162 55.905 2.467 ;
      RECT 55.856 2.15 55.875 2.463 ;
      RECT 55.77 2.122 55.856 2.453 ;
      RECT 55.76 2.097 55.77 2.443 ;
      RECT 55.69 2.065 55.76 2.435 ;
      RECT 55.665 2.025 55.69 2.427 ;
      RECT 55.645 2.007 55.665 2.421 ;
      RECT 55.635 1.997 55.645 2.418 ;
      RECT 55.625 1.99 55.635 2.416 ;
      RECT 55.605 1.977 55.625 2.413 ;
      RECT 55.595 1.967 55.605 2.41 ;
      RECT 55.585 1.96 55.595 2.408 ;
      RECT 55.535 1.952 55.585 2.402 ;
      RECT 55.525 1.95 55.535 2.396 ;
      RECT 55.495 1.95 55.52 2.393 ;
      RECT 55.466 1.95 55.495 2.388 ;
      RECT 55.38 1.95 55.466 2.378 ;
      RECT 55.35 1.95 55.38 2.365 ;
      RECT 55.305 1.95 55.33 2.348 ;
      RECT 55.29 1.95 55.3 2.33 ;
      RECT 55.27 1.957 55.29 2.315 ;
      RECT 55.265 1.972 55.27 2.303 ;
      RECT 55.26 1.977 55.265 2.243 ;
      RECT 55.255 1.982 55.26 2.085 ;
      RECT 55.25 1.985 55.255 2.003 ;
      RECT 55.515 2.67 55.601 2.991 ;
      RECT 55.515 2.67 55.635 2.984 ;
      RECT 55.465 2.67 55.635 2.98 ;
      RECT 55.465 2.672 55.721 2.978 ;
      RECT 55.465 2.674 55.745 2.972 ;
      RECT 55.465 2.681 55.755 2.971 ;
      RECT 55.465 2.69 55.76 2.968 ;
      RECT 55.465 2.696 55.765 2.963 ;
      RECT 55.465 2.74 55.77 2.96 ;
      RECT 55.465 2.832 55.775 2.957 ;
      RECT 54.99 3.275 55.025 3.595 ;
      RECT 55.575 3.46 55.58 3.642 ;
      RECT 55.53 3.342 55.575 3.661 ;
      RECT 55.515 3.319 55.53 3.684 ;
      RECT 55.505 3.309 55.515 3.694 ;
      RECT 55.485 3.304 55.505 3.707 ;
      RECT 55.46 3.302 55.485 3.728 ;
      RECT 55.441 3.301 55.46 3.74 ;
      RECT 55.355 3.298 55.441 3.74 ;
      RECT 55.285 3.293 55.355 3.728 ;
      RECT 55.21 3.289 55.285 3.703 ;
      RECT 55.145 3.285 55.21 3.67 ;
      RECT 55.075 3.282 55.145 3.63 ;
      RECT 55.045 3.278 55.075 3.605 ;
      RECT 55.025 3.276 55.045 3.598 ;
      RECT 54.941 3.274 54.99 3.596 ;
      RECT 54.855 3.271 54.941 3.597 ;
      RECT 54.78 3.27 54.855 3.599 ;
      RECT 54.695 3.27 54.78 3.625 ;
      RECT 54.618 3.271 54.695 3.65 ;
      RECT 54.532 3.272 54.618 3.65 ;
      RECT 54.446 3.272 54.532 3.65 ;
      RECT 54.36 3.273 54.446 3.65 ;
      RECT 54.34 3.274 54.36 3.642 ;
      RECT 54.325 3.28 54.34 3.627 ;
      RECT 54.29 3.3 54.325 3.607 ;
      RECT 54.28 3.32 54.29 3.589 ;
      RECT 55.25 2.625 55.255 2.895 ;
      RECT 55.245 2.616 55.25 2.9 ;
      RECT 55.235 2.606 55.245 2.912 ;
      RECT 55.23 2.595 55.235 2.923 ;
      RECT 55.21 2.589 55.23 2.941 ;
      RECT 55.165 2.586 55.21 2.99 ;
      RECT 55.15 2.585 55.165 3.035 ;
      RECT 55.145 2.585 55.15 3.048 ;
      RECT 55.135 2.585 55.145 3.06 ;
      RECT 55.13 2.586 55.135 3.075 ;
      RECT 55.11 2.594 55.13 3.08 ;
      RECT 55.08 2.61 55.11 3.08 ;
      RECT 55.07 2.622 55.075 3.08 ;
      RECT 55.035 2.637 55.07 3.08 ;
      RECT 55.005 2.657 55.035 3.08 ;
      RECT 54.995 2.682 55.005 3.08 ;
      RECT 54.99 2.71 54.995 3.08 ;
      RECT 54.985 2.74 54.99 3.08 ;
      RECT 54.98 2.757 54.985 3.08 ;
      RECT 54.97 2.785 54.98 3.08 ;
      RECT 54.96 2.82 54.97 3.08 ;
      RECT 54.955 2.855 54.96 3.08 ;
      RECT 55.075 2.62 55.08 3.08 ;
      RECT 54.59 2.722 54.775 2.895 ;
      RECT 54.55 2.64 54.735 2.893 ;
      RECT 54.511 2.645 54.735 2.889 ;
      RECT 54.425 2.654 54.735 2.884 ;
      RECT 54.341 2.67 54.74 2.879 ;
      RECT 54.255 2.69 54.765 2.873 ;
      RECT 54.255 2.71 54.77 2.873 ;
      RECT 54.341 2.68 54.765 2.879 ;
      RECT 54.425 2.655 54.74 2.884 ;
      RECT 54.59 2.637 54.735 2.895 ;
      RECT 54.59 2.632 54.69 2.895 ;
      RECT 54.676 2.626 54.69 2.895 ;
      RECT 54.065 1.95 54.07 2.349 ;
      RECT 53.81 1.95 53.845 2.347 ;
      RECT 53.405 1.985 53.41 2.341 ;
      RECT 54.15 1.988 54.155 2.243 ;
      RECT 54.145 1.986 54.15 2.249 ;
      RECT 54.14 1.985 54.145 2.256 ;
      RECT 54.115 1.978 54.14 2.28 ;
      RECT 54.11 1.971 54.115 2.304 ;
      RECT 54.105 1.967 54.11 2.313 ;
      RECT 54.095 1.962 54.105 2.326 ;
      RECT 54.09 1.959 54.095 2.335 ;
      RECT 54.085 1.957 54.09 2.34 ;
      RECT 54.07 1.953 54.085 2.35 ;
      RECT 54.055 1.947 54.065 2.349 ;
      RECT 54.017 1.945 54.055 2.349 ;
      RECT 53.931 1.947 54.017 2.349 ;
      RECT 53.845 1.949 53.931 2.348 ;
      RECT 53.774 1.95 53.81 2.347 ;
      RECT 53.688 1.952 53.774 2.347 ;
      RECT 53.602 1.954 53.688 2.346 ;
      RECT 53.516 1.956 53.602 2.346 ;
      RECT 53.43 1.959 53.516 2.345 ;
      RECT 53.42 1.965 53.43 2.344 ;
      RECT 53.41 1.977 53.42 2.342 ;
      RECT 53.35 2.012 53.405 2.338 ;
      RECT 53.345 2.042 53.35 2.1 ;
      RECT 54.09 3.122 54.105 3.315 ;
      RECT 54.085 3.09 54.09 3.315 ;
      RECT 54.075 3.065 54.085 3.315 ;
      RECT 54.07 3.037 54.075 3.315 ;
      RECT 54.04 2.96 54.07 3.315 ;
      RECT 54.015 2.842 54.04 3.315 ;
      RECT 54.01 2.78 54.015 3.315 ;
      RECT 54 2.767 54.01 3.315 ;
      RECT 53.98 2.757 54 3.315 ;
      RECT 53.965 2.74 53.98 3.315 ;
      RECT 53.935 2.728 53.965 3.315 ;
      RECT 53.93 2.727 53.935 3.26 ;
      RECT 53.925 2.727 53.93 3.218 ;
      RECT 53.91 2.726 53.925 3.17 ;
      RECT 53.895 2.726 53.91 3.108 ;
      RECT 53.875 2.726 53.895 3.068 ;
      RECT 53.87 2.726 53.875 3.053 ;
      RECT 53.845 2.725 53.87 3.048 ;
      RECT 53.775 2.724 53.845 3.035 ;
      RECT 53.76 2.723 53.775 3.02 ;
      RECT 53.73 2.722 53.76 3.003 ;
      RECT 53.725 2.722 53.73 2.988 ;
      RECT 53.675 2.721 53.725 2.968 ;
      RECT 53.61 2.72 53.675 2.923 ;
      RECT 53.605 2.72 53.61 2.895 ;
      RECT 53.69 3.257 53.695 3.514 ;
      RECT 53.67 3.176 53.69 3.531 ;
      RECT 53.65 3.17 53.67 3.56 ;
      RECT 53.59 3.157 53.65 3.58 ;
      RECT 53.545 3.141 53.59 3.581 ;
      RECT 53.461 3.129 53.545 3.569 ;
      RECT 53.375 3.116 53.461 3.553 ;
      RECT 53.365 3.109 53.375 3.545 ;
      RECT 53.32 3.106 53.365 3.485 ;
      RECT 53.3 3.102 53.32 3.4 ;
      RECT 53.285 3.1 53.3 3.353 ;
      RECT 53.255 3.097 53.285 3.323 ;
      RECT 53.22 3.093 53.255 3.3 ;
      RECT 53.177 3.088 53.22 3.288 ;
      RECT 53.091 3.079 53.177 3.297 ;
      RECT 53.005 3.068 53.091 3.309 ;
      RECT 52.94 3.059 53.005 3.318 ;
      RECT 52.92 3.05 52.94 3.323 ;
      RECT 52.915 3.043 52.92 3.325 ;
      RECT 52.875 3.028 52.915 3.322 ;
      RECT 52.855 3.007 52.875 3.317 ;
      RECT 52.84 2.995 52.855 3.31 ;
      RECT 52.835 2.987 52.84 3.303 ;
      RECT 52.82 2.967 52.835 3.296 ;
      RECT 52.815 2.83 52.82 3.29 ;
      RECT 52.735 2.719 52.815 3.262 ;
      RECT 52.726 2.712 52.735 3.228 ;
      RECT 52.64 2.706 52.726 3.153 ;
      RECT 52.615 2.697 52.64 3.065 ;
      RECT 52.585 2.692 52.615 3.04 ;
      RECT 52.52 2.701 52.585 3.025 ;
      RECT 52.5 2.717 52.52 3 ;
      RECT 52.49 2.723 52.5 2.948 ;
      RECT 52.47 2.745 52.49 2.83 ;
      RECT 53.125 2.71 53.295 2.895 ;
      RECT 53.125 2.71 53.33 2.893 ;
      RECT 53.175 2.62 53.345 2.884 ;
      RECT 53.125 2.777 53.35 2.877 ;
      RECT 53.14 2.655 53.345 2.884 ;
      RECT 52.34 3.388 52.405 3.831 ;
      RECT 52.28 3.413 52.405 3.829 ;
      RECT 52.28 3.413 52.46 3.823 ;
      RECT 52.265 3.438 52.46 3.822 ;
      RECT 52.405 3.375 52.48 3.819 ;
      RECT 52.34 3.4 52.56 3.813 ;
      RECT 52.265 3.439 52.605 3.807 ;
      RECT 52.25 3.466 52.605 3.798 ;
      RECT 52.265 3.459 52.625 3.79 ;
      RECT 52.25 3.468 52.63 3.773 ;
      RECT 52.245 3.485 52.63 3.6 ;
      RECT 52.25 2.207 52.285 2.445 ;
      RECT 52.25 2.207 52.315 2.444 ;
      RECT 52.25 2.207 52.43 2.44 ;
      RECT 52.25 2.207 52.485 2.418 ;
      RECT 52.26 2.15 52.54 2.318 ;
      RECT 52.365 1.99 52.395 2.441 ;
      RECT 52.395 1.985 52.575 2.198 ;
      RECT 52.265 2.126 52.575 2.198 ;
      RECT 52.315 2.022 52.365 2.442 ;
      RECT 52.285 2.078 52.575 2.198 ;
      RECT 50.79 1.74 50.96 2.935 ;
      RECT 50.79 1.74 51.255 1.91 ;
      RECT 50.79 6.97 51.255 7.14 ;
      RECT 50.79 5.945 50.96 7.14 ;
      RECT 49.8 1.74 49.97 2.935 ;
      RECT 49.8 1.74 50.265 1.91 ;
      RECT 49.8 6.97 50.265 7.14 ;
      RECT 49.8 5.945 49.97 7.14 ;
      RECT 47.945 2.635 48.115 3.865 ;
      RECT 48 0.855 48.17 2.805 ;
      RECT 47.945 0.575 48.115 1.025 ;
      RECT 47.945 7.855 48.115 8.305 ;
      RECT 48 6.075 48.17 8.025 ;
      RECT 47.945 5.015 48.115 6.245 ;
      RECT 47.425 0.575 47.595 3.865 ;
      RECT 47.425 2.075 47.83 2.405 ;
      RECT 47.425 1.235 47.83 1.565 ;
      RECT 47.425 5.015 47.595 8.305 ;
      RECT 47.425 7.315 47.83 7.645 ;
      RECT 47.425 6.475 47.83 6.805 ;
      RECT 45.525 3.392 45.54 3.443 ;
      RECT 45.52 3.372 45.525 3.49 ;
      RECT 45.505 3.362 45.52 3.558 ;
      RECT 45.48 3.342 45.505 3.613 ;
      RECT 45.44 3.327 45.48 3.633 ;
      RECT 45.395 3.321 45.44 3.661 ;
      RECT 45.325 3.311 45.395 3.678 ;
      RECT 45.305 3.303 45.325 3.678 ;
      RECT 45.245 3.297 45.305 3.67 ;
      RECT 45.186 3.288 45.245 3.658 ;
      RECT 45.1 3.277 45.186 3.641 ;
      RECT 45.078 3.268 45.1 3.629 ;
      RECT 44.992 3.261 45.078 3.616 ;
      RECT 44.906 3.248 44.992 3.597 ;
      RECT 44.82 3.236 44.906 3.577 ;
      RECT 44.79 3.225 44.82 3.564 ;
      RECT 44.74 3.211 44.79 3.556 ;
      RECT 44.72 3.2 44.74 3.548 ;
      RECT 44.671 3.189 44.72 3.54 ;
      RECT 44.585 3.168 44.671 3.525 ;
      RECT 44.54 3.155 44.585 3.51 ;
      RECT 44.495 3.155 44.54 3.49 ;
      RECT 44.44 3.155 44.495 3.425 ;
      RECT 44.415 3.155 44.44 3.348 ;
      RECT 44.94 2.892 45.11 3.075 ;
      RECT 44.94 2.892 45.125 3.033 ;
      RECT 44.94 2.892 45.13 2.975 ;
      RECT 45 2.66 45.135 2.951 ;
      RECT 45 2.664 45.14 2.934 ;
      RECT 44.945 2.827 45.14 2.934 ;
      RECT 44.97 2.672 45.11 3.075 ;
      RECT 44.97 2.676 45.15 2.875 ;
      RECT 44.955 2.762 45.15 2.875 ;
      RECT 44.965 2.692 45.11 3.075 ;
      RECT 44.965 2.695 45.16 2.788 ;
      RECT 44.96 2.712 45.16 2.788 ;
      RECT 44.73 1.932 44.9 2.415 ;
      RECT 44.725 1.927 44.875 2.405 ;
      RECT 44.725 1.934 44.905 2.399 ;
      RECT 44.715 1.928 44.875 2.378 ;
      RECT 44.715 1.944 44.92 2.337 ;
      RECT 44.685 1.929 44.875 2.3 ;
      RECT 44.685 1.959 44.93 2.24 ;
      RECT 44.68 1.931 44.875 2.238 ;
      RECT 44.66 1.94 44.905 2.195 ;
      RECT 44.635 1.956 44.92 2.107 ;
      RECT 44.635 1.975 44.945 2.098 ;
      RECT 44.63 2.012 44.945 2.05 ;
      RECT 44.635 1.992 44.95 2.018 ;
      RECT 44.73 1.926 44.84 2.415 ;
      RECT 44.816 1.925 44.84 2.415 ;
      RECT 44.05 2.71 44.055 2.921 ;
      RECT 44.65 2.71 44.655 2.895 ;
      RECT 44.715 2.75 44.72 2.863 ;
      RECT 44.71 2.742 44.715 2.869 ;
      RECT 44.705 2.732 44.71 2.877 ;
      RECT 44.7 2.722 44.705 2.886 ;
      RECT 44.695 2.712 44.7 2.89 ;
      RECT 44.655 2.71 44.695 2.893 ;
      RECT 44.627 2.709 44.65 2.897 ;
      RECT 44.541 2.706 44.627 2.904 ;
      RECT 44.455 2.702 44.541 2.915 ;
      RECT 44.435 2.7 44.455 2.921 ;
      RECT 44.417 2.699 44.435 2.924 ;
      RECT 44.331 2.697 44.417 2.931 ;
      RECT 44.245 2.692 44.331 2.944 ;
      RECT 44.226 2.689 44.245 2.949 ;
      RECT 44.14 2.687 44.226 2.94 ;
      RECT 44.13 2.687 44.14 2.933 ;
      RECT 44.055 2.7 44.13 2.927 ;
      RECT 44.04 2.711 44.05 2.921 ;
      RECT 44.03 2.713 44.04 2.92 ;
      RECT 44.02 2.717 44.03 2.916 ;
      RECT 44.015 2.72 44.02 2.91 ;
      RECT 44.005 2.722 44.015 2.904 ;
      RECT 44 2.725 44.005 2.898 ;
      RECT 43.98 3.311 43.985 3.515 ;
      RECT 43.965 3.298 43.98 3.608 ;
      RECT 43.95 3.279 43.965 3.885 ;
      RECT 43.915 3.245 43.95 3.885 ;
      RECT 43.911 3.215 43.915 3.885 ;
      RECT 43.825 3.097 43.911 3.885 ;
      RECT 43.815 2.972 43.825 3.885 ;
      RECT 43.8 2.94 43.815 3.885 ;
      RECT 43.795 2.915 43.8 3.885 ;
      RECT 43.79 2.905 43.795 3.841 ;
      RECT 43.775 2.877 43.79 3.746 ;
      RECT 43.76 2.843 43.775 3.645 ;
      RECT 43.755 2.821 43.76 3.598 ;
      RECT 43.75 2.81 43.755 3.568 ;
      RECT 43.745 2.8 43.75 3.534 ;
      RECT 43.735 2.787 43.745 3.502 ;
      RECT 43.71 2.763 43.735 3.428 ;
      RECT 43.705 2.743 43.71 3.353 ;
      RECT 43.7 2.737 43.705 3.328 ;
      RECT 43.695 2.732 43.7 3.293 ;
      RECT 43.69 2.727 43.695 3.268 ;
      RECT 43.685 2.725 43.69 3.248 ;
      RECT 43.68 2.725 43.685 3.233 ;
      RECT 43.675 2.725 43.68 3.193 ;
      RECT 43.665 2.725 43.675 3.165 ;
      RECT 43.655 2.725 43.665 3.11 ;
      RECT 43.64 2.725 43.655 3.048 ;
      RECT 43.635 2.724 43.64 2.993 ;
      RECT 43.62 2.723 43.635 2.973 ;
      RECT 43.56 2.721 43.62 2.947 ;
      RECT 43.525 2.722 43.56 2.927 ;
      RECT 43.52 2.724 43.525 2.917 ;
      RECT 43.51 2.743 43.52 2.907 ;
      RECT 43.505 2.77 43.51 2.838 ;
      RECT 43.62 2.195 43.79 2.44 ;
      RECT 43.655 1.966 43.79 2.44 ;
      RECT 43.655 1.968 43.8 2.435 ;
      RECT 43.655 1.97 43.825 2.423 ;
      RECT 43.655 1.973 43.85 2.405 ;
      RECT 43.655 1.978 43.9 2.378 ;
      RECT 43.655 1.983 43.92 2.343 ;
      RECT 43.635 1.985 43.93 2.318 ;
      RECT 43.625 2.08 43.93 2.318 ;
      RECT 43.655 1.965 43.765 2.44 ;
      RECT 43.665 1.962 43.76 2.44 ;
      RECT 43.185 3.227 43.375 3.585 ;
      RECT 43.185 3.239 43.41 3.584 ;
      RECT 43.185 3.267 43.43 3.582 ;
      RECT 43.185 3.292 43.435 3.581 ;
      RECT 43.185 3.35 43.45 3.58 ;
      RECT 43.17 3.223 43.33 3.565 ;
      RECT 43.15 3.232 43.375 3.518 ;
      RECT 43.125 3.243 43.41 3.455 ;
      RECT 43.125 3.327 43.445 3.455 ;
      RECT 43.125 3.302 43.44 3.455 ;
      RECT 43.185 3.218 43.33 3.585 ;
      RECT 43.271 3.217 43.33 3.585 ;
      RECT 43.271 3.216 43.315 3.585 ;
      RECT 43.185 7.855 43.355 8.305 ;
      RECT 43.24 6.075 43.41 8.025 ;
      RECT 43.185 5.015 43.355 6.245 ;
      RECT 42.665 5.015 42.835 8.305 ;
      RECT 42.665 7.315 43.07 7.645 ;
      RECT 42.665 6.475 43.07 6.805 ;
      RECT 42.97 2.732 42.975 3.11 ;
      RECT 42.965 2.7 42.97 3.11 ;
      RECT 42.96 2.672 42.965 3.11 ;
      RECT 42.955 2.652 42.96 3.11 ;
      RECT 42.9 2.635 42.955 3.11 ;
      RECT 42.86 2.62 42.9 3.11 ;
      RECT 42.805 2.607 42.86 3.11 ;
      RECT 42.77 2.598 42.805 3.11 ;
      RECT 42.766 2.596 42.77 3.109 ;
      RECT 42.68 2.592 42.766 3.092 ;
      RECT 42.595 2.584 42.68 3.055 ;
      RECT 42.585 2.58 42.595 3.028 ;
      RECT 42.575 2.58 42.585 3.01 ;
      RECT 42.565 2.582 42.575 2.993 ;
      RECT 42.56 2.587 42.565 2.979 ;
      RECT 42.555 2.591 42.56 2.966 ;
      RECT 42.545 2.596 42.555 2.95 ;
      RECT 42.53 2.61 42.545 2.925 ;
      RECT 42.525 2.616 42.53 2.905 ;
      RECT 42.52 2.618 42.525 2.898 ;
      RECT 42.515 2.622 42.52 2.773 ;
      RECT 42.695 3.422 42.94 3.885 ;
      RECT 42.615 3.395 42.935 3.881 ;
      RECT 42.545 3.43 42.94 3.874 ;
      RECT 42.335 3.685 42.94 3.87 ;
      RECT 42.515 3.453 42.94 3.87 ;
      RECT 42.355 3.645 42.94 3.87 ;
      RECT 42.505 3.465 42.94 3.87 ;
      RECT 42.39 3.582 42.94 3.87 ;
      RECT 42.445 3.507 42.94 3.87 ;
      RECT 42.695 3.372 42.935 3.885 ;
      RECT 42.725 3.365 42.935 3.885 ;
      RECT 42.715 3.367 42.935 3.885 ;
      RECT 42.725 3.362 42.855 3.885 ;
      RECT 42.28 1.925 42.366 2.364 ;
      RECT 42.275 1.925 42.366 2.362 ;
      RECT 42.275 1.925 42.435 2.361 ;
      RECT 42.275 1.925 42.465 2.358 ;
      RECT 42.26 1.932 42.465 2.349 ;
      RECT 42.26 1.932 42.47 2.345 ;
      RECT 42.255 1.942 42.47 2.338 ;
      RECT 42.25 1.947 42.47 2.313 ;
      RECT 42.25 1.947 42.485 2.295 ;
      RECT 42.275 1.925 42.505 2.21 ;
      RECT 42.245 1.952 42.505 2.208 ;
      RECT 42.255 1.945 42.51 2.146 ;
      RECT 42.245 2.067 42.515 2.129 ;
      RECT 42.23 1.962 42.51 2.08 ;
      RECT 42.225 1.972 42.51 1.98 ;
      RECT 42.305 2.743 42.31 2.82 ;
      RECT 42.295 2.737 42.305 3.01 ;
      RECT 42.285 2.729 42.295 3.031 ;
      RECT 42.275 2.72 42.285 3.053 ;
      RECT 42.27 2.715 42.275 3.07 ;
      RECT 42.23 2.715 42.27 3.11 ;
      RECT 42.21 2.715 42.23 3.165 ;
      RECT 42.205 2.715 42.21 3.193 ;
      RECT 42.195 2.715 42.205 3.208 ;
      RECT 42.16 2.715 42.195 3.25 ;
      RECT 42.155 2.715 42.16 3.293 ;
      RECT 42.145 2.715 42.155 3.308 ;
      RECT 42.13 2.715 42.145 3.328 ;
      RECT 42.115 2.715 42.13 3.355 ;
      RECT 42.11 2.716 42.115 3.373 ;
      RECT 42.09 2.717 42.11 3.38 ;
      RECT 42.035 2.718 42.09 3.4 ;
      RECT 42.025 2.719 42.035 3.414 ;
      RECT 42.02 2.722 42.025 3.413 ;
      RECT 41.98 2.795 42.02 3.411 ;
      RECT 41.965 2.875 41.98 3.409 ;
      RECT 41.94 2.93 41.965 3.407 ;
      RECT 41.925 2.995 41.94 3.406 ;
      RECT 41.88 3.027 41.925 3.403 ;
      RECT 41.795 3.05 41.88 3.398 ;
      RECT 41.77 3.07 41.795 3.393 ;
      RECT 41.7 3.075 41.77 3.389 ;
      RECT 41.68 3.077 41.7 3.386 ;
      RECT 41.595 3.088 41.68 3.38 ;
      RECT 41.59 3.099 41.595 3.375 ;
      RECT 41.58 3.101 41.59 3.375 ;
      RECT 41.545 3.105 41.58 3.373 ;
      RECT 41.495 3.115 41.545 3.36 ;
      RECT 41.475 3.123 41.495 3.345 ;
      RECT 41.395 3.135 41.475 3.328 ;
      RECT 41.56 2.685 41.73 2.895 ;
      RECT 41.676 2.681 41.73 2.895 ;
      RECT 41.481 2.685 41.73 2.886 ;
      RECT 41.481 2.685 41.735 2.875 ;
      RECT 41.395 2.685 41.735 2.866 ;
      RECT 41.395 2.693 41.745 2.81 ;
      RECT 41.395 2.705 41.75 2.723 ;
      RECT 41.395 2.712 41.755 2.715 ;
      RECT 41.59 2.683 41.73 2.895 ;
      RECT 41.345 3.628 41.59 3.96 ;
      RECT 41.34 3.62 41.345 3.957 ;
      RECT 41.31 3.64 41.59 3.938 ;
      RECT 41.29 3.672 41.59 3.911 ;
      RECT 41.34 3.625 41.517 3.957 ;
      RECT 41.34 3.622 41.431 3.957 ;
      RECT 41.28 1.97 41.45 2.39 ;
      RECT 41.275 1.97 41.45 2.388 ;
      RECT 41.275 1.97 41.475 2.378 ;
      RECT 41.275 1.97 41.495 2.353 ;
      RECT 41.27 1.97 41.495 2.348 ;
      RECT 41.27 1.97 41.505 2.338 ;
      RECT 41.27 1.97 41.51 2.333 ;
      RECT 41.27 1.975 41.515 2.328 ;
      RECT 41.27 2.007 41.53 2.318 ;
      RECT 41.27 2.077 41.555 2.301 ;
      RECT 41.25 2.077 41.555 2.293 ;
      RECT 41.25 2.137 41.565 2.27 ;
      RECT 41.25 2.177 41.575 2.215 ;
      RECT 41.235 1.97 41.51 2.195 ;
      RECT 41.225 1.985 41.515 2.093 ;
      RECT 40.815 3.375 40.985 3.9 ;
      RECT 40.81 3.375 40.985 3.893 ;
      RECT 40.8 3.375 40.99 3.858 ;
      RECT 40.795 3.385 40.99 3.83 ;
      RECT 40.79 3.405 40.99 3.813 ;
      RECT 40.8 3.38 40.995 3.803 ;
      RECT 40.785 3.425 40.995 3.795 ;
      RECT 40.78 3.445 40.995 3.78 ;
      RECT 40.775 3.475 40.995 3.77 ;
      RECT 40.765 3.52 40.995 3.745 ;
      RECT 40.795 3.39 41 3.728 ;
      RECT 40.76 3.572 41 3.723 ;
      RECT 40.795 3.4 41.005 3.693 ;
      RECT 40.755 3.605 41.005 3.69 ;
      RECT 40.75 3.63 41.005 3.67 ;
      RECT 40.79 3.417 41.015 3.61 ;
      RECT 40.785 3.439 41.025 3.503 ;
      RECT 40.735 2.686 40.75 2.955 ;
      RECT 40.69 2.67 40.735 3 ;
      RECT 40.685 2.658 40.69 3.05 ;
      RECT 40.675 2.654 40.685 3.083 ;
      RECT 40.67 2.651 40.675 3.111 ;
      RECT 40.655 2.653 40.67 3.153 ;
      RECT 40.65 2.657 40.655 3.193 ;
      RECT 40.63 2.662 40.65 3.245 ;
      RECT 40.626 2.667 40.63 3.302 ;
      RECT 40.54 2.686 40.626 3.339 ;
      RECT 40.53 2.707 40.54 3.375 ;
      RECT 40.525 2.715 40.53 3.376 ;
      RECT 40.52 2.757 40.525 3.377 ;
      RECT 40.505 2.845 40.52 3.378 ;
      RECT 40.495 2.995 40.505 3.38 ;
      RECT 40.49 3.04 40.495 3.382 ;
      RECT 40.455 3.082 40.49 3.385 ;
      RECT 40.45 3.1 40.455 3.388 ;
      RECT 40.373 3.106 40.45 3.394 ;
      RECT 40.287 3.12 40.373 3.407 ;
      RECT 40.201 3.134 40.287 3.421 ;
      RECT 40.115 3.148 40.201 3.434 ;
      RECT 40.055 3.16 40.115 3.446 ;
      RECT 40.03 3.167 40.055 3.453 ;
      RECT 40.016 3.17 40.03 3.458 ;
      RECT 39.93 3.178 40.016 3.474 ;
      RECT 39.925 3.185 39.93 3.489 ;
      RECT 39.901 3.185 39.925 3.496 ;
      RECT 39.815 3.188 39.901 3.524 ;
      RECT 39.73 3.192 39.815 3.568 ;
      RECT 39.665 3.196 39.73 3.605 ;
      RECT 39.64 3.199 39.665 3.621 ;
      RECT 39.565 3.212 39.64 3.625 ;
      RECT 39.54 3.23 39.565 3.629 ;
      RECT 39.53 3.237 39.54 3.631 ;
      RECT 39.515 3.24 39.53 3.632 ;
      RECT 39.455 3.252 39.515 3.636 ;
      RECT 39.445 3.266 39.455 3.64 ;
      RECT 39.39 3.276 39.445 3.628 ;
      RECT 39.365 3.297 39.39 3.611 ;
      RECT 39.345 3.317 39.365 3.602 ;
      RECT 39.34 3.33 39.345 3.597 ;
      RECT 39.325 3.342 39.34 3.593 ;
      RECT 40.56 1.997 40.565 2.02 ;
      RECT 40.555 1.988 40.56 2.06 ;
      RECT 40.55 1.986 40.555 2.103 ;
      RECT 40.545 1.977 40.55 2.138 ;
      RECT 40.54 1.967 40.545 2.21 ;
      RECT 40.535 1.957 40.54 2.275 ;
      RECT 40.53 1.954 40.535 2.315 ;
      RECT 40.505 1.948 40.53 2.405 ;
      RECT 40.47 1.936 40.505 2.43 ;
      RECT 40.46 1.927 40.47 2.43 ;
      RECT 40.325 1.925 40.335 2.413 ;
      RECT 40.315 1.925 40.325 2.38 ;
      RECT 40.31 1.925 40.315 2.355 ;
      RECT 40.305 1.925 40.31 2.343 ;
      RECT 40.3 1.925 40.305 2.325 ;
      RECT 40.29 1.925 40.3 2.29 ;
      RECT 40.285 1.927 40.29 2.268 ;
      RECT 40.28 1.933 40.285 2.253 ;
      RECT 40.275 1.939 40.28 2.238 ;
      RECT 40.26 1.951 40.275 2.211 ;
      RECT 40.255 1.962 40.26 2.179 ;
      RECT 40.25 1.972 40.255 2.163 ;
      RECT 40.24 1.98 40.25 2.132 ;
      RECT 40.235 1.99 40.24 2.106 ;
      RECT 40.23 2.047 40.235 2.089 ;
      RECT 40.335 1.925 40.46 2.43 ;
      RECT 40.05 2.612 40.31 2.91 ;
      RECT 40.045 2.619 40.31 2.908 ;
      RECT 40.05 2.614 40.325 2.903 ;
      RECT 40.04 2.627 40.325 2.9 ;
      RECT 40.04 2.632 40.33 2.893 ;
      RECT 40.035 2.64 40.33 2.89 ;
      RECT 40.035 2.657 40.335 2.688 ;
      RECT 40.05 2.609 40.281 2.91 ;
      RECT 40.105 2.608 40.281 2.91 ;
      RECT 40.105 2.605 40.195 2.91 ;
      RECT 40.105 2.602 40.191 2.91 ;
      RECT 39.795 2.875 39.8 2.888 ;
      RECT 39.79 2.842 39.795 2.893 ;
      RECT 39.785 2.797 39.79 2.9 ;
      RECT 39.78 2.752 39.785 2.908 ;
      RECT 39.775 2.72 39.78 2.916 ;
      RECT 39.77 2.68 39.775 2.917 ;
      RECT 39.755 2.66 39.77 2.919 ;
      RECT 39.68 2.642 39.755 2.931 ;
      RECT 39.67 2.635 39.68 2.942 ;
      RECT 39.665 2.635 39.67 2.944 ;
      RECT 39.635 2.641 39.665 2.948 ;
      RECT 39.595 2.654 39.635 2.948 ;
      RECT 39.57 2.665 39.595 2.934 ;
      RECT 39.555 2.671 39.57 2.917 ;
      RECT 39.545 2.673 39.555 2.908 ;
      RECT 39.54 2.674 39.545 2.903 ;
      RECT 39.535 2.675 39.54 2.898 ;
      RECT 39.53 2.676 39.535 2.895 ;
      RECT 39.505 2.681 39.53 2.885 ;
      RECT 39.495 2.697 39.505 2.872 ;
      RECT 39.49 2.717 39.495 2.867 ;
      RECT 39.5 2.11 39.505 2.306 ;
      RECT 39.485 2.074 39.5 2.308 ;
      RECT 39.475 2.056 39.485 2.313 ;
      RECT 39.465 2.042 39.475 2.317 ;
      RECT 39.42 2.026 39.465 2.327 ;
      RECT 39.415 2.016 39.42 2.336 ;
      RECT 39.37 2.005 39.415 2.342 ;
      RECT 39.365 1.993 39.37 2.349 ;
      RECT 39.35 1.988 39.365 2.353 ;
      RECT 39.335 1.98 39.35 2.358 ;
      RECT 39.325 1.973 39.335 2.363 ;
      RECT 39.315 1.97 39.325 2.368 ;
      RECT 39.305 1.97 39.315 2.369 ;
      RECT 39.3 1.967 39.305 2.368 ;
      RECT 39.265 1.962 39.29 2.367 ;
      RECT 39.241 1.958 39.265 2.366 ;
      RECT 39.155 1.949 39.241 2.363 ;
      RECT 39.14 1.941 39.155 2.36 ;
      RECT 39.118 1.94 39.14 2.359 ;
      RECT 39.032 1.94 39.118 2.357 ;
      RECT 38.946 1.94 39.032 2.355 ;
      RECT 38.86 1.94 38.946 2.352 ;
      RECT 38.85 1.94 38.86 2.343 ;
      RECT 38.82 1.94 38.85 2.303 ;
      RECT 38.81 1.95 38.82 2.258 ;
      RECT 38.805 1.99 38.81 2.243 ;
      RECT 38.8 2.005 38.805 2.23 ;
      RECT 38.77 2.085 38.8 2.192 ;
      RECT 39.29 1.965 39.3 2.368 ;
      RECT 39.115 2.73 39.13 3.335 ;
      RECT 39.12 2.725 39.13 3.335 ;
      RECT 39.285 2.725 39.29 2.908 ;
      RECT 39.275 2.725 39.285 2.938 ;
      RECT 39.26 2.725 39.275 2.998 ;
      RECT 39.255 2.725 39.26 3.043 ;
      RECT 39.25 2.725 39.255 3.073 ;
      RECT 39.245 2.725 39.25 3.093 ;
      RECT 39.235 2.725 39.245 3.128 ;
      RECT 39.22 2.725 39.235 3.16 ;
      RECT 39.175 2.725 39.22 3.188 ;
      RECT 39.17 2.725 39.175 3.218 ;
      RECT 39.165 2.725 39.17 3.23 ;
      RECT 39.16 2.725 39.165 3.238 ;
      RECT 39.15 2.725 39.16 3.253 ;
      RECT 39.145 2.725 39.15 3.275 ;
      RECT 39.135 2.725 39.145 3.298 ;
      RECT 39.13 2.725 39.135 3.318 ;
      RECT 39.095 2.74 39.115 3.335 ;
      RECT 39.07 2.757 39.095 3.335 ;
      RECT 39.065 2.767 39.07 3.335 ;
      RECT 39.035 2.782 39.065 3.335 ;
      RECT 38.96 2.824 39.035 3.335 ;
      RECT 38.955 2.855 38.96 3.318 ;
      RECT 38.95 2.859 38.955 3.3 ;
      RECT 38.945 2.863 38.95 3.263 ;
      RECT 38.94 3.047 38.945 3.23 ;
      RECT 38.425 3.236 38.511 3.801 ;
      RECT 38.38 3.238 38.545 3.795 ;
      RECT 38.511 3.235 38.545 3.795 ;
      RECT 38.425 3.237 38.63 3.789 ;
      RECT 38.38 3.247 38.64 3.785 ;
      RECT 38.355 3.239 38.63 3.781 ;
      RECT 38.35 3.242 38.63 3.776 ;
      RECT 38.325 3.257 38.64 3.77 ;
      RECT 38.325 3.282 38.68 3.765 ;
      RECT 38.285 3.29 38.68 3.74 ;
      RECT 38.285 3.317 38.695 3.738 ;
      RECT 38.285 3.347 38.705 3.725 ;
      RECT 38.28 3.492 38.705 3.713 ;
      RECT 38.285 3.421 38.725 3.71 ;
      RECT 38.285 3.478 38.73 3.518 ;
      RECT 38.475 2.757 38.645 2.935 ;
      RECT 38.425 2.696 38.475 2.92 ;
      RECT 38.16 2.676 38.425 2.905 ;
      RECT 38.12 2.74 38.595 2.905 ;
      RECT 38.12 2.73 38.55 2.905 ;
      RECT 38.12 2.727 38.54 2.905 ;
      RECT 38.12 2.715 38.53 2.905 ;
      RECT 38.12 2.7 38.475 2.905 ;
      RECT 38.16 2.672 38.361 2.905 ;
      RECT 38.17 2.65 38.361 2.905 ;
      RECT 38.195 2.635 38.275 2.905 ;
      RECT 37.95 3.165 38.07 3.61 ;
      RECT 37.935 3.165 38.07 3.609 ;
      RECT 37.89 3.187 38.07 3.604 ;
      RECT 37.85 3.236 38.07 3.598 ;
      RECT 37.85 3.236 38.075 3.573 ;
      RECT 37.85 3.236 38.095 3.463 ;
      RECT 37.845 3.266 38.095 3.46 ;
      RECT 37.935 3.165 38.105 3.355 ;
      RECT 37.595 1.95 37.6 2.395 ;
      RECT 37.405 1.95 37.425 2.36 ;
      RECT 37.375 1.95 37.38 2.335 ;
      RECT 38.055 2.257 38.07 2.445 ;
      RECT 38.05 2.242 38.055 2.451 ;
      RECT 38.03 2.215 38.05 2.454 ;
      RECT 37.98 2.182 38.03 2.463 ;
      RECT 37.95 2.162 37.98 2.467 ;
      RECT 37.931 2.15 37.95 2.463 ;
      RECT 37.845 2.122 37.931 2.453 ;
      RECT 37.835 2.097 37.845 2.443 ;
      RECT 37.765 2.065 37.835 2.435 ;
      RECT 37.74 2.025 37.765 2.427 ;
      RECT 37.72 2.007 37.74 2.421 ;
      RECT 37.71 1.997 37.72 2.418 ;
      RECT 37.7 1.99 37.71 2.416 ;
      RECT 37.68 1.977 37.7 2.413 ;
      RECT 37.67 1.967 37.68 2.41 ;
      RECT 37.66 1.96 37.67 2.408 ;
      RECT 37.61 1.952 37.66 2.402 ;
      RECT 37.6 1.95 37.61 2.396 ;
      RECT 37.57 1.95 37.595 2.393 ;
      RECT 37.541 1.95 37.57 2.388 ;
      RECT 37.455 1.95 37.541 2.378 ;
      RECT 37.425 1.95 37.455 2.365 ;
      RECT 37.38 1.95 37.405 2.348 ;
      RECT 37.365 1.95 37.375 2.33 ;
      RECT 37.345 1.957 37.365 2.315 ;
      RECT 37.34 1.972 37.345 2.303 ;
      RECT 37.335 1.977 37.34 2.243 ;
      RECT 37.33 1.982 37.335 2.085 ;
      RECT 37.325 1.985 37.33 2.003 ;
      RECT 37.59 2.67 37.676 2.991 ;
      RECT 37.59 2.67 37.71 2.984 ;
      RECT 37.54 2.67 37.71 2.98 ;
      RECT 37.54 2.672 37.796 2.978 ;
      RECT 37.54 2.674 37.82 2.972 ;
      RECT 37.54 2.681 37.83 2.971 ;
      RECT 37.54 2.69 37.835 2.968 ;
      RECT 37.54 2.696 37.84 2.963 ;
      RECT 37.54 2.74 37.845 2.96 ;
      RECT 37.54 2.832 37.85 2.957 ;
      RECT 37.065 3.275 37.1 3.595 ;
      RECT 37.65 3.46 37.655 3.642 ;
      RECT 37.605 3.342 37.65 3.661 ;
      RECT 37.59 3.319 37.605 3.684 ;
      RECT 37.58 3.309 37.59 3.694 ;
      RECT 37.56 3.304 37.58 3.707 ;
      RECT 37.535 3.302 37.56 3.728 ;
      RECT 37.516 3.301 37.535 3.74 ;
      RECT 37.43 3.298 37.516 3.74 ;
      RECT 37.36 3.293 37.43 3.728 ;
      RECT 37.285 3.289 37.36 3.703 ;
      RECT 37.22 3.285 37.285 3.67 ;
      RECT 37.15 3.282 37.22 3.63 ;
      RECT 37.12 3.278 37.15 3.605 ;
      RECT 37.1 3.276 37.12 3.598 ;
      RECT 37.016 3.274 37.065 3.596 ;
      RECT 36.93 3.271 37.016 3.597 ;
      RECT 36.855 3.27 36.93 3.599 ;
      RECT 36.77 3.27 36.855 3.625 ;
      RECT 36.693 3.271 36.77 3.65 ;
      RECT 36.607 3.272 36.693 3.65 ;
      RECT 36.521 3.272 36.607 3.65 ;
      RECT 36.435 3.273 36.521 3.65 ;
      RECT 36.415 3.274 36.435 3.642 ;
      RECT 36.4 3.28 36.415 3.627 ;
      RECT 36.365 3.3 36.4 3.607 ;
      RECT 36.355 3.32 36.365 3.589 ;
      RECT 37.325 2.625 37.33 2.895 ;
      RECT 37.32 2.616 37.325 2.9 ;
      RECT 37.31 2.606 37.32 2.912 ;
      RECT 37.305 2.595 37.31 2.923 ;
      RECT 37.285 2.589 37.305 2.941 ;
      RECT 37.24 2.586 37.285 2.99 ;
      RECT 37.225 2.585 37.24 3.035 ;
      RECT 37.22 2.585 37.225 3.048 ;
      RECT 37.21 2.585 37.22 3.06 ;
      RECT 37.205 2.586 37.21 3.075 ;
      RECT 37.185 2.594 37.205 3.08 ;
      RECT 37.155 2.61 37.185 3.08 ;
      RECT 37.145 2.622 37.15 3.08 ;
      RECT 37.11 2.637 37.145 3.08 ;
      RECT 37.08 2.657 37.11 3.08 ;
      RECT 37.07 2.682 37.08 3.08 ;
      RECT 37.065 2.71 37.07 3.08 ;
      RECT 37.06 2.74 37.065 3.08 ;
      RECT 37.055 2.757 37.06 3.08 ;
      RECT 37.045 2.785 37.055 3.08 ;
      RECT 37.035 2.82 37.045 3.08 ;
      RECT 37.03 2.855 37.035 3.08 ;
      RECT 37.15 2.62 37.155 3.08 ;
      RECT 36.665 2.722 36.85 2.895 ;
      RECT 36.625 2.64 36.81 2.893 ;
      RECT 36.586 2.645 36.81 2.889 ;
      RECT 36.5 2.654 36.81 2.884 ;
      RECT 36.416 2.67 36.815 2.879 ;
      RECT 36.33 2.69 36.84 2.873 ;
      RECT 36.33 2.71 36.845 2.873 ;
      RECT 36.416 2.68 36.84 2.879 ;
      RECT 36.5 2.655 36.815 2.884 ;
      RECT 36.665 2.637 36.81 2.895 ;
      RECT 36.665 2.632 36.765 2.895 ;
      RECT 36.751 2.626 36.765 2.895 ;
      RECT 36.14 1.95 36.145 2.349 ;
      RECT 35.885 1.95 35.92 2.347 ;
      RECT 35.48 1.985 35.485 2.341 ;
      RECT 36.225 1.988 36.23 2.243 ;
      RECT 36.22 1.986 36.225 2.249 ;
      RECT 36.215 1.985 36.22 2.256 ;
      RECT 36.19 1.978 36.215 2.28 ;
      RECT 36.185 1.971 36.19 2.304 ;
      RECT 36.18 1.967 36.185 2.313 ;
      RECT 36.17 1.962 36.18 2.326 ;
      RECT 36.165 1.959 36.17 2.335 ;
      RECT 36.16 1.957 36.165 2.34 ;
      RECT 36.145 1.953 36.16 2.35 ;
      RECT 36.13 1.947 36.14 2.349 ;
      RECT 36.092 1.945 36.13 2.349 ;
      RECT 36.006 1.947 36.092 2.349 ;
      RECT 35.92 1.949 36.006 2.348 ;
      RECT 35.849 1.95 35.885 2.347 ;
      RECT 35.763 1.952 35.849 2.347 ;
      RECT 35.677 1.954 35.763 2.346 ;
      RECT 35.591 1.956 35.677 2.346 ;
      RECT 35.505 1.959 35.591 2.345 ;
      RECT 35.495 1.965 35.505 2.344 ;
      RECT 35.485 1.977 35.495 2.342 ;
      RECT 35.425 2.012 35.48 2.338 ;
      RECT 35.42 2.042 35.425 2.1 ;
      RECT 36.165 3.122 36.18 3.315 ;
      RECT 36.16 3.09 36.165 3.315 ;
      RECT 36.15 3.065 36.16 3.315 ;
      RECT 36.145 3.037 36.15 3.315 ;
      RECT 36.115 2.96 36.145 3.315 ;
      RECT 36.09 2.842 36.115 3.315 ;
      RECT 36.085 2.78 36.09 3.315 ;
      RECT 36.075 2.767 36.085 3.315 ;
      RECT 36.055 2.757 36.075 3.315 ;
      RECT 36.04 2.74 36.055 3.315 ;
      RECT 36.01 2.728 36.04 3.315 ;
      RECT 36.005 2.727 36.01 3.26 ;
      RECT 36 2.727 36.005 3.218 ;
      RECT 35.985 2.726 36 3.17 ;
      RECT 35.97 2.726 35.985 3.108 ;
      RECT 35.95 2.726 35.97 3.068 ;
      RECT 35.945 2.726 35.95 3.053 ;
      RECT 35.92 2.725 35.945 3.048 ;
      RECT 35.85 2.724 35.92 3.035 ;
      RECT 35.835 2.723 35.85 3.02 ;
      RECT 35.805 2.722 35.835 3.003 ;
      RECT 35.8 2.722 35.805 2.988 ;
      RECT 35.75 2.721 35.8 2.968 ;
      RECT 35.685 2.72 35.75 2.923 ;
      RECT 35.68 2.72 35.685 2.895 ;
      RECT 35.765 3.257 35.77 3.514 ;
      RECT 35.745 3.176 35.765 3.531 ;
      RECT 35.725 3.17 35.745 3.56 ;
      RECT 35.665 3.157 35.725 3.58 ;
      RECT 35.62 3.141 35.665 3.581 ;
      RECT 35.536 3.129 35.62 3.569 ;
      RECT 35.45 3.116 35.536 3.553 ;
      RECT 35.44 3.109 35.45 3.545 ;
      RECT 35.395 3.106 35.44 3.485 ;
      RECT 35.375 3.102 35.395 3.4 ;
      RECT 35.36 3.1 35.375 3.353 ;
      RECT 35.33 3.097 35.36 3.323 ;
      RECT 35.295 3.093 35.33 3.3 ;
      RECT 35.252 3.088 35.295 3.288 ;
      RECT 35.166 3.079 35.252 3.297 ;
      RECT 35.08 3.068 35.166 3.309 ;
      RECT 35.015 3.059 35.08 3.318 ;
      RECT 34.995 3.05 35.015 3.323 ;
      RECT 34.99 3.043 34.995 3.325 ;
      RECT 34.95 3.028 34.99 3.322 ;
      RECT 34.93 3.007 34.95 3.317 ;
      RECT 34.915 2.995 34.93 3.31 ;
      RECT 34.91 2.987 34.915 3.303 ;
      RECT 34.895 2.967 34.91 3.296 ;
      RECT 34.89 2.83 34.895 3.29 ;
      RECT 34.81 2.719 34.89 3.262 ;
      RECT 34.801 2.712 34.81 3.228 ;
      RECT 34.715 2.706 34.801 3.153 ;
      RECT 34.69 2.697 34.715 3.065 ;
      RECT 34.66 2.692 34.69 3.04 ;
      RECT 34.595 2.701 34.66 3.025 ;
      RECT 34.575 2.717 34.595 3 ;
      RECT 34.565 2.723 34.575 2.948 ;
      RECT 34.545 2.745 34.565 2.83 ;
      RECT 35.2 2.71 35.37 2.895 ;
      RECT 35.2 2.71 35.405 2.893 ;
      RECT 35.25 2.62 35.42 2.884 ;
      RECT 35.2 2.777 35.425 2.877 ;
      RECT 35.215 2.655 35.42 2.884 ;
      RECT 34.415 3.388 34.48 3.831 ;
      RECT 34.355 3.413 34.48 3.829 ;
      RECT 34.355 3.413 34.535 3.823 ;
      RECT 34.34 3.438 34.535 3.822 ;
      RECT 34.48 3.375 34.555 3.819 ;
      RECT 34.415 3.4 34.635 3.813 ;
      RECT 34.34 3.439 34.68 3.807 ;
      RECT 34.325 3.466 34.68 3.798 ;
      RECT 34.34 3.459 34.7 3.79 ;
      RECT 34.325 3.468 34.705 3.773 ;
      RECT 34.32 3.485 34.705 3.6 ;
      RECT 34.325 2.207 34.36 2.445 ;
      RECT 34.325 2.207 34.39 2.444 ;
      RECT 34.325 2.207 34.505 2.44 ;
      RECT 34.325 2.207 34.56 2.418 ;
      RECT 34.335 2.15 34.615 2.318 ;
      RECT 34.44 1.99 34.47 2.441 ;
      RECT 34.47 1.985 34.65 2.198 ;
      RECT 34.34 2.126 34.65 2.198 ;
      RECT 34.39 2.022 34.44 2.442 ;
      RECT 34.36 2.078 34.65 2.198 ;
      RECT 32.865 1.74 33.035 2.935 ;
      RECT 32.865 1.74 33.33 1.91 ;
      RECT 32.865 6.97 33.33 7.14 ;
      RECT 32.865 5.945 33.035 7.14 ;
      RECT 31.875 1.74 32.045 2.935 ;
      RECT 31.875 1.74 32.34 1.91 ;
      RECT 31.875 6.97 32.34 7.14 ;
      RECT 31.875 5.945 32.045 7.14 ;
      RECT 30.02 2.635 30.19 3.865 ;
      RECT 30.075 0.855 30.245 2.805 ;
      RECT 30.02 0.575 30.19 1.025 ;
      RECT 30.02 7.855 30.19 8.305 ;
      RECT 30.075 6.075 30.245 8.025 ;
      RECT 30.02 5.015 30.19 6.245 ;
      RECT 29.5 0.575 29.67 3.865 ;
      RECT 29.5 2.075 29.905 2.405 ;
      RECT 29.5 1.235 29.905 1.565 ;
      RECT 29.5 5.015 29.67 8.305 ;
      RECT 29.5 7.315 29.905 7.645 ;
      RECT 29.5 6.475 29.905 6.805 ;
      RECT 27.6 3.392 27.615 3.443 ;
      RECT 27.595 3.372 27.6 3.49 ;
      RECT 27.58 3.362 27.595 3.558 ;
      RECT 27.555 3.342 27.58 3.613 ;
      RECT 27.515 3.327 27.555 3.633 ;
      RECT 27.47 3.321 27.515 3.661 ;
      RECT 27.4 3.311 27.47 3.678 ;
      RECT 27.38 3.303 27.4 3.678 ;
      RECT 27.32 3.297 27.38 3.67 ;
      RECT 27.261 3.288 27.32 3.658 ;
      RECT 27.175 3.277 27.261 3.641 ;
      RECT 27.153 3.268 27.175 3.629 ;
      RECT 27.067 3.261 27.153 3.616 ;
      RECT 26.981 3.248 27.067 3.597 ;
      RECT 26.895 3.236 26.981 3.577 ;
      RECT 26.865 3.225 26.895 3.564 ;
      RECT 26.815 3.211 26.865 3.556 ;
      RECT 26.795 3.2 26.815 3.548 ;
      RECT 26.746 3.189 26.795 3.54 ;
      RECT 26.66 3.168 26.746 3.525 ;
      RECT 26.615 3.155 26.66 3.51 ;
      RECT 26.57 3.155 26.615 3.49 ;
      RECT 26.515 3.155 26.57 3.425 ;
      RECT 26.49 3.155 26.515 3.348 ;
      RECT 27.015 2.892 27.185 3.075 ;
      RECT 27.015 2.892 27.2 3.033 ;
      RECT 27.015 2.892 27.205 2.975 ;
      RECT 27.075 2.66 27.21 2.951 ;
      RECT 27.075 2.664 27.215 2.934 ;
      RECT 27.02 2.827 27.215 2.934 ;
      RECT 27.045 2.672 27.185 3.075 ;
      RECT 27.045 2.676 27.225 2.875 ;
      RECT 27.03 2.762 27.225 2.875 ;
      RECT 27.04 2.692 27.185 3.075 ;
      RECT 27.04 2.695 27.235 2.788 ;
      RECT 27.035 2.712 27.235 2.788 ;
      RECT 26.805 1.932 26.975 2.415 ;
      RECT 26.8 1.927 26.95 2.405 ;
      RECT 26.8 1.934 26.98 2.399 ;
      RECT 26.79 1.928 26.95 2.378 ;
      RECT 26.79 1.944 26.995 2.337 ;
      RECT 26.76 1.929 26.95 2.3 ;
      RECT 26.76 1.959 27.005 2.24 ;
      RECT 26.755 1.931 26.95 2.238 ;
      RECT 26.735 1.94 26.98 2.195 ;
      RECT 26.71 1.956 26.995 2.107 ;
      RECT 26.71 1.975 27.02 2.098 ;
      RECT 26.705 2.012 27.02 2.05 ;
      RECT 26.71 1.992 27.025 2.018 ;
      RECT 26.805 1.926 26.915 2.415 ;
      RECT 26.891 1.925 26.915 2.415 ;
      RECT 26.125 2.71 26.13 2.921 ;
      RECT 26.725 2.71 26.73 2.895 ;
      RECT 26.79 2.75 26.795 2.863 ;
      RECT 26.785 2.742 26.79 2.869 ;
      RECT 26.78 2.732 26.785 2.877 ;
      RECT 26.775 2.722 26.78 2.886 ;
      RECT 26.77 2.712 26.775 2.89 ;
      RECT 26.73 2.71 26.77 2.893 ;
      RECT 26.702 2.709 26.725 2.897 ;
      RECT 26.616 2.706 26.702 2.904 ;
      RECT 26.53 2.702 26.616 2.915 ;
      RECT 26.51 2.7 26.53 2.921 ;
      RECT 26.492 2.699 26.51 2.924 ;
      RECT 26.406 2.697 26.492 2.931 ;
      RECT 26.32 2.692 26.406 2.944 ;
      RECT 26.301 2.689 26.32 2.949 ;
      RECT 26.215 2.687 26.301 2.94 ;
      RECT 26.205 2.687 26.215 2.933 ;
      RECT 26.13 2.7 26.205 2.927 ;
      RECT 26.115 2.711 26.125 2.921 ;
      RECT 26.105 2.713 26.115 2.92 ;
      RECT 26.095 2.717 26.105 2.916 ;
      RECT 26.09 2.72 26.095 2.91 ;
      RECT 26.08 2.722 26.09 2.904 ;
      RECT 26.075 2.725 26.08 2.898 ;
      RECT 26.055 3.311 26.06 3.515 ;
      RECT 26.04 3.298 26.055 3.608 ;
      RECT 26.025 3.279 26.04 3.885 ;
      RECT 25.99 3.245 26.025 3.885 ;
      RECT 25.986 3.215 25.99 3.885 ;
      RECT 25.9 3.097 25.986 3.885 ;
      RECT 25.89 2.972 25.9 3.885 ;
      RECT 25.875 2.94 25.89 3.885 ;
      RECT 25.87 2.915 25.875 3.885 ;
      RECT 25.865 2.905 25.87 3.841 ;
      RECT 25.85 2.877 25.865 3.746 ;
      RECT 25.835 2.843 25.85 3.645 ;
      RECT 25.83 2.821 25.835 3.598 ;
      RECT 25.825 2.81 25.83 3.568 ;
      RECT 25.82 2.8 25.825 3.534 ;
      RECT 25.81 2.787 25.82 3.502 ;
      RECT 25.785 2.763 25.81 3.428 ;
      RECT 25.78 2.743 25.785 3.353 ;
      RECT 25.775 2.737 25.78 3.328 ;
      RECT 25.77 2.732 25.775 3.293 ;
      RECT 25.765 2.727 25.77 3.268 ;
      RECT 25.76 2.725 25.765 3.248 ;
      RECT 25.755 2.725 25.76 3.233 ;
      RECT 25.75 2.725 25.755 3.193 ;
      RECT 25.74 2.725 25.75 3.165 ;
      RECT 25.73 2.725 25.74 3.11 ;
      RECT 25.715 2.725 25.73 3.048 ;
      RECT 25.71 2.724 25.715 2.993 ;
      RECT 25.695 2.723 25.71 2.973 ;
      RECT 25.635 2.721 25.695 2.947 ;
      RECT 25.6 2.722 25.635 2.927 ;
      RECT 25.595 2.724 25.6 2.917 ;
      RECT 25.585 2.743 25.595 2.907 ;
      RECT 25.58 2.77 25.585 2.838 ;
      RECT 25.695 2.195 25.865 2.44 ;
      RECT 25.73 1.966 25.865 2.44 ;
      RECT 25.73 1.968 25.875 2.435 ;
      RECT 25.73 1.97 25.9 2.423 ;
      RECT 25.73 1.973 25.925 2.405 ;
      RECT 25.73 1.978 25.975 2.378 ;
      RECT 25.73 1.983 25.995 2.343 ;
      RECT 25.71 1.985 26.005 2.318 ;
      RECT 25.7 2.08 26.005 2.318 ;
      RECT 25.73 1.965 25.84 2.44 ;
      RECT 25.74 1.962 25.835 2.44 ;
      RECT 25.26 3.227 25.45 3.585 ;
      RECT 25.26 3.239 25.485 3.584 ;
      RECT 25.26 3.267 25.505 3.582 ;
      RECT 25.26 3.292 25.51 3.581 ;
      RECT 25.26 3.35 25.525 3.58 ;
      RECT 25.245 3.223 25.405 3.565 ;
      RECT 25.225 3.232 25.45 3.518 ;
      RECT 25.2 3.243 25.485 3.455 ;
      RECT 25.2 3.327 25.52 3.455 ;
      RECT 25.2 3.302 25.515 3.455 ;
      RECT 25.26 3.218 25.405 3.585 ;
      RECT 25.346 3.217 25.405 3.585 ;
      RECT 25.346 3.216 25.39 3.585 ;
      RECT 25.26 7.855 25.43 8.305 ;
      RECT 25.315 6.075 25.485 8.025 ;
      RECT 25.26 5.015 25.43 6.245 ;
      RECT 24.74 5.015 24.91 8.305 ;
      RECT 24.74 7.315 25.145 7.645 ;
      RECT 24.74 6.475 25.145 6.805 ;
      RECT 25.045 2.732 25.05 3.11 ;
      RECT 25.04 2.7 25.045 3.11 ;
      RECT 25.035 2.672 25.04 3.11 ;
      RECT 25.03 2.652 25.035 3.11 ;
      RECT 24.975 2.635 25.03 3.11 ;
      RECT 24.935 2.62 24.975 3.11 ;
      RECT 24.88 2.607 24.935 3.11 ;
      RECT 24.845 2.598 24.88 3.11 ;
      RECT 24.841 2.596 24.845 3.109 ;
      RECT 24.755 2.592 24.841 3.092 ;
      RECT 24.67 2.584 24.755 3.055 ;
      RECT 24.66 2.58 24.67 3.028 ;
      RECT 24.65 2.58 24.66 3.01 ;
      RECT 24.64 2.582 24.65 2.993 ;
      RECT 24.635 2.587 24.64 2.979 ;
      RECT 24.63 2.591 24.635 2.966 ;
      RECT 24.62 2.596 24.63 2.95 ;
      RECT 24.605 2.61 24.62 2.925 ;
      RECT 24.6 2.616 24.605 2.905 ;
      RECT 24.595 2.618 24.6 2.898 ;
      RECT 24.59 2.622 24.595 2.773 ;
      RECT 24.77 3.422 25.015 3.885 ;
      RECT 24.69 3.395 25.01 3.881 ;
      RECT 24.62 3.43 25.015 3.874 ;
      RECT 24.41 3.685 25.015 3.87 ;
      RECT 24.59 3.453 25.015 3.87 ;
      RECT 24.43 3.645 25.015 3.87 ;
      RECT 24.58 3.465 25.015 3.87 ;
      RECT 24.465 3.582 25.015 3.87 ;
      RECT 24.52 3.507 25.015 3.87 ;
      RECT 24.77 3.372 25.01 3.885 ;
      RECT 24.8 3.365 25.01 3.885 ;
      RECT 24.79 3.367 25.01 3.885 ;
      RECT 24.8 3.362 24.93 3.885 ;
      RECT 24.355 1.925 24.441 2.364 ;
      RECT 24.35 1.925 24.441 2.362 ;
      RECT 24.35 1.925 24.51 2.361 ;
      RECT 24.35 1.925 24.54 2.358 ;
      RECT 24.335 1.932 24.54 2.349 ;
      RECT 24.335 1.932 24.545 2.345 ;
      RECT 24.33 1.942 24.545 2.338 ;
      RECT 24.325 1.947 24.545 2.313 ;
      RECT 24.325 1.947 24.56 2.295 ;
      RECT 24.35 1.925 24.58 2.21 ;
      RECT 24.32 1.952 24.58 2.208 ;
      RECT 24.33 1.945 24.585 2.146 ;
      RECT 24.32 2.067 24.59 2.129 ;
      RECT 24.305 1.962 24.585 2.08 ;
      RECT 24.3 1.972 24.585 1.98 ;
      RECT 24.38 2.743 24.385 2.82 ;
      RECT 24.37 2.737 24.38 3.01 ;
      RECT 24.36 2.729 24.37 3.031 ;
      RECT 24.35 2.72 24.36 3.053 ;
      RECT 24.345 2.715 24.35 3.07 ;
      RECT 24.305 2.715 24.345 3.11 ;
      RECT 24.285 2.715 24.305 3.165 ;
      RECT 24.28 2.715 24.285 3.193 ;
      RECT 24.27 2.715 24.28 3.208 ;
      RECT 24.235 2.715 24.27 3.25 ;
      RECT 24.23 2.715 24.235 3.293 ;
      RECT 24.22 2.715 24.23 3.308 ;
      RECT 24.205 2.715 24.22 3.328 ;
      RECT 24.19 2.715 24.205 3.355 ;
      RECT 24.185 2.716 24.19 3.373 ;
      RECT 24.165 2.717 24.185 3.38 ;
      RECT 24.11 2.718 24.165 3.4 ;
      RECT 24.1 2.719 24.11 3.414 ;
      RECT 24.095 2.722 24.1 3.413 ;
      RECT 24.055 2.795 24.095 3.411 ;
      RECT 24.04 2.875 24.055 3.409 ;
      RECT 24.015 2.93 24.04 3.407 ;
      RECT 24 2.995 24.015 3.406 ;
      RECT 23.955 3.027 24 3.403 ;
      RECT 23.87 3.05 23.955 3.398 ;
      RECT 23.845 3.07 23.87 3.393 ;
      RECT 23.775 3.075 23.845 3.389 ;
      RECT 23.755 3.077 23.775 3.386 ;
      RECT 23.67 3.088 23.755 3.38 ;
      RECT 23.665 3.099 23.67 3.375 ;
      RECT 23.655 3.101 23.665 3.375 ;
      RECT 23.62 3.105 23.655 3.373 ;
      RECT 23.57 3.115 23.62 3.36 ;
      RECT 23.55 3.123 23.57 3.345 ;
      RECT 23.47 3.135 23.55 3.328 ;
      RECT 23.635 2.685 23.805 2.895 ;
      RECT 23.751 2.681 23.805 2.895 ;
      RECT 23.556 2.685 23.805 2.886 ;
      RECT 23.556 2.685 23.81 2.875 ;
      RECT 23.47 2.685 23.81 2.866 ;
      RECT 23.47 2.693 23.82 2.81 ;
      RECT 23.47 2.705 23.825 2.723 ;
      RECT 23.47 2.712 23.83 2.715 ;
      RECT 23.665 2.683 23.805 2.895 ;
      RECT 23.42 3.628 23.665 3.96 ;
      RECT 23.415 3.62 23.42 3.957 ;
      RECT 23.385 3.64 23.665 3.938 ;
      RECT 23.365 3.672 23.665 3.911 ;
      RECT 23.415 3.625 23.592 3.957 ;
      RECT 23.415 3.622 23.506 3.957 ;
      RECT 23.355 1.97 23.525 2.39 ;
      RECT 23.35 1.97 23.525 2.388 ;
      RECT 23.35 1.97 23.55 2.378 ;
      RECT 23.35 1.97 23.57 2.353 ;
      RECT 23.345 1.97 23.57 2.348 ;
      RECT 23.345 1.97 23.58 2.338 ;
      RECT 23.345 1.97 23.585 2.333 ;
      RECT 23.345 1.975 23.59 2.328 ;
      RECT 23.345 2.007 23.605 2.318 ;
      RECT 23.345 2.077 23.63 2.301 ;
      RECT 23.325 2.077 23.63 2.293 ;
      RECT 23.325 2.137 23.64 2.27 ;
      RECT 23.325 2.177 23.65 2.215 ;
      RECT 23.31 1.97 23.585 2.195 ;
      RECT 23.3 1.985 23.59 2.093 ;
      RECT 22.89 3.375 23.06 3.9 ;
      RECT 22.885 3.375 23.06 3.893 ;
      RECT 22.875 3.375 23.065 3.858 ;
      RECT 22.87 3.385 23.065 3.83 ;
      RECT 22.865 3.405 23.065 3.813 ;
      RECT 22.875 3.38 23.07 3.803 ;
      RECT 22.86 3.425 23.07 3.795 ;
      RECT 22.855 3.445 23.07 3.78 ;
      RECT 22.85 3.475 23.07 3.77 ;
      RECT 22.84 3.52 23.07 3.745 ;
      RECT 22.87 3.39 23.075 3.728 ;
      RECT 22.835 3.572 23.075 3.723 ;
      RECT 22.87 3.4 23.08 3.693 ;
      RECT 22.83 3.605 23.08 3.69 ;
      RECT 22.825 3.63 23.08 3.67 ;
      RECT 22.865 3.417 23.09 3.61 ;
      RECT 22.86 3.439 23.1 3.503 ;
      RECT 22.81 2.686 22.825 2.955 ;
      RECT 22.765 2.67 22.81 3 ;
      RECT 22.76 2.658 22.765 3.05 ;
      RECT 22.75 2.654 22.76 3.083 ;
      RECT 22.745 2.651 22.75 3.111 ;
      RECT 22.73 2.653 22.745 3.153 ;
      RECT 22.725 2.657 22.73 3.193 ;
      RECT 22.705 2.662 22.725 3.245 ;
      RECT 22.701 2.667 22.705 3.302 ;
      RECT 22.615 2.686 22.701 3.339 ;
      RECT 22.605 2.707 22.615 3.375 ;
      RECT 22.6 2.715 22.605 3.376 ;
      RECT 22.595 2.757 22.6 3.377 ;
      RECT 22.58 2.845 22.595 3.378 ;
      RECT 22.57 2.995 22.58 3.38 ;
      RECT 22.565 3.04 22.57 3.382 ;
      RECT 22.53 3.082 22.565 3.385 ;
      RECT 22.525 3.1 22.53 3.388 ;
      RECT 22.448 3.106 22.525 3.394 ;
      RECT 22.362 3.12 22.448 3.407 ;
      RECT 22.276 3.134 22.362 3.421 ;
      RECT 22.19 3.148 22.276 3.434 ;
      RECT 22.13 3.16 22.19 3.446 ;
      RECT 22.105 3.167 22.13 3.453 ;
      RECT 22.091 3.17 22.105 3.458 ;
      RECT 22.005 3.178 22.091 3.474 ;
      RECT 22 3.185 22.005 3.489 ;
      RECT 21.976 3.185 22 3.496 ;
      RECT 21.89 3.188 21.976 3.524 ;
      RECT 21.805 3.192 21.89 3.568 ;
      RECT 21.74 3.196 21.805 3.605 ;
      RECT 21.715 3.199 21.74 3.621 ;
      RECT 21.64 3.212 21.715 3.625 ;
      RECT 21.615 3.23 21.64 3.629 ;
      RECT 21.605 3.237 21.615 3.631 ;
      RECT 21.59 3.24 21.605 3.632 ;
      RECT 21.53 3.252 21.59 3.636 ;
      RECT 21.52 3.266 21.53 3.64 ;
      RECT 21.465 3.276 21.52 3.628 ;
      RECT 21.44 3.297 21.465 3.611 ;
      RECT 21.42 3.317 21.44 3.602 ;
      RECT 21.415 3.33 21.42 3.597 ;
      RECT 21.4 3.342 21.415 3.593 ;
      RECT 22.635 1.997 22.64 2.02 ;
      RECT 22.63 1.988 22.635 2.06 ;
      RECT 22.625 1.986 22.63 2.103 ;
      RECT 22.62 1.977 22.625 2.138 ;
      RECT 22.615 1.967 22.62 2.21 ;
      RECT 22.61 1.957 22.615 2.275 ;
      RECT 22.605 1.954 22.61 2.315 ;
      RECT 22.58 1.948 22.605 2.405 ;
      RECT 22.545 1.936 22.58 2.43 ;
      RECT 22.535 1.927 22.545 2.43 ;
      RECT 22.4 1.925 22.41 2.413 ;
      RECT 22.39 1.925 22.4 2.38 ;
      RECT 22.385 1.925 22.39 2.355 ;
      RECT 22.38 1.925 22.385 2.343 ;
      RECT 22.375 1.925 22.38 2.325 ;
      RECT 22.365 1.925 22.375 2.29 ;
      RECT 22.36 1.927 22.365 2.268 ;
      RECT 22.355 1.933 22.36 2.253 ;
      RECT 22.35 1.939 22.355 2.238 ;
      RECT 22.335 1.951 22.35 2.211 ;
      RECT 22.33 1.962 22.335 2.179 ;
      RECT 22.325 1.972 22.33 2.163 ;
      RECT 22.315 1.98 22.325 2.132 ;
      RECT 22.31 1.99 22.315 2.106 ;
      RECT 22.305 2.047 22.31 2.089 ;
      RECT 22.41 1.925 22.535 2.43 ;
      RECT 22.125 2.612 22.385 2.91 ;
      RECT 22.12 2.619 22.385 2.908 ;
      RECT 22.125 2.614 22.4 2.903 ;
      RECT 22.115 2.627 22.4 2.9 ;
      RECT 22.115 2.632 22.405 2.893 ;
      RECT 22.11 2.64 22.405 2.89 ;
      RECT 22.11 2.657 22.41 2.688 ;
      RECT 22.125 2.609 22.356 2.91 ;
      RECT 22.18 2.608 22.356 2.91 ;
      RECT 22.18 2.605 22.27 2.91 ;
      RECT 22.18 2.602 22.266 2.91 ;
      RECT 21.87 2.875 21.875 2.888 ;
      RECT 21.865 2.842 21.87 2.893 ;
      RECT 21.86 2.797 21.865 2.9 ;
      RECT 21.855 2.752 21.86 2.908 ;
      RECT 21.85 2.72 21.855 2.916 ;
      RECT 21.845 2.68 21.85 2.917 ;
      RECT 21.83 2.66 21.845 2.919 ;
      RECT 21.755 2.642 21.83 2.931 ;
      RECT 21.745 2.635 21.755 2.942 ;
      RECT 21.74 2.635 21.745 2.944 ;
      RECT 21.71 2.641 21.74 2.948 ;
      RECT 21.67 2.654 21.71 2.948 ;
      RECT 21.645 2.665 21.67 2.934 ;
      RECT 21.63 2.671 21.645 2.917 ;
      RECT 21.62 2.673 21.63 2.908 ;
      RECT 21.615 2.674 21.62 2.903 ;
      RECT 21.61 2.675 21.615 2.898 ;
      RECT 21.605 2.676 21.61 2.895 ;
      RECT 21.58 2.681 21.605 2.885 ;
      RECT 21.57 2.697 21.58 2.872 ;
      RECT 21.565 2.717 21.57 2.867 ;
      RECT 21.575 2.11 21.58 2.306 ;
      RECT 21.56 2.074 21.575 2.308 ;
      RECT 21.55 2.056 21.56 2.313 ;
      RECT 21.54 2.042 21.55 2.317 ;
      RECT 21.495 2.026 21.54 2.327 ;
      RECT 21.49 2.016 21.495 2.336 ;
      RECT 21.445 2.005 21.49 2.342 ;
      RECT 21.44 1.993 21.445 2.349 ;
      RECT 21.425 1.988 21.44 2.353 ;
      RECT 21.41 1.98 21.425 2.358 ;
      RECT 21.4 1.973 21.41 2.363 ;
      RECT 21.39 1.97 21.4 2.368 ;
      RECT 21.38 1.97 21.39 2.369 ;
      RECT 21.375 1.967 21.38 2.368 ;
      RECT 21.34 1.962 21.365 2.367 ;
      RECT 21.316 1.958 21.34 2.366 ;
      RECT 21.23 1.949 21.316 2.363 ;
      RECT 21.215 1.941 21.23 2.36 ;
      RECT 21.193 1.94 21.215 2.359 ;
      RECT 21.107 1.94 21.193 2.357 ;
      RECT 21.021 1.94 21.107 2.355 ;
      RECT 20.935 1.94 21.021 2.352 ;
      RECT 20.925 1.94 20.935 2.343 ;
      RECT 20.895 1.94 20.925 2.303 ;
      RECT 20.885 1.95 20.895 2.258 ;
      RECT 20.88 1.99 20.885 2.243 ;
      RECT 20.875 2.005 20.88 2.23 ;
      RECT 20.845 2.085 20.875 2.192 ;
      RECT 21.365 1.965 21.375 2.368 ;
      RECT 21.19 2.73 21.205 3.335 ;
      RECT 21.195 2.725 21.205 3.335 ;
      RECT 21.36 2.725 21.365 2.908 ;
      RECT 21.35 2.725 21.36 2.938 ;
      RECT 21.335 2.725 21.35 2.998 ;
      RECT 21.33 2.725 21.335 3.043 ;
      RECT 21.325 2.725 21.33 3.073 ;
      RECT 21.32 2.725 21.325 3.093 ;
      RECT 21.31 2.725 21.32 3.128 ;
      RECT 21.295 2.725 21.31 3.16 ;
      RECT 21.25 2.725 21.295 3.188 ;
      RECT 21.245 2.725 21.25 3.218 ;
      RECT 21.24 2.725 21.245 3.23 ;
      RECT 21.235 2.725 21.24 3.238 ;
      RECT 21.225 2.725 21.235 3.253 ;
      RECT 21.22 2.725 21.225 3.275 ;
      RECT 21.21 2.725 21.22 3.298 ;
      RECT 21.205 2.725 21.21 3.318 ;
      RECT 21.17 2.74 21.19 3.335 ;
      RECT 21.145 2.757 21.17 3.335 ;
      RECT 21.14 2.767 21.145 3.335 ;
      RECT 21.11 2.782 21.14 3.335 ;
      RECT 21.035 2.824 21.11 3.335 ;
      RECT 21.03 2.855 21.035 3.318 ;
      RECT 21.025 2.859 21.03 3.3 ;
      RECT 21.02 2.863 21.025 3.263 ;
      RECT 21.015 3.047 21.02 3.23 ;
      RECT 20.5 3.236 20.586 3.801 ;
      RECT 20.455 3.238 20.62 3.795 ;
      RECT 20.586 3.235 20.62 3.795 ;
      RECT 20.5 3.237 20.705 3.789 ;
      RECT 20.455 3.247 20.715 3.785 ;
      RECT 20.43 3.239 20.705 3.781 ;
      RECT 20.425 3.242 20.705 3.776 ;
      RECT 20.4 3.257 20.715 3.77 ;
      RECT 20.4 3.282 20.755 3.765 ;
      RECT 20.36 3.29 20.755 3.74 ;
      RECT 20.36 3.317 20.77 3.738 ;
      RECT 20.36 3.347 20.78 3.725 ;
      RECT 20.355 3.492 20.78 3.713 ;
      RECT 20.36 3.421 20.8 3.71 ;
      RECT 20.36 3.478 20.805 3.518 ;
      RECT 20.55 2.757 20.72 2.935 ;
      RECT 20.5 2.696 20.55 2.92 ;
      RECT 20.235 2.676 20.5 2.905 ;
      RECT 20.195 2.74 20.67 2.905 ;
      RECT 20.195 2.73 20.625 2.905 ;
      RECT 20.195 2.727 20.615 2.905 ;
      RECT 20.195 2.715 20.605 2.905 ;
      RECT 20.195 2.7 20.55 2.905 ;
      RECT 20.235 2.672 20.436 2.905 ;
      RECT 20.245 2.65 20.436 2.905 ;
      RECT 20.27 2.635 20.35 2.905 ;
      RECT 20.025 3.165 20.145 3.61 ;
      RECT 20.01 3.165 20.145 3.609 ;
      RECT 19.965 3.187 20.145 3.604 ;
      RECT 19.925 3.236 20.145 3.598 ;
      RECT 19.925 3.236 20.15 3.573 ;
      RECT 19.925 3.236 20.17 3.463 ;
      RECT 19.92 3.266 20.17 3.46 ;
      RECT 20.01 3.165 20.18 3.355 ;
      RECT 19.67 1.95 19.675 2.395 ;
      RECT 19.48 1.95 19.5 2.36 ;
      RECT 19.45 1.95 19.455 2.335 ;
      RECT 20.13 2.257 20.145 2.445 ;
      RECT 20.125 2.242 20.13 2.451 ;
      RECT 20.105 2.215 20.125 2.454 ;
      RECT 20.055 2.182 20.105 2.463 ;
      RECT 20.025 2.162 20.055 2.467 ;
      RECT 20.006 2.15 20.025 2.463 ;
      RECT 19.92 2.122 20.006 2.453 ;
      RECT 19.91 2.097 19.92 2.443 ;
      RECT 19.84 2.065 19.91 2.435 ;
      RECT 19.815 2.025 19.84 2.427 ;
      RECT 19.795 2.007 19.815 2.421 ;
      RECT 19.785 1.997 19.795 2.418 ;
      RECT 19.775 1.99 19.785 2.416 ;
      RECT 19.755 1.977 19.775 2.413 ;
      RECT 19.745 1.967 19.755 2.41 ;
      RECT 19.735 1.96 19.745 2.408 ;
      RECT 19.685 1.952 19.735 2.402 ;
      RECT 19.675 1.95 19.685 2.396 ;
      RECT 19.645 1.95 19.67 2.393 ;
      RECT 19.616 1.95 19.645 2.388 ;
      RECT 19.53 1.95 19.616 2.378 ;
      RECT 19.5 1.95 19.53 2.365 ;
      RECT 19.455 1.95 19.48 2.348 ;
      RECT 19.44 1.95 19.45 2.33 ;
      RECT 19.42 1.957 19.44 2.315 ;
      RECT 19.415 1.972 19.42 2.303 ;
      RECT 19.41 1.977 19.415 2.243 ;
      RECT 19.405 1.982 19.41 2.085 ;
      RECT 19.4 1.985 19.405 2.003 ;
      RECT 19.665 2.67 19.751 2.991 ;
      RECT 19.665 2.67 19.785 2.984 ;
      RECT 19.615 2.67 19.785 2.98 ;
      RECT 19.615 2.672 19.871 2.978 ;
      RECT 19.615 2.674 19.895 2.972 ;
      RECT 19.615 2.681 19.905 2.971 ;
      RECT 19.615 2.69 19.91 2.968 ;
      RECT 19.615 2.696 19.915 2.963 ;
      RECT 19.615 2.74 19.92 2.96 ;
      RECT 19.615 2.832 19.925 2.957 ;
      RECT 19.14 3.275 19.175 3.595 ;
      RECT 19.725 3.46 19.73 3.642 ;
      RECT 19.68 3.342 19.725 3.661 ;
      RECT 19.665 3.319 19.68 3.684 ;
      RECT 19.655 3.309 19.665 3.694 ;
      RECT 19.635 3.304 19.655 3.707 ;
      RECT 19.61 3.302 19.635 3.728 ;
      RECT 19.591 3.301 19.61 3.74 ;
      RECT 19.505 3.298 19.591 3.74 ;
      RECT 19.435 3.293 19.505 3.728 ;
      RECT 19.36 3.289 19.435 3.703 ;
      RECT 19.295 3.285 19.36 3.67 ;
      RECT 19.225 3.282 19.295 3.63 ;
      RECT 19.195 3.278 19.225 3.605 ;
      RECT 19.175 3.276 19.195 3.598 ;
      RECT 19.091 3.274 19.14 3.596 ;
      RECT 19.005 3.271 19.091 3.597 ;
      RECT 18.93 3.27 19.005 3.599 ;
      RECT 18.845 3.27 18.93 3.625 ;
      RECT 18.768 3.271 18.845 3.65 ;
      RECT 18.682 3.272 18.768 3.65 ;
      RECT 18.596 3.272 18.682 3.65 ;
      RECT 18.51 3.273 18.596 3.65 ;
      RECT 18.49 3.274 18.51 3.642 ;
      RECT 18.475 3.28 18.49 3.627 ;
      RECT 18.44 3.3 18.475 3.607 ;
      RECT 18.43 3.32 18.44 3.589 ;
      RECT 19.4 2.625 19.405 2.895 ;
      RECT 19.395 2.616 19.4 2.9 ;
      RECT 19.385 2.606 19.395 2.912 ;
      RECT 19.38 2.595 19.385 2.923 ;
      RECT 19.36 2.589 19.38 2.941 ;
      RECT 19.315 2.586 19.36 2.99 ;
      RECT 19.3 2.585 19.315 3.035 ;
      RECT 19.295 2.585 19.3 3.048 ;
      RECT 19.285 2.585 19.295 3.06 ;
      RECT 19.28 2.586 19.285 3.075 ;
      RECT 19.26 2.594 19.28 3.08 ;
      RECT 19.23 2.61 19.26 3.08 ;
      RECT 19.22 2.622 19.225 3.08 ;
      RECT 19.185 2.637 19.22 3.08 ;
      RECT 19.155 2.657 19.185 3.08 ;
      RECT 19.145 2.682 19.155 3.08 ;
      RECT 19.14 2.71 19.145 3.08 ;
      RECT 19.135 2.74 19.14 3.08 ;
      RECT 19.13 2.757 19.135 3.08 ;
      RECT 19.12 2.785 19.13 3.08 ;
      RECT 19.11 2.82 19.12 3.08 ;
      RECT 19.105 2.855 19.11 3.08 ;
      RECT 19.225 2.62 19.23 3.08 ;
      RECT 18.74 2.722 18.925 2.895 ;
      RECT 18.7 2.64 18.885 2.893 ;
      RECT 18.661 2.645 18.885 2.889 ;
      RECT 18.575 2.654 18.885 2.884 ;
      RECT 18.491 2.67 18.89 2.879 ;
      RECT 18.405 2.69 18.915 2.873 ;
      RECT 18.405 2.71 18.92 2.873 ;
      RECT 18.491 2.68 18.915 2.879 ;
      RECT 18.575 2.655 18.89 2.884 ;
      RECT 18.74 2.637 18.885 2.895 ;
      RECT 18.74 2.632 18.84 2.895 ;
      RECT 18.826 2.626 18.84 2.895 ;
      RECT 18.215 1.95 18.22 2.349 ;
      RECT 17.96 1.95 17.995 2.347 ;
      RECT 17.555 1.985 17.56 2.341 ;
      RECT 18.3 1.988 18.305 2.243 ;
      RECT 18.295 1.986 18.3 2.249 ;
      RECT 18.29 1.985 18.295 2.256 ;
      RECT 18.265 1.978 18.29 2.28 ;
      RECT 18.26 1.971 18.265 2.304 ;
      RECT 18.255 1.967 18.26 2.313 ;
      RECT 18.245 1.962 18.255 2.326 ;
      RECT 18.24 1.959 18.245 2.335 ;
      RECT 18.235 1.957 18.24 2.34 ;
      RECT 18.22 1.953 18.235 2.35 ;
      RECT 18.205 1.947 18.215 2.349 ;
      RECT 18.167 1.945 18.205 2.349 ;
      RECT 18.081 1.947 18.167 2.349 ;
      RECT 17.995 1.949 18.081 2.348 ;
      RECT 17.924 1.95 17.96 2.347 ;
      RECT 17.838 1.952 17.924 2.347 ;
      RECT 17.752 1.954 17.838 2.346 ;
      RECT 17.666 1.956 17.752 2.346 ;
      RECT 17.58 1.959 17.666 2.345 ;
      RECT 17.57 1.965 17.58 2.344 ;
      RECT 17.56 1.977 17.57 2.342 ;
      RECT 17.5 2.012 17.555 2.338 ;
      RECT 17.495 2.042 17.5 2.1 ;
      RECT 18.24 3.122 18.255 3.315 ;
      RECT 18.235 3.09 18.24 3.315 ;
      RECT 18.225 3.065 18.235 3.315 ;
      RECT 18.22 3.037 18.225 3.315 ;
      RECT 18.19 2.96 18.22 3.315 ;
      RECT 18.165 2.842 18.19 3.315 ;
      RECT 18.16 2.78 18.165 3.315 ;
      RECT 18.15 2.767 18.16 3.315 ;
      RECT 18.13 2.757 18.15 3.315 ;
      RECT 18.115 2.74 18.13 3.315 ;
      RECT 18.085 2.728 18.115 3.315 ;
      RECT 18.08 2.727 18.085 3.26 ;
      RECT 18.075 2.727 18.08 3.218 ;
      RECT 18.06 2.726 18.075 3.17 ;
      RECT 18.045 2.726 18.06 3.108 ;
      RECT 18.025 2.726 18.045 3.068 ;
      RECT 18.02 2.726 18.025 3.053 ;
      RECT 17.995 2.725 18.02 3.048 ;
      RECT 17.925 2.724 17.995 3.035 ;
      RECT 17.91 2.723 17.925 3.02 ;
      RECT 17.88 2.722 17.91 3.003 ;
      RECT 17.875 2.722 17.88 2.988 ;
      RECT 17.825 2.721 17.875 2.968 ;
      RECT 17.76 2.72 17.825 2.923 ;
      RECT 17.755 2.72 17.76 2.895 ;
      RECT 17.84 3.257 17.845 3.514 ;
      RECT 17.82 3.176 17.84 3.531 ;
      RECT 17.8 3.17 17.82 3.56 ;
      RECT 17.74 3.157 17.8 3.58 ;
      RECT 17.695 3.141 17.74 3.581 ;
      RECT 17.611 3.129 17.695 3.569 ;
      RECT 17.525 3.116 17.611 3.553 ;
      RECT 17.515 3.109 17.525 3.545 ;
      RECT 17.47 3.106 17.515 3.485 ;
      RECT 17.45 3.102 17.47 3.4 ;
      RECT 17.435 3.1 17.45 3.353 ;
      RECT 17.405 3.097 17.435 3.323 ;
      RECT 17.37 3.093 17.405 3.3 ;
      RECT 17.327 3.088 17.37 3.288 ;
      RECT 17.241 3.079 17.327 3.297 ;
      RECT 17.155 3.068 17.241 3.309 ;
      RECT 17.09 3.059 17.155 3.318 ;
      RECT 17.07 3.05 17.09 3.323 ;
      RECT 17.065 3.043 17.07 3.325 ;
      RECT 17.025 3.028 17.065 3.322 ;
      RECT 17.005 3.007 17.025 3.317 ;
      RECT 16.99 2.995 17.005 3.31 ;
      RECT 16.985 2.987 16.99 3.303 ;
      RECT 16.97 2.967 16.985 3.296 ;
      RECT 16.965 2.83 16.97 3.29 ;
      RECT 16.885 2.719 16.965 3.262 ;
      RECT 16.876 2.712 16.885 3.228 ;
      RECT 16.79 2.706 16.876 3.153 ;
      RECT 16.765 2.697 16.79 3.065 ;
      RECT 16.735 2.692 16.765 3.04 ;
      RECT 16.67 2.701 16.735 3.025 ;
      RECT 16.65 2.717 16.67 3 ;
      RECT 16.64 2.723 16.65 2.948 ;
      RECT 16.62 2.745 16.64 2.83 ;
      RECT 17.275 2.71 17.445 2.895 ;
      RECT 17.275 2.71 17.48 2.893 ;
      RECT 17.325 2.62 17.495 2.884 ;
      RECT 17.275 2.777 17.5 2.877 ;
      RECT 17.29 2.655 17.495 2.884 ;
      RECT 16.49 3.388 16.555 3.831 ;
      RECT 16.43 3.413 16.555 3.829 ;
      RECT 16.43 3.413 16.61 3.823 ;
      RECT 16.415 3.438 16.61 3.822 ;
      RECT 16.555 3.375 16.63 3.819 ;
      RECT 16.49 3.4 16.71 3.813 ;
      RECT 16.415 3.439 16.755 3.807 ;
      RECT 16.4 3.466 16.755 3.798 ;
      RECT 16.415 3.459 16.775 3.79 ;
      RECT 16.4 3.468 16.78 3.773 ;
      RECT 16.395 3.485 16.78 3.6 ;
      RECT 16.4 2.207 16.435 2.445 ;
      RECT 16.4 2.207 16.465 2.444 ;
      RECT 16.4 2.207 16.58 2.44 ;
      RECT 16.4 2.207 16.635 2.418 ;
      RECT 16.41 2.15 16.69 2.318 ;
      RECT 16.515 1.99 16.545 2.441 ;
      RECT 16.545 1.985 16.725 2.198 ;
      RECT 16.415 2.126 16.725 2.198 ;
      RECT 16.465 2.022 16.515 2.442 ;
      RECT 16.435 2.078 16.725 2.198 ;
      RECT 14.94 1.74 15.11 2.935 ;
      RECT 14.94 1.74 15.405 1.91 ;
      RECT 14.94 6.97 15.405 7.14 ;
      RECT 14.94 5.945 15.11 7.14 ;
      RECT 13.95 1.74 14.12 2.935 ;
      RECT 13.95 1.74 14.415 1.91 ;
      RECT 13.95 6.97 14.415 7.14 ;
      RECT 13.95 5.945 14.12 7.14 ;
      RECT 12.095 2.635 12.265 3.865 ;
      RECT 12.15 0.855 12.32 2.805 ;
      RECT 12.095 0.575 12.265 1.025 ;
      RECT 12.095 7.855 12.265 8.305 ;
      RECT 12.15 6.075 12.32 8.025 ;
      RECT 12.095 5.015 12.265 6.245 ;
      RECT 11.575 0.575 11.745 3.865 ;
      RECT 11.575 2.075 11.98 2.405 ;
      RECT 11.575 1.235 11.98 1.565 ;
      RECT 11.575 5.015 11.745 8.305 ;
      RECT 11.575 7.315 11.98 7.645 ;
      RECT 11.575 6.475 11.98 6.805 ;
      RECT 9.675 3.392 9.69 3.443 ;
      RECT 9.67 3.372 9.675 3.49 ;
      RECT 9.655 3.362 9.67 3.558 ;
      RECT 9.63 3.342 9.655 3.613 ;
      RECT 9.59 3.327 9.63 3.633 ;
      RECT 9.545 3.321 9.59 3.661 ;
      RECT 9.475 3.311 9.545 3.678 ;
      RECT 9.455 3.303 9.475 3.678 ;
      RECT 9.395 3.297 9.455 3.67 ;
      RECT 9.336 3.288 9.395 3.658 ;
      RECT 9.25 3.277 9.336 3.641 ;
      RECT 9.228 3.268 9.25 3.629 ;
      RECT 9.142 3.261 9.228 3.616 ;
      RECT 9.056 3.248 9.142 3.597 ;
      RECT 8.97 3.236 9.056 3.577 ;
      RECT 8.94 3.225 8.97 3.564 ;
      RECT 8.89 3.211 8.94 3.556 ;
      RECT 8.87 3.2 8.89 3.548 ;
      RECT 8.821 3.189 8.87 3.54 ;
      RECT 8.735 3.168 8.821 3.525 ;
      RECT 8.69 3.155 8.735 3.51 ;
      RECT 8.645 3.155 8.69 3.49 ;
      RECT 8.59 3.155 8.645 3.425 ;
      RECT 8.565 3.155 8.59 3.348 ;
      RECT 9.09 2.892 9.26 3.075 ;
      RECT 9.09 2.892 9.275 3.033 ;
      RECT 9.09 2.892 9.28 2.975 ;
      RECT 9.15 2.66 9.285 2.951 ;
      RECT 9.15 2.664 9.29 2.934 ;
      RECT 9.095 2.827 9.29 2.934 ;
      RECT 9.12 2.672 9.26 3.075 ;
      RECT 9.12 2.676 9.3 2.875 ;
      RECT 9.105 2.762 9.3 2.875 ;
      RECT 9.115 2.692 9.26 3.075 ;
      RECT 9.115 2.695 9.31 2.788 ;
      RECT 9.11 2.712 9.31 2.788 ;
      RECT 8.88 1.932 9.05 2.415 ;
      RECT 8.875 1.927 9.025 2.405 ;
      RECT 8.875 1.934 9.055 2.399 ;
      RECT 8.865 1.928 9.025 2.378 ;
      RECT 8.865 1.944 9.07 2.337 ;
      RECT 8.835 1.929 9.025 2.3 ;
      RECT 8.835 1.959 9.08 2.24 ;
      RECT 8.83 1.931 9.025 2.238 ;
      RECT 8.81 1.94 9.055 2.195 ;
      RECT 8.785 1.956 9.07 2.107 ;
      RECT 8.785 1.975 9.095 2.098 ;
      RECT 8.78 2.012 9.095 2.05 ;
      RECT 8.785 1.992 9.1 2.018 ;
      RECT 8.88 1.926 8.99 2.415 ;
      RECT 8.966 1.925 8.99 2.415 ;
      RECT 8.2 2.71 8.205 2.921 ;
      RECT 8.8 2.71 8.805 2.895 ;
      RECT 8.865 2.75 8.87 2.863 ;
      RECT 8.86 2.742 8.865 2.869 ;
      RECT 8.855 2.732 8.86 2.877 ;
      RECT 8.85 2.722 8.855 2.886 ;
      RECT 8.845 2.712 8.85 2.89 ;
      RECT 8.805 2.71 8.845 2.893 ;
      RECT 8.777 2.709 8.8 2.897 ;
      RECT 8.691 2.706 8.777 2.904 ;
      RECT 8.605 2.702 8.691 2.915 ;
      RECT 8.585 2.7 8.605 2.921 ;
      RECT 8.567 2.699 8.585 2.924 ;
      RECT 8.481 2.697 8.567 2.931 ;
      RECT 8.395 2.692 8.481 2.944 ;
      RECT 8.376 2.689 8.395 2.949 ;
      RECT 8.29 2.687 8.376 2.94 ;
      RECT 8.28 2.687 8.29 2.933 ;
      RECT 8.205 2.7 8.28 2.927 ;
      RECT 8.19 2.711 8.2 2.921 ;
      RECT 8.18 2.713 8.19 2.92 ;
      RECT 8.17 2.717 8.18 2.916 ;
      RECT 8.165 2.72 8.17 2.91 ;
      RECT 8.155 2.722 8.165 2.904 ;
      RECT 8.15 2.725 8.155 2.898 ;
      RECT 8.13 3.311 8.135 3.515 ;
      RECT 8.115 3.298 8.13 3.608 ;
      RECT 8.1 3.279 8.115 3.885 ;
      RECT 8.065 3.245 8.1 3.885 ;
      RECT 8.061 3.215 8.065 3.885 ;
      RECT 7.975 3.097 8.061 3.885 ;
      RECT 7.965 2.972 7.975 3.885 ;
      RECT 7.95 2.94 7.965 3.885 ;
      RECT 7.945 2.915 7.95 3.885 ;
      RECT 7.94 2.905 7.945 3.841 ;
      RECT 7.925 2.877 7.94 3.746 ;
      RECT 7.91 2.843 7.925 3.645 ;
      RECT 7.905 2.821 7.91 3.598 ;
      RECT 7.9 2.81 7.905 3.568 ;
      RECT 7.895 2.8 7.9 3.534 ;
      RECT 7.885 2.787 7.895 3.502 ;
      RECT 7.86 2.763 7.885 3.428 ;
      RECT 7.855 2.743 7.86 3.353 ;
      RECT 7.85 2.737 7.855 3.328 ;
      RECT 7.845 2.732 7.85 3.293 ;
      RECT 7.84 2.727 7.845 3.268 ;
      RECT 7.835 2.725 7.84 3.248 ;
      RECT 7.83 2.725 7.835 3.233 ;
      RECT 7.825 2.725 7.83 3.193 ;
      RECT 7.815 2.725 7.825 3.165 ;
      RECT 7.805 2.725 7.815 3.11 ;
      RECT 7.79 2.725 7.805 3.048 ;
      RECT 7.785 2.724 7.79 2.993 ;
      RECT 7.77 2.723 7.785 2.973 ;
      RECT 7.71 2.721 7.77 2.947 ;
      RECT 7.675 2.722 7.71 2.927 ;
      RECT 7.67 2.724 7.675 2.917 ;
      RECT 7.66 2.743 7.67 2.907 ;
      RECT 7.655 2.77 7.66 2.838 ;
      RECT 7.77 2.195 7.94 2.44 ;
      RECT 7.805 1.966 7.94 2.44 ;
      RECT 7.805 1.968 7.95 2.435 ;
      RECT 7.805 1.97 7.975 2.423 ;
      RECT 7.805 1.973 8 2.405 ;
      RECT 7.805 1.978 8.05 2.378 ;
      RECT 7.805 1.983 8.07 2.343 ;
      RECT 7.785 1.985 8.08 2.318 ;
      RECT 7.775 2.08 8.08 2.318 ;
      RECT 7.805 1.965 7.915 2.44 ;
      RECT 7.815 1.962 7.91 2.44 ;
      RECT 7.335 3.227 7.525 3.585 ;
      RECT 7.335 3.239 7.56 3.584 ;
      RECT 7.335 3.267 7.58 3.582 ;
      RECT 7.335 3.292 7.585 3.581 ;
      RECT 7.335 3.35 7.6 3.58 ;
      RECT 7.32 3.223 7.48 3.565 ;
      RECT 7.3 3.232 7.525 3.518 ;
      RECT 7.275 3.243 7.56 3.455 ;
      RECT 7.275 3.327 7.595 3.455 ;
      RECT 7.275 3.302 7.59 3.455 ;
      RECT 7.335 3.218 7.48 3.585 ;
      RECT 7.421 3.217 7.48 3.585 ;
      RECT 7.421 3.216 7.465 3.585 ;
      RECT 7.335 7.855 7.505 8.305 ;
      RECT 7.39 6.075 7.56 8.025 ;
      RECT 7.335 5.015 7.505 6.245 ;
      RECT 6.815 5.015 6.985 8.305 ;
      RECT 6.815 7.315 7.22 7.645 ;
      RECT 6.815 6.475 7.22 6.805 ;
      RECT 7.12 2.732 7.125 3.11 ;
      RECT 7.115 2.7 7.12 3.11 ;
      RECT 7.11 2.672 7.115 3.11 ;
      RECT 7.105 2.652 7.11 3.11 ;
      RECT 7.05 2.635 7.105 3.11 ;
      RECT 7.01 2.62 7.05 3.11 ;
      RECT 6.955 2.607 7.01 3.11 ;
      RECT 6.92 2.598 6.955 3.11 ;
      RECT 6.916 2.596 6.92 3.109 ;
      RECT 6.83 2.592 6.916 3.092 ;
      RECT 6.745 2.584 6.83 3.055 ;
      RECT 6.735 2.58 6.745 3.028 ;
      RECT 6.725 2.58 6.735 3.01 ;
      RECT 6.715 2.582 6.725 2.993 ;
      RECT 6.71 2.587 6.715 2.979 ;
      RECT 6.705 2.591 6.71 2.966 ;
      RECT 6.695 2.596 6.705 2.95 ;
      RECT 6.68 2.61 6.695 2.925 ;
      RECT 6.675 2.616 6.68 2.905 ;
      RECT 6.67 2.618 6.675 2.898 ;
      RECT 6.665 2.622 6.67 2.773 ;
      RECT 6.845 3.422 7.09 3.885 ;
      RECT 6.765 3.395 7.085 3.881 ;
      RECT 6.695 3.43 7.09 3.874 ;
      RECT 6.485 3.685 7.09 3.87 ;
      RECT 6.665 3.453 7.09 3.87 ;
      RECT 6.505 3.645 7.09 3.87 ;
      RECT 6.655 3.465 7.09 3.87 ;
      RECT 6.54 3.582 7.09 3.87 ;
      RECT 6.595 3.507 7.09 3.87 ;
      RECT 6.845 3.372 7.085 3.885 ;
      RECT 6.875 3.365 7.085 3.885 ;
      RECT 6.865 3.367 7.085 3.885 ;
      RECT 6.875 3.362 7.005 3.885 ;
      RECT 6.43 1.925 6.516 2.364 ;
      RECT 6.425 1.925 6.516 2.362 ;
      RECT 6.425 1.925 6.585 2.361 ;
      RECT 6.425 1.925 6.615 2.358 ;
      RECT 6.41 1.932 6.615 2.349 ;
      RECT 6.41 1.932 6.62 2.345 ;
      RECT 6.405 1.942 6.62 2.338 ;
      RECT 6.4 1.947 6.62 2.313 ;
      RECT 6.4 1.947 6.635 2.295 ;
      RECT 6.425 1.925 6.655 2.21 ;
      RECT 6.395 1.952 6.655 2.208 ;
      RECT 6.405 1.945 6.66 2.146 ;
      RECT 6.395 2.067 6.665 2.129 ;
      RECT 6.38 1.962 6.66 2.08 ;
      RECT 6.375 1.972 6.66 1.98 ;
      RECT 6.455 2.743 6.46 2.82 ;
      RECT 6.445 2.737 6.455 3.01 ;
      RECT 6.435 2.729 6.445 3.031 ;
      RECT 6.425 2.72 6.435 3.053 ;
      RECT 6.42 2.715 6.425 3.07 ;
      RECT 6.38 2.715 6.42 3.11 ;
      RECT 6.36 2.715 6.38 3.165 ;
      RECT 6.355 2.715 6.36 3.193 ;
      RECT 6.345 2.715 6.355 3.208 ;
      RECT 6.31 2.715 6.345 3.25 ;
      RECT 6.305 2.715 6.31 3.293 ;
      RECT 6.295 2.715 6.305 3.308 ;
      RECT 6.28 2.715 6.295 3.328 ;
      RECT 6.265 2.715 6.28 3.355 ;
      RECT 6.26 2.716 6.265 3.373 ;
      RECT 6.24 2.717 6.26 3.38 ;
      RECT 6.185 2.718 6.24 3.4 ;
      RECT 6.175 2.719 6.185 3.414 ;
      RECT 6.17 2.722 6.175 3.413 ;
      RECT 6.13 2.795 6.17 3.411 ;
      RECT 6.115 2.875 6.13 3.409 ;
      RECT 6.09 2.93 6.115 3.407 ;
      RECT 6.075 2.995 6.09 3.406 ;
      RECT 6.03 3.027 6.075 3.403 ;
      RECT 5.945 3.05 6.03 3.398 ;
      RECT 5.92 3.07 5.945 3.393 ;
      RECT 5.85 3.075 5.92 3.389 ;
      RECT 5.83 3.077 5.85 3.386 ;
      RECT 5.745 3.088 5.83 3.38 ;
      RECT 5.74 3.099 5.745 3.375 ;
      RECT 5.73 3.101 5.74 3.375 ;
      RECT 5.695 3.105 5.73 3.373 ;
      RECT 5.645 3.115 5.695 3.36 ;
      RECT 5.625 3.123 5.645 3.345 ;
      RECT 5.545 3.135 5.625 3.328 ;
      RECT 5.71 2.685 5.88 2.895 ;
      RECT 5.826 2.681 5.88 2.895 ;
      RECT 5.631 2.685 5.88 2.886 ;
      RECT 5.631 2.685 5.885 2.875 ;
      RECT 5.545 2.685 5.885 2.866 ;
      RECT 5.545 2.693 5.895 2.81 ;
      RECT 5.545 2.705 5.9 2.723 ;
      RECT 5.545 2.712 5.905 2.715 ;
      RECT 5.74 2.683 5.88 2.895 ;
      RECT 5.495 3.628 5.74 3.96 ;
      RECT 5.49 3.62 5.495 3.957 ;
      RECT 5.46 3.64 5.74 3.938 ;
      RECT 5.44 3.672 5.74 3.911 ;
      RECT 5.49 3.625 5.667 3.957 ;
      RECT 5.49 3.622 5.581 3.957 ;
      RECT 5.43 1.97 5.6 2.39 ;
      RECT 5.425 1.97 5.6 2.388 ;
      RECT 5.425 1.97 5.625 2.378 ;
      RECT 5.425 1.97 5.645 2.353 ;
      RECT 5.42 1.97 5.645 2.348 ;
      RECT 5.42 1.97 5.655 2.338 ;
      RECT 5.42 1.97 5.66 2.333 ;
      RECT 5.42 1.975 5.665 2.328 ;
      RECT 5.42 2.007 5.68 2.318 ;
      RECT 5.42 2.077 5.705 2.301 ;
      RECT 5.4 2.077 5.705 2.293 ;
      RECT 5.4 2.137 5.715 2.27 ;
      RECT 5.4 2.177 5.725 2.215 ;
      RECT 5.385 1.97 5.66 2.195 ;
      RECT 5.375 1.985 5.665 2.093 ;
      RECT 4.965 3.375 5.135 3.9 ;
      RECT 4.96 3.375 5.135 3.893 ;
      RECT 4.95 3.375 5.14 3.858 ;
      RECT 4.945 3.385 5.14 3.83 ;
      RECT 4.94 3.405 5.14 3.813 ;
      RECT 4.95 3.38 5.145 3.803 ;
      RECT 4.935 3.425 5.145 3.795 ;
      RECT 4.93 3.445 5.145 3.78 ;
      RECT 4.925 3.475 5.145 3.77 ;
      RECT 4.915 3.52 5.145 3.745 ;
      RECT 4.945 3.39 5.15 3.728 ;
      RECT 4.91 3.572 5.15 3.723 ;
      RECT 4.945 3.4 5.155 3.693 ;
      RECT 4.905 3.605 5.155 3.69 ;
      RECT 4.9 3.63 5.155 3.67 ;
      RECT 4.94 3.417 5.165 3.61 ;
      RECT 4.935 3.439 5.175 3.503 ;
      RECT 4.885 2.686 4.9 2.955 ;
      RECT 4.84 2.67 4.885 3 ;
      RECT 4.835 2.658 4.84 3.05 ;
      RECT 4.825 2.654 4.835 3.083 ;
      RECT 4.82 2.651 4.825 3.111 ;
      RECT 4.805 2.653 4.82 3.153 ;
      RECT 4.8 2.657 4.805 3.193 ;
      RECT 4.78 2.662 4.8 3.245 ;
      RECT 4.776 2.667 4.78 3.302 ;
      RECT 4.69 2.686 4.776 3.339 ;
      RECT 4.68 2.707 4.69 3.375 ;
      RECT 4.675 2.715 4.68 3.376 ;
      RECT 4.67 2.757 4.675 3.377 ;
      RECT 4.655 2.845 4.67 3.378 ;
      RECT 4.645 2.995 4.655 3.38 ;
      RECT 4.64 3.04 4.645 3.382 ;
      RECT 4.605 3.082 4.64 3.385 ;
      RECT 4.6 3.1 4.605 3.388 ;
      RECT 4.523 3.106 4.6 3.394 ;
      RECT 4.437 3.12 4.523 3.407 ;
      RECT 4.351 3.134 4.437 3.421 ;
      RECT 4.265 3.148 4.351 3.434 ;
      RECT 4.205 3.16 4.265 3.446 ;
      RECT 4.18 3.167 4.205 3.453 ;
      RECT 4.166 3.17 4.18 3.458 ;
      RECT 4.08 3.178 4.166 3.474 ;
      RECT 4.075 3.185 4.08 3.489 ;
      RECT 4.051 3.185 4.075 3.496 ;
      RECT 3.965 3.188 4.051 3.524 ;
      RECT 3.88 3.192 3.965 3.568 ;
      RECT 3.815 3.196 3.88 3.605 ;
      RECT 3.79 3.199 3.815 3.621 ;
      RECT 3.715 3.212 3.79 3.625 ;
      RECT 3.69 3.23 3.715 3.629 ;
      RECT 3.68 3.237 3.69 3.631 ;
      RECT 3.665 3.24 3.68 3.632 ;
      RECT 3.605 3.252 3.665 3.636 ;
      RECT 3.595 3.266 3.605 3.64 ;
      RECT 3.54 3.276 3.595 3.628 ;
      RECT 3.515 3.297 3.54 3.611 ;
      RECT 3.495 3.317 3.515 3.602 ;
      RECT 3.49 3.33 3.495 3.597 ;
      RECT 3.475 3.342 3.49 3.593 ;
      RECT 4.71 1.997 4.715 2.02 ;
      RECT 4.705 1.988 4.71 2.06 ;
      RECT 4.7 1.986 4.705 2.103 ;
      RECT 4.695 1.977 4.7 2.138 ;
      RECT 4.69 1.967 4.695 2.21 ;
      RECT 4.685 1.957 4.69 2.275 ;
      RECT 4.68 1.954 4.685 2.315 ;
      RECT 4.655 1.948 4.68 2.405 ;
      RECT 4.62 1.936 4.655 2.43 ;
      RECT 4.61 1.927 4.62 2.43 ;
      RECT 4.475 1.925 4.485 2.413 ;
      RECT 4.465 1.925 4.475 2.38 ;
      RECT 4.46 1.925 4.465 2.355 ;
      RECT 4.455 1.925 4.46 2.343 ;
      RECT 4.45 1.925 4.455 2.325 ;
      RECT 4.44 1.925 4.45 2.29 ;
      RECT 4.435 1.927 4.44 2.268 ;
      RECT 4.43 1.933 4.435 2.253 ;
      RECT 4.425 1.939 4.43 2.238 ;
      RECT 4.41 1.951 4.425 2.211 ;
      RECT 4.405 1.962 4.41 2.179 ;
      RECT 4.4 1.972 4.405 2.163 ;
      RECT 4.39 1.98 4.4 2.132 ;
      RECT 4.385 1.99 4.39 2.106 ;
      RECT 4.38 2.047 4.385 2.089 ;
      RECT 4.485 1.925 4.61 2.43 ;
      RECT 4.2 2.612 4.46 2.91 ;
      RECT 4.195 2.619 4.46 2.908 ;
      RECT 4.2 2.614 4.475 2.903 ;
      RECT 4.19 2.627 4.475 2.9 ;
      RECT 4.19 2.632 4.48 2.893 ;
      RECT 4.185 2.64 4.48 2.89 ;
      RECT 4.185 2.657 4.485 2.688 ;
      RECT 4.2 2.609 4.431 2.91 ;
      RECT 4.255 2.608 4.431 2.91 ;
      RECT 4.255 2.605 4.345 2.91 ;
      RECT 4.255 2.602 4.341 2.91 ;
      RECT 3.945 2.875 3.95 2.888 ;
      RECT 3.94 2.842 3.945 2.893 ;
      RECT 3.935 2.797 3.94 2.9 ;
      RECT 3.93 2.752 3.935 2.908 ;
      RECT 3.925 2.72 3.93 2.916 ;
      RECT 3.92 2.68 3.925 2.917 ;
      RECT 3.905 2.66 3.92 2.919 ;
      RECT 3.83 2.642 3.905 2.931 ;
      RECT 3.82 2.635 3.83 2.942 ;
      RECT 3.815 2.635 3.82 2.944 ;
      RECT 3.785 2.641 3.815 2.948 ;
      RECT 3.745 2.654 3.785 2.948 ;
      RECT 3.72 2.665 3.745 2.934 ;
      RECT 3.705 2.671 3.72 2.917 ;
      RECT 3.695 2.673 3.705 2.908 ;
      RECT 3.69 2.674 3.695 2.903 ;
      RECT 3.685 2.675 3.69 2.898 ;
      RECT 3.68 2.676 3.685 2.895 ;
      RECT 3.655 2.681 3.68 2.885 ;
      RECT 3.645 2.697 3.655 2.872 ;
      RECT 3.64 2.717 3.645 2.867 ;
      RECT 3.65 2.11 3.655 2.306 ;
      RECT 3.635 2.074 3.65 2.308 ;
      RECT 3.625 2.056 3.635 2.313 ;
      RECT 3.615 2.042 3.625 2.317 ;
      RECT 3.57 2.026 3.615 2.327 ;
      RECT 3.565 2.016 3.57 2.336 ;
      RECT 3.52 2.005 3.565 2.342 ;
      RECT 3.515 1.993 3.52 2.349 ;
      RECT 3.5 1.988 3.515 2.353 ;
      RECT 3.485 1.98 3.5 2.358 ;
      RECT 3.475 1.973 3.485 2.363 ;
      RECT 3.465 1.97 3.475 2.368 ;
      RECT 3.455 1.97 3.465 2.369 ;
      RECT 3.45 1.967 3.455 2.368 ;
      RECT 3.415 1.962 3.44 2.367 ;
      RECT 3.391 1.958 3.415 2.366 ;
      RECT 3.305 1.949 3.391 2.363 ;
      RECT 3.29 1.941 3.305 2.36 ;
      RECT 3.268 1.94 3.29 2.359 ;
      RECT 3.182 1.94 3.268 2.357 ;
      RECT 3.096 1.94 3.182 2.355 ;
      RECT 3.01 1.94 3.096 2.352 ;
      RECT 3 1.94 3.01 2.343 ;
      RECT 2.97 1.94 3 2.303 ;
      RECT 2.96 1.95 2.97 2.258 ;
      RECT 2.955 1.99 2.96 2.243 ;
      RECT 2.95 2.005 2.955 2.23 ;
      RECT 2.92 2.085 2.95 2.192 ;
      RECT 3.44 1.965 3.45 2.368 ;
      RECT 3.265 2.73 3.28 3.335 ;
      RECT 3.27 2.725 3.28 3.335 ;
      RECT 3.435 2.725 3.44 2.908 ;
      RECT 3.425 2.725 3.435 2.938 ;
      RECT 3.41 2.725 3.425 2.998 ;
      RECT 3.405 2.725 3.41 3.043 ;
      RECT 3.4 2.725 3.405 3.073 ;
      RECT 3.395 2.725 3.4 3.093 ;
      RECT 3.385 2.725 3.395 3.128 ;
      RECT 3.37 2.725 3.385 3.16 ;
      RECT 3.325 2.725 3.37 3.188 ;
      RECT 3.32 2.725 3.325 3.218 ;
      RECT 3.315 2.725 3.32 3.23 ;
      RECT 3.31 2.725 3.315 3.238 ;
      RECT 3.3 2.725 3.31 3.253 ;
      RECT 3.295 2.725 3.3 3.275 ;
      RECT 3.285 2.725 3.295 3.298 ;
      RECT 3.28 2.725 3.285 3.318 ;
      RECT 3.245 2.74 3.265 3.335 ;
      RECT 3.22 2.757 3.245 3.335 ;
      RECT 3.215 2.767 3.22 3.335 ;
      RECT 3.185 2.782 3.215 3.335 ;
      RECT 3.11 2.824 3.185 3.335 ;
      RECT 3.105 2.855 3.11 3.318 ;
      RECT 3.1 2.859 3.105 3.3 ;
      RECT 3.095 2.863 3.1 3.263 ;
      RECT 3.09 3.047 3.095 3.23 ;
      RECT 2.575 3.236 2.661 3.801 ;
      RECT 2.53 3.238 2.695 3.795 ;
      RECT 2.661 3.235 2.695 3.795 ;
      RECT 2.575 3.237 2.78 3.789 ;
      RECT 2.53 3.247 2.79 3.785 ;
      RECT 2.505 3.239 2.78 3.781 ;
      RECT 2.5 3.242 2.78 3.776 ;
      RECT 2.475 3.257 2.79 3.77 ;
      RECT 2.475 3.282 2.83 3.765 ;
      RECT 2.435 3.29 2.83 3.74 ;
      RECT 2.435 3.317 2.845 3.738 ;
      RECT 2.435 3.347 2.855 3.725 ;
      RECT 2.43 3.492 2.855 3.713 ;
      RECT 2.435 3.421 2.875 3.71 ;
      RECT 2.435 3.478 2.88 3.518 ;
      RECT 2.625 2.757 2.795 2.935 ;
      RECT 2.575 2.696 2.625 2.92 ;
      RECT 2.31 2.676 2.575 2.905 ;
      RECT 2.27 2.74 2.745 2.905 ;
      RECT 2.27 2.73 2.7 2.905 ;
      RECT 2.27 2.727 2.69 2.905 ;
      RECT 2.27 2.715 2.68 2.905 ;
      RECT 2.27 2.7 2.625 2.905 ;
      RECT 2.31 2.672 2.511 2.905 ;
      RECT 2.32 2.65 2.511 2.905 ;
      RECT 2.345 2.635 2.425 2.905 ;
      RECT 2.1 3.165 2.22 3.61 ;
      RECT 2.085 3.165 2.22 3.609 ;
      RECT 2.04 3.187 2.22 3.604 ;
      RECT 2 3.236 2.22 3.598 ;
      RECT 2 3.236 2.225 3.573 ;
      RECT 2 3.236 2.245 3.463 ;
      RECT 1.995 3.266 2.245 3.46 ;
      RECT 2.085 3.165 2.255 3.355 ;
      RECT 1.745 1.95 1.75 2.395 ;
      RECT 1.555 1.95 1.575 2.36 ;
      RECT 1.525 1.95 1.53 2.335 ;
      RECT 2.205 2.257 2.22 2.445 ;
      RECT 2.2 2.242 2.205 2.451 ;
      RECT 2.18 2.215 2.2 2.454 ;
      RECT 2.13 2.182 2.18 2.463 ;
      RECT 2.1 2.162 2.13 2.467 ;
      RECT 2.081 2.15 2.1 2.463 ;
      RECT 1.995 2.122 2.081 2.453 ;
      RECT 1.985 2.097 1.995 2.443 ;
      RECT 1.915 2.065 1.985 2.435 ;
      RECT 1.89 2.025 1.915 2.427 ;
      RECT 1.87 2.007 1.89 2.421 ;
      RECT 1.86 1.997 1.87 2.418 ;
      RECT 1.85 1.99 1.86 2.416 ;
      RECT 1.83 1.977 1.85 2.413 ;
      RECT 1.82 1.967 1.83 2.41 ;
      RECT 1.81 1.96 1.82 2.408 ;
      RECT 1.76 1.952 1.81 2.402 ;
      RECT 1.75 1.95 1.76 2.396 ;
      RECT 1.72 1.95 1.745 2.393 ;
      RECT 1.691 1.95 1.72 2.388 ;
      RECT 1.605 1.95 1.691 2.378 ;
      RECT 1.575 1.95 1.605 2.365 ;
      RECT 1.53 1.95 1.555 2.348 ;
      RECT 1.515 1.95 1.525 2.33 ;
      RECT 1.495 1.957 1.515 2.315 ;
      RECT 1.49 1.972 1.495 2.303 ;
      RECT 1.485 1.977 1.49 2.243 ;
      RECT 1.48 1.982 1.485 2.085 ;
      RECT 1.475 1.985 1.48 2.003 ;
      RECT 1.74 2.67 1.826 2.991 ;
      RECT 1.74 2.67 1.86 2.984 ;
      RECT 1.69 2.67 1.86 2.98 ;
      RECT 1.69 2.672 1.946 2.978 ;
      RECT 1.69 2.674 1.97 2.972 ;
      RECT 1.69 2.681 1.98 2.971 ;
      RECT 1.69 2.69 1.985 2.968 ;
      RECT 1.69 2.696 1.99 2.963 ;
      RECT 1.69 2.74 1.995 2.96 ;
      RECT 1.69 2.832 2 2.957 ;
      RECT 1.215 3.275 1.25 3.595 ;
      RECT 1.8 3.46 1.805 3.642 ;
      RECT 1.755 3.342 1.8 3.661 ;
      RECT 1.74 3.319 1.755 3.684 ;
      RECT 1.73 3.309 1.74 3.694 ;
      RECT 1.71 3.304 1.73 3.707 ;
      RECT 1.685 3.302 1.71 3.728 ;
      RECT 1.666 3.301 1.685 3.74 ;
      RECT 1.58 3.298 1.666 3.74 ;
      RECT 1.51 3.293 1.58 3.728 ;
      RECT 1.435 3.289 1.51 3.703 ;
      RECT 1.37 3.285 1.435 3.67 ;
      RECT 1.3 3.282 1.37 3.63 ;
      RECT 1.27 3.278 1.3 3.605 ;
      RECT 1.25 3.276 1.27 3.598 ;
      RECT 1.166 3.274 1.215 3.596 ;
      RECT 1.08 3.271 1.166 3.597 ;
      RECT 1.005 3.27 1.08 3.599 ;
      RECT 0.92 3.27 1.005 3.625 ;
      RECT 0.843 3.271 0.92 3.65 ;
      RECT 0.757 3.272 0.843 3.65 ;
      RECT 0.671 3.272 0.757 3.65 ;
      RECT 0.585 3.273 0.671 3.65 ;
      RECT 0.565 3.274 0.585 3.642 ;
      RECT 0.55 3.28 0.565 3.627 ;
      RECT 0.515 3.3 0.55 3.607 ;
      RECT 0.505 3.32 0.515 3.589 ;
      RECT 1.475 2.625 1.48 2.895 ;
      RECT 1.47 2.616 1.475 2.9 ;
      RECT 1.46 2.606 1.47 2.912 ;
      RECT 1.455 2.595 1.46 2.923 ;
      RECT 1.435 2.589 1.455 2.941 ;
      RECT 1.39 2.586 1.435 2.99 ;
      RECT 1.375 2.585 1.39 3.035 ;
      RECT 1.37 2.585 1.375 3.048 ;
      RECT 1.36 2.585 1.37 3.06 ;
      RECT 1.355 2.586 1.36 3.075 ;
      RECT 1.335 2.594 1.355 3.08 ;
      RECT 1.305 2.61 1.335 3.08 ;
      RECT 1.295 2.622 1.3 3.08 ;
      RECT 1.26 2.637 1.295 3.08 ;
      RECT 1.23 2.657 1.26 3.08 ;
      RECT 1.22 2.682 1.23 3.08 ;
      RECT 1.215 2.71 1.22 3.08 ;
      RECT 1.21 2.74 1.215 3.08 ;
      RECT 1.205 2.757 1.21 3.08 ;
      RECT 1.195 2.785 1.205 3.08 ;
      RECT 1.185 2.82 1.195 3.08 ;
      RECT 1.18 2.855 1.185 3.08 ;
      RECT 1.3 2.62 1.305 3.08 ;
      RECT 0.815 2.722 1 2.895 ;
      RECT 0.775 2.64 0.96 2.893 ;
      RECT 0.736 2.645 0.96 2.889 ;
      RECT 0.65 2.654 0.96 2.884 ;
      RECT 0.566 2.67 0.965 2.879 ;
      RECT 0.48 2.69 0.99 2.873 ;
      RECT 0.48 2.71 0.995 2.873 ;
      RECT 0.566 2.68 0.99 2.879 ;
      RECT 0.65 2.655 0.965 2.884 ;
      RECT 0.815 2.637 0.96 2.895 ;
      RECT 0.815 2.632 0.915 2.895 ;
      RECT 0.901 2.626 0.915 2.895 ;
      RECT 0.29 1.95 0.295 2.349 ;
      RECT 0.035 1.95 0.07 2.347 ;
      RECT -0.37 1.985 -0.365 2.341 ;
      RECT 0.375 1.988 0.38 2.243 ;
      RECT 0.37 1.986 0.375 2.249 ;
      RECT 0.365 1.985 0.37 2.256 ;
      RECT 0.34 1.978 0.365 2.28 ;
      RECT 0.335 1.971 0.34 2.304 ;
      RECT 0.33 1.967 0.335 2.313 ;
      RECT 0.32 1.962 0.33 2.326 ;
      RECT 0.315 1.959 0.32 2.335 ;
      RECT 0.31 1.957 0.315 2.34 ;
      RECT 0.295 1.953 0.31 2.35 ;
      RECT 0.28 1.947 0.29 2.349 ;
      RECT 0.242 1.945 0.28 2.349 ;
      RECT 0.156 1.947 0.242 2.349 ;
      RECT 0.07 1.949 0.156 2.348 ;
      RECT -0.001 1.95 0.035 2.347 ;
      RECT -0.087 1.952 -0.001 2.347 ;
      RECT -0.173 1.954 -0.087 2.346 ;
      RECT -0.259 1.956 -0.173 2.346 ;
      RECT -0.345 1.959 -0.259 2.345 ;
      RECT -0.355 1.965 -0.345 2.344 ;
      RECT -0.365 1.977 -0.355 2.342 ;
      RECT -0.425 2.012 -0.37 2.338 ;
      RECT -0.43 2.042 -0.425 2.1 ;
      RECT 0.315 3.122 0.33 3.315 ;
      RECT 0.31 3.09 0.315 3.315 ;
      RECT 0.3 3.065 0.31 3.315 ;
      RECT 0.295 3.037 0.3 3.315 ;
      RECT 0.265 2.96 0.295 3.315 ;
      RECT 0.24 2.842 0.265 3.315 ;
      RECT 0.235 2.78 0.24 3.315 ;
      RECT 0.225 2.767 0.235 3.315 ;
      RECT 0.205 2.757 0.225 3.315 ;
      RECT 0.19 2.74 0.205 3.315 ;
      RECT 0.16 2.728 0.19 3.315 ;
      RECT 0.155 2.727 0.16 3.26 ;
      RECT 0.15 2.727 0.155 3.218 ;
      RECT 0.135 2.726 0.15 3.17 ;
      RECT 0.12 2.726 0.135 3.108 ;
      RECT 0.1 2.726 0.12 3.068 ;
      RECT 0.095 2.726 0.1 3.053 ;
      RECT 0.07 2.725 0.095 3.048 ;
      RECT 0 2.724 0.07 3.035 ;
      RECT -0.015 2.723 0 3.02 ;
      RECT -0.045 2.722 -0.015 3.003 ;
      RECT -0.05 2.722 -0.045 2.988 ;
      RECT -0.1 2.721 -0.05 2.968 ;
      RECT -0.165 2.72 -0.1 2.923 ;
      RECT -0.17 2.72 -0.165 2.895 ;
      RECT -0.085 3.257 -0.08 3.514 ;
      RECT -0.105 3.176 -0.085 3.531 ;
      RECT -0.125 3.17 -0.105 3.56 ;
      RECT -0.185 3.157 -0.125 3.58 ;
      RECT -0.23 3.141 -0.185 3.581 ;
      RECT -0.314 3.129 -0.23 3.569 ;
      RECT -0.4 3.116 -0.314 3.553 ;
      RECT -0.41 3.109 -0.4 3.545 ;
      RECT -0.455 3.106 -0.41 3.485 ;
      RECT -0.475 3.102 -0.455 3.4 ;
      RECT -0.49 3.1 -0.475 3.353 ;
      RECT -0.52 3.097 -0.49 3.323 ;
      RECT -0.555 3.093 -0.52 3.3 ;
      RECT -0.598 3.088 -0.555 3.288 ;
      RECT -0.684 3.079 -0.598 3.297 ;
      RECT -0.77 3.068 -0.684 3.309 ;
      RECT -0.835 3.059 -0.77 3.318 ;
      RECT -0.855 3.05 -0.835 3.323 ;
      RECT -0.86 3.043 -0.855 3.325 ;
      RECT -0.9 3.028 -0.86 3.322 ;
      RECT -0.92 3.007 -0.9 3.317 ;
      RECT -0.935 2.995 -0.92 3.31 ;
      RECT -0.94 2.987 -0.935 3.303 ;
      RECT -0.955 2.967 -0.94 3.296 ;
      RECT -0.96 2.83 -0.955 3.29 ;
      RECT -1.04 2.719 -0.96 3.262 ;
      RECT -1.049 2.712 -1.04 3.228 ;
      RECT -1.135 2.706 -1.049 3.153 ;
      RECT -1.16 2.697 -1.135 3.065 ;
      RECT -1.19 2.692 -1.16 3.04 ;
      RECT -1.255 2.701 -1.19 3.025 ;
      RECT -1.275 2.717 -1.255 3 ;
      RECT -1.285 2.723 -1.275 2.948 ;
      RECT -1.305 2.745 -1.285 2.83 ;
      RECT -0.65 2.71 -0.48 2.895 ;
      RECT -0.65 2.71 -0.445 2.893 ;
      RECT -0.6 2.62 -0.43 2.884 ;
      RECT -0.65 2.777 -0.425 2.877 ;
      RECT -0.635 2.655 -0.43 2.884 ;
      RECT -1.435 3.388 -1.37 3.831 ;
      RECT -1.495 3.413 -1.37 3.829 ;
      RECT -1.495 3.413 -1.315 3.823 ;
      RECT -1.51 3.438 -1.315 3.822 ;
      RECT -1.37 3.375 -1.295 3.819 ;
      RECT -1.435 3.4 -1.215 3.813 ;
      RECT -1.51 3.439 -1.17 3.807 ;
      RECT -1.525 3.466 -1.17 3.798 ;
      RECT -1.51 3.459 -1.15 3.79 ;
      RECT -1.525 3.468 -1.145 3.773 ;
      RECT -1.53 3.485 -1.145 3.6 ;
      RECT -1.525 2.207 -1.49 2.445 ;
      RECT -1.525 2.207 -1.46 2.444 ;
      RECT -1.525 2.207 -1.345 2.44 ;
      RECT -1.525 2.207 -1.29 2.418 ;
      RECT -1.515 2.15 -1.235 2.318 ;
      RECT -1.41 1.99 -1.38 2.441 ;
      RECT -1.38 1.985 -1.2 2.198 ;
      RECT -1.51 2.126 -1.2 2.198 ;
      RECT -1.46 2.022 -1.41 2.442 ;
      RECT -1.49 2.078 -1.2 2.198 ;
      RECT -3.695 7.855 -3.525 8.305 ;
      RECT -3.64 6.075 -3.47 8.025 ;
      RECT -3.695 5.015 -3.525 6.245 ;
      RECT -4.215 5.015 -4.045 8.305 ;
      RECT -4.215 7.315 -3.81 7.645 ;
      RECT -4.215 6.475 -3.81 6.805 ;
      RECT 87.01 0.575 87.18 1.085 ;
      RECT 87.01 2.395 87.18 3.865 ;
      RECT 87.01 5.015 87.18 6.485 ;
      RECT 87.01 7.795 87.18 8.305 ;
      RECT 86.02 0.575 86.19 1.085 ;
      RECT 86.02 2.395 86.19 3.865 ;
      RECT 86.02 5.015 86.19 6.485 ;
      RECT 86.02 7.795 86.19 8.305 ;
      RECT 84.655 0.575 84.825 3.865 ;
      RECT 84.655 5.015 84.825 8.305 ;
      RECT 84.225 0.575 84.395 1.085 ;
      RECT 84.225 1.655 84.395 3.865 ;
      RECT 84.225 5.015 84.395 7.225 ;
      RECT 84.225 7.795 84.395 8.305 ;
      RECT 82.855 1.66 83.025 2.935 ;
      RECT 82.855 5.945 83.025 7.22 ;
      RECT 79.895 5.015 80.065 8.305 ;
      RECT 79.465 5.015 79.635 7.225 ;
      RECT 79.465 7.795 79.635 8.305 ;
      RECT 78.095 5.945 78.265 7.22 ;
      RECT 69.085 0.575 69.255 1.085 ;
      RECT 69.085 2.395 69.255 3.865 ;
      RECT 69.085 5.015 69.255 6.485 ;
      RECT 69.085 7.795 69.255 8.305 ;
      RECT 68.095 0.575 68.265 1.085 ;
      RECT 68.095 2.395 68.265 3.865 ;
      RECT 68.095 5.015 68.265 6.485 ;
      RECT 68.095 7.795 68.265 8.305 ;
      RECT 66.73 0.575 66.9 3.865 ;
      RECT 66.73 5.015 66.9 8.305 ;
      RECT 66.3 0.575 66.47 1.085 ;
      RECT 66.3 1.655 66.47 3.865 ;
      RECT 66.3 5.015 66.47 7.225 ;
      RECT 66.3 7.795 66.47 8.305 ;
      RECT 64.93 1.66 65.1 2.935 ;
      RECT 64.93 5.945 65.1 7.22 ;
      RECT 61.97 5.015 62.14 8.305 ;
      RECT 61.54 5.015 61.71 7.225 ;
      RECT 61.54 7.795 61.71 8.305 ;
      RECT 60.17 5.945 60.34 7.22 ;
      RECT 51.16 0.575 51.33 1.085 ;
      RECT 51.16 2.395 51.33 3.865 ;
      RECT 51.16 5.015 51.33 6.485 ;
      RECT 51.16 7.795 51.33 8.305 ;
      RECT 50.17 0.575 50.34 1.085 ;
      RECT 50.17 2.395 50.34 3.865 ;
      RECT 50.17 5.015 50.34 6.485 ;
      RECT 50.17 7.795 50.34 8.305 ;
      RECT 48.805 0.575 48.975 3.865 ;
      RECT 48.805 5.015 48.975 8.305 ;
      RECT 48.375 0.575 48.545 1.085 ;
      RECT 48.375 1.655 48.545 3.865 ;
      RECT 48.375 5.015 48.545 7.225 ;
      RECT 48.375 7.795 48.545 8.305 ;
      RECT 47.005 1.66 47.175 2.935 ;
      RECT 47.005 5.945 47.175 7.22 ;
      RECT 44.045 5.015 44.215 8.305 ;
      RECT 43.615 5.015 43.785 7.225 ;
      RECT 43.615 7.795 43.785 8.305 ;
      RECT 42.245 5.945 42.415 7.22 ;
      RECT 33.235 0.575 33.405 1.085 ;
      RECT 33.235 2.395 33.405 3.865 ;
      RECT 33.235 5.015 33.405 6.485 ;
      RECT 33.235 7.795 33.405 8.305 ;
      RECT 32.245 0.575 32.415 1.085 ;
      RECT 32.245 2.395 32.415 3.865 ;
      RECT 32.245 5.015 32.415 6.485 ;
      RECT 32.245 7.795 32.415 8.305 ;
      RECT 30.88 0.575 31.05 3.865 ;
      RECT 30.88 5.015 31.05 8.305 ;
      RECT 30.45 0.575 30.62 1.085 ;
      RECT 30.45 1.655 30.62 3.865 ;
      RECT 30.45 5.015 30.62 7.225 ;
      RECT 30.45 7.795 30.62 8.305 ;
      RECT 29.08 1.66 29.25 2.935 ;
      RECT 29.08 5.945 29.25 7.22 ;
      RECT 26.12 5.015 26.29 8.305 ;
      RECT 25.69 5.015 25.86 7.225 ;
      RECT 25.69 7.795 25.86 8.305 ;
      RECT 24.32 5.945 24.49 7.22 ;
      RECT 15.31 0.575 15.48 1.085 ;
      RECT 15.31 2.395 15.48 3.865 ;
      RECT 15.31 5.015 15.48 6.485 ;
      RECT 15.31 7.795 15.48 8.305 ;
      RECT 14.32 0.575 14.49 1.085 ;
      RECT 14.32 2.395 14.49 3.865 ;
      RECT 14.32 5.015 14.49 6.485 ;
      RECT 14.32 7.795 14.49 8.305 ;
      RECT 12.955 0.575 13.125 3.865 ;
      RECT 12.955 5.015 13.125 8.305 ;
      RECT 12.525 0.575 12.695 1.085 ;
      RECT 12.525 1.655 12.695 3.865 ;
      RECT 12.525 5.015 12.695 7.225 ;
      RECT 12.525 7.795 12.695 8.305 ;
      RECT 11.155 1.66 11.325 2.935 ;
      RECT 11.155 5.945 11.325 7.22 ;
      RECT 8.195 5.015 8.365 8.305 ;
      RECT 7.765 5.015 7.935 7.225 ;
      RECT 7.765 7.795 7.935 8.305 ;
      RECT 6.395 5.945 6.565 7.22 ;
      RECT -3.265 5.015 -3.095 7.225 ;
      RECT -3.265 7.795 -3.095 8.305 ;
      RECT -4.635 5.945 -4.465 7.22 ;
  END
END sky130_osu_ring_oscillator_mpr2at_8_b0r1

MACRO sky130_osu_ring_oscillator_mpr2at_8_b0r2
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 92.575 BY 8.88 ;
  SYMMETRY X Y R90 ;
  SITE CoreSite ;
  OBS
    LAYER met3 ;
      RECT 84.38 7.055 84.755 7.425 ;
      RECT 84.415 4.925 84.725 7.425 ;
      RECT 84.415 4.925 87.51 5.235 ;
      RECT 87.2 1.125 87.51 5.235 ;
      RECT 87.2 1.14 87.575 1.51 ;
      RECT 84.33 3.685 84.885 4.015 ;
      RECT 84.33 2.02 84.63 4.015 ;
      RECT 80.395 3.125 80.95 3.455 ;
      RECT 80.65 2.02 80.95 3.455 ;
      RECT 81.445 1.885 81.595 2.535 ;
      RECT 80.65 2.02 84.63 2.32 ;
      RECT 79.165 0.96 79.465 3.91 ;
      RECT 79.155 2.565 79.885 2.895 ;
      RECT 79.12 0.96 79.495 1.33 ;
      RECT 77.715 3.125 78.445 3.455 ;
      RECT 77.73 0.96 78.03 3.455 ;
      RECT 75.605 2.565 76.335 2.895 ;
      RECT 75.76 0.93 76.06 2.895 ;
      RECT 77.685 0.96 78.06 1.33 ;
      RECT 75.715 0.93 76.09 1.3 ;
      RECT 75.715 0.97 78.06 1.27 ;
      RECT 66.455 7.055 66.83 7.425 ;
      RECT 66.49 4.925 66.8 7.425 ;
      RECT 66.49 4.925 69.585 5.235 ;
      RECT 69.275 1.125 69.585 5.235 ;
      RECT 69.275 1.14 69.65 1.51 ;
      RECT 66.405 3.685 66.96 4.015 ;
      RECT 66.405 2.02 66.705 4.015 ;
      RECT 62.47 3.125 63.025 3.455 ;
      RECT 62.725 2.02 63.025 3.455 ;
      RECT 63.52 1.885 63.67 2.535 ;
      RECT 62.725 2.02 66.705 2.32 ;
      RECT 61.24 0.96 61.54 3.91 ;
      RECT 61.23 2.565 61.96 2.895 ;
      RECT 61.195 0.96 61.57 1.33 ;
      RECT 59.79 3.125 60.52 3.455 ;
      RECT 59.805 0.96 60.105 3.455 ;
      RECT 57.68 2.565 58.41 2.895 ;
      RECT 57.835 0.93 58.135 2.895 ;
      RECT 59.76 0.96 60.135 1.33 ;
      RECT 57.79 0.93 58.165 1.3 ;
      RECT 57.79 0.97 60.135 1.27 ;
      RECT 48.53 7.055 48.905 7.425 ;
      RECT 48.565 4.925 48.875 7.425 ;
      RECT 48.565 4.925 51.66 5.235 ;
      RECT 51.35 1.125 51.66 5.235 ;
      RECT 51.35 1.14 51.725 1.51 ;
      RECT 48.48 3.685 49.035 4.015 ;
      RECT 48.48 2.02 48.78 4.015 ;
      RECT 44.545 3.125 45.1 3.455 ;
      RECT 44.8 2.02 45.1 3.455 ;
      RECT 45.595 1.885 45.745 2.535 ;
      RECT 44.8 2.02 48.78 2.32 ;
      RECT 43.315 0.96 43.615 3.91 ;
      RECT 43.305 2.565 44.035 2.895 ;
      RECT 43.27 0.96 43.645 1.33 ;
      RECT 41.865 3.125 42.595 3.455 ;
      RECT 41.88 0.96 42.18 3.455 ;
      RECT 39.755 2.565 40.485 2.895 ;
      RECT 39.91 0.93 40.21 2.895 ;
      RECT 41.835 0.96 42.21 1.33 ;
      RECT 39.865 0.93 40.24 1.3 ;
      RECT 39.865 0.97 42.21 1.27 ;
      RECT 30.605 7.055 30.98 7.425 ;
      RECT 30.64 4.925 30.95 7.425 ;
      RECT 30.64 4.925 33.735 5.235 ;
      RECT 33.425 1.125 33.735 5.235 ;
      RECT 33.425 1.14 33.8 1.51 ;
      RECT 30.555 3.685 31.11 4.015 ;
      RECT 30.555 2.02 30.855 4.015 ;
      RECT 26.62 3.125 27.175 3.455 ;
      RECT 26.875 2.02 27.175 3.455 ;
      RECT 27.67 1.885 27.82 2.535 ;
      RECT 26.875 2.02 30.855 2.32 ;
      RECT 25.39 0.96 25.69 3.91 ;
      RECT 25.38 2.565 26.11 2.895 ;
      RECT 25.345 0.96 25.72 1.33 ;
      RECT 23.94 3.125 24.67 3.455 ;
      RECT 23.955 0.96 24.255 3.455 ;
      RECT 21.83 2.565 22.56 2.895 ;
      RECT 21.985 0.93 22.285 2.895 ;
      RECT 23.91 0.96 24.285 1.33 ;
      RECT 21.94 0.93 22.315 1.3 ;
      RECT 21.94 0.97 24.285 1.27 ;
      RECT 12.68 7.055 13.055 7.425 ;
      RECT 12.715 4.925 13.025 7.425 ;
      RECT 12.715 4.925 15.81 5.235 ;
      RECT 15.5 1.125 15.81 5.235 ;
      RECT 15.5 1.14 15.875 1.51 ;
      RECT 12.63 3.685 13.185 4.015 ;
      RECT 12.63 2.02 12.93 4.015 ;
      RECT 8.695 3.125 9.25 3.455 ;
      RECT 8.95 2.02 9.25 3.455 ;
      RECT 9.745 1.885 9.895 2.535 ;
      RECT 8.95 2.02 12.93 2.32 ;
      RECT 7.465 0.96 7.765 3.91 ;
      RECT 7.455 2.565 8.185 2.895 ;
      RECT 7.42 0.96 7.795 1.33 ;
      RECT 6.015 3.125 6.745 3.455 ;
      RECT 6.03 0.96 6.33 3.455 ;
      RECT 3.905 2.565 4.635 2.895 ;
      RECT 4.06 0.93 4.36 2.895 ;
      RECT 5.985 0.96 6.36 1.33 ;
      RECT 4.015 0.93 4.39 1.3 ;
      RECT 4.015 0.97 6.36 1.27 ;
      RECT 85.515 2.005 86.245 2.335 ;
      RECT 83.295 3.685 84.025 4.015 ;
      RECT 81.595 3.685 82.325 4.015 ;
      RECT 76.64 2.565 77.37 2.895 ;
      RECT 75.275 3.685 76.005 4.015 ;
      RECT 67.59 2.005 68.32 2.335 ;
      RECT 65.37 3.685 66.1 4.015 ;
      RECT 63.67 3.685 64.4 4.015 ;
      RECT 58.715 2.565 59.445 2.895 ;
      RECT 57.35 3.685 58.08 4.015 ;
      RECT 49.665 2.005 50.395 2.335 ;
      RECT 47.445 3.685 48.175 4.015 ;
      RECT 45.745 3.685 46.475 4.015 ;
      RECT 40.79 2.565 41.52 2.895 ;
      RECT 39.425 3.685 40.155 4.015 ;
      RECT 31.74 2.005 32.47 2.335 ;
      RECT 29.52 3.685 30.25 4.015 ;
      RECT 27.82 3.685 28.55 4.015 ;
      RECT 22.865 2.565 23.595 2.895 ;
      RECT 21.5 3.685 22.23 4.015 ;
      RECT 13.815 2.005 14.545 2.335 ;
      RECT 11.595 3.685 12.325 4.015 ;
      RECT 9.895 3.685 10.625 4.015 ;
      RECT 4.94 2.565 5.67 2.895 ;
      RECT 3.575 3.685 4.305 4.015 ;
    LAYER via2 ;
      RECT 87.29 1.225 87.49 1.425 ;
      RECT 85.58 2.07 85.78 2.27 ;
      RECT 84.62 3.75 84.82 3.95 ;
      RECT 84.47 7.14 84.67 7.34 ;
      RECT 83.62 3.75 83.82 3.95 ;
      RECT 81.66 3.75 81.86 3.95 ;
      RECT 80.46 3.19 80.66 3.39 ;
      RECT 79.22 2.63 79.42 2.83 ;
      RECT 79.21 1.045 79.41 1.245 ;
      RECT 77.78 3.19 77.98 3.39 ;
      RECT 77.775 1.04 77.975 1.24 ;
      RECT 77.04 2.63 77.24 2.83 ;
      RECT 75.82 2.63 76.02 2.83 ;
      RECT 75.805 1.015 76.005 1.215 ;
      RECT 75.34 3.75 75.54 3.95 ;
      RECT 69.365 1.225 69.565 1.425 ;
      RECT 67.655 2.07 67.855 2.27 ;
      RECT 66.695 3.75 66.895 3.95 ;
      RECT 66.545 7.14 66.745 7.34 ;
      RECT 65.695 3.75 65.895 3.95 ;
      RECT 63.735 3.75 63.935 3.95 ;
      RECT 62.535 3.19 62.735 3.39 ;
      RECT 61.295 2.63 61.495 2.83 ;
      RECT 61.285 1.045 61.485 1.245 ;
      RECT 59.855 3.19 60.055 3.39 ;
      RECT 59.85 1.04 60.05 1.24 ;
      RECT 59.115 2.63 59.315 2.83 ;
      RECT 57.895 2.63 58.095 2.83 ;
      RECT 57.88 1.015 58.08 1.215 ;
      RECT 57.415 3.75 57.615 3.95 ;
      RECT 51.44 1.225 51.64 1.425 ;
      RECT 49.73 2.07 49.93 2.27 ;
      RECT 48.77 3.75 48.97 3.95 ;
      RECT 48.62 7.14 48.82 7.34 ;
      RECT 47.77 3.75 47.97 3.95 ;
      RECT 45.81 3.75 46.01 3.95 ;
      RECT 44.61 3.19 44.81 3.39 ;
      RECT 43.37 2.63 43.57 2.83 ;
      RECT 43.36 1.045 43.56 1.245 ;
      RECT 41.93 3.19 42.13 3.39 ;
      RECT 41.925 1.04 42.125 1.24 ;
      RECT 41.19 2.63 41.39 2.83 ;
      RECT 39.97 2.63 40.17 2.83 ;
      RECT 39.955 1.015 40.155 1.215 ;
      RECT 39.49 3.75 39.69 3.95 ;
      RECT 33.515 1.225 33.715 1.425 ;
      RECT 31.805 2.07 32.005 2.27 ;
      RECT 30.845 3.75 31.045 3.95 ;
      RECT 30.695 7.14 30.895 7.34 ;
      RECT 29.845 3.75 30.045 3.95 ;
      RECT 27.885 3.75 28.085 3.95 ;
      RECT 26.685 3.19 26.885 3.39 ;
      RECT 25.445 2.63 25.645 2.83 ;
      RECT 25.435 1.045 25.635 1.245 ;
      RECT 24.005 3.19 24.205 3.39 ;
      RECT 24 1.04 24.2 1.24 ;
      RECT 23.265 2.63 23.465 2.83 ;
      RECT 22.045 2.63 22.245 2.83 ;
      RECT 22.03 1.015 22.23 1.215 ;
      RECT 21.565 3.75 21.765 3.95 ;
      RECT 15.59 1.225 15.79 1.425 ;
      RECT 13.88 2.07 14.08 2.27 ;
      RECT 12.92 3.75 13.12 3.95 ;
      RECT 12.77 7.14 12.97 7.34 ;
      RECT 11.92 3.75 12.12 3.95 ;
      RECT 9.96 3.75 10.16 3.95 ;
      RECT 8.76 3.19 8.96 3.39 ;
      RECT 7.52 2.63 7.72 2.83 ;
      RECT 7.51 1.045 7.71 1.245 ;
      RECT 6.08 3.19 6.28 3.39 ;
      RECT 6.075 1.04 6.275 1.24 ;
      RECT 5.34 2.63 5.54 2.83 ;
      RECT 4.12 2.63 4.32 2.83 ;
      RECT 4.105 1.015 4.305 1.215 ;
      RECT 3.64 3.75 3.84 3.95 ;
    LAYER met2 ;
      RECT 1.385 8.4 92.2 8.57 ;
      RECT 92.03 7.275 92.2 8.57 ;
      RECT 1.385 6.255 1.555 8.57 ;
      RECT 92 7.275 92.35 7.625 ;
      RECT 1.325 6.255 1.615 6.605 ;
      RECT 88.845 6.225 89.165 6.545 ;
      RECT 88.875 5.695 89.045 6.545 ;
      RECT 88.875 5.695 89.05 6.045 ;
      RECT 88.875 5.695 89.85 5.87 ;
      RECT 89.675 1.965 89.85 5.87 ;
      RECT 89.62 1.965 89.97 2.315 ;
      RECT 89.645 6.655 89.97 6.98 ;
      RECT 88.53 6.745 89.97 6.915 ;
      RECT 88.53 2.395 88.69 6.915 ;
      RECT 88.845 2.365 89.165 2.685 ;
      RECT 88.53 2.395 89.165 2.565 ;
      RECT 87.79 5.84 88.14 6.19 ;
      RECT 87.865 2.705 88.04 6.19 ;
      RECT 87.8 2.705 88.15 3.055 ;
      RECT 87.2 1.14 87.575 1.51 ;
      RECT 79.12 0.96 79.495 1.33 ;
      RECT 77.685 0.96 78.06 1.33 ;
      RECT 77.685 1.08 87.505 1.25 ;
      RECT 81.805 4.36 87.485 4.53 ;
      RECT 87.315 3.425 87.485 4.53 ;
      RECT 81.615 3.6 81.64 4.53 ;
      RECT 81.87 3.71 81.9 3.99 ;
      RECT 81.575 3.6 81.64 3.86 ;
      RECT 87.225 3.43 87.575 3.78 ;
      RECT 81.405 2.225 81.44 2.485 ;
      RECT 81.18 2.225 81.24 2.485 ;
      RECT 81.86 3.69 81.87 3.99 ;
      RECT 81.855 3.65 81.86 3.99 ;
      RECT 81.84 3.605 81.855 3.99 ;
      RECT 81.835 3.57 81.84 3.99 ;
      RECT 81.83 3.55 81.835 3.99 ;
      RECT 81.805 3.487 81.83 3.99 ;
      RECT 81.8 3.425 81.805 4.53 ;
      RECT 81.78 3.375 81.8 4.53 ;
      RECT 81.77 3.305 81.78 4.53 ;
      RECT 81.725 3.245 81.77 4.53 ;
      RECT 81.64 3.206 81.725 4.53 ;
      RECT 81.635 3.197 81.64 3.57 ;
      RECT 81.625 3.196 81.635 3.553 ;
      RECT 81.6 3.177 81.625 3.523 ;
      RECT 81.595 3.152 81.6 3.502 ;
      RECT 81.585 3.13 81.595 3.493 ;
      RECT 81.58 3.101 81.585 3.483 ;
      RECT 81.54 3.027 81.58 3.455 ;
      RECT 81.52 2.928 81.54 3.42 ;
      RECT 81.505 2.864 81.52 3.403 ;
      RECT 81.475 2.788 81.505 3.375 ;
      RECT 81.455 2.703 81.475 3.348 ;
      RECT 81.415 2.599 81.455 3.255 ;
      RECT 81.41 2.52 81.415 3.163 ;
      RECT 81.405 2.503 81.41 3.14 ;
      RECT 81.4 2.225 81.405 3.12 ;
      RECT 81.37 2.225 81.4 3.058 ;
      RECT 81.365 2.225 81.37 2.99 ;
      RECT 81.355 2.225 81.365 2.955 ;
      RECT 81.345 2.225 81.355 2.92 ;
      RECT 81.28 2.225 81.345 2.775 ;
      RECT 81.275 2.225 81.28 2.645 ;
      RECT 81.245 2.225 81.275 2.578 ;
      RECT 81.24 2.225 81.245 2.503 ;
      RECT 85.575 2.16 85.835 2.42 ;
      RECT 85.57 2.16 85.835 2.368 ;
      RECT 85.565 2.16 85.835 2.338 ;
      RECT 85.54 2.03 85.82 2.31 ;
      RECT 74.055 6.655 74.405 7.005 ;
      RECT 85.3 6.61 85.65 6.96 ;
      RECT 74.055 6.685 85.65 6.885 ;
      RECT 84.58 3.71 84.86 3.99 ;
      RECT 84.62 3.665 84.885 3.925 ;
      RECT 84.61 3.7 84.885 3.925 ;
      RECT 84.615 3.685 84.86 3.99 ;
      RECT 84.62 3.662 84.83 3.99 ;
      RECT 84.62 3.66 84.815 3.99 ;
      RECT 84.66 3.65 84.815 3.99 ;
      RECT 84.63 3.655 84.815 3.99 ;
      RECT 84.66 3.647 84.76 3.99 ;
      RECT 84.685 3.64 84.76 3.99 ;
      RECT 84.665 3.642 84.76 3.99 ;
      RECT 83.995 3.155 84.255 3.415 ;
      RECT 84.045 3.147 84.235 3.415 ;
      RECT 84.05 3.067 84.235 3.415 ;
      RECT 84.17 2.455 84.235 3.415 ;
      RECT 84.075 2.852 84.235 3.415 ;
      RECT 84.15 2.54 84.235 3.415 ;
      RECT 84.185 2.165 84.321 2.893 ;
      RECT 84.13 2.662 84.321 2.893 ;
      RECT 84.145 2.602 84.235 3.415 ;
      RECT 84.185 2.165 84.345 2.558 ;
      RECT 84.185 2.165 84.355 2.455 ;
      RECT 84.175 2.165 84.435 2.425 ;
      RECT 83.58 3.71 83.86 3.99 ;
      RECT 83.6 3.67 83.86 3.99 ;
      RECT 83.24 3.625 83.345 3.885 ;
      RECT 83.095 2.115 83.185 2.375 ;
      RECT 83.635 3.18 83.64 3.22 ;
      RECT 83.63 3.17 83.635 3.305 ;
      RECT 83.625 3.16 83.63 3.398 ;
      RECT 83.615 3.14 83.625 3.454 ;
      RECT 83.535 3.068 83.615 3.534 ;
      RECT 83.57 3.712 83.58 3.937 ;
      RECT 83.565 3.709 83.57 3.932 ;
      RECT 83.55 3.706 83.565 3.925 ;
      RECT 83.515 3.7 83.55 3.907 ;
      RECT 83.53 3.003 83.535 3.608 ;
      RECT 83.51 2.954 83.53 3.623 ;
      RECT 83.5 3.687 83.515 3.89 ;
      RECT 83.505 2.896 83.51 3.638 ;
      RECT 83.5 2.874 83.505 3.648 ;
      RECT 83.465 2.784 83.5 3.885 ;
      RECT 83.45 2.662 83.465 3.885 ;
      RECT 83.445 2.615 83.45 3.885 ;
      RECT 83.42 2.54 83.445 3.885 ;
      RECT 83.405 2.455 83.42 3.885 ;
      RECT 83.4 2.402 83.405 3.885 ;
      RECT 83.395 2.382 83.4 3.885 ;
      RECT 83.39 2.357 83.395 3.119 ;
      RECT 83.375 3.317 83.395 3.885 ;
      RECT 83.385 2.335 83.39 3.096 ;
      RECT 83.375 2.287 83.385 3.061 ;
      RECT 83.37 2.25 83.375 3.027 ;
      RECT 83.37 3.397 83.375 3.885 ;
      RECT 83.355 2.227 83.37 2.982 ;
      RECT 83.35 3.495 83.37 3.885 ;
      RECT 83.3 2.115 83.355 2.824 ;
      RECT 83.345 3.617 83.35 3.885 ;
      RECT 83.285 2.115 83.3 2.663 ;
      RECT 83.28 2.115 83.285 2.615 ;
      RECT 83.275 2.115 83.28 2.603 ;
      RECT 83.23 2.115 83.275 2.54 ;
      RECT 83.205 2.115 83.23 2.458 ;
      RECT 83.19 2.115 83.205 2.41 ;
      RECT 83.185 2.115 83.19 2.38 ;
      RECT 82.51 3.565 82.555 3.825 ;
      RECT 82.415 2.1 82.56 2.36 ;
      RECT 82.92 2.722 82.93 2.813 ;
      RECT 82.905 2.66 82.92 2.869 ;
      RECT 82.9 2.607 82.905 2.915 ;
      RECT 82.85 2.554 82.9 3.041 ;
      RECT 82.845 2.509 82.85 3.188 ;
      RECT 82.835 2.497 82.845 3.23 ;
      RECT 82.8 2.461 82.835 3.335 ;
      RECT 82.795 2.429 82.8 3.441 ;
      RECT 82.78 2.411 82.795 3.486 ;
      RECT 82.775 2.394 82.78 2.72 ;
      RECT 82.77 2.775 82.78 3.543 ;
      RECT 82.765 2.38 82.775 2.693 ;
      RECT 82.76 2.83 82.77 3.825 ;
      RECT 82.755 2.366 82.765 2.678 ;
      RECT 82.755 2.88 82.76 3.825 ;
      RECT 82.74 2.343 82.755 2.658 ;
      RECT 82.72 3.002 82.755 3.825 ;
      RECT 82.735 2.325 82.74 2.64 ;
      RECT 82.73 2.317 82.735 2.63 ;
      RECT 82.7 2.285 82.73 2.594 ;
      RECT 82.71 3.13 82.72 3.825 ;
      RECT 82.705 3.157 82.71 3.825 ;
      RECT 82.7 3.207 82.705 3.825 ;
      RECT 82.69 2.251 82.7 2.559 ;
      RECT 82.65 3.275 82.7 3.825 ;
      RECT 82.675 2.228 82.69 2.535 ;
      RECT 82.65 2.1 82.675 2.498 ;
      RECT 82.645 2.1 82.65 2.47 ;
      RECT 82.615 3.375 82.65 3.825 ;
      RECT 82.64 2.1 82.645 2.463 ;
      RECT 82.635 2.1 82.64 2.453 ;
      RECT 82.62 2.1 82.635 2.438 ;
      RECT 82.605 2.1 82.62 2.41 ;
      RECT 82.57 3.48 82.615 3.825 ;
      RECT 82.59 2.1 82.605 2.383 ;
      RECT 82.56 2.1 82.59 2.368 ;
      RECT 82.555 3.552 82.57 3.825 ;
      RECT 82.48 2.635 82.52 2.895 ;
      RECT 82.255 2.582 82.26 2.84 ;
      RECT 78.21 2.06 78.47 2.32 ;
      RECT 78.21 2.085 78.485 2.3 ;
      RECT 80.6 1.91 80.605 2.055 ;
      RECT 82.47 2.63 82.48 2.895 ;
      RECT 82.45 2.622 82.47 2.895 ;
      RECT 82.432 2.618 82.45 2.895 ;
      RECT 82.346 2.607 82.432 2.895 ;
      RECT 82.26 2.59 82.346 2.895 ;
      RECT 82.205 2.577 82.255 2.825 ;
      RECT 82.171 2.569 82.205 2.8 ;
      RECT 82.085 2.558 82.171 2.765 ;
      RECT 82.05 2.535 82.085 2.73 ;
      RECT 82.04 2.497 82.05 2.716 ;
      RECT 82.035 2.47 82.04 2.712 ;
      RECT 82.03 2.457 82.035 2.709 ;
      RECT 82.02 2.437 82.03 2.705 ;
      RECT 82.015 2.412 82.02 2.701 ;
      RECT 81.99 2.367 82.015 2.695 ;
      RECT 81.98 2.308 81.99 2.687 ;
      RECT 81.97 2.276 81.98 2.678 ;
      RECT 81.95 2.228 81.97 2.658 ;
      RECT 81.945 2.188 81.95 2.628 ;
      RECT 81.93 2.162 81.945 2.602 ;
      RECT 81.925 2.14 81.93 2.578 ;
      RECT 81.91 2.112 81.925 2.554 ;
      RECT 81.895 2.085 81.91 2.518 ;
      RECT 81.88 2.062 81.895 2.48 ;
      RECT 81.875 2.052 81.88 2.455 ;
      RECT 81.865 2.045 81.875 2.438 ;
      RECT 81.85 2.032 81.865 2.408 ;
      RECT 81.845 2.022 81.85 2.383 ;
      RECT 81.84 2.017 81.845 2.37 ;
      RECT 81.83 2.01 81.84 2.35 ;
      RECT 81.825 2.003 81.83 2.335 ;
      RECT 81.8 1.996 81.825 2.293 ;
      RECT 81.785 1.986 81.8 2.243 ;
      RECT 81.775 1.981 81.785 2.213 ;
      RECT 81.765 1.977 81.775 2.188 ;
      RECT 81.75 1.974 81.765 2.178 ;
      RECT 81.7 1.971 81.75 2.163 ;
      RECT 81.68 1.969 81.7 2.148 ;
      RECT 81.631 1.967 81.68 2.143 ;
      RECT 81.545 1.963 81.631 2.138 ;
      RECT 81.506 1.96 81.545 2.134 ;
      RECT 81.42 1.956 81.506 2.129 ;
      RECT 81.37 1.953 81.42 2.123 ;
      RECT 81.321 1.95 81.37 2.118 ;
      RECT 81.235 1.947 81.321 2.113 ;
      RECT 81.231 1.945 81.235 2.11 ;
      RECT 81.145 1.942 81.231 2.105 ;
      RECT 81.096 1.938 81.145 2.098 ;
      RECT 81.01 1.935 81.096 2.093 ;
      RECT 80.986 1.932 81.01 2.089 ;
      RECT 80.9 1.93 80.986 2.084 ;
      RECT 80.835 1.926 80.9 2.077 ;
      RECT 80.832 1.925 80.835 2.074 ;
      RECT 80.746 1.922 80.832 2.071 ;
      RECT 80.66 1.916 80.746 2.064 ;
      RECT 80.63 1.912 80.66 2.06 ;
      RECT 80.605 1.91 80.63 2.058 ;
      RECT 80.55 1.907 80.6 2.055 ;
      RECT 80.47 1.906 80.55 2.055 ;
      RECT 80.415 1.908 80.47 2.058 ;
      RECT 80.4 1.909 80.415 2.062 ;
      RECT 80.345 1.917 80.4 2.072 ;
      RECT 80.315 1.925 80.345 2.085 ;
      RECT 80.296 1.926 80.315 2.091 ;
      RECT 80.21 1.929 80.296 2.096 ;
      RECT 80.14 1.934 80.21 2.105 ;
      RECT 80.121 1.937 80.14 2.111 ;
      RECT 80.035 1.941 80.121 2.116 ;
      RECT 79.995 1.945 80.035 2.123 ;
      RECT 79.986 1.947 79.995 2.126 ;
      RECT 79.9 1.951 79.986 2.131 ;
      RECT 79.897 1.954 79.9 2.135 ;
      RECT 79.811 1.957 79.897 2.139 ;
      RECT 79.725 1.963 79.811 2.147 ;
      RECT 79.701 1.967 79.725 2.151 ;
      RECT 79.615 1.971 79.701 2.156 ;
      RECT 79.57 1.976 79.615 2.163 ;
      RECT 79.49 1.981 79.57 2.17 ;
      RECT 79.41 1.987 79.49 2.185 ;
      RECT 79.385 1.991 79.41 2.198 ;
      RECT 79.32 1.994 79.385 2.21 ;
      RECT 79.265 1.999 79.32 2.225 ;
      RECT 79.235 2.002 79.265 2.243 ;
      RECT 79.225 2.004 79.235 2.256 ;
      RECT 79.165 2.019 79.225 2.266 ;
      RECT 79.15 2.036 79.165 2.275 ;
      RECT 79.145 2.045 79.15 2.275 ;
      RECT 79.135 2.055 79.145 2.275 ;
      RECT 79.125 2.072 79.135 2.275 ;
      RECT 79.105 2.082 79.125 2.276 ;
      RECT 79.06 2.092 79.105 2.277 ;
      RECT 79.025 2.101 79.06 2.279 ;
      RECT 78.96 2.106 79.025 2.281 ;
      RECT 78.88 2.107 78.96 2.284 ;
      RECT 78.876 2.105 78.88 2.285 ;
      RECT 78.79 2.102 78.876 2.287 ;
      RECT 78.743 2.099 78.79 2.289 ;
      RECT 78.657 2.095 78.743 2.292 ;
      RECT 78.571 2.091 78.657 2.295 ;
      RECT 78.485 2.087 78.571 2.299 ;
      RECT 80.42 3.15 80.7 3.43 ;
      RECT 80.46 3.13 80.72 3.39 ;
      RECT 80.45 3.14 80.72 3.39 ;
      RECT 80.46 3.067 80.675 3.43 ;
      RECT 80.515 2.99 80.67 3.43 ;
      RECT 80.52 2.775 80.67 3.43 ;
      RECT 80.51 2.577 80.66 2.828 ;
      RECT 80.5 2.577 80.66 2.695 ;
      RECT 80.495 2.455 80.655 2.598 ;
      RECT 80.48 2.455 80.655 2.503 ;
      RECT 80.475 2.165 80.65 2.48 ;
      RECT 80.46 2.165 80.65 2.45 ;
      RECT 80.42 2.165 80.68 2.425 ;
      RECT 80.33 3.635 80.41 3.895 ;
      RECT 79.735 2.355 79.74 2.62 ;
      RECT 79.615 2.355 79.74 2.615 ;
      RECT 80.29 3.6 80.33 3.895 ;
      RECT 80.245 3.522 80.29 3.895 ;
      RECT 80.225 3.45 80.245 3.895 ;
      RECT 80.215 3.402 80.225 3.895 ;
      RECT 80.18 3.335 80.215 3.895 ;
      RECT 80.15 3.235 80.18 3.895 ;
      RECT 80.13 3.16 80.15 3.695 ;
      RECT 80.12 3.11 80.13 3.65 ;
      RECT 80.115 3.087 80.12 3.623 ;
      RECT 80.11 3.072 80.115 3.61 ;
      RECT 80.105 3.057 80.11 3.588 ;
      RECT 80.1 3.042 80.105 3.57 ;
      RECT 80.075 2.997 80.1 3.525 ;
      RECT 80.065 2.945 80.075 3.468 ;
      RECT 80.055 2.915 80.065 3.435 ;
      RECT 80.045 2.88 80.055 3.403 ;
      RECT 80.01 2.812 80.045 3.335 ;
      RECT 80.005 2.751 80.01 3.27 ;
      RECT 79.995 2.739 80.005 3.25 ;
      RECT 79.99 2.727 79.995 3.23 ;
      RECT 79.985 2.719 79.99 3.218 ;
      RECT 79.98 2.711 79.985 3.198 ;
      RECT 79.97 2.699 79.98 3.17 ;
      RECT 79.96 2.683 79.97 3.14 ;
      RECT 79.935 2.655 79.96 3.078 ;
      RECT 79.925 2.626 79.935 3.023 ;
      RECT 79.91 2.605 79.925 2.983 ;
      RECT 79.905 2.589 79.91 2.955 ;
      RECT 79.9 2.577 79.905 2.945 ;
      RECT 79.895 2.572 79.9 2.918 ;
      RECT 79.89 2.565 79.895 2.905 ;
      RECT 79.875 2.548 79.89 2.878 ;
      RECT 79.865 2.355 79.875 2.838 ;
      RECT 79.855 2.355 79.865 2.805 ;
      RECT 79.845 2.355 79.855 2.78 ;
      RECT 79.775 2.355 79.845 2.715 ;
      RECT 79.765 2.355 79.775 2.663 ;
      RECT 79.75 2.355 79.765 2.645 ;
      RECT 79.74 2.355 79.75 2.63 ;
      RECT 79.57 3.225 79.83 3.485 ;
      RECT 78.105 3.26 78.11 3.467 ;
      RECT 77.74 3.15 77.815 3.465 ;
      RECT 77.555 3.205 77.71 3.465 ;
      RECT 77.74 3.15 77.845 3.43 ;
      RECT 79.555 3.322 79.57 3.483 ;
      RECT 79.53 3.33 79.555 3.488 ;
      RECT 79.505 3.337 79.53 3.493 ;
      RECT 79.442 3.348 79.505 3.502 ;
      RECT 79.356 3.367 79.442 3.519 ;
      RECT 79.27 3.389 79.356 3.538 ;
      RECT 79.255 3.402 79.27 3.549 ;
      RECT 79.215 3.41 79.255 3.556 ;
      RECT 79.195 3.415 79.215 3.563 ;
      RECT 79.157 3.416 79.195 3.566 ;
      RECT 79.071 3.419 79.157 3.567 ;
      RECT 78.985 3.423 79.071 3.568 ;
      RECT 78.936 3.425 78.985 3.57 ;
      RECT 78.85 3.425 78.936 3.572 ;
      RECT 78.81 3.42 78.85 3.574 ;
      RECT 78.8 3.414 78.81 3.575 ;
      RECT 78.76 3.409 78.8 3.572 ;
      RECT 78.75 3.402 78.76 3.568 ;
      RECT 78.735 3.398 78.75 3.566 ;
      RECT 78.718 3.394 78.735 3.564 ;
      RECT 78.632 3.384 78.718 3.556 ;
      RECT 78.546 3.366 78.632 3.542 ;
      RECT 78.46 3.349 78.546 3.528 ;
      RECT 78.435 3.337 78.46 3.519 ;
      RECT 78.365 3.327 78.435 3.512 ;
      RECT 78.32 3.315 78.365 3.503 ;
      RECT 78.26 3.302 78.32 3.495 ;
      RECT 78.255 3.294 78.26 3.49 ;
      RECT 78.22 3.289 78.255 3.488 ;
      RECT 78.165 3.28 78.22 3.481 ;
      RECT 78.125 3.269 78.165 3.473 ;
      RECT 78.11 3.262 78.125 3.469 ;
      RECT 78.09 3.255 78.105 3.466 ;
      RECT 78.075 3.245 78.09 3.464 ;
      RECT 78.06 3.232 78.075 3.461 ;
      RECT 78.035 3.215 78.06 3.457 ;
      RECT 78.02 3.197 78.035 3.454 ;
      RECT 77.995 3.15 78.02 3.452 ;
      RECT 77.971 3.15 77.995 3.449 ;
      RECT 77.885 3.15 77.971 3.441 ;
      RECT 77.845 3.15 77.885 3.433 ;
      RECT 77.71 3.197 77.74 3.465 ;
      RECT 79.39 2.78 79.65 3.04 ;
      RECT 79.35 2.78 79.65 2.918 ;
      RECT 79.315 2.78 79.65 2.903 ;
      RECT 79.26 2.78 79.65 2.883 ;
      RECT 79.18 2.59 79.46 2.87 ;
      RECT 79.18 2.772 79.53 2.87 ;
      RECT 79.18 2.715 79.515 2.87 ;
      RECT 79.18 2.662 79.465 2.87 ;
      RECT 77.01 2.59 77.205 3.375 ;
      RECT 77.09 1.205 77.205 3.375 ;
      RECT 76.945 3.115 77.005 3.375 ;
      RECT 78.315 2.635 78.575 2.895 ;
      RECT 77 2.59 77.205 2.87 ;
      RECT 78.31 2.645 78.575 2.83 ;
      RECT 78.025 2.62 78.035 2.77 ;
      RECT 77.26 1.205 77.34 1.55 ;
      RECT 76.995 1.205 77.205 1.55 ;
      RECT 78.3 2.645 78.31 2.829 ;
      RECT 78.29 2.644 78.3 2.826 ;
      RECT 78.281 2.643 78.29 2.824 ;
      RECT 78.195 2.639 78.281 2.814 ;
      RECT 78.121 2.631 78.195 2.796 ;
      RECT 78.035 2.624 78.121 2.779 ;
      RECT 77.975 2.62 78.025 2.769 ;
      RECT 77.94 2.619 77.975 2.766 ;
      RECT 77.885 2.619 77.94 2.768 ;
      RECT 77.85 2.619 77.885 2.772 ;
      RECT 77.764 2.618 77.85 2.779 ;
      RECT 77.678 2.617 77.764 2.789 ;
      RECT 77.592 2.616 77.678 2.8 ;
      RECT 77.506 2.616 77.592 2.81 ;
      RECT 77.42 2.615 77.506 2.82 ;
      RECT 77.385 2.615 77.42 2.86 ;
      RECT 77.38 2.615 77.385 2.903 ;
      RECT 77.355 2.615 77.38 2.92 ;
      RECT 77.28 2.615 77.355 2.935 ;
      RECT 77.26 2.59 77.28 2.948 ;
      RECT 77.255 1.205 77.26 2.958 ;
      RECT 77.23 1.205 77.255 3 ;
      RECT 77.205 1.205 77.23 3.078 ;
      RECT 77.005 2.997 77.01 3.375 ;
      RECT 76.34 2.949 76.355 3.405 ;
      RECT 76.335 3.021 76.441 3.403 ;
      RECT 76.355 2.115 76.49 3.401 ;
      RECT 76.34 2.965 76.495 3.4 ;
      RECT 76.34 3.015 76.5 3.398 ;
      RECT 76.325 3.08 76.5 3.397 ;
      RECT 76.335 3.072 76.505 3.394 ;
      RECT 76.315 3.12 76.505 3.389 ;
      RECT 76.315 3.12 76.52 3.386 ;
      RECT 76.31 3.12 76.52 3.383 ;
      RECT 76.285 3.12 76.545 3.38 ;
      RECT 76.355 2.115 76.515 2.768 ;
      RECT 76.35 2.115 76.515 2.74 ;
      RECT 76.345 2.115 76.515 2.568 ;
      RECT 76.345 2.115 76.535 2.508 ;
      RECT 76.3 2.115 76.56 2.375 ;
      RECT 75.78 2.59 76.06 2.87 ;
      RECT 75.77 2.605 76.06 2.865 ;
      RECT 75.725 2.667 76.06 2.863 ;
      RECT 75.8 2.582 75.965 2.87 ;
      RECT 75.8 2.567 75.921 2.87 ;
      RECT 75.835 2.56 75.921 2.87 ;
      RECT 75.3 3.71 75.58 3.99 ;
      RECT 75.26 3.672 75.555 3.783 ;
      RECT 75.245 3.622 75.535 3.678 ;
      RECT 75.19 3.385 75.45 3.645 ;
      RECT 75.19 3.587 75.53 3.645 ;
      RECT 75.19 3.527 75.525 3.645 ;
      RECT 75.19 3.477 75.505 3.645 ;
      RECT 75.19 3.457 75.5 3.645 ;
      RECT 75.19 3.435 75.495 3.645 ;
      RECT 75.19 3.42 75.465 3.645 ;
      RECT 70.92 6.225 71.24 6.545 ;
      RECT 70.95 5.695 71.12 6.545 ;
      RECT 70.95 5.695 71.125 6.045 ;
      RECT 70.95 5.695 71.925 5.87 ;
      RECT 71.75 1.965 71.925 5.87 ;
      RECT 71.695 1.965 72.045 2.315 ;
      RECT 71.72 6.655 72.045 6.98 ;
      RECT 70.605 6.745 72.045 6.915 ;
      RECT 70.605 2.395 70.765 6.915 ;
      RECT 70.92 2.365 71.24 2.685 ;
      RECT 70.605 2.395 71.24 2.565 ;
      RECT 69.865 5.84 70.215 6.19 ;
      RECT 69.94 2.705 70.115 6.19 ;
      RECT 69.875 2.705 70.225 3.055 ;
      RECT 69.275 1.14 69.65 1.51 ;
      RECT 61.195 0.96 61.57 1.33 ;
      RECT 59.76 0.96 60.135 1.33 ;
      RECT 59.76 1.08 69.58 1.25 ;
      RECT 63.88 4.36 69.56 4.53 ;
      RECT 69.39 3.425 69.56 4.53 ;
      RECT 63.69 3.6 63.715 4.53 ;
      RECT 63.945 3.71 63.975 3.99 ;
      RECT 63.65 3.6 63.715 3.86 ;
      RECT 69.3 3.43 69.65 3.78 ;
      RECT 63.48 2.225 63.515 2.485 ;
      RECT 63.255 2.225 63.315 2.485 ;
      RECT 63.935 3.69 63.945 3.99 ;
      RECT 63.93 3.65 63.935 3.99 ;
      RECT 63.915 3.605 63.93 3.99 ;
      RECT 63.91 3.57 63.915 3.99 ;
      RECT 63.905 3.55 63.91 3.99 ;
      RECT 63.88 3.487 63.905 3.99 ;
      RECT 63.875 3.425 63.88 4.53 ;
      RECT 63.855 3.375 63.875 4.53 ;
      RECT 63.845 3.305 63.855 4.53 ;
      RECT 63.8 3.245 63.845 4.53 ;
      RECT 63.715 3.206 63.8 4.53 ;
      RECT 63.71 3.197 63.715 3.57 ;
      RECT 63.7 3.196 63.71 3.553 ;
      RECT 63.675 3.177 63.7 3.523 ;
      RECT 63.67 3.152 63.675 3.502 ;
      RECT 63.66 3.13 63.67 3.493 ;
      RECT 63.655 3.101 63.66 3.483 ;
      RECT 63.615 3.027 63.655 3.455 ;
      RECT 63.595 2.928 63.615 3.42 ;
      RECT 63.58 2.864 63.595 3.403 ;
      RECT 63.55 2.788 63.58 3.375 ;
      RECT 63.53 2.703 63.55 3.348 ;
      RECT 63.49 2.599 63.53 3.255 ;
      RECT 63.485 2.52 63.49 3.163 ;
      RECT 63.48 2.503 63.485 3.14 ;
      RECT 63.475 2.225 63.48 3.12 ;
      RECT 63.445 2.225 63.475 3.058 ;
      RECT 63.44 2.225 63.445 2.99 ;
      RECT 63.43 2.225 63.44 2.955 ;
      RECT 63.42 2.225 63.43 2.92 ;
      RECT 63.355 2.225 63.42 2.775 ;
      RECT 63.35 2.225 63.355 2.645 ;
      RECT 63.32 2.225 63.35 2.578 ;
      RECT 63.315 2.225 63.32 2.503 ;
      RECT 67.65 2.16 67.91 2.42 ;
      RECT 67.645 2.16 67.91 2.368 ;
      RECT 67.64 2.16 67.91 2.338 ;
      RECT 67.615 2.03 67.895 2.31 ;
      RECT 56.13 6.655 56.48 7.005 ;
      RECT 67.095 6.61 67.445 6.96 ;
      RECT 56.13 6.685 67.445 6.885 ;
      RECT 66.655 3.71 66.935 3.99 ;
      RECT 66.695 3.665 66.96 3.925 ;
      RECT 66.685 3.7 66.96 3.925 ;
      RECT 66.69 3.685 66.935 3.99 ;
      RECT 66.695 3.662 66.905 3.99 ;
      RECT 66.695 3.66 66.89 3.99 ;
      RECT 66.735 3.65 66.89 3.99 ;
      RECT 66.705 3.655 66.89 3.99 ;
      RECT 66.735 3.647 66.835 3.99 ;
      RECT 66.76 3.64 66.835 3.99 ;
      RECT 66.74 3.642 66.835 3.99 ;
      RECT 66.07 3.155 66.33 3.415 ;
      RECT 66.12 3.147 66.31 3.415 ;
      RECT 66.125 3.067 66.31 3.415 ;
      RECT 66.245 2.455 66.31 3.415 ;
      RECT 66.15 2.852 66.31 3.415 ;
      RECT 66.225 2.54 66.31 3.415 ;
      RECT 66.26 2.165 66.396 2.893 ;
      RECT 66.205 2.662 66.396 2.893 ;
      RECT 66.22 2.602 66.31 3.415 ;
      RECT 66.26 2.165 66.42 2.558 ;
      RECT 66.26 2.165 66.43 2.455 ;
      RECT 66.25 2.165 66.51 2.425 ;
      RECT 65.655 3.71 65.935 3.99 ;
      RECT 65.675 3.67 65.935 3.99 ;
      RECT 65.315 3.625 65.42 3.885 ;
      RECT 65.17 2.115 65.26 2.375 ;
      RECT 65.71 3.18 65.715 3.22 ;
      RECT 65.705 3.17 65.71 3.305 ;
      RECT 65.7 3.16 65.705 3.398 ;
      RECT 65.69 3.14 65.7 3.454 ;
      RECT 65.61 3.068 65.69 3.534 ;
      RECT 65.645 3.712 65.655 3.937 ;
      RECT 65.64 3.709 65.645 3.932 ;
      RECT 65.625 3.706 65.64 3.925 ;
      RECT 65.59 3.7 65.625 3.907 ;
      RECT 65.605 3.003 65.61 3.608 ;
      RECT 65.585 2.954 65.605 3.623 ;
      RECT 65.575 3.687 65.59 3.89 ;
      RECT 65.58 2.896 65.585 3.638 ;
      RECT 65.575 2.874 65.58 3.648 ;
      RECT 65.54 2.784 65.575 3.885 ;
      RECT 65.525 2.662 65.54 3.885 ;
      RECT 65.52 2.615 65.525 3.885 ;
      RECT 65.495 2.54 65.52 3.885 ;
      RECT 65.48 2.455 65.495 3.885 ;
      RECT 65.475 2.402 65.48 3.885 ;
      RECT 65.47 2.382 65.475 3.885 ;
      RECT 65.465 2.357 65.47 3.119 ;
      RECT 65.45 3.317 65.47 3.885 ;
      RECT 65.46 2.335 65.465 3.096 ;
      RECT 65.45 2.287 65.46 3.061 ;
      RECT 65.445 2.25 65.45 3.027 ;
      RECT 65.445 3.397 65.45 3.885 ;
      RECT 65.43 2.227 65.445 2.982 ;
      RECT 65.425 3.495 65.445 3.885 ;
      RECT 65.375 2.115 65.43 2.824 ;
      RECT 65.42 3.617 65.425 3.885 ;
      RECT 65.36 2.115 65.375 2.663 ;
      RECT 65.355 2.115 65.36 2.615 ;
      RECT 65.35 2.115 65.355 2.603 ;
      RECT 65.305 2.115 65.35 2.54 ;
      RECT 65.28 2.115 65.305 2.458 ;
      RECT 65.265 2.115 65.28 2.41 ;
      RECT 65.26 2.115 65.265 2.38 ;
      RECT 64.585 3.565 64.63 3.825 ;
      RECT 64.49 2.1 64.635 2.36 ;
      RECT 64.995 2.722 65.005 2.813 ;
      RECT 64.98 2.66 64.995 2.869 ;
      RECT 64.975 2.607 64.98 2.915 ;
      RECT 64.925 2.554 64.975 3.041 ;
      RECT 64.92 2.509 64.925 3.188 ;
      RECT 64.91 2.497 64.92 3.23 ;
      RECT 64.875 2.461 64.91 3.335 ;
      RECT 64.87 2.429 64.875 3.441 ;
      RECT 64.855 2.411 64.87 3.486 ;
      RECT 64.85 2.394 64.855 2.72 ;
      RECT 64.845 2.775 64.855 3.543 ;
      RECT 64.84 2.38 64.85 2.693 ;
      RECT 64.835 2.83 64.845 3.825 ;
      RECT 64.83 2.366 64.84 2.678 ;
      RECT 64.83 2.88 64.835 3.825 ;
      RECT 64.815 2.343 64.83 2.658 ;
      RECT 64.795 3.002 64.83 3.825 ;
      RECT 64.81 2.325 64.815 2.64 ;
      RECT 64.805 2.317 64.81 2.63 ;
      RECT 64.775 2.285 64.805 2.594 ;
      RECT 64.785 3.13 64.795 3.825 ;
      RECT 64.78 3.157 64.785 3.825 ;
      RECT 64.775 3.207 64.78 3.825 ;
      RECT 64.765 2.251 64.775 2.559 ;
      RECT 64.725 3.275 64.775 3.825 ;
      RECT 64.75 2.228 64.765 2.535 ;
      RECT 64.725 2.1 64.75 2.498 ;
      RECT 64.72 2.1 64.725 2.47 ;
      RECT 64.69 3.375 64.725 3.825 ;
      RECT 64.715 2.1 64.72 2.463 ;
      RECT 64.71 2.1 64.715 2.453 ;
      RECT 64.695 2.1 64.71 2.438 ;
      RECT 64.68 2.1 64.695 2.41 ;
      RECT 64.645 3.48 64.69 3.825 ;
      RECT 64.665 2.1 64.68 2.383 ;
      RECT 64.635 2.1 64.665 2.368 ;
      RECT 64.63 3.552 64.645 3.825 ;
      RECT 64.555 2.635 64.595 2.895 ;
      RECT 64.33 2.582 64.335 2.84 ;
      RECT 60.285 2.06 60.545 2.32 ;
      RECT 60.285 2.085 60.56 2.3 ;
      RECT 62.675 1.91 62.68 2.055 ;
      RECT 64.545 2.63 64.555 2.895 ;
      RECT 64.525 2.622 64.545 2.895 ;
      RECT 64.507 2.618 64.525 2.895 ;
      RECT 64.421 2.607 64.507 2.895 ;
      RECT 64.335 2.59 64.421 2.895 ;
      RECT 64.28 2.577 64.33 2.825 ;
      RECT 64.246 2.569 64.28 2.8 ;
      RECT 64.16 2.558 64.246 2.765 ;
      RECT 64.125 2.535 64.16 2.73 ;
      RECT 64.115 2.497 64.125 2.716 ;
      RECT 64.11 2.47 64.115 2.712 ;
      RECT 64.105 2.457 64.11 2.709 ;
      RECT 64.095 2.437 64.105 2.705 ;
      RECT 64.09 2.412 64.095 2.701 ;
      RECT 64.065 2.367 64.09 2.695 ;
      RECT 64.055 2.308 64.065 2.687 ;
      RECT 64.045 2.276 64.055 2.678 ;
      RECT 64.025 2.228 64.045 2.658 ;
      RECT 64.02 2.188 64.025 2.628 ;
      RECT 64.005 2.162 64.02 2.602 ;
      RECT 64 2.14 64.005 2.578 ;
      RECT 63.985 2.112 64 2.554 ;
      RECT 63.97 2.085 63.985 2.518 ;
      RECT 63.955 2.062 63.97 2.48 ;
      RECT 63.95 2.052 63.955 2.455 ;
      RECT 63.94 2.045 63.95 2.438 ;
      RECT 63.925 2.032 63.94 2.408 ;
      RECT 63.92 2.022 63.925 2.383 ;
      RECT 63.915 2.017 63.92 2.37 ;
      RECT 63.905 2.01 63.915 2.35 ;
      RECT 63.9 2.003 63.905 2.335 ;
      RECT 63.875 1.996 63.9 2.293 ;
      RECT 63.86 1.986 63.875 2.243 ;
      RECT 63.85 1.981 63.86 2.213 ;
      RECT 63.84 1.977 63.85 2.188 ;
      RECT 63.825 1.974 63.84 2.178 ;
      RECT 63.775 1.971 63.825 2.163 ;
      RECT 63.755 1.969 63.775 2.148 ;
      RECT 63.706 1.967 63.755 2.143 ;
      RECT 63.62 1.963 63.706 2.138 ;
      RECT 63.581 1.96 63.62 2.134 ;
      RECT 63.495 1.956 63.581 2.129 ;
      RECT 63.445 1.953 63.495 2.123 ;
      RECT 63.396 1.95 63.445 2.118 ;
      RECT 63.31 1.947 63.396 2.113 ;
      RECT 63.306 1.945 63.31 2.11 ;
      RECT 63.22 1.942 63.306 2.105 ;
      RECT 63.171 1.938 63.22 2.098 ;
      RECT 63.085 1.935 63.171 2.093 ;
      RECT 63.061 1.932 63.085 2.089 ;
      RECT 62.975 1.93 63.061 2.084 ;
      RECT 62.91 1.926 62.975 2.077 ;
      RECT 62.907 1.925 62.91 2.074 ;
      RECT 62.821 1.922 62.907 2.071 ;
      RECT 62.735 1.916 62.821 2.064 ;
      RECT 62.705 1.912 62.735 2.06 ;
      RECT 62.68 1.91 62.705 2.058 ;
      RECT 62.625 1.907 62.675 2.055 ;
      RECT 62.545 1.906 62.625 2.055 ;
      RECT 62.49 1.908 62.545 2.058 ;
      RECT 62.475 1.909 62.49 2.062 ;
      RECT 62.42 1.917 62.475 2.072 ;
      RECT 62.39 1.925 62.42 2.085 ;
      RECT 62.371 1.926 62.39 2.091 ;
      RECT 62.285 1.929 62.371 2.096 ;
      RECT 62.215 1.934 62.285 2.105 ;
      RECT 62.196 1.937 62.215 2.111 ;
      RECT 62.11 1.941 62.196 2.116 ;
      RECT 62.07 1.945 62.11 2.123 ;
      RECT 62.061 1.947 62.07 2.126 ;
      RECT 61.975 1.951 62.061 2.131 ;
      RECT 61.972 1.954 61.975 2.135 ;
      RECT 61.886 1.957 61.972 2.139 ;
      RECT 61.8 1.963 61.886 2.147 ;
      RECT 61.776 1.967 61.8 2.151 ;
      RECT 61.69 1.971 61.776 2.156 ;
      RECT 61.645 1.976 61.69 2.163 ;
      RECT 61.565 1.981 61.645 2.17 ;
      RECT 61.485 1.987 61.565 2.185 ;
      RECT 61.46 1.991 61.485 2.198 ;
      RECT 61.395 1.994 61.46 2.21 ;
      RECT 61.34 1.999 61.395 2.225 ;
      RECT 61.31 2.002 61.34 2.243 ;
      RECT 61.3 2.004 61.31 2.256 ;
      RECT 61.24 2.019 61.3 2.266 ;
      RECT 61.225 2.036 61.24 2.275 ;
      RECT 61.22 2.045 61.225 2.275 ;
      RECT 61.21 2.055 61.22 2.275 ;
      RECT 61.2 2.072 61.21 2.275 ;
      RECT 61.18 2.082 61.2 2.276 ;
      RECT 61.135 2.092 61.18 2.277 ;
      RECT 61.1 2.101 61.135 2.279 ;
      RECT 61.035 2.106 61.1 2.281 ;
      RECT 60.955 2.107 61.035 2.284 ;
      RECT 60.951 2.105 60.955 2.285 ;
      RECT 60.865 2.102 60.951 2.287 ;
      RECT 60.818 2.099 60.865 2.289 ;
      RECT 60.732 2.095 60.818 2.292 ;
      RECT 60.646 2.091 60.732 2.295 ;
      RECT 60.56 2.087 60.646 2.299 ;
      RECT 62.495 3.15 62.775 3.43 ;
      RECT 62.535 3.13 62.795 3.39 ;
      RECT 62.525 3.14 62.795 3.39 ;
      RECT 62.535 3.067 62.75 3.43 ;
      RECT 62.59 2.99 62.745 3.43 ;
      RECT 62.595 2.775 62.745 3.43 ;
      RECT 62.585 2.577 62.735 2.828 ;
      RECT 62.575 2.577 62.735 2.695 ;
      RECT 62.57 2.455 62.73 2.598 ;
      RECT 62.555 2.455 62.73 2.503 ;
      RECT 62.55 2.165 62.725 2.48 ;
      RECT 62.535 2.165 62.725 2.45 ;
      RECT 62.495 2.165 62.755 2.425 ;
      RECT 62.405 3.635 62.485 3.895 ;
      RECT 61.81 2.355 61.815 2.62 ;
      RECT 61.69 2.355 61.815 2.615 ;
      RECT 62.365 3.6 62.405 3.895 ;
      RECT 62.32 3.522 62.365 3.895 ;
      RECT 62.3 3.45 62.32 3.895 ;
      RECT 62.29 3.402 62.3 3.895 ;
      RECT 62.255 3.335 62.29 3.895 ;
      RECT 62.225 3.235 62.255 3.895 ;
      RECT 62.205 3.16 62.225 3.695 ;
      RECT 62.195 3.11 62.205 3.65 ;
      RECT 62.19 3.087 62.195 3.623 ;
      RECT 62.185 3.072 62.19 3.61 ;
      RECT 62.18 3.057 62.185 3.588 ;
      RECT 62.175 3.042 62.18 3.57 ;
      RECT 62.15 2.997 62.175 3.525 ;
      RECT 62.14 2.945 62.15 3.468 ;
      RECT 62.13 2.915 62.14 3.435 ;
      RECT 62.12 2.88 62.13 3.403 ;
      RECT 62.085 2.812 62.12 3.335 ;
      RECT 62.08 2.751 62.085 3.27 ;
      RECT 62.07 2.739 62.08 3.25 ;
      RECT 62.065 2.727 62.07 3.23 ;
      RECT 62.06 2.719 62.065 3.218 ;
      RECT 62.055 2.711 62.06 3.198 ;
      RECT 62.045 2.699 62.055 3.17 ;
      RECT 62.035 2.683 62.045 3.14 ;
      RECT 62.01 2.655 62.035 3.078 ;
      RECT 62 2.626 62.01 3.023 ;
      RECT 61.985 2.605 62 2.983 ;
      RECT 61.98 2.589 61.985 2.955 ;
      RECT 61.975 2.577 61.98 2.945 ;
      RECT 61.97 2.572 61.975 2.918 ;
      RECT 61.965 2.565 61.97 2.905 ;
      RECT 61.95 2.548 61.965 2.878 ;
      RECT 61.94 2.355 61.95 2.838 ;
      RECT 61.93 2.355 61.94 2.805 ;
      RECT 61.92 2.355 61.93 2.78 ;
      RECT 61.85 2.355 61.92 2.715 ;
      RECT 61.84 2.355 61.85 2.663 ;
      RECT 61.825 2.355 61.84 2.645 ;
      RECT 61.815 2.355 61.825 2.63 ;
      RECT 61.645 3.225 61.905 3.485 ;
      RECT 60.18 3.26 60.185 3.467 ;
      RECT 59.815 3.15 59.89 3.465 ;
      RECT 59.63 3.205 59.785 3.465 ;
      RECT 59.815 3.15 59.92 3.43 ;
      RECT 61.63 3.322 61.645 3.483 ;
      RECT 61.605 3.33 61.63 3.488 ;
      RECT 61.58 3.337 61.605 3.493 ;
      RECT 61.517 3.348 61.58 3.502 ;
      RECT 61.431 3.367 61.517 3.519 ;
      RECT 61.345 3.389 61.431 3.538 ;
      RECT 61.33 3.402 61.345 3.549 ;
      RECT 61.29 3.41 61.33 3.556 ;
      RECT 61.27 3.415 61.29 3.563 ;
      RECT 61.232 3.416 61.27 3.566 ;
      RECT 61.146 3.419 61.232 3.567 ;
      RECT 61.06 3.423 61.146 3.568 ;
      RECT 61.011 3.425 61.06 3.57 ;
      RECT 60.925 3.425 61.011 3.572 ;
      RECT 60.885 3.42 60.925 3.574 ;
      RECT 60.875 3.414 60.885 3.575 ;
      RECT 60.835 3.409 60.875 3.572 ;
      RECT 60.825 3.402 60.835 3.568 ;
      RECT 60.81 3.398 60.825 3.566 ;
      RECT 60.793 3.394 60.81 3.564 ;
      RECT 60.707 3.384 60.793 3.556 ;
      RECT 60.621 3.366 60.707 3.542 ;
      RECT 60.535 3.349 60.621 3.528 ;
      RECT 60.51 3.337 60.535 3.519 ;
      RECT 60.44 3.327 60.51 3.512 ;
      RECT 60.395 3.315 60.44 3.503 ;
      RECT 60.335 3.302 60.395 3.495 ;
      RECT 60.33 3.294 60.335 3.49 ;
      RECT 60.295 3.289 60.33 3.488 ;
      RECT 60.24 3.28 60.295 3.481 ;
      RECT 60.2 3.269 60.24 3.473 ;
      RECT 60.185 3.262 60.2 3.469 ;
      RECT 60.165 3.255 60.18 3.466 ;
      RECT 60.15 3.245 60.165 3.464 ;
      RECT 60.135 3.232 60.15 3.461 ;
      RECT 60.11 3.215 60.135 3.457 ;
      RECT 60.095 3.197 60.11 3.454 ;
      RECT 60.07 3.15 60.095 3.452 ;
      RECT 60.046 3.15 60.07 3.449 ;
      RECT 59.96 3.15 60.046 3.441 ;
      RECT 59.92 3.15 59.96 3.433 ;
      RECT 59.785 3.197 59.815 3.465 ;
      RECT 61.465 2.78 61.725 3.04 ;
      RECT 61.425 2.78 61.725 2.918 ;
      RECT 61.39 2.78 61.725 2.903 ;
      RECT 61.335 2.78 61.725 2.883 ;
      RECT 61.255 2.59 61.535 2.87 ;
      RECT 61.255 2.772 61.605 2.87 ;
      RECT 61.255 2.715 61.59 2.87 ;
      RECT 61.255 2.662 61.54 2.87 ;
      RECT 59.085 2.59 59.28 3.375 ;
      RECT 59.165 1.205 59.28 3.375 ;
      RECT 59.02 3.115 59.08 3.375 ;
      RECT 60.39 2.635 60.65 2.895 ;
      RECT 59.075 2.59 59.28 2.87 ;
      RECT 60.385 2.645 60.65 2.83 ;
      RECT 60.1 2.62 60.11 2.77 ;
      RECT 59.335 1.205 59.415 1.55 ;
      RECT 59.07 1.205 59.28 1.55 ;
      RECT 60.375 2.645 60.385 2.829 ;
      RECT 60.365 2.644 60.375 2.826 ;
      RECT 60.356 2.643 60.365 2.824 ;
      RECT 60.27 2.639 60.356 2.814 ;
      RECT 60.196 2.631 60.27 2.796 ;
      RECT 60.11 2.624 60.196 2.779 ;
      RECT 60.05 2.62 60.1 2.769 ;
      RECT 60.015 2.619 60.05 2.766 ;
      RECT 59.96 2.619 60.015 2.768 ;
      RECT 59.925 2.619 59.96 2.772 ;
      RECT 59.839 2.618 59.925 2.779 ;
      RECT 59.753 2.617 59.839 2.789 ;
      RECT 59.667 2.616 59.753 2.8 ;
      RECT 59.581 2.616 59.667 2.81 ;
      RECT 59.495 2.615 59.581 2.82 ;
      RECT 59.46 2.615 59.495 2.86 ;
      RECT 59.455 2.615 59.46 2.903 ;
      RECT 59.43 2.615 59.455 2.92 ;
      RECT 59.355 2.615 59.43 2.935 ;
      RECT 59.335 2.59 59.355 2.948 ;
      RECT 59.33 1.205 59.335 2.958 ;
      RECT 59.305 1.205 59.33 3 ;
      RECT 59.28 1.205 59.305 3.078 ;
      RECT 59.08 2.997 59.085 3.375 ;
      RECT 58.415 2.949 58.43 3.405 ;
      RECT 58.41 3.021 58.516 3.403 ;
      RECT 58.43 2.115 58.565 3.401 ;
      RECT 58.415 2.965 58.57 3.4 ;
      RECT 58.415 3.015 58.575 3.398 ;
      RECT 58.4 3.08 58.575 3.397 ;
      RECT 58.41 3.072 58.58 3.394 ;
      RECT 58.39 3.12 58.58 3.389 ;
      RECT 58.39 3.12 58.595 3.386 ;
      RECT 58.385 3.12 58.595 3.383 ;
      RECT 58.36 3.12 58.62 3.38 ;
      RECT 58.43 2.115 58.59 2.768 ;
      RECT 58.425 2.115 58.59 2.74 ;
      RECT 58.42 2.115 58.59 2.568 ;
      RECT 58.42 2.115 58.61 2.508 ;
      RECT 58.375 2.115 58.635 2.375 ;
      RECT 57.855 2.59 58.135 2.87 ;
      RECT 57.845 2.605 58.135 2.865 ;
      RECT 57.8 2.667 58.135 2.863 ;
      RECT 57.875 2.582 58.04 2.87 ;
      RECT 57.875 2.567 57.996 2.87 ;
      RECT 57.91 2.56 57.996 2.87 ;
      RECT 57.375 3.71 57.655 3.99 ;
      RECT 57.335 3.672 57.63 3.783 ;
      RECT 57.32 3.622 57.61 3.678 ;
      RECT 57.265 3.385 57.525 3.645 ;
      RECT 57.265 3.587 57.605 3.645 ;
      RECT 57.265 3.527 57.6 3.645 ;
      RECT 57.265 3.477 57.58 3.645 ;
      RECT 57.265 3.457 57.575 3.645 ;
      RECT 57.265 3.435 57.57 3.645 ;
      RECT 57.265 3.42 57.54 3.645 ;
      RECT 52.995 6.225 53.315 6.545 ;
      RECT 53.025 5.695 53.195 6.545 ;
      RECT 53.025 5.695 53.2 6.045 ;
      RECT 53.025 5.695 54 5.87 ;
      RECT 53.825 1.965 54 5.87 ;
      RECT 53.77 1.965 54.12 2.315 ;
      RECT 53.795 6.655 54.12 6.98 ;
      RECT 52.68 6.745 54.12 6.915 ;
      RECT 52.68 2.395 52.84 6.915 ;
      RECT 52.995 2.365 53.315 2.685 ;
      RECT 52.68 2.395 53.315 2.565 ;
      RECT 51.94 5.84 52.29 6.19 ;
      RECT 52.015 2.705 52.19 6.19 ;
      RECT 51.95 2.705 52.3 3.055 ;
      RECT 51.35 1.14 51.725 1.51 ;
      RECT 43.27 0.96 43.645 1.33 ;
      RECT 41.835 0.96 42.21 1.33 ;
      RECT 41.835 1.08 51.655 1.25 ;
      RECT 45.955 4.36 51.635 4.53 ;
      RECT 51.465 3.425 51.635 4.53 ;
      RECT 45.765 3.6 45.79 4.53 ;
      RECT 46.02 3.71 46.05 3.99 ;
      RECT 45.725 3.6 45.79 3.86 ;
      RECT 51.375 3.43 51.725 3.78 ;
      RECT 45.555 2.225 45.59 2.485 ;
      RECT 45.33 2.225 45.39 2.485 ;
      RECT 46.01 3.69 46.02 3.99 ;
      RECT 46.005 3.65 46.01 3.99 ;
      RECT 45.99 3.605 46.005 3.99 ;
      RECT 45.985 3.57 45.99 3.99 ;
      RECT 45.98 3.55 45.985 3.99 ;
      RECT 45.955 3.487 45.98 3.99 ;
      RECT 45.95 3.425 45.955 4.53 ;
      RECT 45.93 3.375 45.95 4.53 ;
      RECT 45.92 3.305 45.93 4.53 ;
      RECT 45.875 3.245 45.92 4.53 ;
      RECT 45.79 3.206 45.875 4.53 ;
      RECT 45.785 3.197 45.79 3.57 ;
      RECT 45.775 3.196 45.785 3.553 ;
      RECT 45.75 3.177 45.775 3.523 ;
      RECT 45.745 3.152 45.75 3.502 ;
      RECT 45.735 3.13 45.745 3.493 ;
      RECT 45.73 3.101 45.735 3.483 ;
      RECT 45.69 3.027 45.73 3.455 ;
      RECT 45.67 2.928 45.69 3.42 ;
      RECT 45.655 2.864 45.67 3.403 ;
      RECT 45.625 2.788 45.655 3.375 ;
      RECT 45.605 2.703 45.625 3.348 ;
      RECT 45.565 2.599 45.605 3.255 ;
      RECT 45.56 2.52 45.565 3.163 ;
      RECT 45.555 2.503 45.56 3.14 ;
      RECT 45.55 2.225 45.555 3.12 ;
      RECT 45.52 2.225 45.55 3.058 ;
      RECT 45.515 2.225 45.52 2.99 ;
      RECT 45.505 2.225 45.515 2.955 ;
      RECT 45.495 2.225 45.505 2.92 ;
      RECT 45.43 2.225 45.495 2.775 ;
      RECT 45.425 2.225 45.43 2.645 ;
      RECT 45.395 2.225 45.425 2.578 ;
      RECT 45.39 2.225 45.395 2.503 ;
      RECT 49.725 2.16 49.985 2.42 ;
      RECT 49.72 2.16 49.985 2.368 ;
      RECT 49.715 2.16 49.985 2.338 ;
      RECT 49.69 2.03 49.97 2.31 ;
      RECT 38.25 6.66 38.6 7.01 ;
      RECT 49.225 6.615 49.575 6.965 ;
      RECT 38.25 6.69 49.575 6.89 ;
      RECT 48.73 3.71 49.01 3.99 ;
      RECT 48.77 3.665 49.035 3.925 ;
      RECT 48.76 3.7 49.035 3.925 ;
      RECT 48.765 3.685 49.01 3.99 ;
      RECT 48.77 3.662 48.98 3.99 ;
      RECT 48.77 3.66 48.965 3.99 ;
      RECT 48.81 3.65 48.965 3.99 ;
      RECT 48.78 3.655 48.965 3.99 ;
      RECT 48.81 3.647 48.91 3.99 ;
      RECT 48.835 3.64 48.91 3.99 ;
      RECT 48.815 3.642 48.91 3.99 ;
      RECT 48.145 3.155 48.405 3.415 ;
      RECT 48.195 3.147 48.385 3.415 ;
      RECT 48.2 3.067 48.385 3.415 ;
      RECT 48.32 2.455 48.385 3.415 ;
      RECT 48.225 2.852 48.385 3.415 ;
      RECT 48.3 2.54 48.385 3.415 ;
      RECT 48.335 2.165 48.471 2.893 ;
      RECT 48.28 2.662 48.471 2.893 ;
      RECT 48.295 2.602 48.385 3.415 ;
      RECT 48.335 2.165 48.495 2.558 ;
      RECT 48.335 2.165 48.505 2.455 ;
      RECT 48.325 2.165 48.585 2.425 ;
      RECT 47.73 3.71 48.01 3.99 ;
      RECT 47.75 3.67 48.01 3.99 ;
      RECT 47.39 3.625 47.495 3.885 ;
      RECT 47.245 2.115 47.335 2.375 ;
      RECT 47.785 3.18 47.79 3.22 ;
      RECT 47.78 3.17 47.785 3.305 ;
      RECT 47.775 3.16 47.78 3.398 ;
      RECT 47.765 3.14 47.775 3.454 ;
      RECT 47.685 3.068 47.765 3.534 ;
      RECT 47.72 3.712 47.73 3.937 ;
      RECT 47.715 3.709 47.72 3.932 ;
      RECT 47.7 3.706 47.715 3.925 ;
      RECT 47.665 3.7 47.7 3.907 ;
      RECT 47.68 3.003 47.685 3.608 ;
      RECT 47.66 2.954 47.68 3.623 ;
      RECT 47.65 3.687 47.665 3.89 ;
      RECT 47.655 2.896 47.66 3.638 ;
      RECT 47.65 2.874 47.655 3.648 ;
      RECT 47.615 2.784 47.65 3.885 ;
      RECT 47.6 2.662 47.615 3.885 ;
      RECT 47.595 2.615 47.6 3.885 ;
      RECT 47.57 2.54 47.595 3.885 ;
      RECT 47.555 2.455 47.57 3.885 ;
      RECT 47.55 2.402 47.555 3.885 ;
      RECT 47.545 2.382 47.55 3.885 ;
      RECT 47.54 2.357 47.545 3.119 ;
      RECT 47.525 3.317 47.545 3.885 ;
      RECT 47.535 2.335 47.54 3.096 ;
      RECT 47.525 2.287 47.535 3.061 ;
      RECT 47.52 2.25 47.525 3.027 ;
      RECT 47.52 3.397 47.525 3.885 ;
      RECT 47.505 2.227 47.52 2.982 ;
      RECT 47.5 3.495 47.52 3.885 ;
      RECT 47.45 2.115 47.505 2.824 ;
      RECT 47.495 3.617 47.5 3.885 ;
      RECT 47.435 2.115 47.45 2.663 ;
      RECT 47.43 2.115 47.435 2.615 ;
      RECT 47.425 2.115 47.43 2.603 ;
      RECT 47.38 2.115 47.425 2.54 ;
      RECT 47.355 2.115 47.38 2.458 ;
      RECT 47.34 2.115 47.355 2.41 ;
      RECT 47.335 2.115 47.34 2.38 ;
      RECT 46.66 3.565 46.705 3.825 ;
      RECT 46.565 2.1 46.71 2.36 ;
      RECT 47.07 2.722 47.08 2.813 ;
      RECT 47.055 2.66 47.07 2.869 ;
      RECT 47.05 2.607 47.055 2.915 ;
      RECT 47 2.554 47.05 3.041 ;
      RECT 46.995 2.509 47 3.188 ;
      RECT 46.985 2.497 46.995 3.23 ;
      RECT 46.95 2.461 46.985 3.335 ;
      RECT 46.945 2.429 46.95 3.441 ;
      RECT 46.93 2.411 46.945 3.486 ;
      RECT 46.925 2.394 46.93 2.72 ;
      RECT 46.92 2.775 46.93 3.543 ;
      RECT 46.915 2.38 46.925 2.693 ;
      RECT 46.91 2.83 46.92 3.825 ;
      RECT 46.905 2.366 46.915 2.678 ;
      RECT 46.905 2.88 46.91 3.825 ;
      RECT 46.89 2.343 46.905 2.658 ;
      RECT 46.87 3.002 46.905 3.825 ;
      RECT 46.885 2.325 46.89 2.64 ;
      RECT 46.88 2.317 46.885 2.63 ;
      RECT 46.85 2.285 46.88 2.594 ;
      RECT 46.86 3.13 46.87 3.825 ;
      RECT 46.855 3.157 46.86 3.825 ;
      RECT 46.85 3.207 46.855 3.825 ;
      RECT 46.84 2.251 46.85 2.559 ;
      RECT 46.8 3.275 46.85 3.825 ;
      RECT 46.825 2.228 46.84 2.535 ;
      RECT 46.8 2.1 46.825 2.498 ;
      RECT 46.795 2.1 46.8 2.47 ;
      RECT 46.765 3.375 46.8 3.825 ;
      RECT 46.79 2.1 46.795 2.463 ;
      RECT 46.785 2.1 46.79 2.453 ;
      RECT 46.77 2.1 46.785 2.438 ;
      RECT 46.755 2.1 46.77 2.41 ;
      RECT 46.72 3.48 46.765 3.825 ;
      RECT 46.74 2.1 46.755 2.383 ;
      RECT 46.71 2.1 46.74 2.368 ;
      RECT 46.705 3.552 46.72 3.825 ;
      RECT 46.63 2.635 46.67 2.895 ;
      RECT 46.405 2.582 46.41 2.84 ;
      RECT 42.36 2.06 42.62 2.32 ;
      RECT 42.36 2.085 42.635 2.3 ;
      RECT 44.75 1.91 44.755 2.055 ;
      RECT 46.62 2.63 46.63 2.895 ;
      RECT 46.6 2.622 46.62 2.895 ;
      RECT 46.582 2.618 46.6 2.895 ;
      RECT 46.496 2.607 46.582 2.895 ;
      RECT 46.41 2.59 46.496 2.895 ;
      RECT 46.355 2.577 46.405 2.825 ;
      RECT 46.321 2.569 46.355 2.8 ;
      RECT 46.235 2.558 46.321 2.765 ;
      RECT 46.2 2.535 46.235 2.73 ;
      RECT 46.19 2.497 46.2 2.716 ;
      RECT 46.185 2.47 46.19 2.712 ;
      RECT 46.18 2.457 46.185 2.709 ;
      RECT 46.17 2.437 46.18 2.705 ;
      RECT 46.165 2.412 46.17 2.701 ;
      RECT 46.14 2.367 46.165 2.695 ;
      RECT 46.13 2.308 46.14 2.687 ;
      RECT 46.12 2.276 46.13 2.678 ;
      RECT 46.1 2.228 46.12 2.658 ;
      RECT 46.095 2.188 46.1 2.628 ;
      RECT 46.08 2.162 46.095 2.602 ;
      RECT 46.075 2.14 46.08 2.578 ;
      RECT 46.06 2.112 46.075 2.554 ;
      RECT 46.045 2.085 46.06 2.518 ;
      RECT 46.03 2.062 46.045 2.48 ;
      RECT 46.025 2.052 46.03 2.455 ;
      RECT 46.015 2.045 46.025 2.438 ;
      RECT 46 2.032 46.015 2.408 ;
      RECT 45.995 2.022 46 2.383 ;
      RECT 45.99 2.017 45.995 2.37 ;
      RECT 45.98 2.01 45.99 2.35 ;
      RECT 45.975 2.003 45.98 2.335 ;
      RECT 45.95 1.996 45.975 2.293 ;
      RECT 45.935 1.986 45.95 2.243 ;
      RECT 45.925 1.981 45.935 2.213 ;
      RECT 45.915 1.977 45.925 2.188 ;
      RECT 45.9 1.974 45.915 2.178 ;
      RECT 45.85 1.971 45.9 2.163 ;
      RECT 45.83 1.969 45.85 2.148 ;
      RECT 45.781 1.967 45.83 2.143 ;
      RECT 45.695 1.963 45.781 2.138 ;
      RECT 45.656 1.96 45.695 2.134 ;
      RECT 45.57 1.956 45.656 2.129 ;
      RECT 45.52 1.953 45.57 2.123 ;
      RECT 45.471 1.95 45.52 2.118 ;
      RECT 45.385 1.947 45.471 2.113 ;
      RECT 45.381 1.945 45.385 2.11 ;
      RECT 45.295 1.942 45.381 2.105 ;
      RECT 45.246 1.938 45.295 2.098 ;
      RECT 45.16 1.935 45.246 2.093 ;
      RECT 45.136 1.932 45.16 2.089 ;
      RECT 45.05 1.93 45.136 2.084 ;
      RECT 44.985 1.926 45.05 2.077 ;
      RECT 44.982 1.925 44.985 2.074 ;
      RECT 44.896 1.922 44.982 2.071 ;
      RECT 44.81 1.916 44.896 2.064 ;
      RECT 44.78 1.912 44.81 2.06 ;
      RECT 44.755 1.91 44.78 2.058 ;
      RECT 44.7 1.907 44.75 2.055 ;
      RECT 44.62 1.906 44.7 2.055 ;
      RECT 44.565 1.908 44.62 2.058 ;
      RECT 44.55 1.909 44.565 2.062 ;
      RECT 44.495 1.917 44.55 2.072 ;
      RECT 44.465 1.925 44.495 2.085 ;
      RECT 44.446 1.926 44.465 2.091 ;
      RECT 44.36 1.929 44.446 2.096 ;
      RECT 44.29 1.934 44.36 2.105 ;
      RECT 44.271 1.937 44.29 2.111 ;
      RECT 44.185 1.941 44.271 2.116 ;
      RECT 44.145 1.945 44.185 2.123 ;
      RECT 44.136 1.947 44.145 2.126 ;
      RECT 44.05 1.951 44.136 2.131 ;
      RECT 44.047 1.954 44.05 2.135 ;
      RECT 43.961 1.957 44.047 2.139 ;
      RECT 43.875 1.963 43.961 2.147 ;
      RECT 43.851 1.967 43.875 2.151 ;
      RECT 43.765 1.971 43.851 2.156 ;
      RECT 43.72 1.976 43.765 2.163 ;
      RECT 43.64 1.981 43.72 2.17 ;
      RECT 43.56 1.987 43.64 2.185 ;
      RECT 43.535 1.991 43.56 2.198 ;
      RECT 43.47 1.994 43.535 2.21 ;
      RECT 43.415 1.999 43.47 2.225 ;
      RECT 43.385 2.002 43.415 2.243 ;
      RECT 43.375 2.004 43.385 2.256 ;
      RECT 43.315 2.019 43.375 2.266 ;
      RECT 43.3 2.036 43.315 2.275 ;
      RECT 43.295 2.045 43.3 2.275 ;
      RECT 43.285 2.055 43.295 2.275 ;
      RECT 43.275 2.072 43.285 2.275 ;
      RECT 43.255 2.082 43.275 2.276 ;
      RECT 43.21 2.092 43.255 2.277 ;
      RECT 43.175 2.101 43.21 2.279 ;
      RECT 43.11 2.106 43.175 2.281 ;
      RECT 43.03 2.107 43.11 2.284 ;
      RECT 43.026 2.105 43.03 2.285 ;
      RECT 42.94 2.102 43.026 2.287 ;
      RECT 42.893 2.099 42.94 2.289 ;
      RECT 42.807 2.095 42.893 2.292 ;
      RECT 42.721 2.091 42.807 2.295 ;
      RECT 42.635 2.087 42.721 2.299 ;
      RECT 44.57 3.15 44.85 3.43 ;
      RECT 44.61 3.13 44.87 3.39 ;
      RECT 44.6 3.14 44.87 3.39 ;
      RECT 44.61 3.067 44.825 3.43 ;
      RECT 44.665 2.99 44.82 3.43 ;
      RECT 44.67 2.775 44.82 3.43 ;
      RECT 44.66 2.577 44.81 2.828 ;
      RECT 44.65 2.577 44.81 2.695 ;
      RECT 44.645 2.455 44.805 2.598 ;
      RECT 44.63 2.455 44.805 2.503 ;
      RECT 44.625 2.165 44.8 2.48 ;
      RECT 44.61 2.165 44.8 2.45 ;
      RECT 44.57 2.165 44.83 2.425 ;
      RECT 44.48 3.635 44.56 3.895 ;
      RECT 43.885 2.355 43.89 2.62 ;
      RECT 43.765 2.355 43.89 2.615 ;
      RECT 44.44 3.6 44.48 3.895 ;
      RECT 44.395 3.522 44.44 3.895 ;
      RECT 44.375 3.45 44.395 3.895 ;
      RECT 44.365 3.402 44.375 3.895 ;
      RECT 44.33 3.335 44.365 3.895 ;
      RECT 44.3 3.235 44.33 3.895 ;
      RECT 44.28 3.16 44.3 3.695 ;
      RECT 44.27 3.11 44.28 3.65 ;
      RECT 44.265 3.087 44.27 3.623 ;
      RECT 44.26 3.072 44.265 3.61 ;
      RECT 44.255 3.057 44.26 3.588 ;
      RECT 44.25 3.042 44.255 3.57 ;
      RECT 44.225 2.997 44.25 3.525 ;
      RECT 44.215 2.945 44.225 3.468 ;
      RECT 44.205 2.915 44.215 3.435 ;
      RECT 44.195 2.88 44.205 3.403 ;
      RECT 44.16 2.812 44.195 3.335 ;
      RECT 44.155 2.751 44.16 3.27 ;
      RECT 44.145 2.739 44.155 3.25 ;
      RECT 44.14 2.727 44.145 3.23 ;
      RECT 44.135 2.719 44.14 3.218 ;
      RECT 44.13 2.711 44.135 3.198 ;
      RECT 44.12 2.699 44.13 3.17 ;
      RECT 44.11 2.683 44.12 3.14 ;
      RECT 44.085 2.655 44.11 3.078 ;
      RECT 44.075 2.626 44.085 3.023 ;
      RECT 44.06 2.605 44.075 2.983 ;
      RECT 44.055 2.589 44.06 2.955 ;
      RECT 44.05 2.577 44.055 2.945 ;
      RECT 44.045 2.572 44.05 2.918 ;
      RECT 44.04 2.565 44.045 2.905 ;
      RECT 44.025 2.548 44.04 2.878 ;
      RECT 44.015 2.355 44.025 2.838 ;
      RECT 44.005 2.355 44.015 2.805 ;
      RECT 43.995 2.355 44.005 2.78 ;
      RECT 43.925 2.355 43.995 2.715 ;
      RECT 43.915 2.355 43.925 2.663 ;
      RECT 43.9 2.355 43.915 2.645 ;
      RECT 43.89 2.355 43.9 2.63 ;
      RECT 43.72 3.225 43.98 3.485 ;
      RECT 42.255 3.26 42.26 3.467 ;
      RECT 41.89 3.15 41.965 3.465 ;
      RECT 41.705 3.205 41.86 3.465 ;
      RECT 41.89 3.15 41.995 3.43 ;
      RECT 43.705 3.322 43.72 3.483 ;
      RECT 43.68 3.33 43.705 3.488 ;
      RECT 43.655 3.337 43.68 3.493 ;
      RECT 43.592 3.348 43.655 3.502 ;
      RECT 43.506 3.367 43.592 3.519 ;
      RECT 43.42 3.389 43.506 3.538 ;
      RECT 43.405 3.402 43.42 3.549 ;
      RECT 43.365 3.41 43.405 3.556 ;
      RECT 43.345 3.415 43.365 3.563 ;
      RECT 43.307 3.416 43.345 3.566 ;
      RECT 43.221 3.419 43.307 3.567 ;
      RECT 43.135 3.423 43.221 3.568 ;
      RECT 43.086 3.425 43.135 3.57 ;
      RECT 43 3.425 43.086 3.572 ;
      RECT 42.96 3.42 43 3.574 ;
      RECT 42.95 3.414 42.96 3.575 ;
      RECT 42.91 3.409 42.95 3.572 ;
      RECT 42.9 3.402 42.91 3.568 ;
      RECT 42.885 3.398 42.9 3.566 ;
      RECT 42.868 3.394 42.885 3.564 ;
      RECT 42.782 3.384 42.868 3.556 ;
      RECT 42.696 3.366 42.782 3.542 ;
      RECT 42.61 3.349 42.696 3.528 ;
      RECT 42.585 3.337 42.61 3.519 ;
      RECT 42.515 3.327 42.585 3.512 ;
      RECT 42.47 3.315 42.515 3.503 ;
      RECT 42.41 3.302 42.47 3.495 ;
      RECT 42.405 3.294 42.41 3.49 ;
      RECT 42.37 3.289 42.405 3.488 ;
      RECT 42.315 3.28 42.37 3.481 ;
      RECT 42.275 3.269 42.315 3.473 ;
      RECT 42.26 3.262 42.275 3.469 ;
      RECT 42.24 3.255 42.255 3.466 ;
      RECT 42.225 3.245 42.24 3.464 ;
      RECT 42.21 3.232 42.225 3.461 ;
      RECT 42.185 3.215 42.21 3.457 ;
      RECT 42.17 3.197 42.185 3.454 ;
      RECT 42.145 3.15 42.17 3.452 ;
      RECT 42.121 3.15 42.145 3.449 ;
      RECT 42.035 3.15 42.121 3.441 ;
      RECT 41.995 3.15 42.035 3.433 ;
      RECT 41.86 3.197 41.89 3.465 ;
      RECT 43.54 2.78 43.8 3.04 ;
      RECT 43.5 2.78 43.8 2.918 ;
      RECT 43.465 2.78 43.8 2.903 ;
      RECT 43.41 2.78 43.8 2.883 ;
      RECT 43.33 2.59 43.61 2.87 ;
      RECT 43.33 2.772 43.68 2.87 ;
      RECT 43.33 2.715 43.665 2.87 ;
      RECT 43.33 2.662 43.615 2.87 ;
      RECT 41.16 2.59 41.355 3.375 ;
      RECT 41.24 1.205 41.355 3.375 ;
      RECT 41.095 3.115 41.155 3.375 ;
      RECT 42.465 2.635 42.725 2.895 ;
      RECT 41.15 2.59 41.355 2.87 ;
      RECT 42.46 2.645 42.725 2.83 ;
      RECT 42.175 2.62 42.185 2.77 ;
      RECT 41.41 1.205 41.49 1.55 ;
      RECT 41.145 1.205 41.355 1.55 ;
      RECT 42.45 2.645 42.46 2.829 ;
      RECT 42.44 2.644 42.45 2.826 ;
      RECT 42.431 2.643 42.44 2.824 ;
      RECT 42.345 2.639 42.431 2.814 ;
      RECT 42.271 2.631 42.345 2.796 ;
      RECT 42.185 2.624 42.271 2.779 ;
      RECT 42.125 2.62 42.175 2.769 ;
      RECT 42.09 2.619 42.125 2.766 ;
      RECT 42.035 2.619 42.09 2.768 ;
      RECT 42 2.619 42.035 2.772 ;
      RECT 41.914 2.618 42 2.779 ;
      RECT 41.828 2.617 41.914 2.789 ;
      RECT 41.742 2.616 41.828 2.8 ;
      RECT 41.656 2.616 41.742 2.81 ;
      RECT 41.57 2.615 41.656 2.82 ;
      RECT 41.535 2.615 41.57 2.86 ;
      RECT 41.53 2.615 41.535 2.903 ;
      RECT 41.505 2.615 41.53 2.92 ;
      RECT 41.43 2.615 41.505 2.935 ;
      RECT 41.41 2.59 41.43 2.948 ;
      RECT 41.405 1.205 41.41 2.958 ;
      RECT 41.38 1.205 41.405 3 ;
      RECT 41.355 1.205 41.38 3.078 ;
      RECT 41.155 2.997 41.16 3.375 ;
      RECT 40.49 2.949 40.505 3.405 ;
      RECT 40.485 3.021 40.591 3.403 ;
      RECT 40.505 2.115 40.64 3.401 ;
      RECT 40.49 2.965 40.645 3.4 ;
      RECT 40.49 3.015 40.65 3.398 ;
      RECT 40.475 3.08 40.65 3.397 ;
      RECT 40.485 3.072 40.655 3.394 ;
      RECT 40.465 3.12 40.655 3.389 ;
      RECT 40.465 3.12 40.67 3.386 ;
      RECT 40.46 3.12 40.67 3.383 ;
      RECT 40.435 3.12 40.695 3.38 ;
      RECT 40.505 2.115 40.665 2.768 ;
      RECT 40.5 2.115 40.665 2.74 ;
      RECT 40.495 2.115 40.665 2.568 ;
      RECT 40.495 2.115 40.685 2.508 ;
      RECT 40.45 2.115 40.71 2.375 ;
      RECT 39.93 2.59 40.21 2.87 ;
      RECT 39.92 2.605 40.21 2.865 ;
      RECT 39.875 2.667 40.21 2.863 ;
      RECT 39.95 2.582 40.115 2.87 ;
      RECT 39.95 2.567 40.071 2.87 ;
      RECT 39.985 2.56 40.071 2.87 ;
      RECT 39.45 3.71 39.73 3.99 ;
      RECT 39.41 3.672 39.705 3.783 ;
      RECT 39.395 3.622 39.685 3.678 ;
      RECT 39.34 3.385 39.6 3.645 ;
      RECT 39.34 3.587 39.68 3.645 ;
      RECT 39.34 3.527 39.675 3.645 ;
      RECT 39.34 3.477 39.655 3.645 ;
      RECT 39.34 3.457 39.65 3.645 ;
      RECT 39.34 3.435 39.645 3.645 ;
      RECT 39.34 3.42 39.615 3.645 ;
      RECT 35.07 6.225 35.39 6.545 ;
      RECT 35.1 5.695 35.27 6.545 ;
      RECT 35.1 5.695 35.275 6.045 ;
      RECT 35.1 5.695 36.075 5.87 ;
      RECT 35.9 1.965 36.075 5.87 ;
      RECT 35.845 1.965 36.195 2.315 ;
      RECT 35.87 6.655 36.195 6.98 ;
      RECT 34.755 6.745 36.195 6.915 ;
      RECT 34.755 2.395 34.915 6.915 ;
      RECT 35.07 2.365 35.39 2.685 ;
      RECT 34.755 2.395 35.39 2.565 ;
      RECT 34.015 5.84 34.365 6.19 ;
      RECT 34.09 2.705 34.265 6.19 ;
      RECT 34.025 2.705 34.375 3.055 ;
      RECT 33.425 1.14 33.8 1.51 ;
      RECT 25.345 0.96 25.72 1.33 ;
      RECT 23.91 0.96 24.285 1.33 ;
      RECT 23.91 1.08 33.73 1.25 ;
      RECT 28.03 4.36 33.71 4.53 ;
      RECT 33.54 3.425 33.71 4.53 ;
      RECT 27.84 3.6 27.865 4.53 ;
      RECT 28.095 3.71 28.125 3.99 ;
      RECT 27.8 3.6 27.865 3.86 ;
      RECT 33.45 3.43 33.8 3.78 ;
      RECT 27.63 2.225 27.665 2.485 ;
      RECT 27.405 2.225 27.465 2.485 ;
      RECT 28.085 3.69 28.095 3.99 ;
      RECT 28.08 3.65 28.085 3.99 ;
      RECT 28.065 3.605 28.08 3.99 ;
      RECT 28.06 3.57 28.065 3.99 ;
      RECT 28.055 3.55 28.06 3.99 ;
      RECT 28.03 3.487 28.055 3.99 ;
      RECT 28.025 3.425 28.03 4.53 ;
      RECT 28.005 3.375 28.025 4.53 ;
      RECT 27.995 3.305 28.005 4.53 ;
      RECT 27.95 3.245 27.995 4.53 ;
      RECT 27.865 3.206 27.95 4.53 ;
      RECT 27.86 3.197 27.865 3.57 ;
      RECT 27.85 3.196 27.86 3.553 ;
      RECT 27.825 3.177 27.85 3.523 ;
      RECT 27.82 3.152 27.825 3.502 ;
      RECT 27.81 3.13 27.82 3.493 ;
      RECT 27.805 3.101 27.81 3.483 ;
      RECT 27.765 3.027 27.805 3.455 ;
      RECT 27.745 2.928 27.765 3.42 ;
      RECT 27.73 2.864 27.745 3.403 ;
      RECT 27.7 2.788 27.73 3.375 ;
      RECT 27.68 2.703 27.7 3.348 ;
      RECT 27.64 2.599 27.68 3.255 ;
      RECT 27.635 2.52 27.64 3.163 ;
      RECT 27.63 2.503 27.635 3.14 ;
      RECT 27.625 2.225 27.63 3.12 ;
      RECT 27.595 2.225 27.625 3.058 ;
      RECT 27.59 2.225 27.595 2.99 ;
      RECT 27.58 2.225 27.59 2.955 ;
      RECT 27.57 2.225 27.58 2.92 ;
      RECT 27.505 2.225 27.57 2.775 ;
      RECT 27.5 2.225 27.505 2.645 ;
      RECT 27.47 2.225 27.5 2.578 ;
      RECT 27.465 2.225 27.47 2.503 ;
      RECT 31.8 2.16 32.06 2.42 ;
      RECT 31.795 2.16 32.06 2.368 ;
      RECT 31.79 2.16 32.06 2.338 ;
      RECT 31.765 2.03 32.045 2.31 ;
      RECT 20.325 6.655 20.675 7.005 ;
      RECT 31.295 6.61 31.645 6.96 ;
      RECT 20.325 6.685 31.645 6.885 ;
      RECT 30.805 3.71 31.085 3.99 ;
      RECT 30.845 3.665 31.11 3.925 ;
      RECT 30.835 3.7 31.11 3.925 ;
      RECT 30.84 3.685 31.085 3.99 ;
      RECT 30.845 3.662 31.055 3.99 ;
      RECT 30.845 3.66 31.04 3.99 ;
      RECT 30.885 3.65 31.04 3.99 ;
      RECT 30.855 3.655 31.04 3.99 ;
      RECT 30.885 3.647 30.985 3.99 ;
      RECT 30.91 3.64 30.985 3.99 ;
      RECT 30.89 3.642 30.985 3.99 ;
      RECT 30.22 3.155 30.48 3.415 ;
      RECT 30.27 3.147 30.46 3.415 ;
      RECT 30.275 3.067 30.46 3.415 ;
      RECT 30.395 2.455 30.46 3.415 ;
      RECT 30.3 2.852 30.46 3.415 ;
      RECT 30.375 2.54 30.46 3.415 ;
      RECT 30.41 2.165 30.546 2.893 ;
      RECT 30.355 2.662 30.546 2.893 ;
      RECT 30.37 2.602 30.46 3.415 ;
      RECT 30.41 2.165 30.57 2.558 ;
      RECT 30.41 2.165 30.58 2.455 ;
      RECT 30.4 2.165 30.66 2.425 ;
      RECT 29.805 3.71 30.085 3.99 ;
      RECT 29.825 3.67 30.085 3.99 ;
      RECT 29.465 3.625 29.57 3.885 ;
      RECT 29.32 2.115 29.41 2.375 ;
      RECT 29.86 3.18 29.865 3.22 ;
      RECT 29.855 3.17 29.86 3.305 ;
      RECT 29.85 3.16 29.855 3.398 ;
      RECT 29.84 3.14 29.85 3.454 ;
      RECT 29.76 3.068 29.84 3.534 ;
      RECT 29.795 3.712 29.805 3.937 ;
      RECT 29.79 3.709 29.795 3.932 ;
      RECT 29.775 3.706 29.79 3.925 ;
      RECT 29.74 3.7 29.775 3.907 ;
      RECT 29.755 3.003 29.76 3.608 ;
      RECT 29.735 2.954 29.755 3.623 ;
      RECT 29.725 3.687 29.74 3.89 ;
      RECT 29.73 2.896 29.735 3.638 ;
      RECT 29.725 2.874 29.73 3.648 ;
      RECT 29.69 2.784 29.725 3.885 ;
      RECT 29.675 2.662 29.69 3.885 ;
      RECT 29.67 2.615 29.675 3.885 ;
      RECT 29.645 2.54 29.67 3.885 ;
      RECT 29.63 2.455 29.645 3.885 ;
      RECT 29.625 2.402 29.63 3.885 ;
      RECT 29.62 2.382 29.625 3.885 ;
      RECT 29.615 2.357 29.62 3.119 ;
      RECT 29.6 3.317 29.62 3.885 ;
      RECT 29.61 2.335 29.615 3.096 ;
      RECT 29.6 2.287 29.61 3.061 ;
      RECT 29.595 2.25 29.6 3.027 ;
      RECT 29.595 3.397 29.6 3.885 ;
      RECT 29.58 2.227 29.595 2.982 ;
      RECT 29.575 3.495 29.595 3.885 ;
      RECT 29.525 2.115 29.58 2.824 ;
      RECT 29.57 3.617 29.575 3.885 ;
      RECT 29.51 2.115 29.525 2.663 ;
      RECT 29.505 2.115 29.51 2.615 ;
      RECT 29.5 2.115 29.505 2.603 ;
      RECT 29.455 2.115 29.5 2.54 ;
      RECT 29.43 2.115 29.455 2.458 ;
      RECT 29.415 2.115 29.43 2.41 ;
      RECT 29.41 2.115 29.415 2.38 ;
      RECT 28.735 3.565 28.78 3.825 ;
      RECT 28.64 2.1 28.785 2.36 ;
      RECT 29.145 2.722 29.155 2.813 ;
      RECT 29.13 2.66 29.145 2.869 ;
      RECT 29.125 2.607 29.13 2.915 ;
      RECT 29.075 2.554 29.125 3.041 ;
      RECT 29.07 2.509 29.075 3.188 ;
      RECT 29.06 2.497 29.07 3.23 ;
      RECT 29.025 2.461 29.06 3.335 ;
      RECT 29.02 2.429 29.025 3.441 ;
      RECT 29.005 2.411 29.02 3.486 ;
      RECT 29 2.394 29.005 2.72 ;
      RECT 28.995 2.775 29.005 3.543 ;
      RECT 28.99 2.38 29 2.693 ;
      RECT 28.985 2.83 28.995 3.825 ;
      RECT 28.98 2.366 28.99 2.678 ;
      RECT 28.98 2.88 28.985 3.825 ;
      RECT 28.965 2.343 28.98 2.658 ;
      RECT 28.945 3.002 28.98 3.825 ;
      RECT 28.96 2.325 28.965 2.64 ;
      RECT 28.955 2.317 28.96 2.63 ;
      RECT 28.925 2.285 28.955 2.594 ;
      RECT 28.935 3.13 28.945 3.825 ;
      RECT 28.93 3.157 28.935 3.825 ;
      RECT 28.925 3.207 28.93 3.825 ;
      RECT 28.915 2.251 28.925 2.559 ;
      RECT 28.875 3.275 28.925 3.825 ;
      RECT 28.9 2.228 28.915 2.535 ;
      RECT 28.875 2.1 28.9 2.498 ;
      RECT 28.87 2.1 28.875 2.47 ;
      RECT 28.84 3.375 28.875 3.825 ;
      RECT 28.865 2.1 28.87 2.463 ;
      RECT 28.86 2.1 28.865 2.453 ;
      RECT 28.845 2.1 28.86 2.438 ;
      RECT 28.83 2.1 28.845 2.41 ;
      RECT 28.795 3.48 28.84 3.825 ;
      RECT 28.815 2.1 28.83 2.383 ;
      RECT 28.785 2.1 28.815 2.368 ;
      RECT 28.78 3.552 28.795 3.825 ;
      RECT 28.705 2.635 28.745 2.895 ;
      RECT 28.48 2.582 28.485 2.84 ;
      RECT 24.435 2.06 24.695 2.32 ;
      RECT 24.435 2.085 24.71 2.3 ;
      RECT 26.825 1.91 26.83 2.055 ;
      RECT 28.695 2.63 28.705 2.895 ;
      RECT 28.675 2.622 28.695 2.895 ;
      RECT 28.657 2.618 28.675 2.895 ;
      RECT 28.571 2.607 28.657 2.895 ;
      RECT 28.485 2.59 28.571 2.895 ;
      RECT 28.43 2.577 28.48 2.825 ;
      RECT 28.396 2.569 28.43 2.8 ;
      RECT 28.31 2.558 28.396 2.765 ;
      RECT 28.275 2.535 28.31 2.73 ;
      RECT 28.265 2.497 28.275 2.716 ;
      RECT 28.26 2.47 28.265 2.712 ;
      RECT 28.255 2.457 28.26 2.709 ;
      RECT 28.245 2.437 28.255 2.705 ;
      RECT 28.24 2.412 28.245 2.701 ;
      RECT 28.215 2.367 28.24 2.695 ;
      RECT 28.205 2.308 28.215 2.687 ;
      RECT 28.195 2.276 28.205 2.678 ;
      RECT 28.175 2.228 28.195 2.658 ;
      RECT 28.17 2.188 28.175 2.628 ;
      RECT 28.155 2.162 28.17 2.602 ;
      RECT 28.15 2.14 28.155 2.578 ;
      RECT 28.135 2.112 28.15 2.554 ;
      RECT 28.12 2.085 28.135 2.518 ;
      RECT 28.105 2.062 28.12 2.48 ;
      RECT 28.1 2.052 28.105 2.455 ;
      RECT 28.09 2.045 28.1 2.438 ;
      RECT 28.075 2.032 28.09 2.408 ;
      RECT 28.07 2.022 28.075 2.383 ;
      RECT 28.065 2.017 28.07 2.37 ;
      RECT 28.055 2.01 28.065 2.35 ;
      RECT 28.05 2.003 28.055 2.335 ;
      RECT 28.025 1.996 28.05 2.293 ;
      RECT 28.01 1.986 28.025 2.243 ;
      RECT 28 1.981 28.01 2.213 ;
      RECT 27.99 1.977 28 2.188 ;
      RECT 27.975 1.974 27.99 2.178 ;
      RECT 27.925 1.971 27.975 2.163 ;
      RECT 27.905 1.969 27.925 2.148 ;
      RECT 27.856 1.967 27.905 2.143 ;
      RECT 27.77 1.963 27.856 2.138 ;
      RECT 27.731 1.96 27.77 2.134 ;
      RECT 27.645 1.956 27.731 2.129 ;
      RECT 27.595 1.953 27.645 2.123 ;
      RECT 27.546 1.95 27.595 2.118 ;
      RECT 27.46 1.947 27.546 2.113 ;
      RECT 27.456 1.945 27.46 2.11 ;
      RECT 27.37 1.942 27.456 2.105 ;
      RECT 27.321 1.938 27.37 2.098 ;
      RECT 27.235 1.935 27.321 2.093 ;
      RECT 27.211 1.932 27.235 2.089 ;
      RECT 27.125 1.93 27.211 2.084 ;
      RECT 27.06 1.926 27.125 2.077 ;
      RECT 27.057 1.925 27.06 2.074 ;
      RECT 26.971 1.922 27.057 2.071 ;
      RECT 26.885 1.916 26.971 2.064 ;
      RECT 26.855 1.912 26.885 2.06 ;
      RECT 26.83 1.91 26.855 2.058 ;
      RECT 26.775 1.907 26.825 2.055 ;
      RECT 26.695 1.906 26.775 2.055 ;
      RECT 26.64 1.908 26.695 2.058 ;
      RECT 26.625 1.909 26.64 2.062 ;
      RECT 26.57 1.917 26.625 2.072 ;
      RECT 26.54 1.925 26.57 2.085 ;
      RECT 26.521 1.926 26.54 2.091 ;
      RECT 26.435 1.929 26.521 2.096 ;
      RECT 26.365 1.934 26.435 2.105 ;
      RECT 26.346 1.937 26.365 2.111 ;
      RECT 26.26 1.941 26.346 2.116 ;
      RECT 26.22 1.945 26.26 2.123 ;
      RECT 26.211 1.947 26.22 2.126 ;
      RECT 26.125 1.951 26.211 2.131 ;
      RECT 26.122 1.954 26.125 2.135 ;
      RECT 26.036 1.957 26.122 2.139 ;
      RECT 25.95 1.963 26.036 2.147 ;
      RECT 25.926 1.967 25.95 2.151 ;
      RECT 25.84 1.971 25.926 2.156 ;
      RECT 25.795 1.976 25.84 2.163 ;
      RECT 25.715 1.981 25.795 2.17 ;
      RECT 25.635 1.987 25.715 2.185 ;
      RECT 25.61 1.991 25.635 2.198 ;
      RECT 25.545 1.994 25.61 2.21 ;
      RECT 25.49 1.999 25.545 2.225 ;
      RECT 25.46 2.002 25.49 2.243 ;
      RECT 25.45 2.004 25.46 2.256 ;
      RECT 25.39 2.019 25.45 2.266 ;
      RECT 25.375 2.036 25.39 2.275 ;
      RECT 25.37 2.045 25.375 2.275 ;
      RECT 25.36 2.055 25.37 2.275 ;
      RECT 25.35 2.072 25.36 2.275 ;
      RECT 25.33 2.082 25.35 2.276 ;
      RECT 25.285 2.092 25.33 2.277 ;
      RECT 25.25 2.101 25.285 2.279 ;
      RECT 25.185 2.106 25.25 2.281 ;
      RECT 25.105 2.107 25.185 2.284 ;
      RECT 25.101 2.105 25.105 2.285 ;
      RECT 25.015 2.102 25.101 2.287 ;
      RECT 24.968 2.099 25.015 2.289 ;
      RECT 24.882 2.095 24.968 2.292 ;
      RECT 24.796 2.091 24.882 2.295 ;
      RECT 24.71 2.087 24.796 2.299 ;
      RECT 26.645 3.15 26.925 3.43 ;
      RECT 26.685 3.13 26.945 3.39 ;
      RECT 26.675 3.14 26.945 3.39 ;
      RECT 26.685 3.067 26.9 3.43 ;
      RECT 26.74 2.99 26.895 3.43 ;
      RECT 26.745 2.775 26.895 3.43 ;
      RECT 26.735 2.577 26.885 2.828 ;
      RECT 26.725 2.577 26.885 2.695 ;
      RECT 26.72 2.455 26.88 2.598 ;
      RECT 26.705 2.455 26.88 2.503 ;
      RECT 26.7 2.165 26.875 2.48 ;
      RECT 26.685 2.165 26.875 2.45 ;
      RECT 26.645 2.165 26.905 2.425 ;
      RECT 26.555 3.635 26.635 3.895 ;
      RECT 25.96 2.355 25.965 2.62 ;
      RECT 25.84 2.355 25.965 2.615 ;
      RECT 26.515 3.6 26.555 3.895 ;
      RECT 26.47 3.522 26.515 3.895 ;
      RECT 26.45 3.45 26.47 3.895 ;
      RECT 26.44 3.402 26.45 3.895 ;
      RECT 26.405 3.335 26.44 3.895 ;
      RECT 26.375 3.235 26.405 3.895 ;
      RECT 26.355 3.16 26.375 3.695 ;
      RECT 26.345 3.11 26.355 3.65 ;
      RECT 26.34 3.087 26.345 3.623 ;
      RECT 26.335 3.072 26.34 3.61 ;
      RECT 26.33 3.057 26.335 3.588 ;
      RECT 26.325 3.042 26.33 3.57 ;
      RECT 26.3 2.997 26.325 3.525 ;
      RECT 26.29 2.945 26.3 3.468 ;
      RECT 26.28 2.915 26.29 3.435 ;
      RECT 26.27 2.88 26.28 3.403 ;
      RECT 26.235 2.812 26.27 3.335 ;
      RECT 26.23 2.751 26.235 3.27 ;
      RECT 26.22 2.739 26.23 3.25 ;
      RECT 26.215 2.727 26.22 3.23 ;
      RECT 26.21 2.719 26.215 3.218 ;
      RECT 26.205 2.711 26.21 3.198 ;
      RECT 26.195 2.699 26.205 3.17 ;
      RECT 26.185 2.683 26.195 3.14 ;
      RECT 26.16 2.655 26.185 3.078 ;
      RECT 26.15 2.626 26.16 3.023 ;
      RECT 26.135 2.605 26.15 2.983 ;
      RECT 26.13 2.589 26.135 2.955 ;
      RECT 26.125 2.577 26.13 2.945 ;
      RECT 26.12 2.572 26.125 2.918 ;
      RECT 26.115 2.565 26.12 2.905 ;
      RECT 26.1 2.548 26.115 2.878 ;
      RECT 26.09 2.355 26.1 2.838 ;
      RECT 26.08 2.355 26.09 2.805 ;
      RECT 26.07 2.355 26.08 2.78 ;
      RECT 26 2.355 26.07 2.715 ;
      RECT 25.99 2.355 26 2.663 ;
      RECT 25.975 2.355 25.99 2.645 ;
      RECT 25.965 2.355 25.975 2.63 ;
      RECT 25.795 3.225 26.055 3.485 ;
      RECT 24.33 3.26 24.335 3.467 ;
      RECT 23.965 3.15 24.04 3.465 ;
      RECT 23.78 3.205 23.935 3.465 ;
      RECT 23.965 3.15 24.07 3.43 ;
      RECT 25.78 3.322 25.795 3.483 ;
      RECT 25.755 3.33 25.78 3.488 ;
      RECT 25.73 3.337 25.755 3.493 ;
      RECT 25.667 3.348 25.73 3.502 ;
      RECT 25.581 3.367 25.667 3.519 ;
      RECT 25.495 3.389 25.581 3.538 ;
      RECT 25.48 3.402 25.495 3.549 ;
      RECT 25.44 3.41 25.48 3.556 ;
      RECT 25.42 3.415 25.44 3.563 ;
      RECT 25.382 3.416 25.42 3.566 ;
      RECT 25.296 3.419 25.382 3.567 ;
      RECT 25.21 3.423 25.296 3.568 ;
      RECT 25.161 3.425 25.21 3.57 ;
      RECT 25.075 3.425 25.161 3.572 ;
      RECT 25.035 3.42 25.075 3.574 ;
      RECT 25.025 3.414 25.035 3.575 ;
      RECT 24.985 3.409 25.025 3.572 ;
      RECT 24.975 3.402 24.985 3.568 ;
      RECT 24.96 3.398 24.975 3.566 ;
      RECT 24.943 3.394 24.96 3.564 ;
      RECT 24.857 3.384 24.943 3.556 ;
      RECT 24.771 3.366 24.857 3.542 ;
      RECT 24.685 3.349 24.771 3.528 ;
      RECT 24.66 3.337 24.685 3.519 ;
      RECT 24.59 3.327 24.66 3.512 ;
      RECT 24.545 3.315 24.59 3.503 ;
      RECT 24.485 3.302 24.545 3.495 ;
      RECT 24.48 3.294 24.485 3.49 ;
      RECT 24.445 3.289 24.48 3.488 ;
      RECT 24.39 3.28 24.445 3.481 ;
      RECT 24.35 3.269 24.39 3.473 ;
      RECT 24.335 3.262 24.35 3.469 ;
      RECT 24.315 3.255 24.33 3.466 ;
      RECT 24.3 3.245 24.315 3.464 ;
      RECT 24.285 3.232 24.3 3.461 ;
      RECT 24.26 3.215 24.285 3.457 ;
      RECT 24.245 3.197 24.26 3.454 ;
      RECT 24.22 3.15 24.245 3.452 ;
      RECT 24.196 3.15 24.22 3.449 ;
      RECT 24.11 3.15 24.196 3.441 ;
      RECT 24.07 3.15 24.11 3.433 ;
      RECT 23.935 3.197 23.965 3.465 ;
      RECT 25.615 2.78 25.875 3.04 ;
      RECT 25.575 2.78 25.875 2.918 ;
      RECT 25.54 2.78 25.875 2.903 ;
      RECT 25.485 2.78 25.875 2.883 ;
      RECT 25.405 2.59 25.685 2.87 ;
      RECT 25.405 2.772 25.755 2.87 ;
      RECT 25.405 2.715 25.74 2.87 ;
      RECT 25.405 2.662 25.69 2.87 ;
      RECT 23.235 2.59 23.43 3.375 ;
      RECT 23.315 1.205 23.43 3.375 ;
      RECT 23.17 3.115 23.23 3.375 ;
      RECT 24.54 2.635 24.8 2.895 ;
      RECT 23.225 2.59 23.43 2.87 ;
      RECT 24.535 2.645 24.8 2.83 ;
      RECT 24.25 2.62 24.26 2.77 ;
      RECT 23.485 1.205 23.565 1.55 ;
      RECT 23.22 1.205 23.43 1.55 ;
      RECT 24.525 2.645 24.535 2.829 ;
      RECT 24.515 2.644 24.525 2.826 ;
      RECT 24.506 2.643 24.515 2.824 ;
      RECT 24.42 2.639 24.506 2.814 ;
      RECT 24.346 2.631 24.42 2.796 ;
      RECT 24.26 2.624 24.346 2.779 ;
      RECT 24.2 2.62 24.25 2.769 ;
      RECT 24.165 2.619 24.2 2.766 ;
      RECT 24.11 2.619 24.165 2.768 ;
      RECT 24.075 2.619 24.11 2.772 ;
      RECT 23.989 2.618 24.075 2.779 ;
      RECT 23.903 2.617 23.989 2.789 ;
      RECT 23.817 2.616 23.903 2.8 ;
      RECT 23.731 2.616 23.817 2.81 ;
      RECT 23.645 2.615 23.731 2.82 ;
      RECT 23.61 2.615 23.645 2.86 ;
      RECT 23.605 2.615 23.61 2.903 ;
      RECT 23.58 2.615 23.605 2.92 ;
      RECT 23.505 2.615 23.58 2.935 ;
      RECT 23.485 2.59 23.505 2.948 ;
      RECT 23.48 1.205 23.485 2.958 ;
      RECT 23.455 1.205 23.48 3 ;
      RECT 23.43 1.205 23.455 3.078 ;
      RECT 23.23 2.997 23.235 3.375 ;
      RECT 22.565 2.949 22.58 3.405 ;
      RECT 22.56 3.021 22.666 3.403 ;
      RECT 22.58 2.115 22.715 3.401 ;
      RECT 22.565 2.965 22.72 3.4 ;
      RECT 22.565 3.015 22.725 3.398 ;
      RECT 22.55 3.08 22.725 3.397 ;
      RECT 22.56 3.072 22.73 3.394 ;
      RECT 22.54 3.12 22.73 3.389 ;
      RECT 22.54 3.12 22.745 3.386 ;
      RECT 22.535 3.12 22.745 3.383 ;
      RECT 22.51 3.12 22.77 3.38 ;
      RECT 22.58 2.115 22.74 2.768 ;
      RECT 22.575 2.115 22.74 2.74 ;
      RECT 22.57 2.115 22.74 2.568 ;
      RECT 22.57 2.115 22.76 2.508 ;
      RECT 22.525 2.115 22.785 2.375 ;
      RECT 22.005 2.59 22.285 2.87 ;
      RECT 21.995 2.605 22.285 2.865 ;
      RECT 21.95 2.667 22.285 2.863 ;
      RECT 22.025 2.582 22.19 2.87 ;
      RECT 22.025 2.567 22.146 2.87 ;
      RECT 22.06 2.56 22.146 2.87 ;
      RECT 21.525 3.71 21.805 3.99 ;
      RECT 21.485 3.672 21.78 3.783 ;
      RECT 21.47 3.622 21.76 3.678 ;
      RECT 21.415 3.385 21.675 3.645 ;
      RECT 21.415 3.587 21.755 3.645 ;
      RECT 21.415 3.527 21.75 3.645 ;
      RECT 21.415 3.477 21.73 3.645 ;
      RECT 21.415 3.457 21.725 3.645 ;
      RECT 21.415 3.435 21.72 3.645 ;
      RECT 21.415 3.42 21.69 3.645 ;
      RECT 17.145 6.225 17.465 6.545 ;
      RECT 17.175 5.695 17.345 6.545 ;
      RECT 17.175 5.695 17.35 6.045 ;
      RECT 17.175 5.695 18.15 5.87 ;
      RECT 17.975 1.965 18.15 5.87 ;
      RECT 17.92 1.965 18.27 2.315 ;
      RECT 17.945 6.655 18.27 6.98 ;
      RECT 16.83 6.745 18.27 6.915 ;
      RECT 16.83 2.395 16.99 6.915 ;
      RECT 17.145 2.365 17.465 2.685 ;
      RECT 16.83 2.395 17.465 2.565 ;
      RECT 16.09 5.84 16.44 6.19 ;
      RECT 16.165 2.705 16.34 6.19 ;
      RECT 16.1 2.705 16.45 3.055 ;
      RECT 15.5 1.14 15.875 1.51 ;
      RECT 7.42 0.96 7.795 1.33 ;
      RECT 5.985 0.96 6.36 1.33 ;
      RECT 5.985 1.08 15.805 1.25 ;
      RECT 10.105 4.36 15.785 4.53 ;
      RECT 15.615 3.425 15.785 4.53 ;
      RECT 9.915 3.6 9.94 4.53 ;
      RECT 10.17 3.71 10.2 3.99 ;
      RECT 9.875 3.6 9.94 3.86 ;
      RECT 15.525 3.43 15.875 3.78 ;
      RECT 9.705 2.225 9.74 2.485 ;
      RECT 9.48 2.225 9.54 2.485 ;
      RECT 10.16 3.69 10.17 3.99 ;
      RECT 10.155 3.65 10.16 3.99 ;
      RECT 10.14 3.605 10.155 3.99 ;
      RECT 10.135 3.57 10.14 3.99 ;
      RECT 10.13 3.55 10.135 3.99 ;
      RECT 10.105 3.487 10.13 3.99 ;
      RECT 10.1 3.425 10.105 4.53 ;
      RECT 10.08 3.375 10.1 4.53 ;
      RECT 10.07 3.305 10.08 4.53 ;
      RECT 10.025 3.245 10.07 4.53 ;
      RECT 9.94 3.206 10.025 4.53 ;
      RECT 9.935 3.197 9.94 3.57 ;
      RECT 9.925 3.196 9.935 3.553 ;
      RECT 9.9 3.177 9.925 3.523 ;
      RECT 9.895 3.152 9.9 3.502 ;
      RECT 9.885 3.13 9.895 3.493 ;
      RECT 9.88 3.101 9.885 3.483 ;
      RECT 9.84 3.027 9.88 3.455 ;
      RECT 9.82 2.928 9.84 3.42 ;
      RECT 9.805 2.864 9.82 3.403 ;
      RECT 9.775 2.788 9.805 3.375 ;
      RECT 9.755 2.703 9.775 3.348 ;
      RECT 9.715 2.599 9.755 3.255 ;
      RECT 9.71 2.52 9.715 3.163 ;
      RECT 9.705 2.503 9.71 3.14 ;
      RECT 9.7 2.225 9.705 3.12 ;
      RECT 9.67 2.225 9.7 3.058 ;
      RECT 9.665 2.225 9.67 2.99 ;
      RECT 9.655 2.225 9.665 2.955 ;
      RECT 9.645 2.225 9.655 2.92 ;
      RECT 9.58 2.225 9.645 2.775 ;
      RECT 9.575 2.225 9.58 2.645 ;
      RECT 9.545 2.225 9.575 2.578 ;
      RECT 9.54 2.225 9.545 2.503 ;
      RECT 13.875 2.16 14.135 2.42 ;
      RECT 13.87 2.16 14.135 2.368 ;
      RECT 13.865 2.16 14.135 2.338 ;
      RECT 13.84 2.03 14.12 2.31 ;
      RECT 1.7 6.995 1.99 7.345 ;
      RECT 1.7 7.055 3.01 7.225 ;
      RECT 2.84 6.685 3.01 7.225 ;
      RECT 13.34 6.605 13.69 6.955 ;
      RECT 2.84 6.685 13.69 6.855 ;
      RECT 12.88 3.71 13.16 3.99 ;
      RECT 12.92 3.665 13.185 3.925 ;
      RECT 12.91 3.7 13.185 3.925 ;
      RECT 12.915 3.685 13.16 3.99 ;
      RECT 12.92 3.662 13.13 3.99 ;
      RECT 12.92 3.66 13.115 3.99 ;
      RECT 12.96 3.65 13.115 3.99 ;
      RECT 12.93 3.655 13.115 3.99 ;
      RECT 12.96 3.647 13.06 3.99 ;
      RECT 12.985 3.64 13.06 3.99 ;
      RECT 12.965 3.642 13.06 3.99 ;
      RECT 12.295 3.155 12.555 3.415 ;
      RECT 12.345 3.147 12.535 3.415 ;
      RECT 12.35 3.067 12.535 3.415 ;
      RECT 12.47 2.455 12.535 3.415 ;
      RECT 12.375 2.852 12.535 3.415 ;
      RECT 12.45 2.54 12.535 3.415 ;
      RECT 12.485 2.165 12.621 2.893 ;
      RECT 12.43 2.662 12.621 2.893 ;
      RECT 12.445 2.602 12.535 3.415 ;
      RECT 12.485 2.165 12.645 2.558 ;
      RECT 12.485 2.165 12.655 2.455 ;
      RECT 12.475 2.165 12.735 2.425 ;
      RECT 11.88 3.71 12.16 3.99 ;
      RECT 11.9 3.67 12.16 3.99 ;
      RECT 11.54 3.625 11.645 3.885 ;
      RECT 11.395 2.115 11.485 2.375 ;
      RECT 11.935 3.18 11.94 3.22 ;
      RECT 11.93 3.17 11.935 3.305 ;
      RECT 11.925 3.16 11.93 3.398 ;
      RECT 11.915 3.14 11.925 3.454 ;
      RECT 11.835 3.068 11.915 3.534 ;
      RECT 11.87 3.712 11.88 3.937 ;
      RECT 11.865 3.709 11.87 3.932 ;
      RECT 11.85 3.706 11.865 3.925 ;
      RECT 11.815 3.7 11.85 3.907 ;
      RECT 11.83 3.003 11.835 3.608 ;
      RECT 11.81 2.954 11.83 3.623 ;
      RECT 11.8 3.687 11.815 3.89 ;
      RECT 11.805 2.896 11.81 3.638 ;
      RECT 11.8 2.874 11.805 3.648 ;
      RECT 11.765 2.784 11.8 3.885 ;
      RECT 11.75 2.662 11.765 3.885 ;
      RECT 11.745 2.615 11.75 3.885 ;
      RECT 11.72 2.54 11.745 3.885 ;
      RECT 11.705 2.455 11.72 3.885 ;
      RECT 11.7 2.402 11.705 3.885 ;
      RECT 11.695 2.382 11.7 3.885 ;
      RECT 11.69 2.357 11.695 3.119 ;
      RECT 11.675 3.317 11.695 3.885 ;
      RECT 11.685 2.335 11.69 3.096 ;
      RECT 11.675 2.287 11.685 3.061 ;
      RECT 11.67 2.25 11.675 3.027 ;
      RECT 11.67 3.397 11.675 3.885 ;
      RECT 11.655 2.227 11.67 2.982 ;
      RECT 11.65 3.495 11.67 3.885 ;
      RECT 11.6 2.115 11.655 2.824 ;
      RECT 11.645 3.617 11.65 3.885 ;
      RECT 11.585 2.115 11.6 2.663 ;
      RECT 11.58 2.115 11.585 2.615 ;
      RECT 11.575 2.115 11.58 2.603 ;
      RECT 11.53 2.115 11.575 2.54 ;
      RECT 11.505 2.115 11.53 2.458 ;
      RECT 11.49 2.115 11.505 2.41 ;
      RECT 11.485 2.115 11.49 2.38 ;
      RECT 10.81 3.565 10.855 3.825 ;
      RECT 10.715 2.1 10.86 2.36 ;
      RECT 11.22 2.722 11.23 2.813 ;
      RECT 11.205 2.66 11.22 2.869 ;
      RECT 11.2 2.607 11.205 2.915 ;
      RECT 11.15 2.554 11.2 3.041 ;
      RECT 11.145 2.509 11.15 3.188 ;
      RECT 11.135 2.497 11.145 3.23 ;
      RECT 11.1 2.461 11.135 3.335 ;
      RECT 11.095 2.429 11.1 3.441 ;
      RECT 11.08 2.411 11.095 3.486 ;
      RECT 11.075 2.394 11.08 2.72 ;
      RECT 11.07 2.775 11.08 3.543 ;
      RECT 11.065 2.38 11.075 2.693 ;
      RECT 11.06 2.83 11.07 3.825 ;
      RECT 11.055 2.366 11.065 2.678 ;
      RECT 11.055 2.88 11.06 3.825 ;
      RECT 11.04 2.343 11.055 2.658 ;
      RECT 11.02 3.002 11.055 3.825 ;
      RECT 11.035 2.325 11.04 2.64 ;
      RECT 11.03 2.317 11.035 2.63 ;
      RECT 11 2.285 11.03 2.594 ;
      RECT 11.01 3.13 11.02 3.825 ;
      RECT 11.005 3.157 11.01 3.825 ;
      RECT 11 3.207 11.005 3.825 ;
      RECT 10.99 2.251 11 2.559 ;
      RECT 10.95 3.275 11 3.825 ;
      RECT 10.975 2.228 10.99 2.535 ;
      RECT 10.95 2.1 10.975 2.498 ;
      RECT 10.945 2.1 10.95 2.47 ;
      RECT 10.915 3.375 10.95 3.825 ;
      RECT 10.94 2.1 10.945 2.463 ;
      RECT 10.935 2.1 10.94 2.453 ;
      RECT 10.92 2.1 10.935 2.438 ;
      RECT 10.905 2.1 10.92 2.41 ;
      RECT 10.87 3.48 10.915 3.825 ;
      RECT 10.89 2.1 10.905 2.383 ;
      RECT 10.86 2.1 10.89 2.368 ;
      RECT 10.855 3.552 10.87 3.825 ;
      RECT 10.78 2.635 10.82 2.895 ;
      RECT 10.555 2.582 10.56 2.84 ;
      RECT 6.51 2.06 6.77 2.32 ;
      RECT 6.51 2.085 6.785 2.3 ;
      RECT 8.9 1.91 8.905 2.055 ;
      RECT 10.77 2.63 10.78 2.895 ;
      RECT 10.75 2.622 10.77 2.895 ;
      RECT 10.732 2.618 10.75 2.895 ;
      RECT 10.646 2.607 10.732 2.895 ;
      RECT 10.56 2.59 10.646 2.895 ;
      RECT 10.505 2.577 10.555 2.825 ;
      RECT 10.471 2.569 10.505 2.8 ;
      RECT 10.385 2.558 10.471 2.765 ;
      RECT 10.35 2.535 10.385 2.73 ;
      RECT 10.34 2.497 10.35 2.716 ;
      RECT 10.335 2.47 10.34 2.712 ;
      RECT 10.33 2.457 10.335 2.709 ;
      RECT 10.32 2.437 10.33 2.705 ;
      RECT 10.315 2.412 10.32 2.701 ;
      RECT 10.29 2.367 10.315 2.695 ;
      RECT 10.28 2.308 10.29 2.687 ;
      RECT 10.27 2.276 10.28 2.678 ;
      RECT 10.25 2.228 10.27 2.658 ;
      RECT 10.245 2.188 10.25 2.628 ;
      RECT 10.23 2.162 10.245 2.602 ;
      RECT 10.225 2.14 10.23 2.578 ;
      RECT 10.21 2.112 10.225 2.554 ;
      RECT 10.195 2.085 10.21 2.518 ;
      RECT 10.18 2.062 10.195 2.48 ;
      RECT 10.175 2.052 10.18 2.455 ;
      RECT 10.165 2.045 10.175 2.438 ;
      RECT 10.15 2.032 10.165 2.408 ;
      RECT 10.145 2.022 10.15 2.383 ;
      RECT 10.14 2.017 10.145 2.37 ;
      RECT 10.13 2.01 10.14 2.35 ;
      RECT 10.125 2.003 10.13 2.335 ;
      RECT 10.1 1.996 10.125 2.293 ;
      RECT 10.085 1.986 10.1 2.243 ;
      RECT 10.075 1.981 10.085 2.213 ;
      RECT 10.065 1.977 10.075 2.188 ;
      RECT 10.05 1.974 10.065 2.178 ;
      RECT 10 1.971 10.05 2.163 ;
      RECT 9.98 1.969 10 2.148 ;
      RECT 9.931 1.967 9.98 2.143 ;
      RECT 9.845 1.963 9.931 2.138 ;
      RECT 9.806 1.96 9.845 2.134 ;
      RECT 9.72 1.956 9.806 2.129 ;
      RECT 9.67 1.953 9.72 2.123 ;
      RECT 9.621 1.95 9.67 2.118 ;
      RECT 9.535 1.947 9.621 2.113 ;
      RECT 9.531 1.945 9.535 2.11 ;
      RECT 9.445 1.942 9.531 2.105 ;
      RECT 9.396 1.938 9.445 2.098 ;
      RECT 9.31 1.935 9.396 2.093 ;
      RECT 9.286 1.932 9.31 2.089 ;
      RECT 9.2 1.93 9.286 2.084 ;
      RECT 9.135 1.926 9.2 2.077 ;
      RECT 9.132 1.925 9.135 2.074 ;
      RECT 9.046 1.922 9.132 2.071 ;
      RECT 8.96 1.916 9.046 2.064 ;
      RECT 8.93 1.912 8.96 2.06 ;
      RECT 8.905 1.91 8.93 2.058 ;
      RECT 8.85 1.907 8.9 2.055 ;
      RECT 8.77 1.906 8.85 2.055 ;
      RECT 8.715 1.908 8.77 2.058 ;
      RECT 8.7 1.909 8.715 2.062 ;
      RECT 8.645 1.917 8.7 2.072 ;
      RECT 8.615 1.925 8.645 2.085 ;
      RECT 8.596 1.926 8.615 2.091 ;
      RECT 8.51 1.929 8.596 2.096 ;
      RECT 8.44 1.934 8.51 2.105 ;
      RECT 8.421 1.937 8.44 2.111 ;
      RECT 8.335 1.941 8.421 2.116 ;
      RECT 8.295 1.945 8.335 2.123 ;
      RECT 8.286 1.947 8.295 2.126 ;
      RECT 8.2 1.951 8.286 2.131 ;
      RECT 8.197 1.954 8.2 2.135 ;
      RECT 8.111 1.957 8.197 2.139 ;
      RECT 8.025 1.963 8.111 2.147 ;
      RECT 8.001 1.967 8.025 2.151 ;
      RECT 7.915 1.971 8.001 2.156 ;
      RECT 7.87 1.976 7.915 2.163 ;
      RECT 7.79 1.981 7.87 2.17 ;
      RECT 7.71 1.987 7.79 2.185 ;
      RECT 7.685 1.991 7.71 2.198 ;
      RECT 7.62 1.994 7.685 2.21 ;
      RECT 7.565 1.999 7.62 2.225 ;
      RECT 7.535 2.002 7.565 2.243 ;
      RECT 7.525 2.004 7.535 2.256 ;
      RECT 7.465 2.019 7.525 2.266 ;
      RECT 7.45 2.036 7.465 2.275 ;
      RECT 7.445 2.045 7.45 2.275 ;
      RECT 7.435 2.055 7.445 2.275 ;
      RECT 7.425 2.072 7.435 2.275 ;
      RECT 7.405 2.082 7.425 2.276 ;
      RECT 7.36 2.092 7.405 2.277 ;
      RECT 7.325 2.101 7.36 2.279 ;
      RECT 7.26 2.106 7.325 2.281 ;
      RECT 7.18 2.107 7.26 2.284 ;
      RECT 7.176 2.105 7.18 2.285 ;
      RECT 7.09 2.102 7.176 2.287 ;
      RECT 7.043 2.099 7.09 2.289 ;
      RECT 6.957 2.095 7.043 2.292 ;
      RECT 6.871 2.091 6.957 2.295 ;
      RECT 6.785 2.087 6.871 2.299 ;
      RECT 8.72 3.15 9 3.43 ;
      RECT 8.76 3.13 9.02 3.39 ;
      RECT 8.75 3.14 9.02 3.39 ;
      RECT 8.76 3.067 8.975 3.43 ;
      RECT 8.815 2.99 8.97 3.43 ;
      RECT 8.82 2.775 8.97 3.43 ;
      RECT 8.81 2.577 8.96 2.828 ;
      RECT 8.8 2.577 8.96 2.695 ;
      RECT 8.795 2.455 8.955 2.598 ;
      RECT 8.78 2.455 8.955 2.503 ;
      RECT 8.775 2.165 8.95 2.48 ;
      RECT 8.76 2.165 8.95 2.45 ;
      RECT 8.72 2.165 8.98 2.425 ;
      RECT 8.63 3.635 8.71 3.895 ;
      RECT 8.035 2.355 8.04 2.62 ;
      RECT 7.915 2.355 8.04 2.615 ;
      RECT 8.59 3.6 8.63 3.895 ;
      RECT 8.545 3.522 8.59 3.895 ;
      RECT 8.525 3.45 8.545 3.895 ;
      RECT 8.515 3.402 8.525 3.895 ;
      RECT 8.48 3.335 8.515 3.895 ;
      RECT 8.45 3.235 8.48 3.895 ;
      RECT 8.43 3.16 8.45 3.695 ;
      RECT 8.42 3.11 8.43 3.65 ;
      RECT 8.415 3.087 8.42 3.623 ;
      RECT 8.41 3.072 8.415 3.61 ;
      RECT 8.405 3.057 8.41 3.588 ;
      RECT 8.4 3.042 8.405 3.57 ;
      RECT 8.375 2.997 8.4 3.525 ;
      RECT 8.365 2.945 8.375 3.468 ;
      RECT 8.355 2.915 8.365 3.435 ;
      RECT 8.345 2.88 8.355 3.403 ;
      RECT 8.31 2.812 8.345 3.335 ;
      RECT 8.305 2.751 8.31 3.27 ;
      RECT 8.295 2.739 8.305 3.25 ;
      RECT 8.29 2.727 8.295 3.23 ;
      RECT 8.285 2.719 8.29 3.218 ;
      RECT 8.28 2.711 8.285 3.198 ;
      RECT 8.27 2.699 8.28 3.17 ;
      RECT 8.26 2.683 8.27 3.14 ;
      RECT 8.235 2.655 8.26 3.078 ;
      RECT 8.225 2.626 8.235 3.023 ;
      RECT 8.21 2.605 8.225 2.983 ;
      RECT 8.205 2.589 8.21 2.955 ;
      RECT 8.2 2.577 8.205 2.945 ;
      RECT 8.195 2.572 8.2 2.918 ;
      RECT 8.19 2.565 8.195 2.905 ;
      RECT 8.175 2.548 8.19 2.878 ;
      RECT 8.165 2.355 8.175 2.838 ;
      RECT 8.155 2.355 8.165 2.805 ;
      RECT 8.145 2.355 8.155 2.78 ;
      RECT 8.075 2.355 8.145 2.715 ;
      RECT 8.065 2.355 8.075 2.663 ;
      RECT 8.05 2.355 8.065 2.645 ;
      RECT 8.04 2.355 8.05 2.63 ;
      RECT 7.87 3.225 8.13 3.485 ;
      RECT 6.405 3.26 6.41 3.467 ;
      RECT 6.04 3.15 6.115 3.465 ;
      RECT 5.855 3.205 6.01 3.465 ;
      RECT 6.04 3.15 6.145 3.43 ;
      RECT 7.855 3.322 7.87 3.483 ;
      RECT 7.83 3.33 7.855 3.488 ;
      RECT 7.805 3.337 7.83 3.493 ;
      RECT 7.742 3.348 7.805 3.502 ;
      RECT 7.656 3.367 7.742 3.519 ;
      RECT 7.57 3.389 7.656 3.538 ;
      RECT 7.555 3.402 7.57 3.549 ;
      RECT 7.515 3.41 7.555 3.556 ;
      RECT 7.495 3.415 7.515 3.563 ;
      RECT 7.457 3.416 7.495 3.566 ;
      RECT 7.371 3.419 7.457 3.567 ;
      RECT 7.285 3.423 7.371 3.568 ;
      RECT 7.236 3.425 7.285 3.57 ;
      RECT 7.15 3.425 7.236 3.572 ;
      RECT 7.11 3.42 7.15 3.574 ;
      RECT 7.1 3.414 7.11 3.575 ;
      RECT 7.06 3.409 7.1 3.572 ;
      RECT 7.05 3.402 7.06 3.568 ;
      RECT 7.035 3.398 7.05 3.566 ;
      RECT 7.018 3.394 7.035 3.564 ;
      RECT 6.932 3.384 7.018 3.556 ;
      RECT 6.846 3.366 6.932 3.542 ;
      RECT 6.76 3.349 6.846 3.528 ;
      RECT 6.735 3.337 6.76 3.519 ;
      RECT 6.665 3.327 6.735 3.512 ;
      RECT 6.62 3.315 6.665 3.503 ;
      RECT 6.56 3.302 6.62 3.495 ;
      RECT 6.555 3.294 6.56 3.49 ;
      RECT 6.52 3.289 6.555 3.488 ;
      RECT 6.465 3.28 6.52 3.481 ;
      RECT 6.425 3.269 6.465 3.473 ;
      RECT 6.41 3.262 6.425 3.469 ;
      RECT 6.39 3.255 6.405 3.466 ;
      RECT 6.375 3.245 6.39 3.464 ;
      RECT 6.36 3.232 6.375 3.461 ;
      RECT 6.335 3.215 6.36 3.457 ;
      RECT 6.32 3.197 6.335 3.454 ;
      RECT 6.295 3.15 6.32 3.452 ;
      RECT 6.271 3.15 6.295 3.449 ;
      RECT 6.185 3.15 6.271 3.441 ;
      RECT 6.145 3.15 6.185 3.433 ;
      RECT 6.01 3.197 6.04 3.465 ;
      RECT 7.69 2.78 7.95 3.04 ;
      RECT 7.65 2.78 7.95 2.918 ;
      RECT 7.615 2.78 7.95 2.903 ;
      RECT 7.56 2.78 7.95 2.883 ;
      RECT 7.48 2.59 7.76 2.87 ;
      RECT 7.48 2.772 7.83 2.87 ;
      RECT 7.48 2.715 7.815 2.87 ;
      RECT 7.48 2.662 7.765 2.87 ;
      RECT 5.31 2.59 5.505 3.375 ;
      RECT 5.39 1.205 5.505 3.375 ;
      RECT 5.245 3.115 5.305 3.375 ;
      RECT 6.615 2.635 6.875 2.895 ;
      RECT 5.3 2.59 5.505 2.87 ;
      RECT 6.61 2.645 6.875 2.83 ;
      RECT 6.325 2.62 6.335 2.77 ;
      RECT 5.56 1.205 5.64 1.55 ;
      RECT 5.295 1.205 5.505 1.55 ;
      RECT 6.6 2.645 6.61 2.829 ;
      RECT 6.59 2.644 6.6 2.826 ;
      RECT 6.581 2.643 6.59 2.824 ;
      RECT 6.495 2.639 6.581 2.814 ;
      RECT 6.421 2.631 6.495 2.796 ;
      RECT 6.335 2.624 6.421 2.779 ;
      RECT 6.275 2.62 6.325 2.769 ;
      RECT 6.24 2.619 6.275 2.766 ;
      RECT 6.185 2.619 6.24 2.768 ;
      RECT 6.15 2.619 6.185 2.772 ;
      RECT 6.064 2.618 6.15 2.779 ;
      RECT 5.978 2.617 6.064 2.789 ;
      RECT 5.892 2.616 5.978 2.8 ;
      RECT 5.806 2.616 5.892 2.81 ;
      RECT 5.72 2.615 5.806 2.82 ;
      RECT 5.685 2.615 5.72 2.86 ;
      RECT 5.68 2.615 5.685 2.903 ;
      RECT 5.655 2.615 5.68 2.92 ;
      RECT 5.58 2.615 5.655 2.935 ;
      RECT 5.56 2.59 5.58 2.948 ;
      RECT 5.555 1.205 5.56 2.958 ;
      RECT 5.53 1.205 5.555 3 ;
      RECT 5.505 1.205 5.53 3.078 ;
      RECT 5.305 2.997 5.31 3.375 ;
      RECT 4.64 2.949 4.655 3.405 ;
      RECT 4.635 3.021 4.741 3.403 ;
      RECT 4.655 2.115 4.79 3.401 ;
      RECT 4.64 2.965 4.795 3.4 ;
      RECT 4.64 3.015 4.8 3.398 ;
      RECT 4.625 3.08 4.8 3.397 ;
      RECT 4.635 3.072 4.805 3.394 ;
      RECT 4.615 3.12 4.805 3.389 ;
      RECT 4.615 3.12 4.82 3.386 ;
      RECT 4.61 3.12 4.82 3.383 ;
      RECT 4.585 3.12 4.845 3.38 ;
      RECT 4.655 2.115 4.815 2.768 ;
      RECT 4.65 2.115 4.815 2.74 ;
      RECT 4.645 2.115 4.815 2.568 ;
      RECT 4.645 2.115 4.835 2.508 ;
      RECT 4.6 2.115 4.86 2.375 ;
      RECT 4.08 2.59 4.36 2.87 ;
      RECT 4.07 2.605 4.36 2.865 ;
      RECT 4.025 2.667 4.36 2.863 ;
      RECT 4.1 2.582 4.265 2.87 ;
      RECT 4.1 2.567 4.221 2.87 ;
      RECT 4.135 2.56 4.221 2.87 ;
      RECT 3.6 3.71 3.88 3.99 ;
      RECT 3.56 3.672 3.855 3.783 ;
      RECT 3.545 3.622 3.835 3.678 ;
      RECT 3.49 3.385 3.75 3.645 ;
      RECT 3.49 3.587 3.83 3.645 ;
      RECT 3.49 3.527 3.825 3.645 ;
      RECT 3.49 3.477 3.805 3.645 ;
      RECT 3.49 3.457 3.8 3.645 ;
      RECT 3.49 3.435 3.795 3.645 ;
      RECT 3.49 3.42 3.765 3.645 ;
      RECT 84.38 7.055 84.755 7.425 ;
      RECT 75.715 0.93 76.09 1.3 ;
      RECT 66.455 7.055 66.83 7.425 ;
      RECT 57.79 0.93 58.165 1.3 ;
      RECT 48.53 7.055 48.905 7.425 ;
      RECT 39.865 0.93 40.24 1.3 ;
      RECT 30.605 7.055 30.98 7.425 ;
      RECT 21.94 0.93 22.315 1.3 ;
      RECT 12.68 7.055 13.055 7.425 ;
      RECT 4.015 0.93 4.39 1.3 ;
    LAYER via1 ;
      RECT 92.1 7.375 92.25 7.525 ;
      RECT 89.735 6.74 89.885 6.89 ;
      RECT 89.72 2.065 89.87 2.215 ;
      RECT 88.93 2.45 89.08 2.6 ;
      RECT 88.93 6.325 89.08 6.475 ;
      RECT 87.9 2.805 88.05 2.955 ;
      RECT 87.89 5.94 88.04 6.09 ;
      RECT 87.325 3.53 87.475 3.68 ;
      RECT 87.315 1.25 87.465 1.4 ;
      RECT 85.63 2.215 85.78 2.365 ;
      RECT 85.4 6.71 85.55 6.86 ;
      RECT 84.68 3.72 84.83 3.87 ;
      RECT 84.495 7.165 84.645 7.315 ;
      RECT 84.23 2.22 84.38 2.37 ;
      RECT 84.05 3.21 84.2 3.36 ;
      RECT 83.655 3.725 83.805 3.875 ;
      RECT 83.295 3.68 83.445 3.83 ;
      RECT 83.15 2.17 83.3 2.32 ;
      RECT 82.565 3.62 82.715 3.77 ;
      RECT 82.47 2.155 82.62 2.305 ;
      RECT 82.315 2.69 82.465 2.84 ;
      RECT 81.63 3.655 81.78 3.805 ;
      RECT 81.235 2.28 81.385 2.43 ;
      RECT 80.515 3.185 80.665 3.335 ;
      RECT 80.475 2.22 80.625 2.37 ;
      RECT 80.205 3.69 80.355 3.84 ;
      RECT 79.67 2.41 79.82 2.56 ;
      RECT 79.625 3.28 79.775 3.43 ;
      RECT 79.445 2.835 79.595 2.985 ;
      RECT 78.37 2.69 78.52 2.84 ;
      RECT 78.265 2.115 78.415 2.265 ;
      RECT 77.61 3.26 77.76 3.41 ;
      RECT 77.09 1.3 77.24 1.45 ;
      RECT 77 3.17 77.15 3.32 ;
      RECT 76.355 2.17 76.505 2.32 ;
      RECT 76.34 3.175 76.49 3.325 ;
      RECT 75.825 2.66 75.975 2.81 ;
      RECT 75.245 3.44 75.395 3.59 ;
      RECT 74.155 6.755 74.305 6.905 ;
      RECT 71.81 6.74 71.96 6.89 ;
      RECT 71.795 2.065 71.945 2.215 ;
      RECT 71.005 2.45 71.155 2.6 ;
      RECT 71.005 6.325 71.155 6.475 ;
      RECT 69.975 2.805 70.125 2.955 ;
      RECT 69.965 5.94 70.115 6.09 ;
      RECT 69.4 3.53 69.55 3.68 ;
      RECT 69.39 1.25 69.54 1.4 ;
      RECT 67.705 2.215 67.855 2.365 ;
      RECT 67.195 6.71 67.345 6.86 ;
      RECT 66.755 3.72 66.905 3.87 ;
      RECT 66.57 7.165 66.72 7.315 ;
      RECT 66.305 2.22 66.455 2.37 ;
      RECT 66.125 3.21 66.275 3.36 ;
      RECT 65.73 3.725 65.88 3.875 ;
      RECT 65.37 3.68 65.52 3.83 ;
      RECT 65.225 2.17 65.375 2.32 ;
      RECT 64.64 3.62 64.79 3.77 ;
      RECT 64.545 2.155 64.695 2.305 ;
      RECT 64.39 2.69 64.54 2.84 ;
      RECT 63.705 3.655 63.855 3.805 ;
      RECT 63.31 2.28 63.46 2.43 ;
      RECT 62.59 3.185 62.74 3.335 ;
      RECT 62.55 2.22 62.7 2.37 ;
      RECT 62.28 3.69 62.43 3.84 ;
      RECT 61.745 2.41 61.895 2.56 ;
      RECT 61.7 3.28 61.85 3.43 ;
      RECT 61.52 2.835 61.67 2.985 ;
      RECT 60.445 2.69 60.595 2.84 ;
      RECT 60.34 2.115 60.49 2.265 ;
      RECT 59.685 3.26 59.835 3.41 ;
      RECT 59.165 1.3 59.315 1.45 ;
      RECT 59.075 3.17 59.225 3.32 ;
      RECT 58.43 2.17 58.58 2.32 ;
      RECT 58.415 3.175 58.565 3.325 ;
      RECT 57.9 2.66 58.05 2.81 ;
      RECT 57.32 3.44 57.47 3.59 ;
      RECT 56.23 6.755 56.38 6.905 ;
      RECT 53.885 6.74 54.035 6.89 ;
      RECT 53.87 2.065 54.02 2.215 ;
      RECT 53.08 2.45 53.23 2.6 ;
      RECT 53.08 6.325 53.23 6.475 ;
      RECT 52.05 2.805 52.2 2.955 ;
      RECT 52.04 5.94 52.19 6.09 ;
      RECT 51.475 3.53 51.625 3.68 ;
      RECT 51.465 1.25 51.615 1.4 ;
      RECT 49.78 2.215 49.93 2.365 ;
      RECT 49.325 6.715 49.475 6.865 ;
      RECT 48.83 3.72 48.98 3.87 ;
      RECT 48.645 7.165 48.795 7.315 ;
      RECT 48.38 2.22 48.53 2.37 ;
      RECT 48.2 3.21 48.35 3.36 ;
      RECT 47.805 3.725 47.955 3.875 ;
      RECT 47.445 3.68 47.595 3.83 ;
      RECT 47.3 2.17 47.45 2.32 ;
      RECT 46.715 3.62 46.865 3.77 ;
      RECT 46.62 2.155 46.77 2.305 ;
      RECT 46.465 2.69 46.615 2.84 ;
      RECT 45.78 3.655 45.93 3.805 ;
      RECT 45.385 2.28 45.535 2.43 ;
      RECT 44.665 3.185 44.815 3.335 ;
      RECT 44.625 2.22 44.775 2.37 ;
      RECT 44.355 3.69 44.505 3.84 ;
      RECT 43.82 2.41 43.97 2.56 ;
      RECT 43.775 3.28 43.925 3.43 ;
      RECT 43.595 2.835 43.745 2.985 ;
      RECT 42.52 2.69 42.67 2.84 ;
      RECT 42.415 2.115 42.565 2.265 ;
      RECT 41.76 3.26 41.91 3.41 ;
      RECT 41.24 1.3 41.39 1.45 ;
      RECT 41.15 3.17 41.3 3.32 ;
      RECT 40.505 2.17 40.655 2.32 ;
      RECT 40.49 3.175 40.64 3.325 ;
      RECT 39.975 2.66 40.125 2.81 ;
      RECT 39.395 3.44 39.545 3.59 ;
      RECT 38.35 6.76 38.5 6.91 ;
      RECT 35.96 6.74 36.11 6.89 ;
      RECT 35.945 2.065 36.095 2.215 ;
      RECT 35.155 2.45 35.305 2.6 ;
      RECT 35.155 6.325 35.305 6.475 ;
      RECT 34.125 2.805 34.275 2.955 ;
      RECT 34.115 5.94 34.265 6.09 ;
      RECT 33.55 3.53 33.7 3.68 ;
      RECT 33.54 1.25 33.69 1.4 ;
      RECT 31.855 2.215 32.005 2.365 ;
      RECT 31.395 6.71 31.545 6.86 ;
      RECT 30.905 3.72 31.055 3.87 ;
      RECT 30.72 7.165 30.87 7.315 ;
      RECT 30.455 2.22 30.605 2.37 ;
      RECT 30.275 3.21 30.425 3.36 ;
      RECT 29.88 3.725 30.03 3.875 ;
      RECT 29.52 3.68 29.67 3.83 ;
      RECT 29.375 2.17 29.525 2.32 ;
      RECT 28.79 3.62 28.94 3.77 ;
      RECT 28.695 2.155 28.845 2.305 ;
      RECT 28.54 2.69 28.69 2.84 ;
      RECT 27.855 3.655 28.005 3.805 ;
      RECT 27.46 2.28 27.61 2.43 ;
      RECT 26.74 3.185 26.89 3.335 ;
      RECT 26.7 2.22 26.85 2.37 ;
      RECT 26.43 3.69 26.58 3.84 ;
      RECT 25.895 2.41 26.045 2.56 ;
      RECT 25.85 3.28 26 3.43 ;
      RECT 25.67 2.835 25.82 2.985 ;
      RECT 24.595 2.69 24.745 2.84 ;
      RECT 24.49 2.115 24.64 2.265 ;
      RECT 23.835 3.26 23.985 3.41 ;
      RECT 23.315 1.3 23.465 1.45 ;
      RECT 23.225 3.17 23.375 3.32 ;
      RECT 22.58 2.17 22.73 2.32 ;
      RECT 22.565 3.175 22.715 3.325 ;
      RECT 22.05 2.66 22.2 2.81 ;
      RECT 21.47 3.44 21.62 3.59 ;
      RECT 20.425 6.755 20.575 6.905 ;
      RECT 18.035 6.74 18.185 6.89 ;
      RECT 18.02 2.065 18.17 2.215 ;
      RECT 17.23 2.45 17.38 2.6 ;
      RECT 17.23 6.325 17.38 6.475 ;
      RECT 16.2 2.805 16.35 2.955 ;
      RECT 16.19 5.94 16.34 6.09 ;
      RECT 15.625 3.53 15.775 3.68 ;
      RECT 15.615 1.25 15.765 1.4 ;
      RECT 13.93 2.215 14.08 2.365 ;
      RECT 13.44 6.705 13.59 6.855 ;
      RECT 12.98 3.72 13.13 3.87 ;
      RECT 12.795 7.165 12.945 7.315 ;
      RECT 12.53 2.22 12.68 2.37 ;
      RECT 12.35 3.21 12.5 3.36 ;
      RECT 11.955 3.725 12.105 3.875 ;
      RECT 11.595 3.68 11.745 3.83 ;
      RECT 11.45 2.17 11.6 2.32 ;
      RECT 10.865 3.62 11.015 3.77 ;
      RECT 10.77 2.155 10.92 2.305 ;
      RECT 10.615 2.69 10.765 2.84 ;
      RECT 9.93 3.655 10.08 3.805 ;
      RECT 9.535 2.28 9.685 2.43 ;
      RECT 8.815 3.185 8.965 3.335 ;
      RECT 8.775 2.22 8.925 2.37 ;
      RECT 8.505 3.69 8.655 3.84 ;
      RECT 7.97 2.41 8.12 2.56 ;
      RECT 7.925 3.28 8.075 3.43 ;
      RECT 7.745 2.835 7.895 2.985 ;
      RECT 6.67 2.69 6.82 2.84 ;
      RECT 6.565 2.115 6.715 2.265 ;
      RECT 5.91 3.26 6.06 3.41 ;
      RECT 5.39 1.3 5.54 1.45 ;
      RECT 5.3 3.17 5.45 3.32 ;
      RECT 4.655 2.17 4.805 2.32 ;
      RECT 4.64 3.175 4.79 3.325 ;
      RECT 4.125 2.66 4.275 2.81 ;
      RECT 3.545 3.44 3.695 3.59 ;
      RECT 1.77 7.095 1.92 7.245 ;
      RECT 1.395 6.355 1.545 6.505 ;
    LAYER met1 ;
      RECT 75.025 1.285 86.985 1.89 ;
      RECT 79.45 0 86.985 1.89 ;
      RECT 57.1 1.285 69.06 1.89 ;
      RECT 61.525 0 69.06 1.89 ;
      RECT 39.175 1.285 51.135 1.89 ;
      RECT 43.6 0 51.135 1.89 ;
      RECT 21.25 1.285 33.21 1.89 ;
      RECT 25.675 0 33.21 1.89 ;
      RECT 3.325 1.285 15.285 1.89 ;
      RECT 7.75 0 15.285 1.89 ;
      RECT 75.02 0 75.765 1.68 ;
      RECT 57.095 0 57.84 1.68 ;
      RECT 39.17 0 39.915 1.68 ;
      RECT 21.245 0 21.99 1.68 ;
      RECT 3.32 0 4.065 1.68 ;
      RECT 78.015 0 79.17 1.89 ;
      RECT 75.02 1.255 77.735 1.68 ;
      RECT 76.045 0 77.735 1.89 ;
      RECT 60.09 0 61.245 1.89 ;
      RECT 57.095 1.255 59.81 1.68 ;
      RECT 58.12 0 59.81 1.89 ;
      RECT 42.165 0 43.32 1.89 ;
      RECT 39.17 1.255 41.885 1.68 ;
      RECT 40.195 0 41.885 1.89 ;
      RECT 24.24 0 25.395 1.89 ;
      RECT 21.245 1.255 23.96 1.68 ;
      RECT 22.27 0 23.96 1.89 ;
      RECT 6.315 0 7.47 1.89 ;
      RECT 3.32 1.255 6.035 1.68 ;
      RECT 4.345 0 6.035 1.89 ;
      RECT 76.045 0 86.985 1.005 ;
      RECT 58.12 0 69.06 1.005 ;
      RECT 40.195 0 51.135 1.005 ;
      RECT 22.27 0 33.21 1.005 ;
      RECT 4.345 0 15.285 1.005 ;
      RECT 75.02 0 86.985 0.975 ;
      RECT 57.095 0 69.06 0.975 ;
      RECT 39.17 0 51.135 0.975 ;
      RECT 21.245 0 33.21 0.975 ;
      RECT 3.32 0 15.285 0.975 ;
      RECT 0 0 92.575 0.305 ;
      RECT 0 4.285 92.575 4.745 ;
      RECT 75.025 4.135 92.575 4.745 ;
      RECT 57.1 4.135 74.65 4.745 ;
      RECT 39.175 4.135 56.725 4.745 ;
      RECT 21.25 4.135 38.8 4.745 ;
      RECT 3.325 4.135 20.875 4.745 ;
      RECT 75.025 4.13 86.985 4.745 ;
      RECT 57.1 4.13 69.06 4.745 ;
      RECT 39.175 4.13 51.135 4.745 ;
      RECT 21.25 4.13 33.21 4.745 ;
      RECT 3.325 4.13 15.285 4.745 ;
      RECT 0 8.575 92.575 8.88 ;
      RECT 83.72 6.315 83.89 8.88 ;
      RECT 65.795 6.315 65.965 8.88 ;
      RECT 47.87 6.315 48.04 8.88 ;
      RECT 29.945 6.315 30.115 8.88 ;
      RECT 12.02 6.315 12.19 8.88 ;
      RECT 84.055 6.285 84.345 6.515 ;
      RECT 66.13 6.285 66.42 6.515 ;
      RECT 48.205 6.285 48.495 6.515 ;
      RECT 30.28 6.285 30.57 6.515 ;
      RECT 12.355 6.285 12.645 6.515 ;
      RECT 83.72 6.315 84.345 6.485 ;
      RECT 65.795 6.315 66.42 6.485 ;
      RECT 47.87 6.315 48.495 6.485 ;
      RECT 29.945 6.315 30.57 6.485 ;
      RECT 12.02 6.315 12.645 6.485 ;
      RECT 91.975 7.765 92.265 7.995 ;
      RECT 92.035 6.285 92.205 7.995 ;
      RECT 92 7.275 92.35 7.625 ;
      RECT 91.975 6.285 92.265 6.515 ;
      RECT 91.975 2.365 92.265 2.595 ;
      RECT 92.035 0.885 92.205 2.595 ;
      RECT 91.975 0.885 92.265 1.115 ;
      RECT 91.565 2.735 91.895 2.965 ;
      RECT 91.565 2.765 92.065 2.935 ;
      RECT 91.565 2.395 91.755 2.965 ;
      RECT 90.985 2.365 91.275 2.595 ;
      RECT 90.985 2.395 91.755 2.565 ;
      RECT 91.045 0.885 91.215 2.595 ;
      RECT 90.985 0.885 91.275 1.115 ;
      RECT 90.985 7.765 91.275 7.995 ;
      RECT 91.045 6.285 91.215 7.995 ;
      RECT 90.985 6.285 91.275 6.515 ;
      RECT 90.985 6.325 91.835 6.485 ;
      RECT 91.665 5.915 91.835 6.485 ;
      RECT 90.985 6.32 91.375 6.485 ;
      RECT 91.605 5.915 91.895 6.145 ;
      RECT 91.605 5.945 92.065 6.115 ;
      RECT 90.615 2.735 90.905 2.965 ;
      RECT 90.615 2.765 91.075 2.935 ;
      RECT 90.675 1.655 90.84 2.965 ;
      RECT 89.19 1.625 89.48 1.855 ;
      RECT 89.19 1.655 90.84 1.825 ;
      RECT 89.25 0.885 89.42 1.855 ;
      RECT 89.19 0.885 89.48 1.115 ;
      RECT 89.19 7.765 89.48 7.995 ;
      RECT 89.25 7.025 89.42 7.995 ;
      RECT 89.25 7.12 90.84 7.29 ;
      RECT 90.67 5.915 90.84 7.29 ;
      RECT 89.19 7.025 89.48 7.255 ;
      RECT 90.615 5.915 90.905 6.145 ;
      RECT 90.615 5.945 91.075 6.115 ;
      RECT 87.225 3.43 87.575 3.78 ;
      RECT 87.315 2.025 87.485 3.78 ;
      RECT 89.62 1.965 89.97 2.315 ;
      RECT 87.315 2.025 88.935 2.2 ;
      RECT 87.315 2.025 89.97 2.195 ;
      RECT 89.645 6.655 89.97 6.98 ;
      RECT 85.3 6.61 85.65 6.96 ;
      RECT 89.62 6.655 89.97 6.885 ;
      RECT 84.86 6.655 85.15 6.885 ;
      RECT 84.69 6.685 89.97 6.855 ;
      RECT 88.845 2.365 89.165 2.685 ;
      RECT 88.815 2.365 89.165 2.595 ;
      RECT 88.645 2.395 89.165 2.565 ;
      RECT 88.845 6.225 89.165 6.545 ;
      RECT 88.815 6.285 89.165 6.515 ;
      RECT 88.645 6.315 89.165 6.485 ;
      RECT 87.8 2.705 88.15 3.055 ;
      RECT 87.8 2.765 88.28 2.935 ;
      RECT 87.79 5.84 88.14 6.19 ;
      RECT 83.06 5.915 83.35 6.145 ;
      RECT 83.06 5.945 88.28 6.115 ;
      RECT 84.625 3.665 84.665 3.925 ;
      RECT 84.665 3.645 84.67 3.655 ;
      RECT 85.995 2.89 86.005 3.111 ;
      RECT 85.925 2.885 85.995 3.236 ;
      RECT 85.915 2.885 85.925 3.363 ;
      RECT 85.89 2.885 85.915 3.41 ;
      RECT 85.865 2.885 85.89 3.488 ;
      RECT 85.845 2.885 85.865 3.558 ;
      RECT 85.82 2.885 85.845 3.598 ;
      RECT 85.81 2.885 85.82 3.618 ;
      RECT 85.8 2.887 85.81 3.626 ;
      RECT 85.795 2.892 85.8 3.083 ;
      RECT 85.795 3.092 85.8 3.627 ;
      RECT 85.79 3.137 85.795 3.628 ;
      RECT 85.78 3.202 85.79 3.629 ;
      RECT 85.77 3.297 85.78 3.631 ;
      RECT 85.765 3.35 85.77 3.633 ;
      RECT 85.76 3.37 85.765 3.634 ;
      RECT 85.705 3.395 85.76 3.64 ;
      RECT 85.665 3.43 85.705 3.649 ;
      RECT 85.655 3.447 85.665 3.654 ;
      RECT 85.646 3.453 85.655 3.656 ;
      RECT 85.56 3.491 85.646 3.667 ;
      RECT 85.555 3.53 85.56 3.677 ;
      RECT 85.48 3.537 85.555 3.687 ;
      RECT 85.46 3.547 85.48 3.698 ;
      RECT 85.43 3.554 85.46 3.706 ;
      RECT 85.405 3.561 85.43 3.713 ;
      RECT 85.381 3.567 85.405 3.718 ;
      RECT 85.295 3.58 85.381 3.73 ;
      RECT 85.217 3.587 85.295 3.748 ;
      RECT 85.131 3.582 85.217 3.766 ;
      RECT 85.045 3.577 85.131 3.786 ;
      RECT 84.965 3.571 85.045 3.803 ;
      RECT 84.9 3.567 84.965 3.832 ;
      RECT 84.895 3.281 84.9 3.305 ;
      RECT 84.885 3.557 84.9 3.86 ;
      RECT 84.89 3.275 84.895 3.345 ;
      RECT 84.885 3.269 84.89 3.415 ;
      RECT 84.88 3.263 84.885 3.493 ;
      RECT 84.88 3.54 84.885 3.925 ;
      RECT 84.872 3.26 84.88 3.925 ;
      RECT 84.786 3.258 84.872 3.925 ;
      RECT 84.7 3.256 84.786 3.925 ;
      RECT 84.69 3.257 84.7 3.925 ;
      RECT 84.685 3.262 84.69 3.925 ;
      RECT 84.675 3.275 84.685 3.925 ;
      RECT 84.67 3.297 84.675 3.925 ;
      RECT 84.665 3.657 84.67 3.925 ;
      RECT 85.295 3.125 85.3 3.345 ;
      RECT 85.8 2.16 85.835 2.42 ;
      RECT 85.785 2.16 85.8 2.428 ;
      RECT 85.756 2.16 85.785 2.45 ;
      RECT 85.67 2.16 85.756 2.51 ;
      RECT 85.65 2.16 85.67 2.575 ;
      RECT 85.59 2.16 85.65 2.74 ;
      RECT 85.585 2.16 85.59 2.888 ;
      RECT 85.58 2.16 85.585 2.9 ;
      RECT 85.575 2.16 85.58 2.926 ;
      RECT 85.545 2.346 85.575 3.006 ;
      RECT 85.54 2.394 85.545 3.095 ;
      RECT 85.535 2.408 85.54 3.11 ;
      RECT 85.53 2.427 85.535 3.14 ;
      RECT 85.525 2.442 85.53 3.156 ;
      RECT 85.52 2.457 85.525 3.178 ;
      RECT 85.515 2.477 85.52 3.2 ;
      RECT 85.505 2.497 85.515 3.233 ;
      RECT 85.49 2.539 85.505 3.295 ;
      RECT 85.485 2.57 85.49 3.335 ;
      RECT 85.48 2.582 85.485 3.34 ;
      RECT 85.475 2.594 85.48 3.345 ;
      RECT 85.47 2.607 85.475 3.345 ;
      RECT 85.465 2.625 85.47 3.345 ;
      RECT 85.46 2.645 85.465 3.345 ;
      RECT 85.455 2.657 85.46 3.345 ;
      RECT 85.45 2.67 85.455 3.345 ;
      RECT 85.43 2.705 85.45 3.345 ;
      RECT 85.38 2.807 85.43 3.345 ;
      RECT 85.375 2.892 85.38 3.345 ;
      RECT 85.37 2.9 85.375 3.345 ;
      RECT 85.365 2.917 85.37 3.345 ;
      RECT 85.36 2.932 85.365 3.345 ;
      RECT 85.325 2.997 85.36 3.345 ;
      RECT 85.31 3.062 85.325 3.345 ;
      RECT 85.305 3.092 85.31 3.345 ;
      RECT 85.3 3.117 85.305 3.345 ;
      RECT 85.285 3.127 85.295 3.345 ;
      RECT 85.27 3.14 85.285 3.338 ;
      RECT 85.015 2.73 85.085 2.94 ;
      RECT 84.805 2.707 84.81 2.9 ;
      RECT 82.26 2.635 82.52 2.895 ;
      RECT 85.095 2.917 85.1 2.92 ;
      RECT 85.085 2.735 85.095 2.935 ;
      RECT 84.986 2.728 85.015 2.94 ;
      RECT 84.9 2.72 84.986 2.94 ;
      RECT 84.885 2.714 84.9 2.938 ;
      RECT 84.865 2.713 84.885 2.925 ;
      RECT 84.86 2.712 84.865 2.908 ;
      RECT 84.81 2.709 84.86 2.903 ;
      RECT 84.78 2.706 84.805 2.898 ;
      RECT 84.76 2.704 84.78 2.893 ;
      RECT 84.745 2.702 84.76 2.89 ;
      RECT 84.715 2.7 84.745 2.888 ;
      RECT 84.65 2.696 84.715 2.88 ;
      RECT 84.62 2.691 84.65 2.875 ;
      RECT 84.6 2.689 84.62 2.873 ;
      RECT 84.57 2.686 84.6 2.868 ;
      RECT 84.51 2.682 84.57 2.86 ;
      RECT 84.505 2.679 84.51 2.855 ;
      RECT 84.435 2.677 84.505 2.85 ;
      RECT 84.406 2.673 84.435 2.843 ;
      RECT 84.32 2.668 84.406 2.835 ;
      RECT 84.286 2.663 84.32 2.827 ;
      RECT 84.2 2.655 84.286 2.819 ;
      RECT 84.161 2.648 84.2 2.811 ;
      RECT 84.075 2.643 84.161 2.803 ;
      RECT 84.01 2.637 84.075 2.793 ;
      RECT 83.99 2.632 84.01 2.788 ;
      RECT 83.981 2.629 83.99 2.787 ;
      RECT 83.895 2.625 83.981 2.781 ;
      RECT 83.855 2.621 83.895 2.773 ;
      RECT 83.835 2.617 83.855 2.771 ;
      RECT 83.775 2.617 83.835 2.768 ;
      RECT 83.755 2.62 83.775 2.766 ;
      RECT 83.734 2.62 83.755 2.766 ;
      RECT 83.648 2.622 83.734 2.77 ;
      RECT 83.562 2.624 83.648 2.776 ;
      RECT 83.476 2.626 83.562 2.783 ;
      RECT 83.39 2.629 83.476 2.789 ;
      RECT 83.356 2.63 83.39 2.794 ;
      RECT 83.27 2.633 83.356 2.799 ;
      RECT 83.241 2.64 83.27 2.804 ;
      RECT 83.155 2.64 83.241 2.809 ;
      RECT 83.122 2.64 83.155 2.814 ;
      RECT 83.036 2.642 83.122 2.819 ;
      RECT 82.95 2.644 83.036 2.826 ;
      RECT 82.886 2.646 82.95 2.832 ;
      RECT 82.8 2.648 82.886 2.838 ;
      RECT 82.797 2.65 82.8 2.841 ;
      RECT 82.711 2.651 82.797 2.845 ;
      RECT 82.625 2.654 82.711 2.852 ;
      RECT 82.606 2.656 82.625 2.856 ;
      RECT 82.52 2.658 82.606 2.861 ;
      RECT 82.25 2.67 82.26 2.865 ;
      RECT 84.43 7.765 84.72 7.995 ;
      RECT 84.49 7.025 84.66 7.995 ;
      RECT 84.38 7.055 84.755 7.425 ;
      RECT 84.43 7.025 84.72 7.425 ;
      RECT 84.485 2.25 84.67 2.46 ;
      RECT 84.48 2.251 84.675 2.458 ;
      RECT 84.475 2.256 84.685 2.453 ;
      RECT 84.47 2.232 84.475 2.45 ;
      RECT 84.44 2.229 84.47 2.443 ;
      RECT 84.435 2.225 84.44 2.434 ;
      RECT 84.4 2.256 84.685 2.429 ;
      RECT 84.175 2.165 84.435 2.425 ;
      RECT 84.475 2.234 84.48 2.453 ;
      RECT 84.48 2.235 84.485 2.458 ;
      RECT 84.175 2.247 84.555 2.425 ;
      RECT 84.175 2.245 84.54 2.425 ;
      RECT 84.175 2.24 84.53 2.425 ;
      RECT 84.13 3.155 84.18 3.44 ;
      RECT 84.075 3.125 84.08 3.44 ;
      RECT 84.045 3.105 84.05 3.44 ;
      RECT 84.195 3.155 84.255 3.415 ;
      RECT 84.19 3.155 84.195 3.423 ;
      RECT 84.18 3.155 84.19 3.435 ;
      RECT 84.095 3.145 84.13 3.44 ;
      RECT 84.09 3.132 84.095 3.44 ;
      RECT 84.08 3.127 84.09 3.44 ;
      RECT 84.06 3.117 84.075 3.44 ;
      RECT 84.05 3.11 84.06 3.44 ;
      RECT 84.04 3.102 84.045 3.44 ;
      RECT 84.01 3.092 84.04 3.44 ;
      RECT 83.995 3.08 84.01 3.44 ;
      RECT 83.98 3.07 83.995 3.435 ;
      RECT 83.96 3.06 83.98 3.41 ;
      RECT 83.95 3.052 83.96 3.387 ;
      RECT 83.92 3.035 83.95 3.377 ;
      RECT 83.915 3.012 83.92 3.368 ;
      RECT 83.91 2.999 83.915 3.366 ;
      RECT 83.895 2.975 83.91 3.36 ;
      RECT 83.89 2.951 83.895 3.354 ;
      RECT 83.88 2.94 83.89 3.349 ;
      RECT 83.875 2.93 83.88 3.345 ;
      RECT 83.87 2.922 83.875 3.342 ;
      RECT 83.86 2.917 83.87 3.338 ;
      RECT 83.855 2.912 83.86 3.334 ;
      RECT 83.77 2.91 83.855 3.309 ;
      RECT 83.74 2.91 83.77 3.275 ;
      RECT 83.725 2.91 83.74 3.258 ;
      RECT 83.67 2.91 83.725 3.203 ;
      RECT 83.665 2.915 83.67 3.152 ;
      RECT 83.655 2.92 83.665 3.142 ;
      RECT 83.65 2.93 83.655 3.128 ;
      RECT 83.6 3.67 83.86 3.93 ;
      RECT 83.52 3.685 83.86 3.906 ;
      RECT 83.5 3.685 83.86 3.901 ;
      RECT 83.476 3.685 83.86 3.899 ;
      RECT 83.39 3.685 83.86 3.894 ;
      RECT 83.24 3.625 83.5 3.89 ;
      RECT 83.195 3.685 83.86 3.885 ;
      RECT 83.19 3.692 83.86 3.88 ;
      RECT 83.205 3.68 83.52 3.89 ;
      RECT 83.095 2.115 83.355 2.375 ;
      RECT 83.095 2.172 83.36 2.368 ;
      RECT 83.095 2.202 83.365 2.3 ;
      RECT 83.155 2.633 83.27 2.635 ;
      RECT 83.241 2.63 83.27 2.635 ;
      RECT 82.265 3.634 82.29 3.874 ;
      RECT 82.25 3.637 82.34 3.868 ;
      RECT 82.245 3.642 82.426 3.863 ;
      RECT 82.24 3.65 82.49 3.861 ;
      RECT 82.24 3.65 82.5 3.86 ;
      RECT 82.235 3.657 82.51 3.853 ;
      RECT 82.235 3.657 82.596 3.842 ;
      RECT 82.23 3.692 82.596 3.838 ;
      RECT 82.23 3.692 82.605 3.827 ;
      RECT 82.51 3.565 82.77 3.825 ;
      RECT 82.22 3.742 82.77 3.823 ;
      RECT 82.49 3.61 82.51 3.858 ;
      RECT 82.426 3.613 82.49 3.862 ;
      RECT 82.34 3.618 82.426 3.867 ;
      RECT 82.27 3.629 82.77 3.825 ;
      RECT 82.29 3.623 82.34 3.872 ;
      RECT 82.415 2.1 82.425 2.362 ;
      RECT 82.405 2.157 82.415 2.365 ;
      RECT 82.38 2.162 82.405 2.371 ;
      RECT 82.355 2.166 82.38 2.383 ;
      RECT 82.345 2.169 82.355 2.393 ;
      RECT 82.34 2.17 82.345 2.398 ;
      RECT 82.335 2.171 82.34 2.403 ;
      RECT 82.33 2.172 82.335 2.405 ;
      RECT 82.305 2.175 82.33 2.408 ;
      RECT 82.275 2.181 82.305 2.411 ;
      RECT 82.21 2.192 82.275 2.414 ;
      RECT 82.165 2.2 82.21 2.418 ;
      RECT 82.15 2.2 82.165 2.426 ;
      RECT 82.145 2.201 82.15 2.433 ;
      RECT 82.14 2.203 82.145 2.436 ;
      RECT 82.135 2.207 82.14 2.439 ;
      RECT 82.125 2.215 82.135 2.443 ;
      RECT 82.12 2.228 82.125 2.448 ;
      RECT 82.115 2.236 82.12 2.45 ;
      RECT 82.11 2.242 82.115 2.45 ;
      RECT 82.105 2.246 82.11 2.453 ;
      RECT 82.1 2.248 82.105 2.456 ;
      RECT 82.095 2.251 82.1 2.459 ;
      RECT 82.085 2.256 82.095 2.463 ;
      RECT 82.08 2.262 82.085 2.468 ;
      RECT 82.07 2.268 82.08 2.472 ;
      RECT 82.055 2.275 82.07 2.478 ;
      RECT 82.026 2.289 82.055 2.488 ;
      RECT 81.94 2.324 82.026 2.52 ;
      RECT 81.92 2.357 81.94 2.549 ;
      RECT 81.9 2.37 81.92 2.56 ;
      RECT 81.88 2.382 81.9 2.571 ;
      RECT 81.83 2.404 81.88 2.591 ;
      RECT 81.815 2.422 81.83 2.608 ;
      RECT 81.81 2.428 81.815 2.611 ;
      RECT 81.805 2.432 81.81 2.614 ;
      RECT 81.8 2.436 81.805 2.618 ;
      RECT 81.795 2.438 81.8 2.621 ;
      RECT 81.785 2.445 81.795 2.624 ;
      RECT 81.78 2.45 81.785 2.628 ;
      RECT 81.775 2.452 81.78 2.631 ;
      RECT 81.77 2.456 81.775 2.634 ;
      RECT 81.765 2.458 81.77 2.638 ;
      RECT 81.75 2.463 81.765 2.643 ;
      RECT 81.745 2.468 81.75 2.646 ;
      RECT 81.74 2.476 81.745 2.649 ;
      RECT 81.735 2.478 81.74 2.652 ;
      RECT 81.73 2.48 81.735 2.655 ;
      RECT 81.72 2.482 81.73 2.661 ;
      RECT 81.685 2.496 81.72 2.673 ;
      RECT 81.675 2.511 81.685 2.683 ;
      RECT 81.6 2.54 81.675 2.707 ;
      RECT 81.595 2.565 81.6 2.73 ;
      RECT 81.58 2.569 81.595 2.736 ;
      RECT 81.57 2.577 81.58 2.741 ;
      RECT 81.54 2.59 81.57 2.745 ;
      RECT 81.53 2.605 81.54 2.75 ;
      RECT 81.52 2.61 81.53 2.753 ;
      RECT 81.515 2.612 81.52 2.755 ;
      RECT 81.5 2.615 81.515 2.758 ;
      RECT 81.495 2.617 81.5 2.761 ;
      RECT 81.475 2.622 81.495 2.765 ;
      RECT 81.445 2.627 81.475 2.773 ;
      RECT 81.42 2.634 81.445 2.781 ;
      RECT 81.415 2.639 81.42 2.786 ;
      RECT 81.385 2.642 81.415 2.79 ;
      RECT 81.345 2.645 81.385 2.8 ;
      RECT 81.31 2.642 81.345 2.812 ;
      RECT 81.3 2.638 81.31 2.819 ;
      RECT 81.275 2.634 81.3 2.825 ;
      RECT 81.27 2.63 81.275 2.83 ;
      RECT 81.23 2.627 81.27 2.83 ;
      RECT 81.215 2.612 81.23 2.831 ;
      RECT 81.192 2.6 81.215 2.831 ;
      RECT 81.106 2.6 81.192 2.832 ;
      RECT 81.02 2.6 81.106 2.834 ;
      RECT 81 2.6 81.02 2.831 ;
      RECT 80.995 2.605 81 2.826 ;
      RECT 80.99 2.61 80.995 2.824 ;
      RECT 80.98 2.62 80.99 2.822 ;
      RECT 80.975 2.626 80.98 2.815 ;
      RECT 80.97 2.628 80.975 2.8 ;
      RECT 80.965 2.632 80.97 2.79 ;
      RECT 82.425 2.1 82.675 2.36 ;
      RECT 80.15 3.635 80.41 3.895 ;
      RECT 82.445 3.125 82.45 3.335 ;
      RECT 82.45 3.13 82.46 3.33 ;
      RECT 82.4 3.125 82.445 3.35 ;
      RECT 82.39 3.125 82.4 3.37 ;
      RECT 82.371 3.125 82.39 3.375 ;
      RECT 82.285 3.125 82.371 3.372 ;
      RECT 82.255 3.127 82.285 3.37 ;
      RECT 82.2 3.137 82.255 3.368 ;
      RECT 82.135 3.151 82.2 3.366 ;
      RECT 82.13 3.159 82.135 3.365 ;
      RECT 82.115 3.162 82.13 3.363 ;
      RECT 82.05 3.172 82.115 3.359 ;
      RECT 82.002 3.186 82.05 3.36 ;
      RECT 81.916 3.203 82.002 3.374 ;
      RECT 81.83 3.224 81.916 3.391 ;
      RECT 81.81 3.237 81.83 3.401 ;
      RECT 81.765 3.245 81.81 3.408 ;
      RECT 81.73 3.253 81.765 3.416 ;
      RECT 81.696 3.261 81.73 3.424 ;
      RECT 81.61 3.275 81.696 3.436 ;
      RECT 81.575 3.292 81.61 3.448 ;
      RECT 81.566 3.301 81.575 3.452 ;
      RECT 81.48 3.319 81.566 3.469 ;
      RECT 81.421 3.346 81.48 3.496 ;
      RECT 81.335 3.373 81.421 3.524 ;
      RECT 81.315 3.395 81.335 3.544 ;
      RECT 81.255 3.41 81.315 3.56 ;
      RECT 81.245 3.422 81.255 3.573 ;
      RECT 81.24 3.427 81.245 3.576 ;
      RECT 81.23 3.43 81.24 3.579 ;
      RECT 81.225 3.432 81.23 3.582 ;
      RECT 81.195 3.44 81.225 3.589 ;
      RECT 81.18 3.447 81.195 3.597 ;
      RECT 81.17 3.452 81.18 3.601 ;
      RECT 81.165 3.455 81.17 3.604 ;
      RECT 81.155 3.457 81.165 3.607 ;
      RECT 81.12 3.467 81.155 3.616 ;
      RECT 81.045 3.49 81.12 3.638 ;
      RECT 81.025 3.508 81.045 3.656 ;
      RECT 80.995 3.515 81.025 3.666 ;
      RECT 80.975 3.523 80.995 3.676 ;
      RECT 80.965 3.529 80.975 3.683 ;
      RECT 80.946 3.534 80.965 3.689 ;
      RECT 80.86 3.554 80.946 3.709 ;
      RECT 80.845 3.574 80.86 3.728 ;
      RECT 80.8 3.586 80.845 3.739 ;
      RECT 80.735 3.607 80.8 3.762 ;
      RECT 80.695 3.627 80.735 3.783 ;
      RECT 80.685 3.637 80.695 3.793 ;
      RECT 80.635 3.649 80.685 3.804 ;
      RECT 80.615 3.665 80.635 3.816 ;
      RECT 80.585 3.675 80.615 3.822 ;
      RECT 80.575 3.68 80.585 3.824 ;
      RECT 80.506 3.681 80.575 3.83 ;
      RECT 80.42 3.683 80.506 3.84 ;
      RECT 80.41 3.684 80.42 3.845 ;
      RECT 81.68 3.71 81.87 3.92 ;
      RECT 81.67 3.715 81.88 3.913 ;
      RECT 81.655 3.715 81.88 3.878 ;
      RECT 81.575 3.6 81.835 3.86 ;
      RECT 80.49 3.13 80.675 3.425 ;
      RECT 80.48 3.13 80.675 3.423 ;
      RECT 80.465 3.13 80.68 3.418 ;
      RECT 80.465 3.13 80.685 3.415 ;
      RECT 80.46 3.13 80.685 3.413 ;
      RECT 80.455 3.385 80.685 3.403 ;
      RECT 80.46 3.13 80.72 3.39 ;
      RECT 80.42 2.165 80.68 2.425 ;
      RECT 80.23 2.09 80.316 2.423 ;
      RECT 80.205 2.094 80.36 2.419 ;
      RECT 80.316 2.086 80.36 2.419 ;
      RECT 80.316 2.087 80.365 2.418 ;
      RECT 80.23 2.092 80.38 2.417 ;
      RECT 80.205 2.1 80.42 2.416 ;
      RECT 80.2 2.095 80.38 2.411 ;
      RECT 80.19 2.11 80.42 2.318 ;
      RECT 80.19 2.162 80.62 2.318 ;
      RECT 80.19 2.155 80.6 2.318 ;
      RECT 80.19 2.142 80.57 2.318 ;
      RECT 80.19 2.13 80.51 2.318 ;
      RECT 80.19 2.115 80.485 2.318 ;
      RECT 79.39 2.745 79.525 3.04 ;
      RECT 79.65 2.768 79.655 2.955 ;
      RECT 80.37 2.665 80.515 2.9 ;
      RECT 80.53 2.665 80.535 2.89 ;
      RECT 80.565 2.676 80.57 2.87 ;
      RECT 80.56 2.668 80.565 2.875 ;
      RECT 80.54 2.665 80.56 2.88 ;
      RECT 80.535 2.665 80.54 2.888 ;
      RECT 80.525 2.665 80.53 2.893 ;
      RECT 80.515 2.665 80.525 2.898 ;
      RECT 80.345 2.667 80.37 2.9 ;
      RECT 80.295 2.674 80.345 2.9 ;
      RECT 80.29 2.679 80.295 2.9 ;
      RECT 80.251 2.684 80.29 2.901 ;
      RECT 80.165 2.696 80.251 2.902 ;
      RECT 80.156 2.706 80.165 2.902 ;
      RECT 80.07 2.715 80.156 2.904 ;
      RECT 80.046 2.725 80.07 2.906 ;
      RECT 79.96 2.736 80.046 2.907 ;
      RECT 79.93 2.747 79.96 2.909 ;
      RECT 79.9 2.752 79.93 2.911 ;
      RECT 79.875 2.758 79.9 2.914 ;
      RECT 79.86 2.763 79.875 2.915 ;
      RECT 79.815 2.769 79.86 2.915 ;
      RECT 79.81 2.774 79.815 2.916 ;
      RECT 79.79 2.774 79.81 2.918 ;
      RECT 79.77 2.772 79.79 2.923 ;
      RECT 79.735 2.771 79.77 2.93 ;
      RECT 79.705 2.77 79.735 2.94 ;
      RECT 79.655 2.769 79.705 2.95 ;
      RECT 79.565 2.766 79.65 3.04 ;
      RECT 79.54 2.76 79.565 3.04 ;
      RECT 79.525 2.75 79.54 3.04 ;
      RECT 79.34 2.745 79.39 2.96 ;
      RECT 79.33 2.75 79.34 2.95 ;
      RECT 79.57 3.225 79.83 3.485 ;
      RECT 79.57 3.225 79.86 3.378 ;
      RECT 79.57 3.225 79.895 3.363 ;
      RECT 79.825 3.145 80.015 3.355 ;
      RECT 79.815 3.15 80.025 3.348 ;
      RECT 79.78 3.22 80.025 3.348 ;
      RECT 79.81 3.162 79.83 3.485 ;
      RECT 79.795 3.21 80.025 3.348 ;
      RECT 79.8 3.182 79.83 3.485 ;
      RECT 78.88 2.25 78.95 3.355 ;
      RECT 79.615 2.355 79.875 2.615 ;
      RECT 79.195 2.401 79.21 2.61 ;
      RECT 79.531 2.414 79.615 2.565 ;
      RECT 79.445 2.411 79.531 2.565 ;
      RECT 79.406 2.409 79.445 2.565 ;
      RECT 79.32 2.407 79.406 2.565 ;
      RECT 79.26 2.405 79.32 2.576 ;
      RECT 79.225 2.403 79.26 2.594 ;
      RECT 79.21 2.401 79.225 2.605 ;
      RECT 79.18 2.401 79.195 2.618 ;
      RECT 79.17 2.401 79.18 2.623 ;
      RECT 79.145 2.4 79.17 2.628 ;
      RECT 79.13 2.395 79.145 2.634 ;
      RECT 79.125 2.388 79.13 2.639 ;
      RECT 79.1 2.379 79.125 2.645 ;
      RECT 79.055 2.358 79.1 2.658 ;
      RECT 79.045 2.342 79.055 2.668 ;
      RECT 79.03 2.335 79.045 2.678 ;
      RECT 79.02 2.328 79.03 2.695 ;
      RECT 79.015 2.325 79.02 2.725 ;
      RECT 79.01 2.323 79.015 2.755 ;
      RECT 79.005 2.321 79.01 2.792 ;
      RECT 78.99 2.317 79.005 2.859 ;
      RECT 78.99 3.15 79 3.35 ;
      RECT 78.985 2.313 78.99 2.985 ;
      RECT 78.985 3.137 78.99 3.355 ;
      RECT 78.98 2.311 78.985 3.07 ;
      RECT 78.98 3.127 78.985 3.355 ;
      RECT 78.965 2.282 78.98 3.355 ;
      RECT 78.95 2.255 78.965 3.355 ;
      RECT 78.875 2.25 78.88 2.605 ;
      RECT 78.875 2.66 78.88 3.355 ;
      RECT 78.86 2.25 78.875 2.583 ;
      RECT 78.87 2.682 78.875 3.355 ;
      RECT 78.86 2.722 78.87 3.355 ;
      RECT 78.825 2.25 78.86 2.525 ;
      RECT 78.855 2.757 78.86 3.355 ;
      RECT 78.84 2.812 78.855 3.355 ;
      RECT 78.835 2.877 78.84 3.355 ;
      RECT 78.82 2.925 78.835 3.355 ;
      RECT 78.795 2.25 78.825 2.48 ;
      RECT 78.815 2.98 78.82 3.355 ;
      RECT 78.8 3.04 78.815 3.355 ;
      RECT 78.795 3.088 78.8 3.353 ;
      RECT 78.79 2.25 78.795 2.473 ;
      RECT 78.79 3.12 78.795 3.348 ;
      RECT 78.765 2.25 78.79 2.465 ;
      RECT 78.755 2.255 78.765 2.455 ;
      RECT 78.97 3.53 78.99 3.77 ;
      RECT 78.2 3.46 78.205 3.67 ;
      RECT 79.48 3.533 79.49 3.728 ;
      RECT 79.475 3.523 79.48 3.731 ;
      RECT 79.395 3.52 79.475 3.754 ;
      RECT 79.391 3.52 79.395 3.776 ;
      RECT 79.305 3.52 79.391 3.786 ;
      RECT 79.29 3.52 79.305 3.794 ;
      RECT 79.261 3.521 79.29 3.792 ;
      RECT 79.175 3.526 79.261 3.788 ;
      RECT 79.162 3.53 79.175 3.784 ;
      RECT 79.076 3.53 79.162 3.78 ;
      RECT 78.99 3.53 79.076 3.774 ;
      RECT 78.906 3.53 78.97 3.768 ;
      RECT 78.82 3.53 78.906 3.763 ;
      RECT 78.8 3.53 78.82 3.759 ;
      RECT 78.74 3.525 78.8 3.756 ;
      RECT 78.712 3.519 78.74 3.753 ;
      RECT 78.626 3.514 78.712 3.749 ;
      RECT 78.54 3.508 78.626 3.743 ;
      RECT 78.465 3.49 78.54 3.738 ;
      RECT 78.43 3.467 78.465 3.734 ;
      RECT 78.42 3.457 78.43 3.733 ;
      RECT 78.365 3.455 78.42 3.732 ;
      RECT 78.29 3.455 78.365 3.728 ;
      RECT 78.28 3.455 78.29 3.723 ;
      RECT 78.265 3.455 78.28 3.715 ;
      RECT 78.215 3.457 78.265 3.693 ;
      RECT 78.205 3.46 78.215 3.673 ;
      RECT 78.195 3.465 78.2 3.668 ;
      RECT 78.19 3.47 78.195 3.663 ;
      RECT 78.315 2.635 78.575 2.895 ;
      RECT 78.315 2.65 78.595 2.86 ;
      RECT 78.315 2.655 78.605 2.855 ;
      RECT 76.3 2.115 76.56 2.375 ;
      RECT 76.29 2.145 76.56 2.355 ;
      RECT 78.21 2.06 78.47 2.32 ;
      RECT 78.205 2.135 78.21 2.321 ;
      RECT 78.18 2.14 78.205 2.323 ;
      RECT 78.165 2.147 78.18 2.326 ;
      RECT 78.105 2.165 78.165 2.331 ;
      RECT 78.075 2.185 78.105 2.338 ;
      RECT 78.05 2.193 78.075 2.343 ;
      RECT 78.025 2.201 78.05 2.345 ;
      RECT 78.007 2.205 78.025 2.344 ;
      RECT 77.921 2.203 78.007 2.344 ;
      RECT 77.835 2.201 77.921 2.344 ;
      RECT 77.749 2.199 77.835 2.343 ;
      RECT 77.663 2.197 77.749 2.343 ;
      RECT 77.577 2.195 77.663 2.343 ;
      RECT 77.491 2.193 77.577 2.343 ;
      RECT 77.405 2.191 77.491 2.342 ;
      RECT 77.387 2.19 77.405 2.342 ;
      RECT 77.301 2.189 77.387 2.342 ;
      RECT 77.215 2.187 77.301 2.342 ;
      RECT 77.129 2.186 77.215 2.341 ;
      RECT 77.043 2.185 77.129 2.341 ;
      RECT 76.957 2.183 77.043 2.341 ;
      RECT 76.871 2.182 76.957 2.341 ;
      RECT 76.785 2.18 76.871 2.34 ;
      RECT 76.761 2.178 76.785 2.34 ;
      RECT 76.675 2.171 76.761 2.34 ;
      RECT 76.646 2.163 76.675 2.34 ;
      RECT 76.56 2.155 76.646 2.34 ;
      RECT 76.28 2.152 76.29 2.35 ;
      RECT 77.785 3.115 77.79 3.465 ;
      RECT 77.555 3.205 77.695 3.465 ;
      RECT 78.03 2.89 78.075 3.1 ;
      RECT 78.085 2.901 78.095 3.095 ;
      RECT 78.075 2.893 78.085 3.1 ;
      RECT 78.01 2.89 78.03 3.105 ;
      RECT 77.98 2.89 78.01 3.128 ;
      RECT 77.97 2.89 77.98 3.153 ;
      RECT 77.965 2.89 77.97 3.163 ;
      RECT 77.91 2.89 77.965 3.203 ;
      RECT 77.905 2.89 77.91 3.243 ;
      RECT 77.9 2.892 77.905 3.248 ;
      RECT 77.885 2.902 77.9 3.259 ;
      RECT 77.84 2.96 77.885 3.295 ;
      RECT 77.83 3.015 77.84 3.329 ;
      RECT 77.815 3.042 77.83 3.345 ;
      RECT 77.805 3.069 77.815 3.465 ;
      RECT 77.79 3.092 77.805 3.465 ;
      RECT 77.78 3.132 77.785 3.465 ;
      RECT 77.775 3.142 77.78 3.465 ;
      RECT 77.77 3.157 77.775 3.465 ;
      RECT 77.76 3.162 77.77 3.465 ;
      RECT 77.695 3.185 77.76 3.465 ;
      RECT 77.195 2.68 77.385 2.89 ;
      RECT 75.77 2.605 76.03 2.865 ;
      RECT 76.12 2.6 76.215 2.81 ;
      RECT 76.095 2.615 76.105 2.81 ;
      RECT 77.385 2.687 77.395 2.885 ;
      RECT 77.185 2.687 77.195 2.885 ;
      RECT 77.17 2.702 77.185 2.875 ;
      RECT 77.165 2.71 77.17 2.868 ;
      RECT 77.155 2.713 77.165 2.865 ;
      RECT 77.12 2.712 77.155 2.863 ;
      RECT 77.091 2.708 77.12 2.86 ;
      RECT 77.005 2.703 77.091 2.857 ;
      RECT 76.945 2.697 77.005 2.853 ;
      RECT 76.916 2.693 76.945 2.85 ;
      RECT 76.83 2.685 76.916 2.847 ;
      RECT 76.821 2.679 76.83 2.845 ;
      RECT 76.735 2.674 76.821 2.843 ;
      RECT 76.712 2.669 76.735 2.84 ;
      RECT 76.626 2.663 76.712 2.837 ;
      RECT 76.54 2.654 76.626 2.832 ;
      RECT 76.53 2.649 76.54 2.83 ;
      RECT 76.511 2.648 76.53 2.829 ;
      RECT 76.425 2.643 76.511 2.825 ;
      RECT 76.405 2.638 76.425 2.821 ;
      RECT 76.345 2.633 76.405 2.818 ;
      RECT 76.32 2.623 76.345 2.816 ;
      RECT 76.315 2.616 76.32 2.815 ;
      RECT 76.305 2.607 76.315 2.814 ;
      RECT 76.301 2.6 76.305 2.814 ;
      RECT 76.215 2.6 76.301 2.812 ;
      RECT 76.105 2.607 76.12 2.81 ;
      RECT 76.09 2.617 76.095 2.81 ;
      RECT 76.07 2.62 76.09 2.807 ;
      RECT 76.04 2.62 76.07 2.803 ;
      RECT 76.03 2.62 76.04 2.803 ;
      RECT 76.945 3.115 77.205 3.375 ;
      RECT 76.875 3.125 77.205 3.335 ;
      RECT 76.865 3.132 77.205 3.33 ;
      RECT 76.285 3.12 76.545 3.38 ;
      RECT 76.285 3.16 76.65 3.37 ;
      RECT 76.285 3.162 76.655 3.369 ;
      RECT 76.285 3.17 76.66 3.366 ;
      RECT 75.21 2.245 75.31 3.77 ;
      RECT 75.4 3.385 75.45 3.645 ;
      RECT 75.395 2.258 75.4 2.445 ;
      RECT 75.39 3.366 75.4 3.645 ;
      RECT 75.39 2.255 75.395 2.453 ;
      RECT 75.375 2.249 75.39 2.46 ;
      RECT 75.385 3.354 75.39 3.728 ;
      RECT 75.375 3.342 75.385 3.765 ;
      RECT 75.365 2.245 75.375 2.467 ;
      RECT 75.365 3.327 75.375 3.77 ;
      RECT 75.36 2.245 75.365 2.475 ;
      RECT 75.34 3.297 75.365 3.77 ;
      RECT 75.32 2.245 75.36 2.523 ;
      RECT 75.33 3.257 75.34 3.77 ;
      RECT 75.32 3.212 75.33 3.77 ;
      RECT 75.315 2.245 75.32 2.593 ;
      RECT 75.315 3.17 75.32 3.77 ;
      RECT 75.31 2.245 75.315 3.07 ;
      RECT 75.31 3.152 75.315 3.77 ;
      RECT 75.2 2.248 75.21 3.77 ;
      RECT 75.185 2.255 75.2 3.766 ;
      RECT 75.18 2.265 75.185 3.761 ;
      RECT 75.175 2.465 75.18 3.653 ;
      RECT 75.17 2.55 75.175 3.205 ;
      RECT 74.05 7.765 74.34 7.995 ;
      RECT 74.11 6.285 74.28 7.995 ;
      RECT 74.055 6.655 74.405 7.005 ;
      RECT 74.05 6.285 74.34 6.515 ;
      RECT 74.05 2.365 74.34 2.595 ;
      RECT 74.11 0.885 74.28 2.595 ;
      RECT 74.05 0.885 74.34 1.115 ;
      RECT 73.64 2.735 73.97 2.965 ;
      RECT 73.64 2.765 74.14 2.935 ;
      RECT 73.64 2.395 73.83 2.965 ;
      RECT 73.06 2.365 73.35 2.595 ;
      RECT 73.06 2.395 73.83 2.565 ;
      RECT 73.12 0.885 73.29 2.595 ;
      RECT 73.06 0.885 73.35 1.115 ;
      RECT 73.06 7.765 73.35 7.995 ;
      RECT 73.12 6.285 73.29 7.995 ;
      RECT 73.06 6.285 73.35 6.515 ;
      RECT 73.06 6.325 73.91 6.485 ;
      RECT 73.74 5.915 73.91 6.485 ;
      RECT 73.06 6.32 73.45 6.485 ;
      RECT 73.68 5.915 73.97 6.145 ;
      RECT 73.68 5.945 74.14 6.115 ;
      RECT 72.69 2.735 72.98 2.965 ;
      RECT 72.69 2.765 73.15 2.935 ;
      RECT 72.75 1.655 72.915 2.965 ;
      RECT 71.265 1.625 71.555 1.855 ;
      RECT 71.265 1.655 72.915 1.825 ;
      RECT 71.325 0.885 71.495 1.855 ;
      RECT 71.265 0.885 71.555 1.115 ;
      RECT 71.265 7.765 71.555 7.995 ;
      RECT 71.325 7.025 71.495 7.995 ;
      RECT 71.325 7.12 72.915 7.29 ;
      RECT 72.745 5.915 72.915 7.29 ;
      RECT 71.265 7.025 71.555 7.255 ;
      RECT 72.69 5.915 72.98 6.145 ;
      RECT 72.69 5.945 73.15 6.115 ;
      RECT 69.3 3.43 69.65 3.78 ;
      RECT 69.39 2.025 69.56 3.78 ;
      RECT 71.695 1.965 72.045 2.315 ;
      RECT 69.39 2.025 71.01 2.2 ;
      RECT 69.39 2.025 72.045 2.195 ;
      RECT 71.72 6.655 72.045 6.98 ;
      RECT 67.095 6.61 67.445 6.96 ;
      RECT 71.695 6.655 72.045 6.885 ;
      RECT 66.935 6.655 67.445 6.885 ;
      RECT 66.765 6.685 72.045 6.855 ;
      RECT 70.92 2.365 71.24 2.685 ;
      RECT 70.89 2.365 71.24 2.595 ;
      RECT 70.72 2.395 71.24 2.565 ;
      RECT 70.92 6.225 71.24 6.545 ;
      RECT 70.89 6.285 71.24 6.515 ;
      RECT 70.72 6.315 71.24 6.485 ;
      RECT 69.875 2.705 70.225 3.055 ;
      RECT 69.875 2.765 70.355 2.935 ;
      RECT 69.865 5.84 70.215 6.19 ;
      RECT 65.135 5.915 65.425 6.145 ;
      RECT 65.135 5.945 70.355 6.115 ;
      RECT 66.7 3.665 66.74 3.925 ;
      RECT 66.74 3.645 66.745 3.655 ;
      RECT 68.07 2.89 68.08 3.111 ;
      RECT 68 2.885 68.07 3.236 ;
      RECT 67.99 2.885 68 3.363 ;
      RECT 67.965 2.885 67.99 3.41 ;
      RECT 67.94 2.885 67.965 3.488 ;
      RECT 67.92 2.885 67.94 3.558 ;
      RECT 67.895 2.885 67.92 3.598 ;
      RECT 67.885 2.885 67.895 3.618 ;
      RECT 67.875 2.887 67.885 3.626 ;
      RECT 67.87 2.892 67.875 3.083 ;
      RECT 67.87 3.092 67.875 3.627 ;
      RECT 67.865 3.137 67.87 3.628 ;
      RECT 67.855 3.202 67.865 3.629 ;
      RECT 67.845 3.297 67.855 3.631 ;
      RECT 67.84 3.35 67.845 3.633 ;
      RECT 67.835 3.37 67.84 3.634 ;
      RECT 67.78 3.395 67.835 3.64 ;
      RECT 67.74 3.43 67.78 3.649 ;
      RECT 67.73 3.447 67.74 3.654 ;
      RECT 67.721 3.453 67.73 3.656 ;
      RECT 67.635 3.491 67.721 3.667 ;
      RECT 67.63 3.53 67.635 3.677 ;
      RECT 67.555 3.537 67.63 3.687 ;
      RECT 67.535 3.547 67.555 3.698 ;
      RECT 67.505 3.554 67.535 3.706 ;
      RECT 67.48 3.561 67.505 3.713 ;
      RECT 67.456 3.567 67.48 3.718 ;
      RECT 67.37 3.58 67.456 3.73 ;
      RECT 67.292 3.587 67.37 3.748 ;
      RECT 67.206 3.582 67.292 3.766 ;
      RECT 67.12 3.577 67.206 3.786 ;
      RECT 67.04 3.571 67.12 3.803 ;
      RECT 66.975 3.567 67.04 3.832 ;
      RECT 66.97 3.281 66.975 3.305 ;
      RECT 66.96 3.557 66.975 3.86 ;
      RECT 66.965 3.275 66.97 3.345 ;
      RECT 66.96 3.269 66.965 3.415 ;
      RECT 66.955 3.263 66.96 3.493 ;
      RECT 66.955 3.54 66.96 3.925 ;
      RECT 66.947 3.26 66.955 3.925 ;
      RECT 66.861 3.258 66.947 3.925 ;
      RECT 66.775 3.256 66.861 3.925 ;
      RECT 66.765 3.257 66.775 3.925 ;
      RECT 66.76 3.262 66.765 3.925 ;
      RECT 66.75 3.275 66.76 3.925 ;
      RECT 66.745 3.297 66.75 3.925 ;
      RECT 66.74 3.657 66.745 3.925 ;
      RECT 67.37 3.125 67.375 3.345 ;
      RECT 67.875 2.16 67.91 2.42 ;
      RECT 67.86 2.16 67.875 2.428 ;
      RECT 67.831 2.16 67.86 2.45 ;
      RECT 67.745 2.16 67.831 2.51 ;
      RECT 67.725 2.16 67.745 2.575 ;
      RECT 67.665 2.16 67.725 2.74 ;
      RECT 67.66 2.16 67.665 2.888 ;
      RECT 67.655 2.16 67.66 2.9 ;
      RECT 67.65 2.16 67.655 2.926 ;
      RECT 67.62 2.346 67.65 3.006 ;
      RECT 67.615 2.394 67.62 3.095 ;
      RECT 67.61 2.408 67.615 3.11 ;
      RECT 67.605 2.427 67.61 3.14 ;
      RECT 67.6 2.442 67.605 3.156 ;
      RECT 67.595 2.457 67.6 3.178 ;
      RECT 67.59 2.477 67.595 3.2 ;
      RECT 67.58 2.497 67.59 3.233 ;
      RECT 67.565 2.539 67.58 3.295 ;
      RECT 67.56 2.57 67.565 3.335 ;
      RECT 67.555 2.582 67.56 3.34 ;
      RECT 67.55 2.594 67.555 3.345 ;
      RECT 67.545 2.607 67.55 3.345 ;
      RECT 67.54 2.625 67.545 3.345 ;
      RECT 67.535 2.645 67.54 3.345 ;
      RECT 67.53 2.657 67.535 3.345 ;
      RECT 67.525 2.67 67.53 3.345 ;
      RECT 67.505 2.705 67.525 3.345 ;
      RECT 67.455 2.807 67.505 3.345 ;
      RECT 67.45 2.892 67.455 3.345 ;
      RECT 67.445 2.9 67.45 3.345 ;
      RECT 67.44 2.917 67.445 3.345 ;
      RECT 67.435 2.932 67.44 3.345 ;
      RECT 67.4 2.997 67.435 3.345 ;
      RECT 67.385 3.062 67.4 3.345 ;
      RECT 67.38 3.092 67.385 3.345 ;
      RECT 67.375 3.117 67.38 3.345 ;
      RECT 67.36 3.127 67.37 3.345 ;
      RECT 67.345 3.14 67.36 3.338 ;
      RECT 67.09 2.73 67.16 2.94 ;
      RECT 66.88 2.707 66.885 2.9 ;
      RECT 64.335 2.635 64.595 2.895 ;
      RECT 67.17 2.917 67.175 2.92 ;
      RECT 67.16 2.735 67.17 2.935 ;
      RECT 67.061 2.728 67.09 2.94 ;
      RECT 66.975 2.72 67.061 2.94 ;
      RECT 66.96 2.714 66.975 2.938 ;
      RECT 66.94 2.713 66.96 2.925 ;
      RECT 66.935 2.712 66.94 2.908 ;
      RECT 66.885 2.709 66.935 2.903 ;
      RECT 66.855 2.706 66.88 2.898 ;
      RECT 66.835 2.704 66.855 2.893 ;
      RECT 66.82 2.702 66.835 2.89 ;
      RECT 66.79 2.7 66.82 2.888 ;
      RECT 66.725 2.696 66.79 2.88 ;
      RECT 66.695 2.691 66.725 2.875 ;
      RECT 66.675 2.689 66.695 2.873 ;
      RECT 66.645 2.686 66.675 2.868 ;
      RECT 66.585 2.682 66.645 2.86 ;
      RECT 66.58 2.679 66.585 2.855 ;
      RECT 66.51 2.677 66.58 2.85 ;
      RECT 66.481 2.673 66.51 2.843 ;
      RECT 66.395 2.668 66.481 2.835 ;
      RECT 66.361 2.663 66.395 2.827 ;
      RECT 66.275 2.655 66.361 2.819 ;
      RECT 66.236 2.648 66.275 2.811 ;
      RECT 66.15 2.643 66.236 2.803 ;
      RECT 66.085 2.637 66.15 2.793 ;
      RECT 66.065 2.632 66.085 2.788 ;
      RECT 66.056 2.629 66.065 2.787 ;
      RECT 65.97 2.625 66.056 2.781 ;
      RECT 65.93 2.621 65.97 2.773 ;
      RECT 65.91 2.617 65.93 2.771 ;
      RECT 65.85 2.617 65.91 2.768 ;
      RECT 65.83 2.62 65.85 2.766 ;
      RECT 65.809 2.62 65.83 2.766 ;
      RECT 65.723 2.622 65.809 2.77 ;
      RECT 65.637 2.624 65.723 2.776 ;
      RECT 65.551 2.626 65.637 2.783 ;
      RECT 65.465 2.629 65.551 2.789 ;
      RECT 65.431 2.63 65.465 2.794 ;
      RECT 65.345 2.633 65.431 2.799 ;
      RECT 65.316 2.64 65.345 2.804 ;
      RECT 65.23 2.64 65.316 2.809 ;
      RECT 65.197 2.64 65.23 2.814 ;
      RECT 65.111 2.642 65.197 2.819 ;
      RECT 65.025 2.644 65.111 2.826 ;
      RECT 64.961 2.646 65.025 2.832 ;
      RECT 64.875 2.648 64.961 2.838 ;
      RECT 64.872 2.65 64.875 2.841 ;
      RECT 64.786 2.651 64.872 2.845 ;
      RECT 64.7 2.654 64.786 2.852 ;
      RECT 64.681 2.656 64.7 2.856 ;
      RECT 64.595 2.658 64.681 2.861 ;
      RECT 64.325 2.67 64.335 2.865 ;
      RECT 66.505 7.765 66.795 7.995 ;
      RECT 66.565 7.025 66.735 7.995 ;
      RECT 66.455 7.055 66.83 7.425 ;
      RECT 66.505 7.025 66.795 7.425 ;
      RECT 66.56 2.25 66.745 2.46 ;
      RECT 66.555 2.251 66.75 2.458 ;
      RECT 66.55 2.256 66.76 2.453 ;
      RECT 66.545 2.232 66.55 2.45 ;
      RECT 66.515 2.229 66.545 2.443 ;
      RECT 66.51 2.225 66.515 2.434 ;
      RECT 66.475 2.256 66.76 2.429 ;
      RECT 66.25 2.165 66.51 2.425 ;
      RECT 66.55 2.234 66.555 2.453 ;
      RECT 66.555 2.235 66.56 2.458 ;
      RECT 66.25 2.247 66.63 2.425 ;
      RECT 66.25 2.245 66.615 2.425 ;
      RECT 66.25 2.24 66.605 2.425 ;
      RECT 66.205 3.155 66.255 3.44 ;
      RECT 66.15 3.125 66.155 3.44 ;
      RECT 66.12 3.105 66.125 3.44 ;
      RECT 66.27 3.155 66.33 3.415 ;
      RECT 66.265 3.155 66.27 3.423 ;
      RECT 66.255 3.155 66.265 3.435 ;
      RECT 66.17 3.145 66.205 3.44 ;
      RECT 66.165 3.132 66.17 3.44 ;
      RECT 66.155 3.127 66.165 3.44 ;
      RECT 66.135 3.117 66.15 3.44 ;
      RECT 66.125 3.11 66.135 3.44 ;
      RECT 66.115 3.102 66.12 3.44 ;
      RECT 66.085 3.092 66.115 3.44 ;
      RECT 66.07 3.08 66.085 3.44 ;
      RECT 66.055 3.07 66.07 3.435 ;
      RECT 66.035 3.06 66.055 3.41 ;
      RECT 66.025 3.052 66.035 3.387 ;
      RECT 65.995 3.035 66.025 3.377 ;
      RECT 65.99 3.012 65.995 3.368 ;
      RECT 65.985 2.999 65.99 3.366 ;
      RECT 65.97 2.975 65.985 3.36 ;
      RECT 65.965 2.951 65.97 3.354 ;
      RECT 65.955 2.94 65.965 3.349 ;
      RECT 65.95 2.93 65.955 3.345 ;
      RECT 65.945 2.922 65.95 3.342 ;
      RECT 65.935 2.917 65.945 3.338 ;
      RECT 65.93 2.912 65.935 3.334 ;
      RECT 65.845 2.91 65.93 3.309 ;
      RECT 65.815 2.91 65.845 3.275 ;
      RECT 65.8 2.91 65.815 3.258 ;
      RECT 65.745 2.91 65.8 3.203 ;
      RECT 65.74 2.915 65.745 3.152 ;
      RECT 65.73 2.92 65.74 3.142 ;
      RECT 65.725 2.93 65.73 3.128 ;
      RECT 65.675 3.67 65.935 3.93 ;
      RECT 65.595 3.685 65.935 3.906 ;
      RECT 65.575 3.685 65.935 3.901 ;
      RECT 65.551 3.685 65.935 3.899 ;
      RECT 65.465 3.685 65.935 3.894 ;
      RECT 65.315 3.625 65.575 3.89 ;
      RECT 65.27 3.685 65.935 3.885 ;
      RECT 65.265 3.692 65.935 3.88 ;
      RECT 65.28 3.68 65.595 3.89 ;
      RECT 65.17 2.115 65.43 2.375 ;
      RECT 65.17 2.172 65.435 2.368 ;
      RECT 65.17 2.202 65.44 2.3 ;
      RECT 65.23 2.633 65.345 2.635 ;
      RECT 65.316 2.63 65.345 2.635 ;
      RECT 64.34 3.634 64.365 3.874 ;
      RECT 64.325 3.637 64.415 3.868 ;
      RECT 64.32 3.642 64.501 3.863 ;
      RECT 64.315 3.65 64.565 3.861 ;
      RECT 64.315 3.65 64.575 3.86 ;
      RECT 64.31 3.657 64.585 3.853 ;
      RECT 64.31 3.657 64.671 3.842 ;
      RECT 64.305 3.692 64.671 3.838 ;
      RECT 64.305 3.692 64.68 3.827 ;
      RECT 64.585 3.565 64.845 3.825 ;
      RECT 64.295 3.742 64.845 3.823 ;
      RECT 64.565 3.61 64.585 3.858 ;
      RECT 64.501 3.613 64.565 3.862 ;
      RECT 64.415 3.618 64.501 3.867 ;
      RECT 64.345 3.629 64.845 3.825 ;
      RECT 64.365 3.623 64.415 3.872 ;
      RECT 64.49 2.1 64.5 2.362 ;
      RECT 64.48 2.157 64.49 2.365 ;
      RECT 64.455 2.162 64.48 2.371 ;
      RECT 64.43 2.166 64.455 2.383 ;
      RECT 64.42 2.169 64.43 2.393 ;
      RECT 64.415 2.17 64.42 2.398 ;
      RECT 64.41 2.171 64.415 2.403 ;
      RECT 64.405 2.172 64.41 2.405 ;
      RECT 64.38 2.175 64.405 2.408 ;
      RECT 64.35 2.181 64.38 2.411 ;
      RECT 64.285 2.192 64.35 2.414 ;
      RECT 64.24 2.2 64.285 2.418 ;
      RECT 64.225 2.2 64.24 2.426 ;
      RECT 64.22 2.201 64.225 2.433 ;
      RECT 64.215 2.203 64.22 2.436 ;
      RECT 64.21 2.207 64.215 2.439 ;
      RECT 64.2 2.215 64.21 2.443 ;
      RECT 64.195 2.228 64.2 2.448 ;
      RECT 64.19 2.236 64.195 2.45 ;
      RECT 64.185 2.242 64.19 2.45 ;
      RECT 64.18 2.246 64.185 2.453 ;
      RECT 64.175 2.248 64.18 2.456 ;
      RECT 64.17 2.251 64.175 2.459 ;
      RECT 64.16 2.256 64.17 2.463 ;
      RECT 64.155 2.262 64.16 2.468 ;
      RECT 64.145 2.268 64.155 2.472 ;
      RECT 64.13 2.275 64.145 2.478 ;
      RECT 64.101 2.289 64.13 2.488 ;
      RECT 64.015 2.324 64.101 2.52 ;
      RECT 63.995 2.357 64.015 2.549 ;
      RECT 63.975 2.37 63.995 2.56 ;
      RECT 63.955 2.382 63.975 2.571 ;
      RECT 63.905 2.404 63.955 2.591 ;
      RECT 63.89 2.422 63.905 2.608 ;
      RECT 63.885 2.428 63.89 2.611 ;
      RECT 63.88 2.432 63.885 2.614 ;
      RECT 63.875 2.436 63.88 2.618 ;
      RECT 63.87 2.438 63.875 2.621 ;
      RECT 63.86 2.445 63.87 2.624 ;
      RECT 63.855 2.45 63.86 2.628 ;
      RECT 63.85 2.452 63.855 2.631 ;
      RECT 63.845 2.456 63.85 2.634 ;
      RECT 63.84 2.458 63.845 2.638 ;
      RECT 63.825 2.463 63.84 2.643 ;
      RECT 63.82 2.468 63.825 2.646 ;
      RECT 63.815 2.476 63.82 2.649 ;
      RECT 63.81 2.478 63.815 2.652 ;
      RECT 63.805 2.48 63.81 2.655 ;
      RECT 63.795 2.482 63.805 2.661 ;
      RECT 63.76 2.496 63.795 2.673 ;
      RECT 63.75 2.511 63.76 2.683 ;
      RECT 63.675 2.54 63.75 2.707 ;
      RECT 63.67 2.565 63.675 2.73 ;
      RECT 63.655 2.569 63.67 2.736 ;
      RECT 63.645 2.577 63.655 2.741 ;
      RECT 63.615 2.59 63.645 2.745 ;
      RECT 63.605 2.605 63.615 2.75 ;
      RECT 63.595 2.61 63.605 2.753 ;
      RECT 63.59 2.612 63.595 2.755 ;
      RECT 63.575 2.615 63.59 2.758 ;
      RECT 63.57 2.617 63.575 2.761 ;
      RECT 63.55 2.622 63.57 2.765 ;
      RECT 63.52 2.627 63.55 2.773 ;
      RECT 63.495 2.634 63.52 2.781 ;
      RECT 63.49 2.639 63.495 2.786 ;
      RECT 63.46 2.642 63.49 2.79 ;
      RECT 63.42 2.645 63.46 2.8 ;
      RECT 63.385 2.642 63.42 2.812 ;
      RECT 63.375 2.638 63.385 2.819 ;
      RECT 63.35 2.634 63.375 2.825 ;
      RECT 63.345 2.63 63.35 2.83 ;
      RECT 63.305 2.627 63.345 2.83 ;
      RECT 63.29 2.612 63.305 2.831 ;
      RECT 63.267 2.6 63.29 2.831 ;
      RECT 63.181 2.6 63.267 2.832 ;
      RECT 63.095 2.6 63.181 2.834 ;
      RECT 63.075 2.6 63.095 2.831 ;
      RECT 63.07 2.605 63.075 2.826 ;
      RECT 63.065 2.61 63.07 2.824 ;
      RECT 63.055 2.62 63.065 2.822 ;
      RECT 63.05 2.626 63.055 2.815 ;
      RECT 63.045 2.628 63.05 2.8 ;
      RECT 63.04 2.632 63.045 2.79 ;
      RECT 64.5 2.1 64.75 2.36 ;
      RECT 62.225 3.635 62.485 3.895 ;
      RECT 64.52 3.125 64.525 3.335 ;
      RECT 64.525 3.13 64.535 3.33 ;
      RECT 64.475 3.125 64.52 3.35 ;
      RECT 64.465 3.125 64.475 3.37 ;
      RECT 64.446 3.125 64.465 3.375 ;
      RECT 64.36 3.125 64.446 3.372 ;
      RECT 64.33 3.127 64.36 3.37 ;
      RECT 64.275 3.137 64.33 3.368 ;
      RECT 64.21 3.151 64.275 3.366 ;
      RECT 64.205 3.159 64.21 3.365 ;
      RECT 64.19 3.162 64.205 3.363 ;
      RECT 64.125 3.172 64.19 3.359 ;
      RECT 64.077 3.186 64.125 3.36 ;
      RECT 63.991 3.203 64.077 3.374 ;
      RECT 63.905 3.224 63.991 3.391 ;
      RECT 63.885 3.237 63.905 3.401 ;
      RECT 63.84 3.245 63.885 3.408 ;
      RECT 63.805 3.253 63.84 3.416 ;
      RECT 63.771 3.261 63.805 3.424 ;
      RECT 63.685 3.275 63.771 3.436 ;
      RECT 63.65 3.292 63.685 3.448 ;
      RECT 63.641 3.301 63.65 3.452 ;
      RECT 63.555 3.319 63.641 3.469 ;
      RECT 63.496 3.346 63.555 3.496 ;
      RECT 63.41 3.373 63.496 3.524 ;
      RECT 63.39 3.395 63.41 3.544 ;
      RECT 63.33 3.41 63.39 3.56 ;
      RECT 63.32 3.422 63.33 3.573 ;
      RECT 63.315 3.427 63.32 3.576 ;
      RECT 63.305 3.43 63.315 3.579 ;
      RECT 63.3 3.432 63.305 3.582 ;
      RECT 63.27 3.44 63.3 3.589 ;
      RECT 63.255 3.447 63.27 3.597 ;
      RECT 63.245 3.452 63.255 3.601 ;
      RECT 63.24 3.455 63.245 3.604 ;
      RECT 63.23 3.457 63.24 3.607 ;
      RECT 63.195 3.467 63.23 3.616 ;
      RECT 63.12 3.49 63.195 3.638 ;
      RECT 63.1 3.508 63.12 3.656 ;
      RECT 63.07 3.515 63.1 3.666 ;
      RECT 63.05 3.523 63.07 3.676 ;
      RECT 63.04 3.529 63.05 3.683 ;
      RECT 63.021 3.534 63.04 3.689 ;
      RECT 62.935 3.554 63.021 3.709 ;
      RECT 62.92 3.574 62.935 3.728 ;
      RECT 62.875 3.586 62.92 3.739 ;
      RECT 62.81 3.607 62.875 3.762 ;
      RECT 62.77 3.627 62.81 3.783 ;
      RECT 62.76 3.637 62.77 3.793 ;
      RECT 62.71 3.649 62.76 3.804 ;
      RECT 62.69 3.665 62.71 3.816 ;
      RECT 62.66 3.675 62.69 3.822 ;
      RECT 62.65 3.68 62.66 3.824 ;
      RECT 62.581 3.681 62.65 3.83 ;
      RECT 62.495 3.683 62.581 3.84 ;
      RECT 62.485 3.684 62.495 3.845 ;
      RECT 63.755 3.71 63.945 3.92 ;
      RECT 63.745 3.715 63.955 3.913 ;
      RECT 63.73 3.715 63.955 3.878 ;
      RECT 63.65 3.6 63.91 3.86 ;
      RECT 62.565 3.13 62.75 3.425 ;
      RECT 62.555 3.13 62.75 3.423 ;
      RECT 62.54 3.13 62.755 3.418 ;
      RECT 62.54 3.13 62.76 3.415 ;
      RECT 62.535 3.13 62.76 3.413 ;
      RECT 62.53 3.385 62.76 3.403 ;
      RECT 62.535 3.13 62.795 3.39 ;
      RECT 62.495 2.165 62.755 2.425 ;
      RECT 62.305 2.09 62.391 2.423 ;
      RECT 62.28 2.094 62.435 2.419 ;
      RECT 62.391 2.086 62.435 2.419 ;
      RECT 62.391 2.087 62.44 2.418 ;
      RECT 62.305 2.092 62.455 2.417 ;
      RECT 62.28 2.1 62.495 2.416 ;
      RECT 62.275 2.095 62.455 2.411 ;
      RECT 62.265 2.11 62.495 2.318 ;
      RECT 62.265 2.162 62.695 2.318 ;
      RECT 62.265 2.155 62.675 2.318 ;
      RECT 62.265 2.142 62.645 2.318 ;
      RECT 62.265 2.13 62.585 2.318 ;
      RECT 62.265 2.115 62.56 2.318 ;
      RECT 61.465 2.745 61.6 3.04 ;
      RECT 61.725 2.768 61.73 2.955 ;
      RECT 62.445 2.665 62.59 2.9 ;
      RECT 62.605 2.665 62.61 2.89 ;
      RECT 62.64 2.676 62.645 2.87 ;
      RECT 62.635 2.668 62.64 2.875 ;
      RECT 62.615 2.665 62.635 2.88 ;
      RECT 62.61 2.665 62.615 2.888 ;
      RECT 62.6 2.665 62.605 2.893 ;
      RECT 62.59 2.665 62.6 2.898 ;
      RECT 62.42 2.667 62.445 2.9 ;
      RECT 62.37 2.674 62.42 2.9 ;
      RECT 62.365 2.679 62.37 2.9 ;
      RECT 62.326 2.684 62.365 2.901 ;
      RECT 62.24 2.696 62.326 2.902 ;
      RECT 62.231 2.706 62.24 2.902 ;
      RECT 62.145 2.715 62.231 2.904 ;
      RECT 62.121 2.725 62.145 2.906 ;
      RECT 62.035 2.736 62.121 2.907 ;
      RECT 62.005 2.747 62.035 2.909 ;
      RECT 61.975 2.752 62.005 2.911 ;
      RECT 61.95 2.758 61.975 2.914 ;
      RECT 61.935 2.763 61.95 2.915 ;
      RECT 61.89 2.769 61.935 2.915 ;
      RECT 61.885 2.774 61.89 2.916 ;
      RECT 61.865 2.774 61.885 2.918 ;
      RECT 61.845 2.772 61.865 2.923 ;
      RECT 61.81 2.771 61.845 2.93 ;
      RECT 61.78 2.77 61.81 2.94 ;
      RECT 61.73 2.769 61.78 2.95 ;
      RECT 61.64 2.766 61.725 3.04 ;
      RECT 61.615 2.76 61.64 3.04 ;
      RECT 61.6 2.75 61.615 3.04 ;
      RECT 61.415 2.745 61.465 2.96 ;
      RECT 61.405 2.75 61.415 2.95 ;
      RECT 61.645 3.225 61.905 3.485 ;
      RECT 61.645 3.225 61.935 3.378 ;
      RECT 61.645 3.225 61.97 3.363 ;
      RECT 61.9 3.145 62.09 3.355 ;
      RECT 61.89 3.15 62.1 3.348 ;
      RECT 61.855 3.22 62.1 3.348 ;
      RECT 61.885 3.162 61.905 3.485 ;
      RECT 61.87 3.21 62.1 3.348 ;
      RECT 61.875 3.182 61.905 3.485 ;
      RECT 60.955 2.25 61.025 3.355 ;
      RECT 61.69 2.355 61.95 2.615 ;
      RECT 61.27 2.401 61.285 2.61 ;
      RECT 61.606 2.414 61.69 2.565 ;
      RECT 61.52 2.411 61.606 2.565 ;
      RECT 61.481 2.409 61.52 2.565 ;
      RECT 61.395 2.407 61.481 2.565 ;
      RECT 61.335 2.405 61.395 2.576 ;
      RECT 61.3 2.403 61.335 2.594 ;
      RECT 61.285 2.401 61.3 2.605 ;
      RECT 61.255 2.401 61.27 2.618 ;
      RECT 61.245 2.401 61.255 2.623 ;
      RECT 61.22 2.4 61.245 2.628 ;
      RECT 61.205 2.395 61.22 2.634 ;
      RECT 61.2 2.388 61.205 2.639 ;
      RECT 61.175 2.379 61.2 2.645 ;
      RECT 61.13 2.358 61.175 2.658 ;
      RECT 61.12 2.342 61.13 2.668 ;
      RECT 61.105 2.335 61.12 2.678 ;
      RECT 61.095 2.328 61.105 2.695 ;
      RECT 61.09 2.325 61.095 2.725 ;
      RECT 61.085 2.323 61.09 2.755 ;
      RECT 61.08 2.321 61.085 2.792 ;
      RECT 61.065 2.317 61.08 2.859 ;
      RECT 61.065 3.15 61.075 3.35 ;
      RECT 61.06 2.313 61.065 2.985 ;
      RECT 61.06 3.137 61.065 3.355 ;
      RECT 61.055 2.311 61.06 3.07 ;
      RECT 61.055 3.127 61.06 3.355 ;
      RECT 61.04 2.282 61.055 3.355 ;
      RECT 61.025 2.255 61.04 3.355 ;
      RECT 60.95 2.25 60.955 2.605 ;
      RECT 60.95 2.66 60.955 3.355 ;
      RECT 60.935 2.25 60.95 2.583 ;
      RECT 60.945 2.682 60.95 3.355 ;
      RECT 60.935 2.722 60.945 3.355 ;
      RECT 60.9 2.25 60.935 2.525 ;
      RECT 60.93 2.757 60.935 3.355 ;
      RECT 60.915 2.812 60.93 3.355 ;
      RECT 60.91 2.877 60.915 3.355 ;
      RECT 60.895 2.925 60.91 3.355 ;
      RECT 60.87 2.25 60.9 2.48 ;
      RECT 60.89 2.98 60.895 3.355 ;
      RECT 60.875 3.04 60.89 3.355 ;
      RECT 60.87 3.088 60.875 3.353 ;
      RECT 60.865 2.25 60.87 2.473 ;
      RECT 60.865 3.12 60.87 3.348 ;
      RECT 60.84 2.25 60.865 2.465 ;
      RECT 60.83 2.255 60.84 2.455 ;
      RECT 61.045 3.53 61.065 3.77 ;
      RECT 60.275 3.46 60.28 3.67 ;
      RECT 61.555 3.533 61.565 3.728 ;
      RECT 61.55 3.523 61.555 3.731 ;
      RECT 61.47 3.52 61.55 3.754 ;
      RECT 61.466 3.52 61.47 3.776 ;
      RECT 61.38 3.52 61.466 3.786 ;
      RECT 61.365 3.52 61.38 3.794 ;
      RECT 61.336 3.521 61.365 3.792 ;
      RECT 61.25 3.526 61.336 3.788 ;
      RECT 61.237 3.53 61.25 3.784 ;
      RECT 61.151 3.53 61.237 3.78 ;
      RECT 61.065 3.53 61.151 3.774 ;
      RECT 60.981 3.53 61.045 3.768 ;
      RECT 60.895 3.53 60.981 3.763 ;
      RECT 60.875 3.53 60.895 3.759 ;
      RECT 60.815 3.525 60.875 3.756 ;
      RECT 60.787 3.519 60.815 3.753 ;
      RECT 60.701 3.514 60.787 3.749 ;
      RECT 60.615 3.508 60.701 3.743 ;
      RECT 60.54 3.49 60.615 3.738 ;
      RECT 60.505 3.467 60.54 3.734 ;
      RECT 60.495 3.457 60.505 3.733 ;
      RECT 60.44 3.455 60.495 3.732 ;
      RECT 60.365 3.455 60.44 3.728 ;
      RECT 60.355 3.455 60.365 3.723 ;
      RECT 60.34 3.455 60.355 3.715 ;
      RECT 60.29 3.457 60.34 3.693 ;
      RECT 60.28 3.46 60.29 3.673 ;
      RECT 60.27 3.465 60.275 3.668 ;
      RECT 60.265 3.47 60.27 3.663 ;
      RECT 60.39 2.635 60.65 2.895 ;
      RECT 60.39 2.65 60.67 2.86 ;
      RECT 60.39 2.655 60.68 2.855 ;
      RECT 58.375 2.115 58.635 2.375 ;
      RECT 58.365 2.145 58.635 2.355 ;
      RECT 60.285 2.06 60.545 2.32 ;
      RECT 60.28 2.135 60.285 2.321 ;
      RECT 60.255 2.14 60.28 2.323 ;
      RECT 60.24 2.147 60.255 2.326 ;
      RECT 60.18 2.165 60.24 2.331 ;
      RECT 60.15 2.185 60.18 2.338 ;
      RECT 60.125 2.193 60.15 2.343 ;
      RECT 60.1 2.201 60.125 2.345 ;
      RECT 60.082 2.205 60.1 2.344 ;
      RECT 59.996 2.203 60.082 2.344 ;
      RECT 59.91 2.201 59.996 2.344 ;
      RECT 59.824 2.199 59.91 2.343 ;
      RECT 59.738 2.197 59.824 2.343 ;
      RECT 59.652 2.195 59.738 2.343 ;
      RECT 59.566 2.193 59.652 2.343 ;
      RECT 59.48 2.191 59.566 2.342 ;
      RECT 59.462 2.19 59.48 2.342 ;
      RECT 59.376 2.189 59.462 2.342 ;
      RECT 59.29 2.187 59.376 2.342 ;
      RECT 59.204 2.186 59.29 2.341 ;
      RECT 59.118 2.185 59.204 2.341 ;
      RECT 59.032 2.183 59.118 2.341 ;
      RECT 58.946 2.182 59.032 2.341 ;
      RECT 58.86 2.18 58.946 2.34 ;
      RECT 58.836 2.178 58.86 2.34 ;
      RECT 58.75 2.171 58.836 2.34 ;
      RECT 58.721 2.163 58.75 2.34 ;
      RECT 58.635 2.155 58.721 2.34 ;
      RECT 58.355 2.152 58.365 2.35 ;
      RECT 59.86 3.115 59.865 3.465 ;
      RECT 59.63 3.205 59.77 3.465 ;
      RECT 60.105 2.89 60.15 3.1 ;
      RECT 60.16 2.901 60.17 3.095 ;
      RECT 60.15 2.893 60.16 3.1 ;
      RECT 60.085 2.89 60.105 3.105 ;
      RECT 60.055 2.89 60.085 3.128 ;
      RECT 60.045 2.89 60.055 3.153 ;
      RECT 60.04 2.89 60.045 3.163 ;
      RECT 59.985 2.89 60.04 3.203 ;
      RECT 59.98 2.89 59.985 3.243 ;
      RECT 59.975 2.892 59.98 3.248 ;
      RECT 59.96 2.902 59.975 3.259 ;
      RECT 59.915 2.96 59.96 3.295 ;
      RECT 59.905 3.015 59.915 3.329 ;
      RECT 59.89 3.042 59.905 3.345 ;
      RECT 59.88 3.069 59.89 3.465 ;
      RECT 59.865 3.092 59.88 3.465 ;
      RECT 59.855 3.132 59.86 3.465 ;
      RECT 59.85 3.142 59.855 3.465 ;
      RECT 59.845 3.157 59.85 3.465 ;
      RECT 59.835 3.162 59.845 3.465 ;
      RECT 59.77 3.185 59.835 3.465 ;
      RECT 59.27 2.68 59.46 2.89 ;
      RECT 57.845 2.605 58.105 2.865 ;
      RECT 58.195 2.6 58.29 2.81 ;
      RECT 58.17 2.615 58.18 2.81 ;
      RECT 59.46 2.687 59.47 2.885 ;
      RECT 59.26 2.687 59.27 2.885 ;
      RECT 59.245 2.702 59.26 2.875 ;
      RECT 59.24 2.71 59.245 2.868 ;
      RECT 59.23 2.713 59.24 2.865 ;
      RECT 59.195 2.712 59.23 2.863 ;
      RECT 59.166 2.708 59.195 2.86 ;
      RECT 59.08 2.703 59.166 2.857 ;
      RECT 59.02 2.697 59.08 2.853 ;
      RECT 58.991 2.693 59.02 2.85 ;
      RECT 58.905 2.685 58.991 2.847 ;
      RECT 58.896 2.679 58.905 2.845 ;
      RECT 58.81 2.674 58.896 2.843 ;
      RECT 58.787 2.669 58.81 2.84 ;
      RECT 58.701 2.663 58.787 2.837 ;
      RECT 58.615 2.654 58.701 2.832 ;
      RECT 58.605 2.649 58.615 2.83 ;
      RECT 58.586 2.648 58.605 2.829 ;
      RECT 58.5 2.643 58.586 2.825 ;
      RECT 58.48 2.638 58.5 2.821 ;
      RECT 58.42 2.633 58.48 2.818 ;
      RECT 58.395 2.623 58.42 2.816 ;
      RECT 58.39 2.616 58.395 2.815 ;
      RECT 58.38 2.607 58.39 2.814 ;
      RECT 58.376 2.6 58.38 2.814 ;
      RECT 58.29 2.6 58.376 2.812 ;
      RECT 58.18 2.607 58.195 2.81 ;
      RECT 58.165 2.617 58.17 2.81 ;
      RECT 58.145 2.62 58.165 2.807 ;
      RECT 58.115 2.62 58.145 2.803 ;
      RECT 58.105 2.62 58.115 2.803 ;
      RECT 59.02 3.115 59.28 3.375 ;
      RECT 58.95 3.125 59.28 3.335 ;
      RECT 58.94 3.132 59.28 3.33 ;
      RECT 58.36 3.12 58.62 3.38 ;
      RECT 58.36 3.16 58.725 3.37 ;
      RECT 58.36 3.162 58.73 3.369 ;
      RECT 58.36 3.17 58.735 3.366 ;
      RECT 57.285 2.245 57.385 3.77 ;
      RECT 57.475 3.385 57.525 3.645 ;
      RECT 57.47 2.258 57.475 2.445 ;
      RECT 57.465 3.366 57.475 3.645 ;
      RECT 57.465 2.255 57.47 2.453 ;
      RECT 57.45 2.249 57.465 2.46 ;
      RECT 57.46 3.354 57.465 3.728 ;
      RECT 57.45 3.342 57.46 3.765 ;
      RECT 57.44 2.245 57.45 2.467 ;
      RECT 57.44 3.327 57.45 3.77 ;
      RECT 57.435 2.245 57.44 2.475 ;
      RECT 57.415 3.297 57.44 3.77 ;
      RECT 57.395 2.245 57.435 2.523 ;
      RECT 57.405 3.257 57.415 3.77 ;
      RECT 57.395 3.212 57.405 3.77 ;
      RECT 57.39 2.245 57.395 2.593 ;
      RECT 57.39 3.17 57.395 3.77 ;
      RECT 57.385 2.245 57.39 3.07 ;
      RECT 57.385 3.152 57.39 3.77 ;
      RECT 57.275 2.248 57.285 3.77 ;
      RECT 57.26 2.255 57.275 3.766 ;
      RECT 57.255 2.265 57.26 3.761 ;
      RECT 57.25 2.465 57.255 3.653 ;
      RECT 57.245 2.55 57.25 3.205 ;
      RECT 56.125 7.765 56.415 7.995 ;
      RECT 56.185 6.285 56.355 7.995 ;
      RECT 56.13 6.655 56.48 7.005 ;
      RECT 56.125 6.285 56.415 6.515 ;
      RECT 56.125 2.365 56.415 2.595 ;
      RECT 56.185 0.885 56.355 2.595 ;
      RECT 56.125 0.885 56.415 1.115 ;
      RECT 55.715 2.735 56.045 2.965 ;
      RECT 55.715 2.765 56.215 2.935 ;
      RECT 55.715 2.395 55.905 2.965 ;
      RECT 55.135 2.365 55.425 2.595 ;
      RECT 55.135 2.395 55.905 2.565 ;
      RECT 55.195 0.885 55.365 2.595 ;
      RECT 55.135 0.885 55.425 1.115 ;
      RECT 55.135 7.765 55.425 7.995 ;
      RECT 55.195 6.285 55.365 7.995 ;
      RECT 55.135 6.285 55.425 6.515 ;
      RECT 55.135 6.325 55.985 6.485 ;
      RECT 55.815 5.915 55.985 6.485 ;
      RECT 55.135 6.32 55.525 6.485 ;
      RECT 55.755 5.915 56.045 6.145 ;
      RECT 55.755 5.945 56.215 6.115 ;
      RECT 54.765 2.735 55.055 2.965 ;
      RECT 54.765 2.765 55.225 2.935 ;
      RECT 54.825 1.655 54.99 2.965 ;
      RECT 53.34 1.625 53.63 1.855 ;
      RECT 53.34 1.655 54.99 1.825 ;
      RECT 53.4 0.885 53.57 1.855 ;
      RECT 53.34 0.885 53.63 1.115 ;
      RECT 53.34 7.765 53.63 7.995 ;
      RECT 53.4 7.025 53.57 7.995 ;
      RECT 53.4 7.12 54.99 7.29 ;
      RECT 54.82 5.915 54.99 7.29 ;
      RECT 53.34 7.025 53.63 7.255 ;
      RECT 54.765 5.915 55.055 6.145 ;
      RECT 54.765 5.945 55.225 6.115 ;
      RECT 51.375 3.43 51.725 3.78 ;
      RECT 51.465 2.025 51.635 3.78 ;
      RECT 53.77 1.965 54.12 2.315 ;
      RECT 51.465 2.025 53.085 2.2 ;
      RECT 51.465 2.025 54.12 2.195 ;
      RECT 53.795 6.655 54.12 6.98 ;
      RECT 49.225 6.615 49.575 6.965 ;
      RECT 53.77 6.655 54.12 6.885 ;
      RECT 49.01 6.655 49.575 6.885 ;
      RECT 48.84 6.685 54.12 6.855 ;
      RECT 52.995 2.365 53.315 2.685 ;
      RECT 52.965 2.365 53.315 2.595 ;
      RECT 52.795 2.395 53.315 2.565 ;
      RECT 52.995 6.225 53.315 6.545 ;
      RECT 52.965 6.285 53.315 6.515 ;
      RECT 52.795 6.315 53.315 6.485 ;
      RECT 51.95 2.705 52.3 3.055 ;
      RECT 51.95 2.765 52.43 2.935 ;
      RECT 51.94 5.84 52.29 6.19 ;
      RECT 47.21 5.915 47.5 6.145 ;
      RECT 47.21 5.945 52.43 6.115 ;
      RECT 48.775 3.665 48.815 3.925 ;
      RECT 48.815 3.645 48.82 3.655 ;
      RECT 50.145 2.89 50.155 3.111 ;
      RECT 50.075 2.885 50.145 3.236 ;
      RECT 50.065 2.885 50.075 3.363 ;
      RECT 50.04 2.885 50.065 3.41 ;
      RECT 50.015 2.885 50.04 3.488 ;
      RECT 49.995 2.885 50.015 3.558 ;
      RECT 49.97 2.885 49.995 3.598 ;
      RECT 49.96 2.885 49.97 3.618 ;
      RECT 49.95 2.887 49.96 3.626 ;
      RECT 49.945 2.892 49.95 3.083 ;
      RECT 49.945 3.092 49.95 3.627 ;
      RECT 49.94 3.137 49.945 3.628 ;
      RECT 49.93 3.202 49.94 3.629 ;
      RECT 49.92 3.297 49.93 3.631 ;
      RECT 49.915 3.35 49.92 3.633 ;
      RECT 49.91 3.37 49.915 3.634 ;
      RECT 49.855 3.395 49.91 3.64 ;
      RECT 49.815 3.43 49.855 3.649 ;
      RECT 49.805 3.447 49.815 3.654 ;
      RECT 49.796 3.453 49.805 3.656 ;
      RECT 49.71 3.491 49.796 3.667 ;
      RECT 49.705 3.53 49.71 3.677 ;
      RECT 49.63 3.537 49.705 3.687 ;
      RECT 49.61 3.547 49.63 3.698 ;
      RECT 49.58 3.554 49.61 3.706 ;
      RECT 49.555 3.561 49.58 3.713 ;
      RECT 49.531 3.567 49.555 3.718 ;
      RECT 49.445 3.58 49.531 3.73 ;
      RECT 49.367 3.587 49.445 3.748 ;
      RECT 49.281 3.582 49.367 3.766 ;
      RECT 49.195 3.577 49.281 3.786 ;
      RECT 49.115 3.571 49.195 3.803 ;
      RECT 49.05 3.567 49.115 3.832 ;
      RECT 49.045 3.281 49.05 3.305 ;
      RECT 49.035 3.557 49.05 3.86 ;
      RECT 49.04 3.275 49.045 3.345 ;
      RECT 49.035 3.269 49.04 3.415 ;
      RECT 49.03 3.263 49.035 3.493 ;
      RECT 49.03 3.54 49.035 3.925 ;
      RECT 49.022 3.26 49.03 3.925 ;
      RECT 48.936 3.258 49.022 3.925 ;
      RECT 48.85 3.256 48.936 3.925 ;
      RECT 48.84 3.257 48.85 3.925 ;
      RECT 48.835 3.262 48.84 3.925 ;
      RECT 48.825 3.275 48.835 3.925 ;
      RECT 48.82 3.297 48.825 3.925 ;
      RECT 48.815 3.657 48.82 3.925 ;
      RECT 49.445 3.125 49.45 3.345 ;
      RECT 49.95 2.16 49.985 2.42 ;
      RECT 49.935 2.16 49.95 2.428 ;
      RECT 49.906 2.16 49.935 2.45 ;
      RECT 49.82 2.16 49.906 2.51 ;
      RECT 49.8 2.16 49.82 2.575 ;
      RECT 49.74 2.16 49.8 2.74 ;
      RECT 49.735 2.16 49.74 2.888 ;
      RECT 49.73 2.16 49.735 2.9 ;
      RECT 49.725 2.16 49.73 2.926 ;
      RECT 49.695 2.346 49.725 3.006 ;
      RECT 49.69 2.394 49.695 3.095 ;
      RECT 49.685 2.408 49.69 3.11 ;
      RECT 49.68 2.427 49.685 3.14 ;
      RECT 49.675 2.442 49.68 3.156 ;
      RECT 49.67 2.457 49.675 3.178 ;
      RECT 49.665 2.477 49.67 3.2 ;
      RECT 49.655 2.497 49.665 3.233 ;
      RECT 49.64 2.539 49.655 3.295 ;
      RECT 49.635 2.57 49.64 3.335 ;
      RECT 49.63 2.582 49.635 3.34 ;
      RECT 49.625 2.594 49.63 3.345 ;
      RECT 49.62 2.607 49.625 3.345 ;
      RECT 49.615 2.625 49.62 3.345 ;
      RECT 49.61 2.645 49.615 3.345 ;
      RECT 49.605 2.657 49.61 3.345 ;
      RECT 49.6 2.67 49.605 3.345 ;
      RECT 49.58 2.705 49.6 3.345 ;
      RECT 49.53 2.807 49.58 3.345 ;
      RECT 49.525 2.892 49.53 3.345 ;
      RECT 49.52 2.9 49.525 3.345 ;
      RECT 49.515 2.917 49.52 3.345 ;
      RECT 49.51 2.932 49.515 3.345 ;
      RECT 49.475 2.997 49.51 3.345 ;
      RECT 49.46 3.062 49.475 3.345 ;
      RECT 49.455 3.092 49.46 3.345 ;
      RECT 49.45 3.117 49.455 3.345 ;
      RECT 49.435 3.127 49.445 3.345 ;
      RECT 49.42 3.14 49.435 3.338 ;
      RECT 49.165 2.73 49.235 2.94 ;
      RECT 48.955 2.707 48.96 2.9 ;
      RECT 46.41 2.635 46.67 2.895 ;
      RECT 49.245 2.917 49.25 2.92 ;
      RECT 49.235 2.735 49.245 2.935 ;
      RECT 49.136 2.728 49.165 2.94 ;
      RECT 49.05 2.72 49.136 2.94 ;
      RECT 49.035 2.714 49.05 2.938 ;
      RECT 49.015 2.713 49.035 2.925 ;
      RECT 49.01 2.712 49.015 2.908 ;
      RECT 48.96 2.709 49.01 2.903 ;
      RECT 48.93 2.706 48.955 2.898 ;
      RECT 48.91 2.704 48.93 2.893 ;
      RECT 48.895 2.702 48.91 2.89 ;
      RECT 48.865 2.7 48.895 2.888 ;
      RECT 48.8 2.696 48.865 2.88 ;
      RECT 48.77 2.691 48.8 2.875 ;
      RECT 48.75 2.689 48.77 2.873 ;
      RECT 48.72 2.686 48.75 2.868 ;
      RECT 48.66 2.682 48.72 2.86 ;
      RECT 48.655 2.679 48.66 2.855 ;
      RECT 48.585 2.677 48.655 2.85 ;
      RECT 48.556 2.673 48.585 2.843 ;
      RECT 48.47 2.668 48.556 2.835 ;
      RECT 48.436 2.663 48.47 2.827 ;
      RECT 48.35 2.655 48.436 2.819 ;
      RECT 48.311 2.648 48.35 2.811 ;
      RECT 48.225 2.643 48.311 2.803 ;
      RECT 48.16 2.637 48.225 2.793 ;
      RECT 48.14 2.632 48.16 2.788 ;
      RECT 48.131 2.629 48.14 2.787 ;
      RECT 48.045 2.625 48.131 2.781 ;
      RECT 48.005 2.621 48.045 2.773 ;
      RECT 47.985 2.617 48.005 2.771 ;
      RECT 47.925 2.617 47.985 2.768 ;
      RECT 47.905 2.62 47.925 2.766 ;
      RECT 47.884 2.62 47.905 2.766 ;
      RECT 47.798 2.622 47.884 2.77 ;
      RECT 47.712 2.624 47.798 2.776 ;
      RECT 47.626 2.626 47.712 2.783 ;
      RECT 47.54 2.629 47.626 2.789 ;
      RECT 47.506 2.63 47.54 2.794 ;
      RECT 47.42 2.633 47.506 2.799 ;
      RECT 47.391 2.64 47.42 2.804 ;
      RECT 47.305 2.64 47.391 2.809 ;
      RECT 47.272 2.64 47.305 2.814 ;
      RECT 47.186 2.642 47.272 2.819 ;
      RECT 47.1 2.644 47.186 2.826 ;
      RECT 47.036 2.646 47.1 2.832 ;
      RECT 46.95 2.648 47.036 2.838 ;
      RECT 46.947 2.65 46.95 2.841 ;
      RECT 46.861 2.651 46.947 2.845 ;
      RECT 46.775 2.654 46.861 2.852 ;
      RECT 46.756 2.656 46.775 2.856 ;
      RECT 46.67 2.658 46.756 2.861 ;
      RECT 46.4 2.67 46.41 2.865 ;
      RECT 48.58 7.765 48.87 7.995 ;
      RECT 48.64 7.025 48.81 7.995 ;
      RECT 48.53 7.055 48.905 7.425 ;
      RECT 48.58 7.025 48.87 7.425 ;
      RECT 48.635 2.25 48.82 2.46 ;
      RECT 48.63 2.251 48.825 2.458 ;
      RECT 48.625 2.256 48.835 2.453 ;
      RECT 48.62 2.232 48.625 2.45 ;
      RECT 48.59 2.229 48.62 2.443 ;
      RECT 48.585 2.225 48.59 2.434 ;
      RECT 48.55 2.256 48.835 2.429 ;
      RECT 48.325 2.165 48.585 2.425 ;
      RECT 48.625 2.234 48.63 2.453 ;
      RECT 48.63 2.235 48.635 2.458 ;
      RECT 48.325 2.247 48.705 2.425 ;
      RECT 48.325 2.245 48.69 2.425 ;
      RECT 48.325 2.24 48.68 2.425 ;
      RECT 48.28 3.155 48.33 3.44 ;
      RECT 48.225 3.125 48.23 3.44 ;
      RECT 48.195 3.105 48.2 3.44 ;
      RECT 48.345 3.155 48.405 3.415 ;
      RECT 48.34 3.155 48.345 3.423 ;
      RECT 48.33 3.155 48.34 3.435 ;
      RECT 48.245 3.145 48.28 3.44 ;
      RECT 48.24 3.132 48.245 3.44 ;
      RECT 48.23 3.127 48.24 3.44 ;
      RECT 48.21 3.117 48.225 3.44 ;
      RECT 48.2 3.11 48.21 3.44 ;
      RECT 48.19 3.102 48.195 3.44 ;
      RECT 48.16 3.092 48.19 3.44 ;
      RECT 48.145 3.08 48.16 3.44 ;
      RECT 48.13 3.07 48.145 3.435 ;
      RECT 48.11 3.06 48.13 3.41 ;
      RECT 48.1 3.052 48.11 3.387 ;
      RECT 48.07 3.035 48.1 3.377 ;
      RECT 48.065 3.012 48.07 3.368 ;
      RECT 48.06 2.999 48.065 3.366 ;
      RECT 48.045 2.975 48.06 3.36 ;
      RECT 48.04 2.951 48.045 3.354 ;
      RECT 48.03 2.94 48.04 3.349 ;
      RECT 48.025 2.93 48.03 3.345 ;
      RECT 48.02 2.922 48.025 3.342 ;
      RECT 48.01 2.917 48.02 3.338 ;
      RECT 48.005 2.912 48.01 3.334 ;
      RECT 47.92 2.91 48.005 3.309 ;
      RECT 47.89 2.91 47.92 3.275 ;
      RECT 47.875 2.91 47.89 3.258 ;
      RECT 47.82 2.91 47.875 3.203 ;
      RECT 47.815 2.915 47.82 3.152 ;
      RECT 47.805 2.92 47.815 3.142 ;
      RECT 47.8 2.93 47.805 3.128 ;
      RECT 47.75 3.67 48.01 3.93 ;
      RECT 47.67 3.685 48.01 3.906 ;
      RECT 47.65 3.685 48.01 3.901 ;
      RECT 47.626 3.685 48.01 3.899 ;
      RECT 47.54 3.685 48.01 3.894 ;
      RECT 47.39 3.625 47.65 3.89 ;
      RECT 47.345 3.685 48.01 3.885 ;
      RECT 47.34 3.692 48.01 3.88 ;
      RECT 47.355 3.68 47.67 3.89 ;
      RECT 47.245 2.115 47.505 2.375 ;
      RECT 47.245 2.172 47.51 2.368 ;
      RECT 47.245 2.202 47.515 2.3 ;
      RECT 47.305 2.633 47.42 2.635 ;
      RECT 47.391 2.63 47.42 2.635 ;
      RECT 46.415 3.634 46.44 3.874 ;
      RECT 46.4 3.637 46.49 3.868 ;
      RECT 46.395 3.642 46.576 3.863 ;
      RECT 46.39 3.65 46.64 3.861 ;
      RECT 46.39 3.65 46.65 3.86 ;
      RECT 46.385 3.657 46.66 3.853 ;
      RECT 46.385 3.657 46.746 3.842 ;
      RECT 46.38 3.692 46.746 3.838 ;
      RECT 46.38 3.692 46.755 3.827 ;
      RECT 46.66 3.565 46.92 3.825 ;
      RECT 46.37 3.742 46.92 3.823 ;
      RECT 46.64 3.61 46.66 3.858 ;
      RECT 46.576 3.613 46.64 3.862 ;
      RECT 46.49 3.618 46.576 3.867 ;
      RECT 46.42 3.629 46.92 3.825 ;
      RECT 46.44 3.623 46.49 3.872 ;
      RECT 46.565 2.1 46.575 2.362 ;
      RECT 46.555 2.157 46.565 2.365 ;
      RECT 46.53 2.162 46.555 2.371 ;
      RECT 46.505 2.166 46.53 2.383 ;
      RECT 46.495 2.169 46.505 2.393 ;
      RECT 46.49 2.17 46.495 2.398 ;
      RECT 46.485 2.171 46.49 2.403 ;
      RECT 46.48 2.172 46.485 2.405 ;
      RECT 46.455 2.175 46.48 2.408 ;
      RECT 46.425 2.181 46.455 2.411 ;
      RECT 46.36 2.192 46.425 2.414 ;
      RECT 46.315 2.2 46.36 2.418 ;
      RECT 46.3 2.2 46.315 2.426 ;
      RECT 46.295 2.201 46.3 2.433 ;
      RECT 46.29 2.203 46.295 2.436 ;
      RECT 46.285 2.207 46.29 2.439 ;
      RECT 46.275 2.215 46.285 2.443 ;
      RECT 46.27 2.228 46.275 2.448 ;
      RECT 46.265 2.236 46.27 2.45 ;
      RECT 46.26 2.242 46.265 2.45 ;
      RECT 46.255 2.246 46.26 2.453 ;
      RECT 46.25 2.248 46.255 2.456 ;
      RECT 46.245 2.251 46.25 2.459 ;
      RECT 46.235 2.256 46.245 2.463 ;
      RECT 46.23 2.262 46.235 2.468 ;
      RECT 46.22 2.268 46.23 2.472 ;
      RECT 46.205 2.275 46.22 2.478 ;
      RECT 46.176 2.289 46.205 2.488 ;
      RECT 46.09 2.324 46.176 2.52 ;
      RECT 46.07 2.357 46.09 2.549 ;
      RECT 46.05 2.37 46.07 2.56 ;
      RECT 46.03 2.382 46.05 2.571 ;
      RECT 45.98 2.404 46.03 2.591 ;
      RECT 45.965 2.422 45.98 2.608 ;
      RECT 45.96 2.428 45.965 2.611 ;
      RECT 45.955 2.432 45.96 2.614 ;
      RECT 45.95 2.436 45.955 2.618 ;
      RECT 45.945 2.438 45.95 2.621 ;
      RECT 45.935 2.445 45.945 2.624 ;
      RECT 45.93 2.45 45.935 2.628 ;
      RECT 45.925 2.452 45.93 2.631 ;
      RECT 45.92 2.456 45.925 2.634 ;
      RECT 45.915 2.458 45.92 2.638 ;
      RECT 45.9 2.463 45.915 2.643 ;
      RECT 45.895 2.468 45.9 2.646 ;
      RECT 45.89 2.476 45.895 2.649 ;
      RECT 45.885 2.478 45.89 2.652 ;
      RECT 45.88 2.48 45.885 2.655 ;
      RECT 45.87 2.482 45.88 2.661 ;
      RECT 45.835 2.496 45.87 2.673 ;
      RECT 45.825 2.511 45.835 2.683 ;
      RECT 45.75 2.54 45.825 2.707 ;
      RECT 45.745 2.565 45.75 2.73 ;
      RECT 45.73 2.569 45.745 2.736 ;
      RECT 45.72 2.577 45.73 2.741 ;
      RECT 45.69 2.59 45.72 2.745 ;
      RECT 45.68 2.605 45.69 2.75 ;
      RECT 45.67 2.61 45.68 2.753 ;
      RECT 45.665 2.612 45.67 2.755 ;
      RECT 45.65 2.615 45.665 2.758 ;
      RECT 45.645 2.617 45.65 2.761 ;
      RECT 45.625 2.622 45.645 2.765 ;
      RECT 45.595 2.627 45.625 2.773 ;
      RECT 45.57 2.634 45.595 2.781 ;
      RECT 45.565 2.639 45.57 2.786 ;
      RECT 45.535 2.642 45.565 2.79 ;
      RECT 45.495 2.645 45.535 2.8 ;
      RECT 45.46 2.642 45.495 2.812 ;
      RECT 45.45 2.638 45.46 2.819 ;
      RECT 45.425 2.634 45.45 2.825 ;
      RECT 45.42 2.63 45.425 2.83 ;
      RECT 45.38 2.627 45.42 2.83 ;
      RECT 45.365 2.612 45.38 2.831 ;
      RECT 45.342 2.6 45.365 2.831 ;
      RECT 45.256 2.6 45.342 2.832 ;
      RECT 45.17 2.6 45.256 2.834 ;
      RECT 45.15 2.6 45.17 2.831 ;
      RECT 45.145 2.605 45.15 2.826 ;
      RECT 45.14 2.61 45.145 2.824 ;
      RECT 45.13 2.62 45.14 2.822 ;
      RECT 45.125 2.626 45.13 2.815 ;
      RECT 45.12 2.628 45.125 2.8 ;
      RECT 45.115 2.632 45.12 2.79 ;
      RECT 46.575 2.1 46.825 2.36 ;
      RECT 44.3 3.635 44.56 3.895 ;
      RECT 46.595 3.125 46.6 3.335 ;
      RECT 46.6 3.13 46.61 3.33 ;
      RECT 46.55 3.125 46.595 3.35 ;
      RECT 46.54 3.125 46.55 3.37 ;
      RECT 46.521 3.125 46.54 3.375 ;
      RECT 46.435 3.125 46.521 3.372 ;
      RECT 46.405 3.127 46.435 3.37 ;
      RECT 46.35 3.137 46.405 3.368 ;
      RECT 46.285 3.151 46.35 3.366 ;
      RECT 46.28 3.159 46.285 3.365 ;
      RECT 46.265 3.162 46.28 3.363 ;
      RECT 46.2 3.172 46.265 3.359 ;
      RECT 46.152 3.186 46.2 3.36 ;
      RECT 46.066 3.203 46.152 3.374 ;
      RECT 45.98 3.224 46.066 3.391 ;
      RECT 45.96 3.237 45.98 3.401 ;
      RECT 45.915 3.245 45.96 3.408 ;
      RECT 45.88 3.253 45.915 3.416 ;
      RECT 45.846 3.261 45.88 3.424 ;
      RECT 45.76 3.275 45.846 3.436 ;
      RECT 45.725 3.292 45.76 3.448 ;
      RECT 45.716 3.301 45.725 3.452 ;
      RECT 45.63 3.319 45.716 3.469 ;
      RECT 45.571 3.346 45.63 3.496 ;
      RECT 45.485 3.373 45.571 3.524 ;
      RECT 45.465 3.395 45.485 3.544 ;
      RECT 45.405 3.41 45.465 3.56 ;
      RECT 45.395 3.422 45.405 3.573 ;
      RECT 45.39 3.427 45.395 3.576 ;
      RECT 45.38 3.43 45.39 3.579 ;
      RECT 45.375 3.432 45.38 3.582 ;
      RECT 45.345 3.44 45.375 3.589 ;
      RECT 45.33 3.447 45.345 3.597 ;
      RECT 45.32 3.452 45.33 3.601 ;
      RECT 45.315 3.455 45.32 3.604 ;
      RECT 45.305 3.457 45.315 3.607 ;
      RECT 45.27 3.467 45.305 3.616 ;
      RECT 45.195 3.49 45.27 3.638 ;
      RECT 45.175 3.508 45.195 3.656 ;
      RECT 45.145 3.515 45.175 3.666 ;
      RECT 45.125 3.523 45.145 3.676 ;
      RECT 45.115 3.529 45.125 3.683 ;
      RECT 45.096 3.534 45.115 3.689 ;
      RECT 45.01 3.554 45.096 3.709 ;
      RECT 44.995 3.574 45.01 3.728 ;
      RECT 44.95 3.586 44.995 3.739 ;
      RECT 44.885 3.607 44.95 3.762 ;
      RECT 44.845 3.627 44.885 3.783 ;
      RECT 44.835 3.637 44.845 3.793 ;
      RECT 44.785 3.649 44.835 3.804 ;
      RECT 44.765 3.665 44.785 3.816 ;
      RECT 44.735 3.675 44.765 3.822 ;
      RECT 44.725 3.68 44.735 3.824 ;
      RECT 44.656 3.681 44.725 3.83 ;
      RECT 44.57 3.683 44.656 3.84 ;
      RECT 44.56 3.684 44.57 3.845 ;
      RECT 45.83 3.71 46.02 3.92 ;
      RECT 45.82 3.715 46.03 3.913 ;
      RECT 45.805 3.715 46.03 3.878 ;
      RECT 45.725 3.6 45.985 3.86 ;
      RECT 44.64 3.13 44.825 3.425 ;
      RECT 44.63 3.13 44.825 3.423 ;
      RECT 44.615 3.13 44.83 3.418 ;
      RECT 44.615 3.13 44.835 3.415 ;
      RECT 44.61 3.13 44.835 3.413 ;
      RECT 44.605 3.385 44.835 3.403 ;
      RECT 44.61 3.13 44.87 3.39 ;
      RECT 44.57 2.165 44.83 2.425 ;
      RECT 44.38 2.09 44.466 2.423 ;
      RECT 44.355 2.094 44.51 2.419 ;
      RECT 44.466 2.086 44.51 2.419 ;
      RECT 44.466 2.087 44.515 2.418 ;
      RECT 44.38 2.092 44.53 2.417 ;
      RECT 44.355 2.1 44.57 2.416 ;
      RECT 44.35 2.095 44.53 2.411 ;
      RECT 44.34 2.11 44.57 2.318 ;
      RECT 44.34 2.162 44.77 2.318 ;
      RECT 44.34 2.155 44.75 2.318 ;
      RECT 44.34 2.142 44.72 2.318 ;
      RECT 44.34 2.13 44.66 2.318 ;
      RECT 44.34 2.115 44.635 2.318 ;
      RECT 43.54 2.745 43.675 3.04 ;
      RECT 43.8 2.768 43.805 2.955 ;
      RECT 44.52 2.665 44.665 2.9 ;
      RECT 44.68 2.665 44.685 2.89 ;
      RECT 44.715 2.676 44.72 2.87 ;
      RECT 44.71 2.668 44.715 2.875 ;
      RECT 44.69 2.665 44.71 2.88 ;
      RECT 44.685 2.665 44.69 2.888 ;
      RECT 44.675 2.665 44.68 2.893 ;
      RECT 44.665 2.665 44.675 2.898 ;
      RECT 44.495 2.667 44.52 2.9 ;
      RECT 44.445 2.674 44.495 2.9 ;
      RECT 44.44 2.679 44.445 2.9 ;
      RECT 44.401 2.684 44.44 2.901 ;
      RECT 44.315 2.696 44.401 2.902 ;
      RECT 44.306 2.706 44.315 2.902 ;
      RECT 44.22 2.715 44.306 2.904 ;
      RECT 44.196 2.725 44.22 2.906 ;
      RECT 44.11 2.736 44.196 2.907 ;
      RECT 44.08 2.747 44.11 2.909 ;
      RECT 44.05 2.752 44.08 2.911 ;
      RECT 44.025 2.758 44.05 2.914 ;
      RECT 44.01 2.763 44.025 2.915 ;
      RECT 43.965 2.769 44.01 2.915 ;
      RECT 43.96 2.774 43.965 2.916 ;
      RECT 43.94 2.774 43.96 2.918 ;
      RECT 43.92 2.772 43.94 2.923 ;
      RECT 43.885 2.771 43.92 2.93 ;
      RECT 43.855 2.77 43.885 2.94 ;
      RECT 43.805 2.769 43.855 2.95 ;
      RECT 43.715 2.766 43.8 3.04 ;
      RECT 43.69 2.76 43.715 3.04 ;
      RECT 43.675 2.75 43.69 3.04 ;
      RECT 43.49 2.745 43.54 2.96 ;
      RECT 43.48 2.75 43.49 2.95 ;
      RECT 43.72 3.225 43.98 3.485 ;
      RECT 43.72 3.225 44.01 3.378 ;
      RECT 43.72 3.225 44.045 3.363 ;
      RECT 43.975 3.145 44.165 3.355 ;
      RECT 43.965 3.15 44.175 3.348 ;
      RECT 43.93 3.22 44.175 3.348 ;
      RECT 43.96 3.162 43.98 3.485 ;
      RECT 43.945 3.21 44.175 3.348 ;
      RECT 43.95 3.182 43.98 3.485 ;
      RECT 43.03 2.25 43.1 3.355 ;
      RECT 43.765 2.355 44.025 2.615 ;
      RECT 43.345 2.401 43.36 2.61 ;
      RECT 43.681 2.414 43.765 2.565 ;
      RECT 43.595 2.411 43.681 2.565 ;
      RECT 43.556 2.409 43.595 2.565 ;
      RECT 43.47 2.407 43.556 2.565 ;
      RECT 43.41 2.405 43.47 2.576 ;
      RECT 43.375 2.403 43.41 2.594 ;
      RECT 43.36 2.401 43.375 2.605 ;
      RECT 43.33 2.401 43.345 2.618 ;
      RECT 43.32 2.401 43.33 2.623 ;
      RECT 43.295 2.4 43.32 2.628 ;
      RECT 43.28 2.395 43.295 2.634 ;
      RECT 43.275 2.388 43.28 2.639 ;
      RECT 43.25 2.379 43.275 2.645 ;
      RECT 43.205 2.358 43.25 2.658 ;
      RECT 43.195 2.342 43.205 2.668 ;
      RECT 43.18 2.335 43.195 2.678 ;
      RECT 43.17 2.328 43.18 2.695 ;
      RECT 43.165 2.325 43.17 2.725 ;
      RECT 43.16 2.323 43.165 2.755 ;
      RECT 43.155 2.321 43.16 2.792 ;
      RECT 43.14 2.317 43.155 2.859 ;
      RECT 43.14 3.15 43.15 3.35 ;
      RECT 43.135 2.313 43.14 2.985 ;
      RECT 43.135 3.137 43.14 3.355 ;
      RECT 43.13 2.311 43.135 3.07 ;
      RECT 43.13 3.127 43.135 3.355 ;
      RECT 43.115 2.282 43.13 3.355 ;
      RECT 43.1 2.255 43.115 3.355 ;
      RECT 43.025 2.25 43.03 2.605 ;
      RECT 43.025 2.66 43.03 3.355 ;
      RECT 43.01 2.25 43.025 2.583 ;
      RECT 43.02 2.682 43.025 3.355 ;
      RECT 43.01 2.722 43.02 3.355 ;
      RECT 42.975 2.25 43.01 2.525 ;
      RECT 43.005 2.757 43.01 3.355 ;
      RECT 42.99 2.812 43.005 3.355 ;
      RECT 42.985 2.877 42.99 3.355 ;
      RECT 42.97 2.925 42.985 3.355 ;
      RECT 42.945 2.25 42.975 2.48 ;
      RECT 42.965 2.98 42.97 3.355 ;
      RECT 42.95 3.04 42.965 3.355 ;
      RECT 42.945 3.088 42.95 3.353 ;
      RECT 42.94 2.25 42.945 2.473 ;
      RECT 42.94 3.12 42.945 3.348 ;
      RECT 42.915 2.25 42.94 2.465 ;
      RECT 42.905 2.255 42.915 2.455 ;
      RECT 43.12 3.53 43.14 3.77 ;
      RECT 42.35 3.46 42.355 3.67 ;
      RECT 43.63 3.533 43.64 3.728 ;
      RECT 43.625 3.523 43.63 3.731 ;
      RECT 43.545 3.52 43.625 3.754 ;
      RECT 43.541 3.52 43.545 3.776 ;
      RECT 43.455 3.52 43.541 3.786 ;
      RECT 43.44 3.52 43.455 3.794 ;
      RECT 43.411 3.521 43.44 3.792 ;
      RECT 43.325 3.526 43.411 3.788 ;
      RECT 43.312 3.53 43.325 3.784 ;
      RECT 43.226 3.53 43.312 3.78 ;
      RECT 43.14 3.53 43.226 3.774 ;
      RECT 43.056 3.53 43.12 3.768 ;
      RECT 42.97 3.53 43.056 3.763 ;
      RECT 42.95 3.53 42.97 3.759 ;
      RECT 42.89 3.525 42.95 3.756 ;
      RECT 42.862 3.519 42.89 3.753 ;
      RECT 42.776 3.514 42.862 3.749 ;
      RECT 42.69 3.508 42.776 3.743 ;
      RECT 42.615 3.49 42.69 3.738 ;
      RECT 42.58 3.467 42.615 3.734 ;
      RECT 42.57 3.457 42.58 3.733 ;
      RECT 42.515 3.455 42.57 3.732 ;
      RECT 42.44 3.455 42.515 3.728 ;
      RECT 42.43 3.455 42.44 3.723 ;
      RECT 42.415 3.455 42.43 3.715 ;
      RECT 42.365 3.457 42.415 3.693 ;
      RECT 42.355 3.46 42.365 3.673 ;
      RECT 42.345 3.465 42.35 3.668 ;
      RECT 42.34 3.47 42.345 3.663 ;
      RECT 42.465 2.635 42.725 2.895 ;
      RECT 42.465 2.65 42.745 2.86 ;
      RECT 42.465 2.655 42.755 2.855 ;
      RECT 40.45 2.115 40.71 2.375 ;
      RECT 40.44 2.145 40.71 2.355 ;
      RECT 42.36 2.06 42.62 2.32 ;
      RECT 42.355 2.135 42.36 2.321 ;
      RECT 42.33 2.14 42.355 2.323 ;
      RECT 42.315 2.147 42.33 2.326 ;
      RECT 42.255 2.165 42.315 2.331 ;
      RECT 42.225 2.185 42.255 2.338 ;
      RECT 42.2 2.193 42.225 2.343 ;
      RECT 42.175 2.201 42.2 2.345 ;
      RECT 42.157 2.205 42.175 2.344 ;
      RECT 42.071 2.203 42.157 2.344 ;
      RECT 41.985 2.201 42.071 2.344 ;
      RECT 41.899 2.199 41.985 2.343 ;
      RECT 41.813 2.197 41.899 2.343 ;
      RECT 41.727 2.195 41.813 2.343 ;
      RECT 41.641 2.193 41.727 2.343 ;
      RECT 41.555 2.191 41.641 2.342 ;
      RECT 41.537 2.19 41.555 2.342 ;
      RECT 41.451 2.189 41.537 2.342 ;
      RECT 41.365 2.187 41.451 2.342 ;
      RECT 41.279 2.186 41.365 2.341 ;
      RECT 41.193 2.185 41.279 2.341 ;
      RECT 41.107 2.183 41.193 2.341 ;
      RECT 41.021 2.182 41.107 2.341 ;
      RECT 40.935 2.18 41.021 2.34 ;
      RECT 40.911 2.178 40.935 2.34 ;
      RECT 40.825 2.171 40.911 2.34 ;
      RECT 40.796 2.163 40.825 2.34 ;
      RECT 40.71 2.155 40.796 2.34 ;
      RECT 40.43 2.152 40.44 2.35 ;
      RECT 41.935 3.115 41.94 3.465 ;
      RECT 41.705 3.205 41.845 3.465 ;
      RECT 42.18 2.89 42.225 3.1 ;
      RECT 42.235 2.901 42.245 3.095 ;
      RECT 42.225 2.893 42.235 3.1 ;
      RECT 42.16 2.89 42.18 3.105 ;
      RECT 42.13 2.89 42.16 3.128 ;
      RECT 42.12 2.89 42.13 3.153 ;
      RECT 42.115 2.89 42.12 3.163 ;
      RECT 42.06 2.89 42.115 3.203 ;
      RECT 42.055 2.89 42.06 3.243 ;
      RECT 42.05 2.892 42.055 3.248 ;
      RECT 42.035 2.902 42.05 3.259 ;
      RECT 41.99 2.96 42.035 3.295 ;
      RECT 41.98 3.015 41.99 3.329 ;
      RECT 41.965 3.042 41.98 3.345 ;
      RECT 41.955 3.069 41.965 3.465 ;
      RECT 41.94 3.092 41.955 3.465 ;
      RECT 41.93 3.132 41.935 3.465 ;
      RECT 41.925 3.142 41.93 3.465 ;
      RECT 41.92 3.157 41.925 3.465 ;
      RECT 41.91 3.162 41.92 3.465 ;
      RECT 41.845 3.185 41.91 3.465 ;
      RECT 41.345 2.68 41.535 2.89 ;
      RECT 39.92 2.605 40.18 2.865 ;
      RECT 40.27 2.6 40.365 2.81 ;
      RECT 40.245 2.615 40.255 2.81 ;
      RECT 41.535 2.687 41.545 2.885 ;
      RECT 41.335 2.687 41.345 2.885 ;
      RECT 41.32 2.702 41.335 2.875 ;
      RECT 41.315 2.71 41.32 2.868 ;
      RECT 41.305 2.713 41.315 2.865 ;
      RECT 41.27 2.712 41.305 2.863 ;
      RECT 41.241 2.708 41.27 2.86 ;
      RECT 41.155 2.703 41.241 2.857 ;
      RECT 41.095 2.697 41.155 2.853 ;
      RECT 41.066 2.693 41.095 2.85 ;
      RECT 40.98 2.685 41.066 2.847 ;
      RECT 40.971 2.679 40.98 2.845 ;
      RECT 40.885 2.674 40.971 2.843 ;
      RECT 40.862 2.669 40.885 2.84 ;
      RECT 40.776 2.663 40.862 2.837 ;
      RECT 40.69 2.654 40.776 2.832 ;
      RECT 40.68 2.649 40.69 2.83 ;
      RECT 40.661 2.648 40.68 2.829 ;
      RECT 40.575 2.643 40.661 2.825 ;
      RECT 40.555 2.638 40.575 2.821 ;
      RECT 40.495 2.633 40.555 2.818 ;
      RECT 40.47 2.623 40.495 2.816 ;
      RECT 40.465 2.616 40.47 2.815 ;
      RECT 40.455 2.607 40.465 2.814 ;
      RECT 40.451 2.6 40.455 2.814 ;
      RECT 40.365 2.6 40.451 2.812 ;
      RECT 40.255 2.607 40.27 2.81 ;
      RECT 40.24 2.617 40.245 2.81 ;
      RECT 40.22 2.62 40.24 2.807 ;
      RECT 40.19 2.62 40.22 2.803 ;
      RECT 40.18 2.62 40.19 2.803 ;
      RECT 41.095 3.115 41.355 3.375 ;
      RECT 41.025 3.125 41.355 3.335 ;
      RECT 41.015 3.132 41.355 3.33 ;
      RECT 40.435 3.12 40.695 3.38 ;
      RECT 40.435 3.16 40.8 3.37 ;
      RECT 40.435 3.162 40.805 3.369 ;
      RECT 40.435 3.17 40.81 3.366 ;
      RECT 39.36 2.245 39.46 3.77 ;
      RECT 39.55 3.385 39.6 3.645 ;
      RECT 39.545 2.258 39.55 2.445 ;
      RECT 39.54 3.366 39.55 3.645 ;
      RECT 39.54 2.255 39.545 2.453 ;
      RECT 39.525 2.249 39.54 2.46 ;
      RECT 39.535 3.354 39.54 3.728 ;
      RECT 39.525 3.342 39.535 3.765 ;
      RECT 39.515 2.245 39.525 2.467 ;
      RECT 39.515 3.327 39.525 3.77 ;
      RECT 39.51 2.245 39.515 2.475 ;
      RECT 39.49 3.297 39.515 3.77 ;
      RECT 39.47 2.245 39.51 2.523 ;
      RECT 39.48 3.257 39.49 3.77 ;
      RECT 39.47 3.212 39.48 3.77 ;
      RECT 39.465 2.245 39.47 2.593 ;
      RECT 39.465 3.17 39.47 3.77 ;
      RECT 39.46 2.245 39.465 3.07 ;
      RECT 39.46 3.152 39.465 3.77 ;
      RECT 39.35 2.248 39.36 3.77 ;
      RECT 39.335 2.255 39.35 3.766 ;
      RECT 39.33 2.265 39.335 3.761 ;
      RECT 39.325 2.465 39.33 3.653 ;
      RECT 39.32 2.55 39.325 3.205 ;
      RECT 38.2 7.765 38.49 7.995 ;
      RECT 38.26 6.285 38.43 7.995 ;
      RECT 38.245 6.66 38.6 7.015 ;
      RECT 38.2 6.285 38.49 6.515 ;
      RECT 38.2 2.365 38.49 2.595 ;
      RECT 38.26 0.885 38.43 2.595 ;
      RECT 38.2 0.885 38.49 1.115 ;
      RECT 37.79 2.735 38.12 2.965 ;
      RECT 37.79 2.765 38.29 2.935 ;
      RECT 37.79 2.395 37.98 2.965 ;
      RECT 37.21 2.365 37.5 2.595 ;
      RECT 37.21 2.395 37.98 2.565 ;
      RECT 37.27 0.885 37.44 2.595 ;
      RECT 37.21 0.885 37.5 1.115 ;
      RECT 37.21 7.765 37.5 7.995 ;
      RECT 37.27 6.285 37.44 7.995 ;
      RECT 37.21 6.285 37.5 6.515 ;
      RECT 37.21 6.325 38.06 6.485 ;
      RECT 37.89 5.915 38.06 6.485 ;
      RECT 37.21 6.32 37.6 6.485 ;
      RECT 37.83 5.915 38.12 6.145 ;
      RECT 37.83 5.945 38.29 6.115 ;
      RECT 36.84 2.735 37.13 2.965 ;
      RECT 36.84 2.765 37.3 2.935 ;
      RECT 36.9 1.655 37.065 2.965 ;
      RECT 35.415 1.625 35.705 1.855 ;
      RECT 35.415 1.655 37.065 1.825 ;
      RECT 35.475 0.885 35.645 1.855 ;
      RECT 35.415 0.885 35.705 1.115 ;
      RECT 35.415 7.765 35.705 7.995 ;
      RECT 35.475 7.025 35.645 7.995 ;
      RECT 35.475 7.12 37.065 7.29 ;
      RECT 36.895 5.915 37.065 7.29 ;
      RECT 35.415 7.025 35.705 7.255 ;
      RECT 36.84 5.915 37.13 6.145 ;
      RECT 36.84 5.945 37.3 6.115 ;
      RECT 33.45 3.43 33.8 3.78 ;
      RECT 33.54 2.025 33.71 3.78 ;
      RECT 35.845 1.965 36.195 2.315 ;
      RECT 33.54 2.025 35.16 2.2 ;
      RECT 33.54 2.025 36.195 2.195 ;
      RECT 35.87 6.655 36.195 6.98 ;
      RECT 31.295 6.61 31.645 6.96 ;
      RECT 35.845 6.655 36.195 6.885 ;
      RECT 31.085 6.655 31.645 6.885 ;
      RECT 30.915 6.685 36.195 6.855 ;
      RECT 35.07 2.365 35.39 2.685 ;
      RECT 35.04 2.365 35.39 2.595 ;
      RECT 34.87 2.395 35.39 2.565 ;
      RECT 35.07 6.225 35.39 6.545 ;
      RECT 35.04 6.285 35.39 6.515 ;
      RECT 34.87 6.315 35.39 6.485 ;
      RECT 34.025 2.705 34.375 3.055 ;
      RECT 34.025 2.765 34.505 2.935 ;
      RECT 34.015 5.84 34.365 6.19 ;
      RECT 29.285 5.915 29.575 6.145 ;
      RECT 29.285 5.945 34.505 6.115 ;
      RECT 30.85 3.665 30.89 3.925 ;
      RECT 30.89 3.645 30.895 3.655 ;
      RECT 32.22 2.89 32.23 3.111 ;
      RECT 32.15 2.885 32.22 3.236 ;
      RECT 32.14 2.885 32.15 3.363 ;
      RECT 32.115 2.885 32.14 3.41 ;
      RECT 32.09 2.885 32.115 3.488 ;
      RECT 32.07 2.885 32.09 3.558 ;
      RECT 32.045 2.885 32.07 3.598 ;
      RECT 32.035 2.885 32.045 3.618 ;
      RECT 32.025 2.887 32.035 3.626 ;
      RECT 32.02 2.892 32.025 3.083 ;
      RECT 32.02 3.092 32.025 3.627 ;
      RECT 32.015 3.137 32.02 3.628 ;
      RECT 32.005 3.202 32.015 3.629 ;
      RECT 31.995 3.297 32.005 3.631 ;
      RECT 31.99 3.35 31.995 3.633 ;
      RECT 31.985 3.37 31.99 3.634 ;
      RECT 31.93 3.395 31.985 3.64 ;
      RECT 31.89 3.43 31.93 3.649 ;
      RECT 31.88 3.447 31.89 3.654 ;
      RECT 31.871 3.453 31.88 3.656 ;
      RECT 31.785 3.491 31.871 3.667 ;
      RECT 31.78 3.53 31.785 3.677 ;
      RECT 31.705 3.537 31.78 3.687 ;
      RECT 31.685 3.547 31.705 3.698 ;
      RECT 31.655 3.554 31.685 3.706 ;
      RECT 31.63 3.561 31.655 3.713 ;
      RECT 31.606 3.567 31.63 3.718 ;
      RECT 31.52 3.58 31.606 3.73 ;
      RECT 31.442 3.587 31.52 3.748 ;
      RECT 31.356 3.582 31.442 3.766 ;
      RECT 31.27 3.577 31.356 3.786 ;
      RECT 31.19 3.571 31.27 3.803 ;
      RECT 31.125 3.567 31.19 3.832 ;
      RECT 31.12 3.281 31.125 3.305 ;
      RECT 31.11 3.557 31.125 3.86 ;
      RECT 31.115 3.275 31.12 3.345 ;
      RECT 31.11 3.269 31.115 3.415 ;
      RECT 31.105 3.263 31.11 3.493 ;
      RECT 31.105 3.54 31.11 3.925 ;
      RECT 31.097 3.26 31.105 3.925 ;
      RECT 31.011 3.258 31.097 3.925 ;
      RECT 30.925 3.256 31.011 3.925 ;
      RECT 30.915 3.257 30.925 3.925 ;
      RECT 30.91 3.262 30.915 3.925 ;
      RECT 30.9 3.275 30.91 3.925 ;
      RECT 30.895 3.297 30.9 3.925 ;
      RECT 30.89 3.657 30.895 3.925 ;
      RECT 31.52 3.125 31.525 3.345 ;
      RECT 32.025 2.16 32.06 2.42 ;
      RECT 32.01 2.16 32.025 2.428 ;
      RECT 31.981 2.16 32.01 2.45 ;
      RECT 31.895 2.16 31.981 2.51 ;
      RECT 31.875 2.16 31.895 2.575 ;
      RECT 31.815 2.16 31.875 2.74 ;
      RECT 31.81 2.16 31.815 2.888 ;
      RECT 31.805 2.16 31.81 2.9 ;
      RECT 31.8 2.16 31.805 2.926 ;
      RECT 31.77 2.346 31.8 3.006 ;
      RECT 31.765 2.394 31.77 3.095 ;
      RECT 31.76 2.408 31.765 3.11 ;
      RECT 31.755 2.427 31.76 3.14 ;
      RECT 31.75 2.442 31.755 3.156 ;
      RECT 31.745 2.457 31.75 3.178 ;
      RECT 31.74 2.477 31.745 3.2 ;
      RECT 31.73 2.497 31.74 3.233 ;
      RECT 31.715 2.539 31.73 3.295 ;
      RECT 31.71 2.57 31.715 3.335 ;
      RECT 31.705 2.582 31.71 3.34 ;
      RECT 31.7 2.594 31.705 3.345 ;
      RECT 31.695 2.607 31.7 3.345 ;
      RECT 31.69 2.625 31.695 3.345 ;
      RECT 31.685 2.645 31.69 3.345 ;
      RECT 31.68 2.657 31.685 3.345 ;
      RECT 31.675 2.67 31.68 3.345 ;
      RECT 31.655 2.705 31.675 3.345 ;
      RECT 31.605 2.807 31.655 3.345 ;
      RECT 31.6 2.892 31.605 3.345 ;
      RECT 31.595 2.9 31.6 3.345 ;
      RECT 31.59 2.917 31.595 3.345 ;
      RECT 31.585 2.932 31.59 3.345 ;
      RECT 31.55 2.997 31.585 3.345 ;
      RECT 31.535 3.062 31.55 3.345 ;
      RECT 31.53 3.092 31.535 3.345 ;
      RECT 31.525 3.117 31.53 3.345 ;
      RECT 31.51 3.127 31.52 3.345 ;
      RECT 31.495 3.14 31.51 3.338 ;
      RECT 31.24 2.73 31.31 2.94 ;
      RECT 31.03 2.707 31.035 2.9 ;
      RECT 28.485 2.635 28.745 2.895 ;
      RECT 31.32 2.917 31.325 2.92 ;
      RECT 31.31 2.735 31.32 2.935 ;
      RECT 31.211 2.728 31.24 2.94 ;
      RECT 31.125 2.72 31.211 2.94 ;
      RECT 31.11 2.714 31.125 2.938 ;
      RECT 31.09 2.713 31.11 2.925 ;
      RECT 31.085 2.712 31.09 2.908 ;
      RECT 31.035 2.709 31.085 2.903 ;
      RECT 31.005 2.706 31.03 2.898 ;
      RECT 30.985 2.704 31.005 2.893 ;
      RECT 30.97 2.702 30.985 2.89 ;
      RECT 30.94 2.7 30.97 2.888 ;
      RECT 30.875 2.696 30.94 2.88 ;
      RECT 30.845 2.691 30.875 2.875 ;
      RECT 30.825 2.689 30.845 2.873 ;
      RECT 30.795 2.686 30.825 2.868 ;
      RECT 30.735 2.682 30.795 2.86 ;
      RECT 30.73 2.679 30.735 2.855 ;
      RECT 30.66 2.677 30.73 2.85 ;
      RECT 30.631 2.673 30.66 2.843 ;
      RECT 30.545 2.668 30.631 2.835 ;
      RECT 30.511 2.663 30.545 2.827 ;
      RECT 30.425 2.655 30.511 2.819 ;
      RECT 30.386 2.648 30.425 2.811 ;
      RECT 30.3 2.643 30.386 2.803 ;
      RECT 30.235 2.637 30.3 2.793 ;
      RECT 30.215 2.632 30.235 2.788 ;
      RECT 30.206 2.629 30.215 2.787 ;
      RECT 30.12 2.625 30.206 2.781 ;
      RECT 30.08 2.621 30.12 2.773 ;
      RECT 30.06 2.617 30.08 2.771 ;
      RECT 30 2.617 30.06 2.768 ;
      RECT 29.98 2.62 30 2.766 ;
      RECT 29.959 2.62 29.98 2.766 ;
      RECT 29.873 2.622 29.959 2.77 ;
      RECT 29.787 2.624 29.873 2.776 ;
      RECT 29.701 2.626 29.787 2.783 ;
      RECT 29.615 2.629 29.701 2.789 ;
      RECT 29.581 2.63 29.615 2.794 ;
      RECT 29.495 2.633 29.581 2.799 ;
      RECT 29.466 2.64 29.495 2.804 ;
      RECT 29.38 2.64 29.466 2.809 ;
      RECT 29.347 2.64 29.38 2.814 ;
      RECT 29.261 2.642 29.347 2.819 ;
      RECT 29.175 2.644 29.261 2.826 ;
      RECT 29.111 2.646 29.175 2.832 ;
      RECT 29.025 2.648 29.111 2.838 ;
      RECT 29.022 2.65 29.025 2.841 ;
      RECT 28.936 2.651 29.022 2.845 ;
      RECT 28.85 2.654 28.936 2.852 ;
      RECT 28.831 2.656 28.85 2.856 ;
      RECT 28.745 2.658 28.831 2.861 ;
      RECT 28.475 2.67 28.485 2.865 ;
      RECT 30.655 7.765 30.945 7.995 ;
      RECT 30.715 7.025 30.885 7.995 ;
      RECT 30.605 7.055 30.98 7.425 ;
      RECT 30.655 7.025 30.945 7.425 ;
      RECT 30.71 2.25 30.895 2.46 ;
      RECT 30.705 2.251 30.9 2.458 ;
      RECT 30.7 2.256 30.91 2.453 ;
      RECT 30.695 2.232 30.7 2.45 ;
      RECT 30.665 2.229 30.695 2.443 ;
      RECT 30.66 2.225 30.665 2.434 ;
      RECT 30.625 2.256 30.91 2.429 ;
      RECT 30.4 2.165 30.66 2.425 ;
      RECT 30.7 2.234 30.705 2.453 ;
      RECT 30.705 2.235 30.71 2.458 ;
      RECT 30.4 2.247 30.78 2.425 ;
      RECT 30.4 2.245 30.765 2.425 ;
      RECT 30.4 2.24 30.755 2.425 ;
      RECT 30.355 3.155 30.405 3.44 ;
      RECT 30.3 3.125 30.305 3.44 ;
      RECT 30.27 3.105 30.275 3.44 ;
      RECT 30.42 3.155 30.48 3.415 ;
      RECT 30.415 3.155 30.42 3.423 ;
      RECT 30.405 3.155 30.415 3.435 ;
      RECT 30.32 3.145 30.355 3.44 ;
      RECT 30.315 3.132 30.32 3.44 ;
      RECT 30.305 3.127 30.315 3.44 ;
      RECT 30.285 3.117 30.3 3.44 ;
      RECT 30.275 3.11 30.285 3.44 ;
      RECT 30.265 3.102 30.27 3.44 ;
      RECT 30.235 3.092 30.265 3.44 ;
      RECT 30.22 3.08 30.235 3.44 ;
      RECT 30.205 3.07 30.22 3.435 ;
      RECT 30.185 3.06 30.205 3.41 ;
      RECT 30.175 3.052 30.185 3.387 ;
      RECT 30.145 3.035 30.175 3.377 ;
      RECT 30.14 3.012 30.145 3.368 ;
      RECT 30.135 2.999 30.14 3.366 ;
      RECT 30.12 2.975 30.135 3.36 ;
      RECT 30.115 2.951 30.12 3.354 ;
      RECT 30.105 2.94 30.115 3.349 ;
      RECT 30.1 2.93 30.105 3.345 ;
      RECT 30.095 2.922 30.1 3.342 ;
      RECT 30.085 2.917 30.095 3.338 ;
      RECT 30.08 2.912 30.085 3.334 ;
      RECT 29.995 2.91 30.08 3.309 ;
      RECT 29.965 2.91 29.995 3.275 ;
      RECT 29.95 2.91 29.965 3.258 ;
      RECT 29.895 2.91 29.95 3.203 ;
      RECT 29.89 2.915 29.895 3.152 ;
      RECT 29.88 2.92 29.89 3.142 ;
      RECT 29.875 2.93 29.88 3.128 ;
      RECT 29.825 3.67 30.085 3.93 ;
      RECT 29.745 3.685 30.085 3.906 ;
      RECT 29.725 3.685 30.085 3.901 ;
      RECT 29.701 3.685 30.085 3.899 ;
      RECT 29.615 3.685 30.085 3.894 ;
      RECT 29.465 3.625 29.725 3.89 ;
      RECT 29.42 3.685 30.085 3.885 ;
      RECT 29.415 3.692 30.085 3.88 ;
      RECT 29.43 3.68 29.745 3.89 ;
      RECT 29.32 2.115 29.58 2.375 ;
      RECT 29.32 2.172 29.585 2.368 ;
      RECT 29.32 2.202 29.59 2.3 ;
      RECT 29.38 2.633 29.495 2.635 ;
      RECT 29.466 2.63 29.495 2.635 ;
      RECT 28.49 3.634 28.515 3.874 ;
      RECT 28.475 3.637 28.565 3.868 ;
      RECT 28.47 3.642 28.651 3.863 ;
      RECT 28.465 3.65 28.715 3.861 ;
      RECT 28.465 3.65 28.725 3.86 ;
      RECT 28.46 3.657 28.735 3.853 ;
      RECT 28.46 3.657 28.821 3.842 ;
      RECT 28.455 3.692 28.821 3.838 ;
      RECT 28.455 3.692 28.83 3.827 ;
      RECT 28.735 3.565 28.995 3.825 ;
      RECT 28.445 3.742 28.995 3.823 ;
      RECT 28.715 3.61 28.735 3.858 ;
      RECT 28.651 3.613 28.715 3.862 ;
      RECT 28.565 3.618 28.651 3.867 ;
      RECT 28.495 3.629 28.995 3.825 ;
      RECT 28.515 3.623 28.565 3.872 ;
      RECT 28.64 2.1 28.65 2.362 ;
      RECT 28.63 2.157 28.64 2.365 ;
      RECT 28.605 2.162 28.63 2.371 ;
      RECT 28.58 2.166 28.605 2.383 ;
      RECT 28.57 2.169 28.58 2.393 ;
      RECT 28.565 2.17 28.57 2.398 ;
      RECT 28.56 2.171 28.565 2.403 ;
      RECT 28.555 2.172 28.56 2.405 ;
      RECT 28.53 2.175 28.555 2.408 ;
      RECT 28.5 2.181 28.53 2.411 ;
      RECT 28.435 2.192 28.5 2.414 ;
      RECT 28.39 2.2 28.435 2.418 ;
      RECT 28.375 2.2 28.39 2.426 ;
      RECT 28.37 2.201 28.375 2.433 ;
      RECT 28.365 2.203 28.37 2.436 ;
      RECT 28.36 2.207 28.365 2.439 ;
      RECT 28.35 2.215 28.36 2.443 ;
      RECT 28.345 2.228 28.35 2.448 ;
      RECT 28.34 2.236 28.345 2.45 ;
      RECT 28.335 2.242 28.34 2.45 ;
      RECT 28.33 2.246 28.335 2.453 ;
      RECT 28.325 2.248 28.33 2.456 ;
      RECT 28.32 2.251 28.325 2.459 ;
      RECT 28.31 2.256 28.32 2.463 ;
      RECT 28.305 2.262 28.31 2.468 ;
      RECT 28.295 2.268 28.305 2.472 ;
      RECT 28.28 2.275 28.295 2.478 ;
      RECT 28.251 2.289 28.28 2.488 ;
      RECT 28.165 2.324 28.251 2.52 ;
      RECT 28.145 2.357 28.165 2.549 ;
      RECT 28.125 2.37 28.145 2.56 ;
      RECT 28.105 2.382 28.125 2.571 ;
      RECT 28.055 2.404 28.105 2.591 ;
      RECT 28.04 2.422 28.055 2.608 ;
      RECT 28.035 2.428 28.04 2.611 ;
      RECT 28.03 2.432 28.035 2.614 ;
      RECT 28.025 2.436 28.03 2.618 ;
      RECT 28.02 2.438 28.025 2.621 ;
      RECT 28.01 2.445 28.02 2.624 ;
      RECT 28.005 2.45 28.01 2.628 ;
      RECT 28 2.452 28.005 2.631 ;
      RECT 27.995 2.456 28 2.634 ;
      RECT 27.99 2.458 27.995 2.638 ;
      RECT 27.975 2.463 27.99 2.643 ;
      RECT 27.97 2.468 27.975 2.646 ;
      RECT 27.965 2.476 27.97 2.649 ;
      RECT 27.96 2.478 27.965 2.652 ;
      RECT 27.955 2.48 27.96 2.655 ;
      RECT 27.945 2.482 27.955 2.661 ;
      RECT 27.91 2.496 27.945 2.673 ;
      RECT 27.9 2.511 27.91 2.683 ;
      RECT 27.825 2.54 27.9 2.707 ;
      RECT 27.82 2.565 27.825 2.73 ;
      RECT 27.805 2.569 27.82 2.736 ;
      RECT 27.795 2.577 27.805 2.741 ;
      RECT 27.765 2.59 27.795 2.745 ;
      RECT 27.755 2.605 27.765 2.75 ;
      RECT 27.745 2.61 27.755 2.753 ;
      RECT 27.74 2.612 27.745 2.755 ;
      RECT 27.725 2.615 27.74 2.758 ;
      RECT 27.72 2.617 27.725 2.761 ;
      RECT 27.7 2.622 27.72 2.765 ;
      RECT 27.67 2.627 27.7 2.773 ;
      RECT 27.645 2.634 27.67 2.781 ;
      RECT 27.64 2.639 27.645 2.786 ;
      RECT 27.61 2.642 27.64 2.79 ;
      RECT 27.57 2.645 27.61 2.8 ;
      RECT 27.535 2.642 27.57 2.812 ;
      RECT 27.525 2.638 27.535 2.819 ;
      RECT 27.5 2.634 27.525 2.825 ;
      RECT 27.495 2.63 27.5 2.83 ;
      RECT 27.455 2.627 27.495 2.83 ;
      RECT 27.44 2.612 27.455 2.831 ;
      RECT 27.417 2.6 27.44 2.831 ;
      RECT 27.331 2.6 27.417 2.832 ;
      RECT 27.245 2.6 27.331 2.834 ;
      RECT 27.225 2.6 27.245 2.831 ;
      RECT 27.22 2.605 27.225 2.826 ;
      RECT 27.215 2.61 27.22 2.824 ;
      RECT 27.205 2.62 27.215 2.822 ;
      RECT 27.2 2.626 27.205 2.815 ;
      RECT 27.195 2.628 27.2 2.8 ;
      RECT 27.19 2.632 27.195 2.79 ;
      RECT 28.65 2.1 28.9 2.36 ;
      RECT 26.375 3.635 26.635 3.895 ;
      RECT 28.67 3.125 28.675 3.335 ;
      RECT 28.675 3.13 28.685 3.33 ;
      RECT 28.625 3.125 28.67 3.35 ;
      RECT 28.615 3.125 28.625 3.37 ;
      RECT 28.596 3.125 28.615 3.375 ;
      RECT 28.51 3.125 28.596 3.372 ;
      RECT 28.48 3.127 28.51 3.37 ;
      RECT 28.425 3.137 28.48 3.368 ;
      RECT 28.36 3.151 28.425 3.366 ;
      RECT 28.355 3.159 28.36 3.365 ;
      RECT 28.34 3.162 28.355 3.363 ;
      RECT 28.275 3.172 28.34 3.359 ;
      RECT 28.227 3.186 28.275 3.36 ;
      RECT 28.141 3.203 28.227 3.374 ;
      RECT 28.055 3.224 28.141 3.391 ;
      RECT 28.035 3.237 28.055 3.401 ;
      RECT 27.99 3.245 28.035 3.408 ;
      RECT 27.955 3.253 27.99 3.416 ;
      RECT 27.921 3.261 27.955 3.424 ;
      RECT 27.835 3.275 27.921 3.436 ;
      RECT 27.8 3.292 27.835 3.448 ;
      RECT 27.791 3.301 27.8 3.452 ;
      RECT 27.705 3.319 27.791 3.469 ;
      RECT 27.646 3.346 27.705 3.496 ;
      RECT 27.56 3.373 27.646 3.524 ;
      RECT 27.54 3.395 27.56 3.544 ;
      RECT 27.48 3.41 27.54 3.56 ;
      RECT 27.47 3.422 27.48 3.573 ;
      RECT 27.465 3.427 27.47 3.576 ;
      RECT 27.455 3.43 27.465 3.579 ;
      RECT 27.45 3.432 27.455 3.582 ;
      RECT 27.42 3.44 27.45 3.589 ;
      RECT 27.405 3.447 27.42 3.597 ;
      RECT 27.395 3.452 27.405 3.601 ;
      RECT 27.39 3.455 27.395 3.604 ;
      RECT 27.38 3.457 27.39 3.607 ;
      RECT 27.345 3.467 27.38 3.616 ;
      RECT 27.27 3.49 27.345 3.638 ;
      RECT 27.25 3.508 27.27 3.656 ;
      RECT 27.22 3.515 27.25 3.666 ;
      RECT 27.2 3.523 27.22 3.676 ;
      RECT 27.19 3.529 27.2 3.683 ;
      RECT 27.171 3.534 27.19 3.689 ;
      RECT 27.085 3.554 27.171 3.709 ;
      RECT 27.07 3.574 27.085 3.728 ;
      RECT 27.025 3.586 27.07 3.739 ;
      RECT 26.96 3.607 27.025 3.762 ;
      RECT 26.92 3.627 26.96 3.783 ;
      RECT 26.91 3.637 26.92 3.793 ;
      RECT 26.86 3.649 26.91 3.804 ;
      RECT 26.84 3.665 26.86 3.816 ;
      RECT 26.81 3.675 26.84 3.822 ;
      RECT 26.8 3.68 26.81 3.824 ;
      RECT 26.731 3.681 26.8 3.83 ;
      RECT 26.645 3.683 26.731 3.84 ;
      RECT 26.635 3.684 26.645 3.845 ;
      RECT 27.905 3.71 28.095 3.92 ;
      RECT 27.895 3.715 28.105 3.913 ;
      RECT 27.88 3.715 28.105 3.878 ;
      RECT 27.8 3.6 28.06 3.86 ;
      RECT 26.715 3.13 26.9 3.425 ;
      RECT 26.705 3.13 26.9 3.423 ;
      RECT 26.69 3.13 26.905 3.418 ;
      RECT 26.69 3.13 26.91 3.415 ;
      RECT 26.685 3.13 26.91 3.413 ;
      RECT 26.68 3.385 26.91 3.403 ;
      RECT 26.685 3.13 26.945 3.39 ;
      RECT 26.645 2.165 26.905 2.425 ;
      RECT 26.455 2.09 26.541 2.423 ;
      RECT 26.43 2.094 26.585 2.419 ;
      RECT 26.541 2.086 26.585 2.419 ;
      RECT 26.541 2.087 26.59 2.418 ;
      RECT 26.455 2.092 26.605 2.417 ;
      RECT 26.43 2.1 26.645 2.416 ;
      RECT 26.425 2.095 26.605 2.411 ;
      RECT 26.415 2.11 26.645 2.318 ;
      RECT 26.415 2.162 26.845 2.318 ;
      RECT 26.415 2.155 26.825 2.318 ;
      RECT 26.415 2.142 26.795 2.318 ;
      RECT 26.415 2.13 26.735 2.318 ;
      RECT 26.415 2.115 26.71 2.318 ;
      RECT 25.615 2.745 25.75 3.04 ;
      RECT 25.875 2.768 25.88 2.955 ;
      RECT 26.595 2.665 26.74 2.9 ;
      RECT 26.755 2.665 26.76 2.89 ;
      RECT 26.79 2.676 26.795 2.87 ;
      RECT 26.785 2.668 26.79 2.875 ;
      RECT 26.765 2.665 26.785 2.88 ;
      RECT 26.76 2.665 26.765 2.888 ;
      RECT 26.75 2.665 26.755 2.893 ;
      RECT 26.74 2.665 26.75 2.898 ;
      RECT 26.57 2.667 26.595 2.9 ;
      RECT 26.52 2.674 26.57 2.9 ;
      RECT 26.515 2.679 26.52 2.9 ;
      RECT 26.476 2.684 26.515 2.901 ;
      RECT 26.39 2.696 26.476 2.902 ;
      RECT 26.381 2.706 26.39 2.902 ;
      RECT 26.295 2.715 26.381 2.904 ;
      RECT 26.271 2.725 26.295 2.906 ;
      RECT 26.185 2.736 26.271 2.907 ;
      RECT 26.155 2.747 26.185 2.909 ;
      RECT 26.125 2.752 26.155 2.911 ;
      RECT 26.1 2.758 26.125 2.914 ;
      RECT 26.085 2.763 26.1 2.915 ;
      RECT 26.04 2.769 26.085 2.915 ;
      RECT 26.035 2.774 26.04 2.916 ;
      RECT 26.015 2.774 26.035 2.918 ;
      RECT 25.995 2.772 26.015 2.923 ;
      RECT 25.96 2.771 25.995 2.93 ;
      RECT 25.93 2.77 25.96 2.94 ;
      RECT 25.88 2.769 25.93 2.95 ;
      RECT 25.79 2.766 25.875 3.04 ;
      RECT 25.765 2.76 25.79 3.04 ;
      RECT 25.75 2.75 25.765 3.04 ;
      RECT 25.565 2.745 25.615 2.96 ;
      RECT 25.555 2.75 25.565 2.95 ;
      RECT 25.795 3.225 26.055 3.485 ;
      RECT 25.795 3.225 26.085 3.378 ;
      RECT 25.795 3.225 26.12 3.363 ;
      RECT 26.05 3.145 26.24 3.355 ;
      RECT 26.04 3.15 26.25 3.348 ;
      RECT 26.005 3.22 26.25 3.348 ;
      RECT 26.035 3.162 26.055 3.485 ;
      RECT 26.02 3.21 26.25 3.348 ;
      RECT 26.025 3.182 26.055 3.485 ;
      RECT 25.105 2.25 25.175 3.355 ;
      RECT 25.84 2.355 26.1 2.615 ;
      RECT 25.42 2.401 25.435 2.61 ;
      RECT 25.756 2.414 25.84 2.565 ;
      RECT 25.67 2.411 25.756 2.565 ;
      RECT 25.631 2.409 25.67 2.565 ;
      RECT 25.545 2.407 25.631 2.565 ;
      RECT 25.485 2.405 25.545 2.576 ;
      RECT 25.45 2.403 25.485 2.594 ;
      RECT 25.435 2.401 25.45 2.605 ;
      RECT 25.405 2.401 25.42 2.618 ;
      RECT 25.395 2.401 25.405 2.623 ;
      RECT 25.37 2.4 25.395 2.628 ;
      RECT 25.355 2.395 25.37 2.634 ;
      RECT 25.35 2.388 25.355 2.639 ;
      RECT 25.325 2.379 25.35 2.645 ;
      RECT 25.28 2.358 25.325 2.658 ;
      RECT 25.27 2.342 25.28 2.668 ;
      RECT 25.255 2.335 25.27 2.678 ;
      RECT 25.245 2.328 25.255 2.695 ;
      RECT 25.24 2.325 25.245 2.725 ;
      RECT 25.235 2.323 25.24 2.755 ;
      RECT 25.23 2.321 25.235 2.792 ;
      RECT 25.215 2.317 25.23 2.859 ;
      RECT 25.215 3.15 25.225 3.35 ;
      RECT 25.21 2.313 25.215 2.985 ;
      RECT 25.21 3.137 25.215 3.355 ;
      RECT 25.205 2.311 25.21 3.07 ;
      RECT 25.205 3.127 25.21 3.355 ;
      RECT 25.19 2.282 25.205 3.355 ;
      RECT 25.175 2.255 25.19 3.355 ;
      RECT 25.1 2.25 25.105 2.605 ;
      RECT 25.1 2.66 25.105 3.355 ;
      RECT 25.085 2.25 25.1 2.583 ;
      RECT 25.095 2.682 25.1 3.355 ;
      RECT 25.085 2.722 25.095 3.355 ;
      RECT 25.05 2.25 25.085 2.525 ;
      RECT 25.08 2.757 25.085 3.355 ;
      RECT 25.065 2.812 25.08 3.355 ;
      RECT 25.06 2.877 25.065 3.355 ;
      RECT 25.045 2.925 25.06 3.355 ;
      RECT 25.02 2.25 25.05 2.48 ;
      RECT 25.04 2.98 25.045 3.355 ;
      RECT 25.025 3.04 25.04 3.355 ;
      RECT 25.02 3.088 25.025 3.353 ;
      RECT 25.015 2.25 25.02 2.473 ;
      RECT 25.015 3.12 25.02 3.348 ;
      RECT 24.99 2.25 25.015 2.465 ;
      RECT 24.98 2.255 24.99 2.455 ;
      RECT 25.195 3.53 25.215 3.77 ;
      RECT 24.425 3.46 24.43 3.67 ;
      RECT 25.705 3.533 25.715 3.728 ;
      RECT 25.7 3.523 25.705 3.731 ;
      RECT 25.62 3.52 25.7 3.754 ;
      RECT 25.616 3.52 25.62 3.776 ;
      RECT 25.53 3.52 25.616 3.786 ;
      RECT 25.515 3.52 25.53 3.794 ;
      RECT 25.486 3.521 25.515 3.792 ;
      RECT 25.4 3.526 25.486 3.788 ;
      RECT 25.387 3.53 25.4 3.784 ;
      RECT 25.301 3.53 25.387 3.78 ;
      RECT 25.215 3.53 25.301 3.774 ;
      RECT 25.131 3.53 25.195 3.768 ;
      RECT 25.045 3.53 25.131 3.763 ;
      RECT 25.025 3.53 25.045 3.759 ;
      RECT 24.965 3.525 25.025 3.756 ;
      RECT 24.937 3.519 24.965 3.753 ;
      RECT 24.851 3.514 24.937 3.749 ;
      RECT 24.765 3.508 24.851 3.743 ;
      RECT 24.69 3.49 24.765 3.738 ;
      RECT 24.655 3.467 24.69 3.734 ;
      RECT 24.645 3.457 24.655 3.733 ;
      RECT 24.59 3.455 24.645 3.732 ;
      RECT 24.515 3.455 24.59 3.728 ;
      RECT 24.505 3.455 24.515 3.723 ;
      RECT 24.49 3.455 24.505 3.715 ;
      RECT 24.44 3.457 24.49 3.693 ;
      RECT 24.43 3.46 24.44 3.673 ;
      RECT 24.42 3.465 24.425 3.668 ;
      RECT 24.415 3.47 24.42 3.663 ;
      RECT 24.54 2.635 24.8 2.895 ;
      RECT 24.54 2.65 24.82 2.86 ;
      RECT 24.54 2.655 24.83 2.855 ;
      RECT 22.525 2.115 22.785 2.375 ;
      RECT 22.515 2.145 22.785 2.355 ;
      RECT 24.435 2.06 24.695 2.32 ;
      RECT 24.43 2.135 24.435 2.321 ;
      RECT 24.405 2.14 24.43 2.323 ;
      RECT 24.39 2.147 24.405 2.326 ;
      RECT 24.33 2.165 24.39 2.331 ;
      RECT 24.3 2.185 24.33 2.338 ;
      RECT 24.275 2.193 24.3 2.343 ;
      RECT 24.25 2.201 24.275 2.345 ;
      RECT 24.232 2.205 24.25 2.344 ;
      RECT 24.146 2.203 24.232 2.344 ;
      RECT 24.06 2.201 24.146 2.344 ;
      RECT 23.974 2.199 24.06 2.343 ;
      RECT 23.888 2.197 23.974 2.343 ;
      RECT 23.802 2.195 23.888 2.343 ;
      RECT 23.716 2.193 23.802 2.343 ;
      RECT 23.63 2.191 23.716 2.342 ;
      RECT 23.612 2.19 23.63 2.342 ;
      RECT 23.526 2.189 23.612 2.342 ;
      RECT 23.44 2.187 23.526 2.342 ;
      RECT 23.354 2.186 23.44 2.341 ;
      RECT 23.268 2.185 23.354 2.341 ;
      RECT 23.182 2.183 23.268 2.341 ;
      RECT 23.096 2.182 23.182 2.341 ;
      RECT 23.01 2.18 23.096 2.34 ;
      RECT 22.986 2.178 23.01 2.34 ;
      RECT 22.9 2.171 22.986 2.34 ;
      RECT 22.871 2.163 22.9 2.34 ;
      RECT 22.785 2.155 22.871 2.34 ;
      RECT 22.505 2.152 22.515 2.35 ;
      RECT 24.01 3.115 24.015 3.465 ;
      RECT 23.78 3.205 23.92 3.465 ;
      RECT 24.255 2.89 24.3 3.1 ;
      RECT 24.31 2.901 24.32 3.095 ;
      RECT 24.3 2.893 24.31 3.1 ;
      RECT 24.235 2.89 24.255 3.105 ;
      RECT 24.205 2.89 24.235 3.128 ;
      RECT 24.195 2.89 24.205 3.153 ;
      RECT 24.19 2.89 24.195 3.163 ;
      RECT 24.135 2.89 24.19 3.203 ;
      RECT 24.13 2.89 24.135 3.243 ;
      RECT 24.125 2.892 24.13 3.248 ;
      RECT 24.11 2.902 24.125 3.259 ;
      RECT 24.065 2.96 24.11 3.295 ;
      RECT 24.055 3.015 24.065 3.329 ;
      RECT 24.04 3.042 24.055 3.345 ;
      RECT 24.03 3.069 24.04 3.465 ;
      RECT 24.015 3.092 24.03 3.465 ;
      RECT 24.005 3.132 24.01 3.465 ;
      RECT 24 3.142 24.005 3.465 ;
      RECT 23.995 3.157 24 3.465 ;
      RECT 23.985 3.162 23.995 3.465 ;
      RECT 23.92 3.185 23.985 3.465 ;
      RECT 23.42 2.68 23.61 2.89 ;
      RECT 21.995 2.605 22.255 2.865 ;
      RECT 22.345 2.6 22.44 2.81 ;
      RECT 22.32 2.615 22.33 2.81 ;
      RECT 23.61 2.687 23.62 2.885 ;
      RECT 23.41 2.687 23.42 2.885 ;
      RECT 23.395 2.702 23.41 2.875 ;
      RECT 23.39 2.71 23.395 2.868 ;
      RECT 23.38 2.713 23.39 2.865 ;
      RECT 23.345 2.712 23.38 2.863 ;
      RECT 23.316 2.708 23.345 2.86 ;
      RECT 23.23 2.703 23.316 2.857 ;
      RECT 23.17 2.697 23.23 2.853 ;
      RECT 23.141 2.693 23.17 2.85 ;
      RECT 23.055 2.685 23.141 2.847 ;
      RECT 23.046 2.679 23.055 2.845 ;
      RECT 22.96 2.674 23.046 2.843 ;
      RECT 22.937 2.669 22.96 2.84 ;
      RECT 22.851 2.663 22.937 2.837 ;
      RECT 22.765 2.654 22.851 2.832 ;
      RECT 22.755 2.649 22.765 2.83 ;
      RECT 22.736 2.648 22.755 2.829 ;
      RECT 22.65 2.643 22.736 2.825 ;
      RECT 22.63 2.638 22.65 2.821 ;
      RECT 22.57 2.633 22.63 2.818 ;
      RECT 22.545 2.623 22.57 2.816 ;
      RECT 22.54 2.616 22.545 2.815 ;
      RECT 22.53 2.607 22.54 2.814 ;
      RECT 22.526 2.6 22.53 2.814 ;
      RECT 22.44 2.6 22.526 2.812 ;
      RECT 22.33 2.607 22.345 2.81 ;
      RECT 22.315 2.617 22.32 2.81 ;
      RECT 22.295 2.62 22.315 2.807 ;
      RECT 22.265 2.62 22.295 2.803 ;
      RECT 22.255 2.62 22.265 2.803 ;
      RECT 23.17 3.115 23.43 3.375 ;
      RECT 23.1 3.125 23.43 3.335 ;
      RECT 23.09 3.132 23.43 3.33 ;
      RECT 22.51 3.12 22.77 3.38 ;
      RECT 22.51 3.16 22.875 3.37 ;
      RECT 22.51 3.162 22.88 3.369 ;
      RECT 22.51 3.17 22.885 3.366 ;
      RECT 21.435 2.245 21.535 3.77 ;
      RECT 21.625 3.385 21.675 3.645 ;
      RECT 21.62 2.258 21.625 2.445 ;
      RECT 21.615 3.366 21.625 3.645 ;
      RECT 21.615 2.255 21.62 2.453 ;
      RECT 21.6 2.249 21.615 2.46 ;
      RECT 21.61 3.354 21.615 3.728 ;
      RECT 21.6 3.342 21.61 3.765 ;
      RECT 21.59 2.245 21.6 2.467 ;
      RECT 21.59 3.327 21.6 3.77 ;
      RECT 21.585 2.245 21.59 2.475 ;
      RECT 21.565 3.297 21.59 3.77 ;
      RECT 21.545 2.245 21.585 2.523 ;
      RECT 21.555 3.257 21.565 3.77 ;
      RECT 21.545 3.212 21.555 3.77 ;
      RECT 21.54 2.245 21.545 2.593 ;
      RECT 21.54 3.17 21.545 3.77 ;
      RECT 21.535 2.245 21.54 3.07 ;
      RECT 21.535 3.152 21.54 3.77 ;
      RECT 21.425 2.248 21.435 3.77 ;
      RECT 21.41 2.255 21.425 3.766 ;
      RECT 21.405 2.265 21.41 3.761 ;
      RECT 21.4 2.465 21.405 3.653 ;
      RECT 21.395 2.55 21.4 3.205 ;
      RECT 20.275 7.765 20.565 7.995 ;
      RECT 20.335 6.285 20.505 7.995 ;
      RECT 20.325 6.655 20.675 7.005 ;
      RECT 20.275 6.285 20.565 6.515 ;
      RECT 20.275 2.365 20.565 2.595 ;
      RECT 20.335 0.885 20.505 2.595 ;
      RECT 20.275 0.885 20.565 1.115 ;
      RECT 19.865 2.735 20.195 2.965 ;
      RECT 19.865 2.765 20.365 2.935 ;
      RECT 19.865 2.395 20.055 2.965 ;
      RECT 19.285 2.365 19.575 2.595 ;
      RECT 19.285 2.395 20.055 2.565 ;
      RECT 19.345 0.885 19.515 2.595 ;
      RECT 19.285 0.885 19.575 1.115 ;
      RECT 19.285 7.765 19.575 7.995 ;
      RECT 19.345 6.285 19.515 7.995 ;
      RECT 19.285 6.285 19.575 6.515 ;
      RECT 19.285 6.325 20.135 6.485 ;
      RECT 19.965 5.915 20.135 6.485 ;
      RECT 19.285 6.32 19.675 6.485 ;
      RECT 19.905 5.915 20.195 6.145 ;
      RECT 19.905 5.945 20.365 6.115 ;
      RECT 18.915 2.735 19.205 2.965 ;
      RECT 18.915 2.765 19.375 2.935 ;
      RECT 18.975 1.655 19.14 2.965 ;
      RECT 17.49 1.625 17.78 1.855 ;
      RECT 17.49 1.655 19.14 1.825 ;
      RECT 17.55 0.885 17.72 1.855 ;
      RECT 17.49 0.885 17.78 1.115 ;
      RECT 17.49 7.765 17.78 7.995 ;
      RECT 17.55 7.025 17.72 7.995 ;
      RECT 17.55 7.12 19.14 7.29 ;
      RECT 18.97 5.915 19.14 7.29 ;
      RECT 17.49 7.025 17.78 7.255 ;
      RECT 18.915 5.915 19.205 6.145 ;
      RECT 18.915 5.945 19.375 6.115 ;
      RECT 15.525 3.43 15.875 3.78 ;
      RECT 15.615 2.025 15.785 3.78 ;
      RECT 17.92 1.965 18.27 2.315 ;
      RECT 15.615 2.025 17.235 2.2 ;
      RECT 15.615 2.025 18.27 2.195 ;
      RECT 17.945 6.655 18.27 6.98 ;
      RECT 13.34 6.605 13.69 6.955 ;
      RECT 17.92 6.655 18.27 6.885 ;
      RECT 13.16 6.655 13.69 6.885 ;
      RECT 12.99 6.685 18.27 6.855 ;
      RECT 17.145 2.365 17.465 2.685 ;
      RECT 17.115 2.365 17.465 2.595 ;
      RECT 16.945 2.395 17.465 2.565 ;
      RECT 17.145 6.225 17.465 6.545 ;
      RECT 17.115 6.285 17.465 6.515 ;
      RECT 16.945 6.315 17.465 6.485 ;
      RECT 16.1 2.705 16.45 3.055 ;
      RECT 16.1 2.765 16.58 2.935 ;
      RECT 16.09 5.84 16.44 6.19 ;
      RECT 11.36 5.915 11.65 6.145 ;
      RECT 11.36 5.945 16.58 6.115 ;
      RECT 12.925 3.665 12.965 3.925 ;
      RECT 12.965 3.645 12.97 3.655 ;
      RECT 14.295 2.89 14.305 3.111 ;
      RECT 14.225 2.885 14.295 3.236 ;
      RECT 14.215 2.885 14.225 3.363 ;
      RECT 14.19 2.885 14.215 3.41 ;
      RECT 14.165 2.885 14.19 3.488 ;
      RECT 14.145 2.885 14.165 3.558 ;
      RECT 14.12 2.885 14.145 3.598 ;
      RECT 14.11 2.885 14.12 3.618 ;
      RECT 14.1 2.887 14.11 3.626 ;
      RECT 14.095 2.892 14.1 3.083 ;
      RECT 14.095 3.092 14.1 3.627 ;
      RECT 14.09 3.137 14.095 3.628 ;
      RECT 14.08 3.202 14.09 3.629 ;
      RECT 14.07 3.297 14.08 3.631 ;
      RECT 14.065 3.35 14.07 3.633 ;
      RECT 14.06 3.37 14.065 3.634 ;
      RECT 14.005 3.395 14.06 3.64 ;
      RECT 13.965 3.43 14.005 3.649 ;
      RECT 13.955 3.447 13.965 3.654 ;
      RECT 13.946 3.453 13.955 3.656 ;
      RECT 13.86 3.491 13.946 3.667 ;
      RECT 13.855 3.53 13.86 3.677 ;
      RECT 13.78 3.537 13.855 3.687 ;
      RECT 13.76 3.547 13.78 3.698 ;
      RECT 13.73 3.554 13.76 3.706 ;
      RECT 13.705 3.561 13.73 3.713 ;
      RECT 13.681 3.567 13.705 3.718 ;
      RECT 13.595 3.58 13.681 3.73 ;
      RECT 13.517 3.587 13.595 3.748 ;
      RECT 13.431 3.582 13.517 3.766 ;
      RECT 13.345 3.577 13.431 3.786 ;
      RECT 13.265 3.571 13.345 3.803 ;
      RECT 13.2 3.567 13.265 3.832 ;
      RECT 13.195 3.281 13.2 3.305 ;
      RECT 13.185 3.557 13.2 3.86 ;
      RECT 13.19 3.275 13.195 3.345 ;
      RECT 13.185 3.269 13.19 3.415 ;
      RECT 13.18 3.263 13.185 3.493 ;
      RECT 13.18 3.54 13.185 3.925 ;
      RECT 13.172 3.26 13.18 3.925 ;
      RECT 13.086 3.258 13.172 3.925 ;
      RECT 13 3.256 13.086 3.925 ;
      RECT 12.99 3.257 13 3.925 ;
      RECT 12.985 3.262 12.99 3.925 ;
      RECT 12.975 3.275 12.985 3.925 ;
      RECT 12.97 3.297 12.975 3.925 ;
      RECT 12.965 3.657 12.97 3.925 ;
      RECT 13.595 3.125 13.6 3.345 ;
      RECT 14.1 2.16 14.135 2.42 ;
      RECT 14.085 2.16 14.1 2.428 ;
      RECT 14.056 2.16 14.085 2.45 ;
      RECT 13.97 2.16 14.056 2.51 ;
      RECT 13.95 2.16 13.97 2.575 ;
      RECT 13.89 2.16 13.95 2.74 ;
      RECT 13.885 2.16 13.89 2.888 ;
      RECT 13.88 2.16 13.885 2.9 ;
      RECT 13.875 2.16 13.88 2.926 ;
      RECT 13.845 2.346 13.875 3.006 ;
      RECT 13.84 2.394 13.845 3.095 ;
      RECT 13.835 2.408 13.84 3.11 ;
      RECT 13.83 2.427 13.835 3.14 ;
      RECT 13.825 2.442 13.83 3.156 ;
      RECT 13.82 2.457 13.825 3.178 ;
      RECT 13.815 2.477 13.82 3.2 ;
      RECT 13.805 2.497 13.815 3.233 ;
      RECT 13.79 2.539 13.805 3.295 ;
      RECT 13.785 2.57 13.79 3.335 ;
      RECT 13.78 2.582 13.785 3.34 ;
      RECT 13.775 2.594 13.78 3.345 ;
      RECT 13.77 2.607 13.775 3.345 ;
      RECT 13.765 2.625 13.77 3.345 ;
      RECT 13.76 2.645 13.765 3.345 ;
      RECT 13.755 2.657 13.76 3.345 ;
      RECT 13.75 2.67 13.755 3.345 ;
      RECT 13.73 2.705 13.75 3.345 ;
      RECT 13.68 2.807 13.73 3.345 ;
      RECT 13.675 2.892 13.68 3.345 ;
      RECT 13.67 2.9 13.675 3.345 ;
      RECT 13.665 2.917 13.67 3.345 ;
      RECT 13.66 2.932 13.665 3.345 ;
      RECT 13.625 2.997 13.66 3.345 ;
      RECT 13.61 3.062 13.625 3.345 ;
      RECT 13.605 3.092 13.61 3.345 ;
      RECT 13.6 3.117 13.605 3.345 ;
      RECT 13.585 3.127 13.595 3.345 ;
      RECT 13.57 3.14 13.585 3.338 ;
      RECT 13.315 2.73 13.385 2.94 ;
      RECT 13.105 2.707 13.11 2.9 ;
      RECT 10.56 2.635 10.82 2.895 ;
      RECT 13.395 2.917 13.4 2.92 ;
      RECT 13.385 2.735 13.395 2.935 ;
      RECT 13.286 2.728 13.315 2.94 ;
      RECT 13.2 2.72 13.286 2.94 ;
      RECT 13.185 2.714 13.2 2.938 ;
      RECT 13.165 2.713 13.185 2.925 ;
      RECT 13.16 2.712 13.165 2.908 ;
      RECT 13.11 2.709 13.16 2.903 ;
      RECT 13.08 2.706 13.105 2.898 ;
      RECT 13.06 2.704 13.08 2.893 ;
      RECT 13.045 2.702 13.06 2.89 ;
      RECT 13.015 2.7 13.045 2.888 ;
      RECT 12.95 2.696 13.015 2.88 ;
      RECT 12.92 2.691 12.95 2.875 ;
      RECT 12.9 2.689 12.92 2.873 ;
      RECT 12.87 2.686 12.9 2.868 ;
      RECT 12.81 2.682 12.87 2.86 ;
      RECT 12.805 2.679 12.81 2.855 ;
      RECT 12.735 2.677 12.805 2.85 ;
      RECT 12.706 2.673 12.735 2.843 ;
      RECT 12.62 2.668 12.706 2.835 ;
      RECT 12.586 2.663 12.62 2.827 ;
      RECT 12.5 2.655 12.586 2.819 ;
      RECT 12.461 2.648 12.5 2.811 ;
      RECT 12.375 2.643 12.461 2.803 ;
      RECT 12.31 2.637 12.375 2.793 ;
      RECT 12.29 2.632 12.31 2.788 ;
      RECT 12.281 2.629 12.29 2.787 ;
      RECT 12.195 2.625 12.281 2.781 ;
      RECT 12.155 2.621 12.195 2.773 ;
      RECT 12.135 2.617 12.155 2.771 ;
      RECT 12.075 2.617 12.135 2.768 ;
      RECT 12.055 2.62 12.075 2.766 ;
      RECT 12.034 2.62 12.055 2.766 ;
      RECT 11.948 2.622 12.034 2.77 ;
      RECT 11.862 2.624 11.948 2.776 ;
      RECT 11.776 2.626 11.862 2.783 ;
      RECT 11.69 2.629 11.776 2.789 ;
      RECT 11.656 2.63 11.69 2.794 ;
      RECT 11.57 2.633 11.656 2.799 ;
      RECT 11.541 2.64 11.57 2.804 ;
      RECT 11.455 2.64 11.541 2.809 ;
      RECT 11.422 2.64 11.455 2.814 ;
      RECT 11.336 2.642 11.422 2.819 ;
      RECT 11.25 2.644 11.336 2.826 ;
      RECT 11.186 2.646 11.25 2.832 ;
      RECT 11.1 2.648 11.186 2.838 ;
      RECT 11.097 2.65 11.1 2.841 ;
      RECT 11.011 2.651 11.097 2.845 ;
      RECT 10.925 2.654 11.011 2.852 ;
      RECT 10.906 2.656 10.925 2.856 ;
      RECT 10.82 2.658 10.906 2.861 ;
      RECT 10.55 2.67 10.56 2.865 ;
      RECT 12.73 7.765 13.02 7.995 ;
      RECT 12.79 7.025 12.96 7.995 ;
      RECT 12.68 7.055 13.055 7.425 ;
      RECT 12.73 7.025 13.02 7.425 ;
      RECT 12.785 2.25 12.97 2.46 ;
      RECT 12.78 2.251 12.975 2.458 ;
      RECT 12.775 2.256 12.985 2.453 ;
      RECT 12.77 2.232 12.775 2.45 ;
      RECT 12.74 2.229 12.77 2.443 ;
      RECT 12.735 2.225 12.74 2.434 ;
      RECT 12.7 2.256 12.985 2.429 ;
      RECT 12.475 2.165 12.735 2.425 ;
      RECT 12.775 2.234 12.78 2.453 ;
      RECT 12.78 2.235 12.785 2.458 ;
      RECT 12.475 2.247 12.855 2.425 ;
      RECT 12.475 2.245 12.84 2.425 ;
      RECT 12.475 2.24 12.83 2.425 ;
      RECT 12.43 3.155 12.48 3.44 ;
      RECT 12.375 3.125 12.38 3.44 ;
      RECT 12.345 3.105 12.35 3.44 ;
      RECT 12.495 3.155 12.555 3.415 ;
      RECT 12.49 3.155 12.495 3.423 ;
      RECT 12.48 3.155 12.49 3.435 ;
      RECT 12.395 3.145 12.43 3.44 ;
      RECT 12.39 3.132 12.395 3.44 ;
      RECT 12.38 3.127 12.39 3.44 ;
      RECT 12.36 3.117 12.375 3.44 ;
      RECT 12.35 3.11 12.36 3.44 ;
      RECT 12.34 3.102 12.345 3.44 ;
      RECT 12.31 3.092 12.34 3.44 ;
      RECT 12.295 3.08 12.31 3.44 ;
      RECT 12.28 3.07 12.295 3.435 ;
      RECT 12.26 3.06 12.28 3.41 ;
      RECT 12.25 3.052 12.26 3.387 ;
      RECT 12.22 3.035 12.25 3.377 ;
      RECT 12.215 3.012 12.22 3.368 ;
      RECT 12.21 2.999 12.215 3.366 ;
      RECT 12.195 2.975 12.21 3.36 ;
      RECT 12.19 2.951 12.195 3.354 ;
      RECT 12.18 2.94 12.19 3.349 ;
      RECT 12.175 2.93 12.18 3.345 ;
      RECT 12.17 2.922 12.175 3.342 ;
      RECT 12.16 2.917 12.17 3.338 ;
      RECT 12.155 2.912 12.16 3.334 ;
      RECT 12.07 2.91 12.155 3.309 ;
      RECT 12.04 2.91 12.07 3.275 ;
      RECT 12.025 2.91 12.04 3.258 ;
      RECT 11.97 2.91 12.025 3.203 ;
      RECT 11.965 2.915 11.97 3.152 ;
      RECT 11.955 2.92 11.965 3.142 ;
      RECT 11.95 2.93 11.955 3.128 ;
      RECT 11.9 3.67 12.16 3.93 ;
      RECT 11.82 3.685 12.16 3.906 ;
      RECT 11.8 3.685 12.16 3.901 ;
      RECT 11.776 3.685 12.16 3.899 ;
      RECT 11.69 3.685 12.16 3.894 ;
      RECT 11.54 3.625 11.8 3.89 ;
      RECT 11.495 3.685 12.16 3.885 ;
      RECT 11.49 3.692 12.16 3.88 ;
      RECT 11.505 3.68 11.82 3.89 ;
      RECT 11.395 2.115 11.655 2.375 ;
      RECT 11.395 2.172 11.66 2.368 ;
      RECT 11.395 2.202 11.665 2.3 ;
      RECT 11.455 2.633 11.57 2.635 ;
      RECT 11.541 2.63 11.57 2.635 ;
      RECT 10.565 3.634 10.59 3.874 ;
      RECT 10.55 3.637 10.64 3.868 ;
      RECT 10.545 3.642 10.726 3.863 ;
      RECT 10.54 3.65 10.79 3.861 ;
      RECT 10.54 3.65 10.8 3.86 ;
      RECT 10.535 3.657 10.81 3.853 ;
      RECT 10.535 3.657 10.896 3.842 ;
      RECT 10.53 3.692 10.896 3.838 ;
      RECT 10.53 3.692 10.905 3.827 ;
      RECT 10.81 3.565 11.07 3.825 ;
      RECT 10.52 3.742 11.07 3.823 ;
      RECT 10.79 3.61 10.81 3.858 ;
      RECT 10.726 3.613 10.79 3.862 ;
      RECT 10.64 3.618 10.726 3.867 ;
      RECT 10.57 3.629 11.07 3.825 ;
      RECT 10.59 3.623 10.64 3.872 ;
      RECT 10.715 2.1 10.725 2.362 ;
      RECT 10.705 2.157 10.715 2.365 ;
      RECT 10.68 2.162 10.705 2.371 ;
      RECT 10.655 2.166 10.68 2.383 ;
      RECT 10.645 2.169 10.655 2.393 ;
      RECT 10.64 2.17 10.645 2.398 ;
      RECT 10.635 2.171 10.64 2.403 ;
      RECT 10.63 2.172 10.635 2.405 ;
      RECT 10.605 2.175 10.63 2.408 ;
      RECT 10.575 2.181 10.605 2.411 ;
      RECT 10.51 2.192 10.575 2.414 ;
      RECT 10.465 2.2 10.51 2.418 ;
      RECT 10.45 2.2 10.465 2.426 ;
      RECT 10.445 2.201 10.45 2.433 ;
      RECT 10.44 2.203 10.445 2.436 ;
      RECT 10.435 2.207 10.44 2.439 ;
      RECT 10.425 2.215 10.435 2.443 ;
      RECT 10.42 2.228 10.425 2.448 ;
      RECT 10.415 2.236 10.42 2.45 ;
      RECT 10.41 2.242 10.415 2.45 ;
      RECT 10.405 2.246 10.41 2.453 ;
      RECT 10.4 2.248 10.405 2.456 ;
      RECT 10.395 2.251 10.4 2.459 ;
      RECT 10.385 2.256 10.395 2.463 ;
      RECT 10.38 2.262 10.385 2.468 ;
      RECT 10.37 2.268 10.38 2.472 ;
      RECT 10.355 2.275 10.37 2.478 ;
      RECT 10.326 2.289 10.355 2.488 ;
      RECT 10.24 2.324 10.326 2.52 ;
      RECT 10.22 2.357 10.24 2.549 ;
      RECT 10.2 2.37 10.22 2.56 ;
      RECT 10.18 2.382 10.2 2.571 ;
      RECT 10.13 2.404 10.18 2.591 ;
      RECT 10.115 2.422 10.13 2.608 ;
      RECT 10.11 2.428 10.115 2.611 ;
      RECT 10.105 2.432 10.11 2.614 ;
      RECT 10.1 2.436 10.105 2.618 ;
      RECT 10.095 2.438 10.1 2.621 ;
      RECT 10.085 2.445 10.095 2.624 ;
      RECT 10.08 2.45 10.085 2.628 ;
      RECT 10.075 2.452 10.08 2.631 ;
      RECT 10.07 2.456 10.075 2.634 ;
      RECT 10.065 2.458 10.07 2.638 ;
      RECT 10.05 2.463 10.065 2.643 ;
      RECT 10.045 2.468 10.05 2.646 ;
      RECT 10.04 2.476 10.045 2.649 ;
      RECT 10.035 2.478 10.04 2.652 ;
      RECT 10.03 2.48 10.035 2.655 ;
      RECT 10.02 2.482 10.03 2.661 ;
      RECT 9.985 2.496 10.02 2.673 ;
      RECT 9.975 2.511 9.985 2.683 ;
      RECT 9.9 2.54 9.975 2.707 ;
      RECT 9.895 2.565 9.9 2.73 ;
      RECT 9.88 2.569 9.895 2.736 ;
      RECT 9.87 2.577 9.88 2.741 ;
      RECT 9.84 2.59 9.87 2.745 ;
      RECT 9.83 2.605 9.84 2.75 ;
      RECT 9.82 2.61 9.83 2.753 ;
      RECT 9.815 2.612 9.82 2.755 ;
      RECT 9.8 2.615 9.815 2.758 ;
      RECT 9.795 2.617 9.8 2.761 ;
      RECT 9.775 2.622 9.795 2.765 ;
      RECT 9.745 2.627 9.775 2.773 ;
      RECT 9.72 2.634 9.745 2.781 ;
      RECT 9.715 2.639 9.72 2.786 ;
      RECT 9.685 2.642 9.715 2.79 ;
      RECT 9.645 2.645 9.685 2.8 ;
      RECT 9.61 2.642 9.645 2.812 ;
      RECT 9.6 2.638 9.61 2.819 ;
      RECT 9.575 2.634 9.6 2.825 ;
      RECT 9.57 2.63 9.575 2.83 ;
      RECT 9.53 2.627 9.57 2.83 ;
      RECT 9.515 2.612 9.53 2.831 ;
      RECT 9.492 2.6 9.515 2.831 ;
      RECT 9.406 2.6 9.492 2.832 ;
      RECT 9.32 2.6 9.406 2.834 ;
      RECT 9.3 2.6 9.32 2.831 ;
      RECT 9.295 2.605 9.3 2.826 ;
      RECT 9.29 2.61 9.295 2.824 ;
      RECT 9.28 2.62 9.29 2.822 ;
      RECT 9.275 2.626 9.28 2.815 ;
      RECT 9.27 2.628 9.275 2.8 ;
      RECT 9.265 2.632 9.27 2.79 ;
      RECT 10.725 2.1 10.975 2.36 ;
      RECT 8.45 3.635 8.71 3.895 ;
      RECT 10.745 3.125 10.75 3.335 ;
      RECT 10.75 3.13 10.76 3.33 ;
      RECT 10.7 3.125 10.745 3.35 ;
      RECT 10.69 3.125 10.7 3.37 ;
      RECT 10.671 3.125 10.69 3.375 ;
      RECT 10.585 3.125 10.671 3.372 ;
      RECT 10.555 3.127 10.585 3.37 ;
      RECT 10.5 3.137 10.555 3.368 ;
      RECT 10.435 3.151 10.5 3.366 ;
      RECT 10.43 3.159 10.435 3.365 ;
      RECT 10.415 3.162 10.43 3.363 ;
      RECT 10.35 3.172 10.415 3.359 ;
      RECT 10.302 3.186 10.35 3.36 ;
      RECT 10.216 3.203 10.302 3.374 ;
      RECT 10.13 3.224 10.216 3.391 ;
      RECT 10.11 3.237 10.13 3.401 ;
      RECT 10.065 3.245 10.11 3.408 ;
      RECT 10.03 3.253 10.065 3.416 ;
      RECT 9.996 3.261 10.03 3.424 ;
      RECT 9.91 3.275 9.996 3.436 ;
      RECT 9.875 3.292 9.91 3.448 ;
      RECT 9.866 3.301 9.875 3.452 ;
      RECT 9.78 3.319 9.866 3.469 ;
      RECT 9.721 3.346 9.78 3.496 ;
      RECT 9.635 3.373 9.721 3.524 ;
      RECT 9.615 3.395 9.635 3.544 ;
      RECT 9.555 3.41 9.615 3.56 ;
      RECT 9.545 3.422 9.555 3.573 ;
      RECT 9.54 3.427 9.545 3.576 ;
      RECT 9.53 3.43 9.54 3.579 ;
      RECT 9.525 3.432 9.53 3.582 ;
      RECT 9.495 3.44 9.525 3.589 ;
      RECT 9.48 3.447 9.495 3.597 ;
      RECT 9.47 3.452 9.48 3.601 ;
      RECT 9.465 3.455 9.47 3.604 ;
      RECT 9.455 3.457 9.465 3.607 ;
      RECT 9.42 3.467 9.455 3.616 ;
      RECT 9.345 3.49 9.42 3.638 ;
      RECT 9.325 3.508 9.345 3.656 ;
      RECT 9.295 3.515 9.325 3.666 ;
      RECT 9.275 3.523 9.295 3.676 ;
      RECT 9.265 3.529 9.275 3.683 ;
      RECT 9.246 3.534 9.265 3.689 ;
      RECT 9.16 3.554 9.246 3.709 ;
      RECT 9.145 3.574 9.16 3.728 ;
      RECT 9.1 3.586 9.145 3.739 ;
      RECT 9.035 3.607 9.1 3.762 ;
      RECT 8.995 3.627 9.035 3.783 ;
      RECT 8.985 3.637 8.995 3.793 ;
      RECT 8.935 3.649 8.985 3.804 ;
      RECT 8.915 3.665 8.935 3.816 ;
      RECT 8.885 3.675 8.915 3.822 ;
      RECT 8.875 3.68 8.885 3.824 ;
      RECT 8.806 3.681 8.875 3.83 ;
      RECT 8.72 3.683 8.806 3.84 ;
      RECT 8.71 3.684 8.72 3.845 ;
      RECT 9.98 3.71 10.17 3.92 ;
      RECT 9.97 3.715 10.18 3.913 ;
      RECT 9.955 3.715 10.18 3.878 ;
      RECT 9.875 3.6 10.135 3.86 ;
      RECT 8.79 3.13 8.975 3.425 ;
      RECT 8.78 3.13 8.975 3.423 ;
      RECT 8.765 3.13 8.98 3.418 ;
      RECT 8.765 3.13 8.985 3.415 ;
      RECT 8.76 3.13 8.985 3.413 ;
      RECT 8.755 3.385 8.985 3.403 ;
      RECT 8.76 3.13 9.02 3.39 ;
      RECT 8.72 2.165 8.98 2.425 ;
      RECT 8.53 2.09 8.616 2.423 ;
      RECT 8.505 2.094 8.66 2.419 ;
      RECT 8.616 2.086 8.66 2.419 ;
      RECT 8.616 2.087 8.665 2.418 ;
      RECT 8.53 2.092 8.68 2.417 ;
      RECT 8.505 2.1 8.72 2.416 ;
      RECT 8.5 2.095 8.68 2.411 ;
      RECT 8.49 2.11 8.72 2.318 ;
      RECT 8.49 2.162 8.92 2.318 ;
      RECT 8.49 2.155 8.9 2.318 ;
      RECT 8.49 2.142 8.87 2.318 ;
      RECT 8.49 2.13 8.81 2.318 ;
      RECT 8.49 2.115 8.785 2.318 ;
      RECT 7.69 2.745 7.825 3.04 ;
      RECT 7.95 2.768 7.955 2.955 ;
      RECT 8.67 2.665 8.815 2.9 ;
      RECT 8.83 2.665 8.835 2.89 ;
      RECT 8.865 2.676 8.87 2.87 ;
      RECT 8.86 2.668 8.865 2.875 ;
      RECT 8.84 2.665 8.86 2.88 ;
      RECT 8.835 2.665 8.84 2.888 ;
      RECT 8.825 2.665 8.83 2.893 ;
      RECT 8.815 2.665 8.825 2.898 ;
      RECT 8.645 2.667 8.67 2.9 ;
      RECT 8.595 2.674 8.645 2.9 ;
      RECT 8.59 2.679 8.595 2.9 ;
      RECT 8.551 2.684 8.59 2.901 ;
      RECT 8.465 2.696 8.551 2.902 ;
      RECT 8.456 2.706 8.465 2.902 ;
      RECT 8.37 2.715 8.456 2.904 ;
      RECT 8.346 2.725 8.37 2.906 ;
      RECT 8.26 2.736 8.346 2.907 ;
      RECT 8.23 2.747 8.26 2.909 ;
      RECT 8.2 2.752 8.23 2.911 ;
      RECT 8.175 2.758 8.2 2.914 ;
      RECT 8.16 2.763 8.175 2.915 ;
      RECT 8.115 2.769 8.16 2.915 ;
      RECT 8.11 2.774 8.115 2.916 ;
      RECT 8.09 2.774 8.11 2.918 ;
      RECT 8.07 2.772 8.09 2.923 ;
      RECT 8.035 2.771 8.07 2.93 ;
      RECT 8.005 2.77 8.035 2.94 ;
      RECT 7.955 2.769 8.005 2.95 ;
      RECT 7.865 2.766 7.95 3.04 ;
      RECT 7.84 2.76 7.865 3.04 ;
      RECT 7.825 2.75 7.84 3.04 ;
      RECT 7.64 2.745 7.69 2.96 ;
      RECT 7.63 2.75 7.64 2.95 ;
      RECT 7.87 3.225 8.13 3.485 ;
      RECT 7.87 3.225 8.16 3.378 ;
      RECT 7.87 3.225 8.195 3.363 ;
      RECT 8.125 3.145 8.315 3.355 ;
      RECT 8.115 3.15 8.325 3.348 ;
      RECT 8.08 3.22 8.325 3.348 ;
      RECT 8.11 3.162 8.13 3.485 ;
      RECT 8.095 3.21 8.325 3.348 ;
      RECT 8.1 3.182 8.13 3.485 ;
      RECT 7.18 2.25 7.25 3.355 ;
      RECT 7.915 2.355 8.175 2.615 ;
      RECT 7.495 2.401 7.51 2.61 ;
      RECT 7.831 2.414 7.915 2.565 ;
      RECT 7.745 2.411 7.831 2.565 ;
      RECT 7.706 2.409 7.745 2.565 ;
      RECT 7.62 2.407 7.706 2.565 ;
      RECT 7.56 2.405 7.62 2.576 ;
      RECT 7.525 2.403 7.56 2.594 ;
      RECT 7.51 2.401 7.525 2.605 ;
      RECT 7.48 2.401 7.495 2.618 ;
      RECT 7.47 2.401 7.48 2.623 ;
      RECT 7.445 2.4 7.47 2.628 ;
      RECT 7.43 2.395 7.445 2.634 ;
      RECT 7.425 2.388 7.43 2.639 ;
      RECT 7.4 2.379 7.425 2.645 ;
      RECT 7.355 2.358 7.4 2.658 ;
      RECT 7.345 2.342 7.355 2.668 ;
      RECT 7.33 2.335 7.345 2.678 ;
      RECT 7.32 2.328 7.33 2.695 ;
      RECT 7.315 2.325 7.32 2.725 ;
      RECT 7.31 2.323 7.315 2.755 ;
      RECT 7.305 2.321 7.31 2.792 ;
      RECT 7.29 2.317 7.305 2.859 ;
      RECT 7.29 3.15 7.3 3.35 ;
      RECT 7.285 2.313 7.29 2.985 ;
      RECT 7.285 3.137 7.29 3.355 ;
      RECT 7.28 2.311 7.285 3.07 ;
      RECT 7.28 3.127 7.285 3.355 ;
      RECT 7.265 2.282 7.28 3.355 ;
      RECT 7.25 2.255 7.265 3.355 ;
      RECT 7.175 2.25 7.18 2.605 ;
      RECT 7.175 2.66 7.18 3.355 ;
      RECT 7.16 2.25 7.175 2.583 ;
      RECT 7.17 2.682 7.175 3.355 ;
      RECT 7.16 2.722 7.17 3.355 ;
      RECT 7.125 2.25 7.16 2.525 ;
      RECT 7.155 2.757 7.16 3.355 ;
      RECT 7.14 2.812 7.155 3.355 ;
      RECT 7.135 2.877 7.14 3.355 ;
      RECT 7.12 2.925 7.135 3.355 ;
      RECT 7.095 2.25 7.125 2.48 ;
      RECT 7.115 2.98 7.12 3.355 ;
      RECT 7.1 3.04 7.115 3.355 ;
      RECT 7.095 3.088 7.1 3.353 ;
      RECT 7.09 2.25 7.095 2.473 ;
      RECT 7.09 3.12 7.095 3.348 ;
      RECT 7.065 2.25 7.09 2.465 ;
      RECT 7.055 2.255 7.065 2.455 ;
      RECT 7.27 3.53 7.29 3.77 ;
      RECT 6.5 3.46 6.505 3.67 ;
      RECT 7.78 3.533 7.79 3.728 ;
      RECT 7.775 3.523 7.78 3.731 ;
      RECT 7.695 3.52 7.775 3.754 ;
      RECT 7.691 3.52 7.695 3.776 ;
      RECT 7.605 3.52 7.691 3.786 ;
      RECT 7.59 3.52 7.605 3.794 ;
      RECT 7.561 3.521 7.59 3.792 ;
      RECT 7.475 3.526 7.561 3.788 ;
      RECT 7.462 3.53 7.475 3.784 ;
      RECT 7.376 3.53 7.462 3.78 ;
      RECT 7.29 3.53 7.376 3.774 ;
      RECT 7.206 3.53 7.27 3.768 ;
      RECT 7.12 3.53 7.206 3.763 ;
      RECT 7.1 3.53 7.12 3.759 ;
      RECT 7.04 3.525 7.1 3.756 ;
      RECT 7.012 3.519 7.04 3.753 ;
      RECT 6.926 3.514 7.012 3.749 ;
      RECT 6.84 3.508 6.926 3.743 ;
      RECT 6.765 3.49 6.84 3.738 ;
      RECT 6.73 3.467 6.765 3.734 ;
      RECT 6.72 3.457 6.73 3.733 ;
      RECT 6.665 3.455 6.72 3.732 ;
      RECT 6.59 3.455 6.665 3.728 ;
      RECT 6.58 3.455 6.59 3.723 ;
      RECT 6.565 3.455 6.58 3.715 ;
      RECT 6.515 3.457 6.565 3.693 ;
      RECT 6.505 3.46 6.515 3.673 ;
      RECT 6.495 3.465 6.5 3.668 ;
      RECT 6.49 3.47 6.495 3.663 ;
      RECT 6.615 2.635 6.875 2.895 ;
      RECT 6.615 2.65 6.895 2.86 ;
      RECT 6.615 2.655 6.905 2.855 ;
      RECT 4.6 2.115 4.86 2.375 ;
      RECT 4.59 2.145 4.86 2.355 ;
      RECT 6.51 2.06 6.77 2.32 ;
      RECT 6.505 2.135 6.51 2.321 ;
      RECT 6.48 2.14 6.505 2.323 ;
      RECT 6.465 2.147 6.48 2.326 ;
      RECT 6.405 2.165 6.465 2.331 ;
      RECT 6.375 2.185 6.405 2.338 ;
      RECT 6.35 2.193 6.375 2.343 ;
      RECT 6.325 2.201 6.35 2.345 ;
      RECT 6.307 2.205 6.325 2.344 ;
      RECT 6.221 2.203 6.307 2.344 ;
      RECT 6.135 2.201 6.221 2.344 ;
      RECT 6.049 2.199 6.135 2.343 ;
      RECT 5.963 2.197 6.049 2.343 ;
      RECT 5.877 2.195 5.963 2.343 ;
      RECT 5.791 2.193 5.877 2.343 ;
      RECT 5.705 2.191 5.791 2.342 ;
      RECT 5.687 2.19 5.705 2.342 ;
      RECT 5.601 2.189 5.687 2.342 ;
      RECT 5.515 2.187 5.601 2.342 ;
      RECT 5.429 2.186 5.515 2.341 ;
      RECT 5.343 2.185 5.429 2.341 ;
      RECT 5.257 2.183 5.343 2.341 ;
      RECT 5.171 2.182 5.257 2.341 ;
      RECT 5.085 2.18 5.171 2.34 ;
      RECT 5.061 2.178 5.085 2.34 ;
      RECT 4.975 2.171 5.061 2.34 ;
      RECT 4.946 2.163 4.975 2.34 ;
      RECT 4.86 2.155 4.946 2.34 ;
      RECT 4.58 2.152 4.59 2.35 ;
      RECT 6.085 3.115 6.09 3.465 ;
      RECT 5.855 3.205 5.995 3.465 ;
      RECT 6.33 2.89 6.375 3.1 ;
      RECT 6.385 2.901 6.395 3.095 ;
      RECT 6.375 2.893 6.385 3.1 ;
      RECT 6.31 2.89 6.33 3.105 ;
      RECT 6.28 2.89 6.31 3.128 ;
      RECT 6.27 2.89 6.28 3.153 ;
      RECT 6.265 2.89 6.27 3.163 ;
      RECT 6.21 2.89 6.265 3.203 ;
      RECT 6.205 2.89 6.21 3.243 ;
      RECT 6.2 2.892 6.205 3.248 ;
      RECT 6.185 2.902 6.2 3.259 ;
      RECT 6.14 2.96 6.185 3.295 ;
      RECT 6.13 3.015 6.14 3.329 ;
      RECT 6.115 3.042 6.13 3.345 ;
      RECT 6.105 3.069 6.115 3.465 ;
      RECT 6.09 3.092 6.105 3.465 ;
      RECT 6.08 3.132 6.085 3.465 ;
      RECT 6.075 3.142 6.08 3.465 ;
      RECT 6.07 3.157 6.075 3.465 ;
      RECT 6.06 3.162 6.07 3.465 ;
      RECT 5.995 3.185 6.06 3.465 ;
      RECT 5.495 2.68 5.685 2.89 ;
      RECT 4.07 2.605 4.33 2.865 ;
      RECT 4.42 2.6 4.515 2.81 ;
      RECT 4.395 2.615 4.405 2.81 ;
      RECT 5.685 2.687 5.695 2.885 ;
      RECT 5.485 2.687 5.495 2.885 ;
      RECT 5.47 2.702 5.485 2.875 ;
      RECT 5.465 2.71 5.47 2.868 ;
      RECT 5.455 2.713 5.465 2.865 ;
      RECT 5.42 2.712 5.455 2.863 ;
      RECT 5.391 2.708 5.42 2.86 ;
      RECT 5.305 2.703 5.391 2.857 ;
      RECT 5.245 2.697 5.305 2.853 ;
      RECT 5.216 2.693 5.245 2.85 ;
      RECT 5.13 2.685 5.216 2.847 ;
      RECT 5.121 2.679 5.13 2.845 ;
      RECT 5.035 2.674 5.121 2.843 ;
      RECT 5.012 2.669 5.035 2.84 ;
      RECT 4.926 2.663 5.012 2.837 ;
      RECT 4.84 2.654 4.926 2.832 ;
      RECT 4.83 2.649 4.84 2.83 ;
      RECT 4.811 2.648 4.83 2.829 ;
      RECT 4.725 2.643 4.811 2.825 ;
      RECT 4.705 2.638 4.725 2.821 ;
      RECT 4.645 2.633 4.705 2.818 ;
      RECT 4.62 2.623 4.645 2.816 ;
      RECT 4.615 2.616 4.62 2.815 ;
      RECT 4.605 2.607 4.615 2.814 ;
      RECT 4.601 2.6 4.605 2.814 ;
      RECT 4.515 2.6 4.601 2.812 ;
      RECT 4.405 2.607 4.42 2.81 ;
      RECT 4.39 2.617 4.395 2.81 ;
      RECT 4.37 2.62 4.39 2.807 ;
      RECT 4.34 2.62 4.37 2.803 ;
      RECT 4.33 2.62 4.34 2.803 ;
      RECT 5.245 3.115 5.505 3.375 ;
      RECT 5.175 3.125 5.505 3.335 ;
      RECT 5.165 3.132 5.505 3.33 ;
      RECT 4.585 3.12 4.845 3.38 ;
      RECT 4.585 3.16 4.95 3.37 ;
      RECT 4.585 3.162 4.955 3.369 ;
      RECT 4.585 3.17 4.96 3.366 ;
      RECT 3.51 2.245 3.61 3.77 ;
      RECT 3.7 3.385 3.75 3.645 ;
      RECT 3.695 2.258 3.7 2.445 ;
      RECT 3.69 3.366 3.7 3.645 ;
      RECT 3.69 2.255 3.695 2.453 ;
      RECT 3.675 2.249 3.69 2.46 ;
      RECT 3.685 3.354 3.69 3.728 ;
      RECT 3.675 3.342 3.685 3.765 ;
      RECT 3.665 2.245 3.675 2.467 ;
      RECT 3.665 3.327 3.675 3.77 ;
      RECT 3.66 2.245 3.665 2.475 ;
      RECT 3.64 3.297 3.665 3.77 ;
      RECT 3.62 2.245 3.66 2.523 ;
      RECT 3.63 3.257 3.64 3.77 ;
      RECT 3.62 3.212 3.63 3.77 ;
      RECT 3.615 2.245 3.62 2.593 ;
      RECT 3.615 3.17 3.62 3.77 ;
      RECT 3.61 2.245 3.615 3.07 ;
      RECT 3.61 3.152 3.615 3.77 ;
      RECT 3.5 2.248 3.51 3.77 ;
      RECT 3.485 2.255 3.5 3.766 ;
      RECT 3.48 2.265 3.485 3.761 ;
      RECT 3.475 2.465 3.48 3.653 ;
      RECT 3.47 2.55 3.475 3.205 ;
      RECT 2.13 6.655 2.42 6.885 ;
      RECT 1.96 6.685 2.42 6.855 ;
      RECT 1.7 7.765 1.99 7.995 ;
      RECT 1.76 7.025 1.93 7.995 ;
      RECT 1.67 7.025 2.02 7.315 ;
      RECT 1.295 6.285 1.645 6.575 ;
      RECT 1.155 6.315 1.645 6.485 ;
      RECT 0.33 5.915 0.62 6.145 ;
      RECT 0.33 5.945 0.79 6.115 ;
      RECT 87.2 1.14 87.575 1.51 ;
      RECT 81.18 2.225 81.44 2.485 ;
      RECT 69.275 1.14 69.65 1.51 ;
      RECT 63.255 2.225 63.515 2.485 ;
      RECT 51.35 1.14 51.725 1.51 ;
      RECT 45.33 2.225 45.59 2.485 ;
      RECT 33.425 1.14 33.8 1.51 ;
      RECT 27.405 2.225 27.665 2.485 ;
      RECT 15.5 1.14 15.875 1.51 ;
      RECT 9.48 2.225 9.74 2.485 ;
    LAYER mcon ;
      RECT 92.035 0.915 92.205 1.085 ;
      RECT 92.035 2.395 92.205 2.565 ;
      RECT 92.035 6.315 92.205 6.485 ;
      RECT 92.035 7.795 92.205 7.965 ;
      RECT 91.685 0.105 91.855 0.275 ;
      RECT 91.685 4.165 91.855 4.335 ;
      RECT 91.685 4.545 91.855 4.715 ;
      RECT 91.685 8.605 91.855 8.775 ;
      RECT 91.665 2.765 91.835 2.935 ;
      RECT 91.665 5.945 91.835 6.115 ;
      RECT 91.045 0.915 91.215 1.085 ;
      RECT 91.045 2.395 91.215 2.565 ;
      RECT 91.045 6.315 91.215 6.485 ;
      RECT 91.045 7.795 91.215 7.965 ;
      RECT 90.695 0.105 90.865 0.275 ;
      RECT 90.695 4.165 90.865 4.335 ;
      RECT 90.695 4.545 90.865 4.715 ;
      RECT 90.695 8.605 90.865 8.775 ;
      RECT 90.675 2.765 90.845 2.935 ;
      RECT 90.675 5.945 90.845 6.115 ;
      RECT 89.99 0.105 90.16 0.275 ;
      RECT 89.99 4.165 90.16 4.335 ;
      RECT 89.99 4.545 90.16 4.715 ;
      RECT 89.99 8.605 90.16 8.775 ;
      RECT 89.68 2.025 89.85 2.195 ;
      RECT 89.68 6.685 89.85 6.855 ;
      RECT 89.31 0.105 89.48 0.275 ;
      RECT 89.31 8.605 89.48 8.775 ;
      RECT 89.25 0.915 89.42 1.085 ;
      RECT 89.25 1.655 89.42 1.825 ;
      RECT 89.25 7.055 89.42 7.225 ;
      RECT 89.25 7.795 89.42 7.965 ;
      RECT 88.875 2.395 89.045 2.565 ;
      RECT 88.875 6.315 89.045 6.485 ;
      RECT 88.63 0.105 88.8 0.275 ;
      RECT 88.63 8.605 88.8 8.775 ;
      RECT 87.95 0.105 88.12 0.275 ;
      RECT 87.95 8.605 88.12 8.775 ;
      RECT 87.88 2.765 88.05 2.935 ;
      RECT 87.88 5.945 88.05 6.115 ;
      RECT 86.67 1.565 86.84 1.735 ;
      RECT 86.67 4.285 86.84 4.455 ;
      RECT 86.21 1.565 86.38 1.735 ;
      RECT 86.21 4.285 86.38 4.455 ;
      RECT 85.815 2.905 85.985 3.075 ;
      RECT 85.75 1.565 85.92 1.735 ;
      RECT 85.75 4.285 85.92 4.455 ;
      RECT 85.605 2.245 85.775 2.415 ;
      RECT 85.29 1.565 85.46 1.735 ;
      RECT 85.29 3.155 85.46 3.325 ;
      RECT 85.29 4.285 85.46 4.455 ;
      RECT 85.23 4.545 85.4 4.715 ;
      RECT 85.23 8.605 85.4 8.775 ;
      RECT 84.92 6.685 85.09 6.855 ;
      RECT 84.905 2.75 85.075 2.92 ;
      RECT 84.83 1.565 85 1.735 ;
      RECT 84.83 4.285 85 4.455 ;
      RECT 84.69 3.315 84.86 3.485 ;
      RECT 84.67 3.715 84.84 3.885 ;
      RECT 84.55 8.605 84.72 8.775 ;
      RECT 84.495 2.27 84.665 2.44 ;
      RECT 84.49 7.055 84.66 7.225 ;
      RECT 84.49 7.795 84.66 7.965 ;
      RECT 84.37 1.565 84.54 1.735 ;
      RECT 84.37 4.285 84.54 4.455 ;
      RECT 84.115 6.315 84.285 6.485 ;
      RECT 84 3.25 84.17 3.42 ;
      RECT 83.91 1.565 84.08 1.735 ;
      RECT 83.91 4.285 84.08 4.455 ;
      RECT 83.87 8.605 84.04 8.775 ;
      RECT 83.675 2.935 83.845 3.105 ;
      RECT 83.61 3.715 83.78 3.885 ;
      RECT 83.45 1.565 83.62 1.735 ;
      RECT 83.45 4.285 83.62 4.455 ;
      RECT 83.21 3.7 83.38 3.87 ;
      RECT 83.19 8.605 83.36 8.775 ;
      RECT 83.17 2.185 83.34 2.355 ;
      RECT 83.12 5.945 83.29 6.115 ;
      RECT 82.99 1.565 83.16 1.735 ;
      RECT 82.99 4.285 83.16 4.455 ;
      RECT 82.53 1.565 82.7 1.735 ;
      RECT 82.53 4.285 82.7 4.455 ;
      RECT 82.27 2.685 82.44 2.855 ;
      RECT 82.27 3.145 82.44 3.315 ;
      RECT 82.27 3.66 82.44 3.83 ;
      RECT 82.155 2.22 82.325 2.39 ;
      RECT 82.07 1.565 82.24 1.735 ;
      RECT 82.07 4.285 82.24 4.455 ;
      RECT 81.69 3.73 81.86 3.9 ;
      RECT 81.61 1.565 81.78 1.735 ;
      RECT 81.61 4.285 81.78 4.455 ;
      RECT 81.21 2.26 81.38 2.43 ;
      RECT 81.15 1.565 81.32 1.735 ;
      RECT 81.15 4.285 81.32 4.455 ;
      RECT 80.995 2.635 81.165 2.805 ;
      RECT 80.69 1.565 80.86 1.735 ;
      RECT 80.69 4.285 80.86 4.455 ;
      RECT 80.495 3.235 80.665 3.405 ;
      RECT 80.38 2.685 80.55 2.855 ;
      RECT 80.23 1.565 80.4 1.735 ;
      RECT 80.23 4.285 80.4 4.455 ;
      RECT 80.21 2.135 80.38 2.305 ;
      RECT 79.835 3.165 80.005 3.335 ;
      RECT 79.77 1.565 79.94 1.735 ;
      RECT 79.77 4.285 79.94 4.455 ;
      RECT 79.35 2.765 79.52 2.935 ;
      RECT 79.31 1.565 79.48 1.735 ;
      RECT 79.31 4.285 79.48 4.455 ;
      RECT 79.3 3.54 79.47 3.71 ;
      RECT 78.85 1.565 79.02 1.735 ;
      RECT 78.85 4.285 79.02 4.455 ;
      RECT 78.81 3.165 78.98 3.335 ;
      RECT 78.775 2.27 78.945 2.44 ;
      RECT 78.415 2.67 78.585 2.84 ;
      RECT 78.39 1.565 78.56 1.735 ;
      RECT 78.39 4.285 78.56 4.455 ;
      RECT 78.21 3.48 78.38 3.65 ;
      RECT 77.93 1.565 78.1 1.735 ;
      RECT 77.93 4.285 78.1 4.455 ;
      RECT 77.905 2.91 78.075 3.08 ;
      RECT 77.47 1.565 77.64 1.735 ;
      RECT 77.47 4.285 77.64 4.455 ;
      RECT 77.205 2.7 77.375 2.87 ;
      RECT 77.01 1.565 77.18 1.735 ;
      RECT 77.01 4.285 77.18 4.455 ;
      RECT 76.885 3.145 77.055 3.315 ;
      RECT 76.55 1.565 76.72 1.735 ;
      RECT 76.55 4.285 76.72 4.455 ;
      RECT 76.47 3.18 76.64 3.35 ;
      RECT 76.3 2.165 76.47 2.335 ;
      RECT 76.125 2.62 76.295 2.79 ;
      RECT 76.09 1.565 76.26 1.735 ;
      RECT 76.09 4.285 76.26 4.455 ;
      RECT 75.63 1.565 75.8 1.735 ;
      RECT 75.63 4.285 75.8 4.455 ;
      RECT 75.205 2.27 75.375 2.44 ;
      RECT 75.2 3.585 75.37 3.755 ;
      RECT 75.17 1.565 75.34 1.735 ;
      RECT 75.17 4.285 75.34 4.455 ;
      RECT 74.11 0.915 74.28 1.085 ;
      RECT 74.11 2.395 74.28 2.565 ;
      RECT 74.11 6.315 74.28 6.485 ;
      RECT 74.11 7.795 74.28 7.965 ;
      RECT 73.76 0.105 73.93 0.275 ;
      RECT 73.76 4.165 73.93 4.335 ;
      RECT 73.76 4.545 73.93 4.715 ;
      RECT 73.76 8.605 73.93 8.775 ;
      RECT 73.74 2.765 73.91 2.935 ;
      RECT 73.74 5.945 73.91 6.115 ;
      RECT 73.12 0.915 73.29 1.085 ;
      RECT 73.12 2.395 73.29 2.565 ;
      RECT 73.12 6.315 73.29 6.485 ;
      RECT 73.12 7.795 73.29 7.965 ;
      RECT 72.77 0.105 72.94 0.275 ;
      RECT 72.77 4.165 72.94 4.335 ;
      RECT 72.77 4.545 72.94 4.715 ;
      RECT 72.77 8.605 72.94 8.775 ;
      RECT 72.75 2.765 72.92 2.935 ;
      RECT 72.75 5.945 72.92 6.115 ;
      RECT 72.065 0.105 72.235 0.275 ;
      RECT 72.065 4.165 72.235 4.335 ;
      RECT 72.065 4.545 72.235 4.715 ;
      RECT 72.065 8.605 72.235 8.775 ;
      RECT 71.755 2.025 71.925 2.195 ;
      RECT 71.755 6.685 71.925 6.855 ;
      RECT 71.385 0.105 71.555 0.275 ;
      RECT 71.385 8.605 71.555 8.775 ;
      RECT 71.325 0.915 71.495 1.085 ;
      RECT 71.325 1.655 71.495 1.825 ;
      RECT 71.325 7.055 71.495 7.225 ;
      RECT 71.325 7.795 71.495 7.965 ;
      RECT 70.95 2.395 71.12 2.565 ;
      RECT 70.95 6.315 71.12 6.485 ;
      RECT 70.705 0.105 70.875 0.275 ;
      RECT 70.705 8.605 70.875 8.775 ;
      RECT 70.025 0.105 70.195 0.275 ;
      RECT 70.025 8.605 70.195 8.775 ;
      RECT 69.955 2.765 70.125 2.935 ;
      RECT 69.955 5.945 70.125 6.115 ;
      RECT 68.745 1.565 68.915 1.735 ;
      RECT 68.745 4.285 68.915 4.455 ;
      RECT 68.285 1.565 68.455 1.735 ;
      RECT 68.285 4.285 68.455 4.455 ;
      RECT 67.89 2.905 68.06 3.075 ;
      RECT 67.825 1.565 67.995 1.735 ;
      RECT 67.825 4.285 67.995 4.455 ;
      RECT 67.68 2.245 67.85 2.415 ;
      RECT 67.365 1.565 67.535 1.735 ;
      RECT 67.365 3.155 67.535 3.325 ;
      RECT 67.365 4.285 67.535 4.455 ;
      RECT 67.305 4.545 67.475 4.715 ;
      RECT 67.305 8.605 67.475 8.775 ;
      RECT 66.995 6.685 67.165 6.855 ;
      RECT 66.98 2.75 67.15 2.92 ;
      RECT 66.905 1.565 67.075 1.735 ;
      RECT 66.905 4.285 67.075 4.455 ;
      RECT 66.765 3.315 66.935 3.485 ;
      RECT 66.745 3.715 66.915 3.885 ;
      RECT 66.625 8.605 66.795 8.775 ;
      RECT 66.57 2.27 66.74 2.44 ;
      RECT 66.565 7.055 66.735 7.225 ;
      RECT 66.565 7.795 66.735 7.965 ;
      RECT 66.445 1.565 66.615 1.735 ;
      RECT 66.445 4.285 66.615 4.455 ;
      RECT 66.19 6.315 66.36 6.485 ;
      RECT 66.075 3.25 66.245 3.42 ;
      RECT 65.985 1.565 66.155 1.735 ;
      RECT 65.985 4.285 66.155 4.455 ;
      RECT 65.945 8.605 66.115 8.775 ;
      RECT 65.75 2.935 65.92 3.105 ;
      RECT 65.685 3.715 65.855 3.885 ;
      RECT 65.525 1.565 65.695 1.735 ;
      RECT 65.525 4.285 65.695 4.455 ;
      RECT 65.285 3.7 65.455 3.87 ;
      RECT 65.265 8.605 65.435 8.775 ;
      RECT 65.245 2.185 65.415 2.355 ;
      RECT 65.195 5.945 65.365 6.115 ;
      RECT 65.065 1.565 65.235 1.735 ;
      RECT 65.065 4.285 65.235 4.455 ;
      RECT 64.605 1.565 64.775 1.735 ;
      RECT 64.605 4.285 64.775 4.455 ;
      RECT 64.345 2.685 64.515 2.855 ;
      RECT 64.345 3.145 64.515 3.315 ;
      RECT 64.345 3.66 64.515 3.83 ;
      RECT 64.23 2.22 64.4 2.39 ;
      RECT 64.145 1.565 64.315 1.735 ;
      RECT 64.145 4.285 64.315 4.455 ;
      RECT 63.765 3.73 63.935 3.9 ;
      RECT 63.685 1.565 63.855 1.735 ;
      RECT 63.685 4.285 63.855 4.455 ;
      RECT 63.285 2.26 63.455 2.43 ;
      RECT 63.225 1.565 63.395 1.735 ;
      RECT 63.225 4.285 63.395 4.455 ;
      RECT 63.07 2.635 63.24 2.805 ;
      RECT 62.765 1.565 62.935 1.735 ;
      RECT 62.765 4.285 62.935 4.455 ;
      RECT 62.57 3.235 62.74 3.405 ;
      RECT 62.455 2.685 62.625 2.855 ;
      RECT 62.305 1.565 62.475 1.735 ;
      RECT 62.305 4.285 62.475 4.455 ;
      RECT 62.285 2.135 62.455 2.305 ;
      RECT 61.91 3.165 62.08 3.335 ;
      RECT 61.845 1.565 62.015 1.735 ;
      RECT 61.845 4.285 62.015 4.455 ;
      RECT 61.425 2.765 61.595 2.935 ;
      RECT 61.385 1.565 61.555 1.735 ;
      RECT 61.385 4.285 61.555 4.455 ;
      RECT 61.375 3.54 61.545 3.71 ;
      RECT 60.925 1.565 61.095 1.735 ;
      RECT 60.925 4.285 61.095 4.455 ;
      RECT 60.885 3.165 61.055 3.335 ;
      RECT 60.85 2.27 61.02 2.44 ;
      RECT 60.49 2.67 60.66 2.84 ;
      RECT 60.465 1.565 60.635 1.735 ;
      RECT 60.465 4.285 60.635 4.455 ;
      RECT 60.285 3.48 60.455 3.65 ;
      RECT 60.005 1.565 60.175 1.735 ;
      RECT 60.005 4.285 60.175 4.455 ;
      RECT 59.98 2.91 60.15 3.08 ;
      RECT 59.545 1.565 59.715 1.735 ;
      RECT 59.545 4.285 59.715 4.455 ;
      RECT 59.28 2.7 59.45 2.87 ;
      RECT 59.085 1.565 59.255 1.735 ;
      RECT 59.085 4.285 59.255 4.455 ;
      RECT 58.96 3.145 59.13 3.315 ;
      RECT 58.625 1.565 58.795 1.735 ;
      RECT 58.625 4.285 58.795 4.455 ;
      RECT 58.545 3.18 58.715 3.35 ;
      RECT 58.375 2.165 58.545 2.335 ;
      RECT 58.2 2.62 58.37 2.79 ;
      RECT 58.165 1.565 58.335 1.735 ;
      RECT 58.165 4.285 58.335 4.455 ;
      RECT 57.705 1.565 57.875 1.735 ;
      RECT 57.705 4.285 57.875 4.455 ;
      RECT 57.28 2.27 57.45 2.44 ;
      RECT 57.275 3.585 57.445 3.755 ;
      RECT 57.245 1.565 57.415 1.735 ;
      RECT 57.245 4.285 57.415 4.455 ;
      RECT 56.185 0.915 56.355 1.085 ;
      RECT 56.185 2.395 56.355 2.565 ;
      RECT 56.185 6.315 56.355 6.485 ;
      RECT 56.185 7.795 56.355 7.965 ;
      RECT 55.835 0.105 56.005 0.275 ;
      RECT 55.835 4.165 56.005 4.335 ;
      RECT 55.835 4.545 56.005 4.715 ;
      RECT 55.835 8.605 56.005 8.775 ;
      RECT 55.815 2.765 55.985 2.935 ;
      RECT 55.815 5.945 55.985 6.115 ;
      RECT 55.195 0.915 55.365 1.085 ;
      RECT 55.195 2.395 55.365 2.565 ;
      RECT 55.195 6.315 55.365 6.485 ;
      RECT 55.195 7.795 55.365 7.965 ;
      RECT 54.845 0.105 55.015 0.275 ;
      RECT 54.845 4.165 55.015 4.335 ;
      RECT 54.845 4.545 55.015 4.715 ;
      RECT 54.845 8.605 55.015 8.775 ;
      RECT 54.825 2.765 54.995 2.935 ;
      RECT 54.825 5.945 54.995 6.115 ;
      RECT 54.14 0.105 54.31 0.275 ;
      RECT 54.14 4.165 54.31 4.335 ;
      RECT 54.14 4.545 54.31 4.715 ;
      RECT 54.14 8.605 54.31 8.775 ;
      RECT 53.83 2.025 54 2.195 ;
      RECT 53.83 6.685 54 6.855 ;
      RECT 53.46 0.105 53.63 0.275 ;
      RECT 53.46 8.605 53.63 8.775 ;
      RECT 53.4 0.915 53.57 1.085 ;
      RECT 53.4 1.655 53.57 1.825 ;
      RECT 53.4 7.055 53.57 7.225 ;
      RECT 53.4 7.795 53.57 7.965 ;
      RECT 53.025 2.395 53.195 2.565 ;
      RECT 53.025 6.315 53.195 6.485 ;
      RECT 52.78 0.105 52.95 0.275 ;
      RECT 52.78 8.605 52.95 8.775 ;
      RECT 52.1 0.105 52.27 0.275 ;
      RECT 52.1 8.605 52.27 8.775 ;
      RECT 52.03 2.765 52.2 2.935 ;
      RECT 52.03 5.945 52.2 6.115 ;
      RECT 50.82 1.565 50.99 1.735 ;
      RECT 50.82 4.285 50.99 4.455 ;
      RECT 50.36 1.565 50.53 1.735 ;
      RECT 50.36 4.285 50.53 4.455 ;
      RECT 49.965 2.905 50.135 3.075 ;
      RECT 49.9 1.565 50.07 1.735 ;
      RECT 49.9 4.285 50.07 4.455 ;
      RECT 49.755 2.245 49.925 2.415 ;
      RECT 49.44 1.565 49.61 1.735 ;
      RECT 49.44 3.155 49.61 3.325 ;
      RECT 49.44 4.285 49.61 4.455 ;
      RECT 49.38 4.545 49.55 4.715 ;
      RECT 49.38 8.605 49.55 8.775 ;
      RECT 49.07 6.685 49.24 6.855 ;
      RECT 49.055 2.75 49.225 2.92 ;
      RECT 48.98 1.565 49.15 1.735 ;
      RECT 48.98 4.285 49.15 4.455 ;
      RECT 48.84 3.315 49.01 3.485 ;
      RECT 48.82 3.715 48.99 3.885 ;
      RECT 48.7 8.605 48.87 8.775 ;
      RECT 48.645 2.27 48.815 2.44 ;
      RECT 48.64 7.055 48.81 7.225 ;
      RECT 48.64 7.795 48.81 7.965 ;
      RECT 48.52 1.565 48.69 1.735 ;
      RECT 48.52 4.285 48.69 4.455 ;
      RECT 48.265 6.315 48.435 6.485 ;
      RECT 48.15 3.25 48.32 3.42 ;
      RECT 48.06 1.565 48.23 1.735 ;
      RECT 48.06 4.285 48.23 4.455 ;
      RECT 48.02 8.605 48.19 8.775 ;
      RECT 47.825 2.935 47.995 3.105 ;
      RECT 47.76 3.715 47.93 3.885 ;
      RECT 47.6 1.565 47.77 1.735 ;
      RECT 47.6 4.285 47.77 4.455 ;
      RECT 47.36 3.7 47.53 3.87 ;
      RECT 47.34 8.605 47.51 8.775 ;
      RECT 47.32 2.185 47.49 2.355 ;
      RECT 47.27 5.945 47.44 6.115 ;
      RECT 47.14 1.565 47.31 1.735 ;
      RECT 47.14 4.285 47.31 4.455 ;
      RECT 46.68 1.565 46.85 1.735 ;
      RECT 46.68 4.285 46.85 4.455 ;
      RECT 46.42 2.685 46.59 2.855 ;
      RECT 46.42 3.145 46.59 3.315 ;
      RECT 46.42 3.66 46.59 3.83 ;
      RECT 46.305 2.22 46.475 2.39 ;
      RECT 46.22 1.565 46.39 1.735 ;
      RECT 46.22 4.285 46.39 4.455 ;
      RECT 45.84 3.73 46.01 3.9 ;
      RECT 45.76 1.565 45.93 1.735 ;
      RECT 45.76 4.285 45.93 4.455 ;
      RECT 45.36 2.26 45.53 2.43 ;
      RECT 45.3 1.565 45.47 1.735 ;
      RECT 45.3 4.285 45.47 4.455 ;
      RECT 45.145 2.635 45.315 2.805 ;
      RECT 44.84 1.565 45.01 1.735 ;
      RECT 44.84 4.285 45.01 4.455 ;
      RECT 44.645 3.235 44.815 3.405 ;
      RECT 44.53 2.685 44.7 2.855 ;
      RECT 44.38 1.565 44.55 1.735 ;
      RECT 44.38 4.285 44.55 4.455 ;
      RECT 44.36 2.135 44.53 2.305 ;
      RECT 43.985 3.165 44.155 3.335 ;
      RECT 43.92 1.565 44.09 1.735 ;
      RECT 43.92 4.285 44.09 4.455 ;
      RECT 43.5 2.765 43.67 2.935 ;
      RECT 43.46 1.565 43.63 1.735 ;
      RECT 43.46 4.285 43.63 4.455 ;
      RECT 43.45 3.54 43.62 3.71 ;
      RECT 43 1.565 43.17 1.735 ;
      RECT 43 4.285 43.17 4.455 ;
      RECT 42.96 3.165 43.13 3.335 ;
      RECT 42.925 2.27 43.095 2.44 ;
      RECT 42.565 2.67 42.735 2.84 ;
      RECT 42.54 1.565 42.71 1.735 ;
      RECT 42.54 4.285 42.71 4.455 ;
      RECT 42.36 3.48 42.53 3.65 ;
      RECT 42.08 1.565 42.25 1.735 ;
      RECT 42.08 4.285 42.25 4.455 ;
      RECT 42.055 2.91 42.225 3.08 ;
      RECT 41.62 1.565 41.79 1.735 ;
      RECT 41.62 4.285 41.79 4.455 ;
      RECT 41.355 2.7 41.525 2.87 ;
      RECT 41.16 1.565 41.33 1.735 ;
      RECT 41.16 4.285 41.33 4.455 ;
      RECT 41.035 3.145 41.205 3.315 ;
      RECT 40.7 1.565 40.87 1.735 ;
      RECT 40.7 4.285 40.87 4.455 ;
      RECT 40.62 3.18 40.79 3.35 ;
      RECT 40.45 2.165 40.62 2.335 ;
      RECT 40.275 2.62 40.445 2.79 ;
      RECT 40.24 1.565 40.41 1.735 ;
      RECT 40.24 4.285 40.41 4.455 ;
      RECT 39.78 1.565 39.95 1.735 ;
      RECT 39.78 4.285 39.95 4.455 ;
      RECT 39.355 2.27 39.525 2.44 ;
      RECT 39.35 3.585 39.52 3.755 ;
      RECT 39.32 1.565 39.49 1.735 ;
      RECT 39.32 4.285 39.49 4.455 ;
      RECT 38.26 0.915 38.43 1.085 ;
      RECT 38.26 2.395 38.43 2.565 ;
      RECT 38.26 6.315 38.43 6.485 ;
      RECT 38.26 7.795 38.43 7.965 ;
      RECT 37.91 0.105 38.08 0.275 ;
      RECT 37.91 4.165 38.08 4.335 ;
      RECT 37.91 4.545 38.08 4.715 ;
      RECT 37.91 8.605 38.08 8.775 ;
      RECT 37.89 2.765 38.06 2.935 ;
      RECT 37.89 5.945 38.06 6.115 ;
      RECT 37.27 0.915 37.44 1.085 ;
      RECT 37.27 2.395 37.44 2.565 ;
      RECT 37.27 6.315 37.44 6.485 ;
      RECT 37.27 7.795 37.44 7.965 ;
      RECT 36.92 0.105 37.09 0.275 ;
      RECT 36.92 4.165 37.09 4.335 ;
      RECT 36.92 4.545 37.09 4.715 ;
      RECT 36.92 8.605 37.09 8.775 ;
      RECT 36.9 2.765 37.07 2.935 ;
      RECT 36.9 5.945 37.07 6.115 ;
      RECT 36.215 0.105 36.385 0.275 ;
      RECT 36.215 4.165 36.385 4.335 ;
      RECT 36.215 4.545 36.385 4.715 ;
      RECT 36.215 8.605 36.385 8.775 ;
      RECT 35.905 2.025 36.075 2.195 ;
      RECT 35.905 6.685 36.075 6.855 ;
      RECT 35.535 0.105 35.705 0.275 ;
      RECT 35.535 8.605 35.705 8.775 ;
      RECT 35.475 0.915 35.645 1.085 ;
      RECT 35.475 1.655 35.645 1.825 ;
      RECT 35.475 7.055 35.645 7.225 ;
      RECT 35.475 7.795 35.645 7.965 ;
      RECT 35.1 2.395 35.27 2.565 ;
      RECT 35.1 6.315 35.27 6.485 ;
      RECT 34.855 0.105 35.025 0.275 ;
      RECT 34.855 8.605 35.025 8.775 ;
      RECT 34.175 0.105 34.345 0.275 ;
      RECT 34.175 8.605 34.345 8.775 ;
      RECT 34.105 2.765 34.275 2.935 ;
      RECT 34.105 5.945 34.275 6.115 ;
      RECT 32.895 1.565 33.065 1.735 ;
      RECT 32.895 4.285 33.065 4.455 ;
      RECT 32.435 1.565 32.605 1.735 ;
      RECT 32.435 4.285 32.605 4.455 ;
      RECT 32.04 2.905 32.21 3.075 ;
      RECT 31.975 1.565 32.145 1.735 ;
      RECT 31.975 4.285 32.145 4.455 ;
      RECT 31.83 2.245 32 2.415 ;
      RECT 31.515 1.565 31.685 1.735 ;
      RECT 31.515 3.155 31.685 3.325 ;
      RECT 31.515 4.285 31.685 4.455 ;
      RECT 31.455 4.545 31.625 4.715 ;
      RECT 31.455 8.605 31.625 8.775 ;
      RECT 31.145 6.685 31.315 6.855 ;
      RECT 31.13 2.75 31.3 2.92 ;
      RECT 31.055 1.565 31.225 1.735 ;
      RECT 31.055 4.285 31.225 4.455 ;
      RECT 30.915 3.315 31.085 3.485 ;
      RECT 30.895 3.715 31.065 3.885 ;
      RECT 30.775 8.605 30.945 8.775 ;
      RECT 30.72 2.27 30.89 2.44 ;
      RECT 30.715 7.055 30.885 7.225 ;
      RECT 30.715 7.795 30.885 7.965 ;
      RECT 30.595 1.565 30.765 1.735 ;
      RECT 30.595 4.285 30.765 4.455 ;
      RECT 30.34 6.315 30.51 6.485 ;
      RECT 30.225 3.25 30.395 3.42 ;
      RECT 30.135 1.565 30.305 1.735 ;
      RECT 30.135 4.285 30.305 4.455 ;
      RECT 30.095 8.605 30.265 8.775 ;
      RECT 29.9 2.935 30.07 3.105 ;
      RECT 29.835 3.715 30.005 3.885 ;
      RECT 29.675 1.565 29.845 1.735 ;
      RECT 29.675 4.285 29.845 4.455 ;
      RECT 29.435 3.7 29.605 3.87 ;
      RECT 29.415 8.605 29.585 8.775 ;
      RECT 29.395 2.185 29.565 2.355 ;
      RECT 29.345 5.945 29.515 6.115 ;
      RECT 29.215 1.565 29.385 1.735 ;
      RECT 29.215 4.285 29.385 4.455 ;
      RECT 28.755 1.565 28.925 1.735 ;
      RECT 28.755 4.285 28.925 4.455 ;
      RECT 28.495 2.685 28.665 2.855 ;
      RECT 28.495 3.145 28.665 3.315 ;
      RECT 28.495 3.66 28.665 3.83 ;
      RECT 28.38 2.22 28.55 2.39 ;
      RECT 28.295 1.565 28.465 1.735 ;
      RECT 28.295 4.285 28.465 4.455 ;
      RECT 27.915 3.73 28.085 3.9 ;
      RECT 27.835 1.565 28.005 1.735 ;
      RECT 27.835 4.285 28.005 4.455 ;
      RECT 27.435 2.26 27.605 2.43 ;
      RECT 27.375 1.565 27.545 1.735 ;
      RECT 27.375 4.285 27.545 4.455 ;
      RECT 27.22 2.635 27.39 2.805 ;
      RECT 26.915 1.565 27.085 1.735 ;
      RECT 26.915 4.285 27.085 4.455 ;
      RECT 26.72 3.235 26.89 3.405 ;
      RECT 26.605 2.685 26.775 2.855 ;
      RECT 26.455 1.565 26.625 1.735 ;
      RECT 26.455 4.285 26.625 4.455 ;
      RECT 26.435 2.135 26.605 2.305 ;
      RECT 26.06 3.165 26.23 3.335 ;
      RECT 25.995 1.565 26.165 1.735 ;
      RECT 25.995 4.285 26.165 4.455 ;
      RECT 25.575 2.765 25.745 2.935 ;
      RECT 25.535 1.565 25.705 1.735 ;
      RECT 25.535 4.285 25.705 4.455 ;
      RECT 25.525 3.54 25.695 3.71 ;
      RECT 25.075 1.565 25.245 1.735 ;
      RECT 25.075 4.285 25.245 4.455 ;
      RECT 25.035 3.165 25.205 3.335 ;
      RECT 25 2.27 25.17 2.44 ;
      RECT 24.64 2.67 24.81 2.84 ;
      RECT 24.615 1.565 24.785 1.735 ;
      RECT 24.615 4.285 24.785 4.455 ;
      RECT 24.435 3.48 24.605 3.65 ;
      RECT 24.155 1.565 24.325 1.735 ;
      RECT 24.155 4.285 24.325 4.455 ;
      RECT 24.13 2.91 24.3 3.08 ;
      RECT 23.695 1.565 23.865 1.735 ;
      RECT 23.695 4.285 23.865 4.455 ;
      RECT 23.43 2.7 23.6 2.87 ;
      RECT 23.235 1.565 23.405 1.735 ;
      RECT 23.235 4.285 23.405 4.455 ;
      RECT 23.11 3.145 23.28 3.315 ;
      RECT 22.775 1.565 22.945 1.735 ;
      RECT 22.775 4.285 22.945 4.455 ;
      RECT 22.695 3.18 22.865 3.35 ;
      RECT 22.525 2.165 22.695 2.335 ;
      RECT 22.35 2.62 22.52 2.79 ;
      RECT 22.315 1.565 22.485 1.735 ;
      RECT 22.315 4.285 22.485 4.455 ;
      RECT 21.855 1.565 22.025 1.735 ;
      RECT 21.855 4.285 22.025 4.455 ;
      RECT 21.43 2.27 21.6 2.44 ;
      RECT 21.425 3.585 21.595 3.755 ;
      RECT 21.395 1.565 21.565 1.735 ;
      RECT 21.395 4.285 21.565 4.455 ;
      RECT 20.335 0.915 20.505 1.085 ;
      RECT 20.335 2.395 20.505 2.565 ;
      RECT 20.335 6.315 20.505 6.485 ;
      RECT 20.335 7.795 20.505 7.965 ;
      RECT 19.985 0.105 20.155 0.275 ;
      RECT 19.985 4.165 20.155 4.335 ;
      RECT 19.985 4.545 20.155 4.715 ;
      RECT 19.985 8.605 20.155 8.775 ;
      RECT 19.965 2.765 20.135 2.935 ;
      RECT 19.965 5.945 20.135 6.115 ;
      RECT 19.345 0.915 19.515 1.085 ;
      RECT 19.345 2.395 19.515 2.565 ;
      RECT 19.345 6.315 19.515 6.485 ;
      RECT 19.345 7.795 19.515 7.965 ;
      RECT 18.995 0.105 19.165 0.275 ;
      RECT 18.995 4.165 19.165 4.335 ;
      RECT 18.995 4.545 19.165 4.715 ;
      RECT 18.995 8.605 19.165 8.775 ;
      RECT 18.975 2.765 19.145 2.935 ;
      RECT 18.975 5.945 19.145 6.115 ;
      RECT 18.29 0.105 18.46 0.275 ;
      RECT 18.29 4.165 18.46 4.335 ;
      RECT 18.29 4.545 18.46 4.715 ;
      RECT 18.29 8.605 18.46 8.775 ;
      RECT 17.98 2.025 18.15 2.195 ;
      RECT 17.98 6.685 18.15 6.855 ;
      RECT 17.61 0.105 17.78 0.275 ;
      RECT 17.61 8.605 17.78 8.775 ;
      RECT 17.55 0.915 17.72 1.085 ;
      RECT 17.55 1.655 17.72 1.825 ;
      RECT 17.55 7.055 17.72 7.225 ;
      RECT 17.55 7.795 17.72 7.965 ;
      RECT 17.175 2.395 17.345 2.565 ;
      RECT 17.175 6.315 17.345 6.485 ;
      RECT 16.93 0.105 17.1 0.275 ;
      RECT 16.93 8.605 17.1 8.775 ;
      RECT 16.25 0.105 16.42 0.275 ;
      RECT 16.25 8.605 16.42 8.775 ;
      RECT 16.18 2.765 16.35 2.935 ;
      RECT 16.18 5.945 16.35 6.115 ;
      RECT 14.97 1.565 15.14 1.735 ;
      RECT 14.97 4.285 15.14 4.455 ;
      RECT 14.51 1.565 14.68 1.735 ;
      RECT 14.51 4.285 14.68 4.455 ;
      RECT 14.115 2.905 14.285 3.075 ;
      RECT 14.05 1.565 14.22 1.735 ;
      RECT 14.05 4.285 14.22 4.455 ;
      RECT 13.905 2.245 14.075 2.415 ;
      RECT 13.59 1.565 13.76 1.735 ;
      RECT 13.59 3.155 13.76 3.325 ;
      RECT 13.59 4.285 13.76 4.455 ;
      RECT 13.53 4.545 13.7 4.715 ;
      RECT 13.53 8.605 13.7 8.775 ;
      RECT 13.22 6.685 13.39 6.855 ;
      RECT 13.205 2.75 13.375 2.92 ;
      RECT 13.13 1.565 13.3 1.735 ;
      RECT 13.13 4.285 13.3 4.455 ;
      RECT 12.99 3.315 13.16 3.485 ;
      RECT 12.97 3.715 13.14 3.885 ;
      RECT 12.85 8.605 13.02 8.775 ;
      RECT 12.795 2.27 12.965 2.44 ;
      RECT 12.79 7.055 12.96 7.225 ;
      RECT 12.79 7.795 12.96 7.965 ;
      RECT 12.67 1.565 12.84 1.735 ;
      RECT 12.67 4.285 12.84 4.455 ;
      RECT 12.415 6.315 12.585 6.485 ;
      RECT 12.3 3.25 12.47 3.42 ;
      RECT 12.21 1.565 12.38 1.735 ;
      RECT 12.21 4.285 12.38 4.455 ;
      RECT 12.17 8.605 12.34 8.775 ;
      RECT 11.975 2.935 12.145 3.105 ;
      RECT 11.91 3.715 12.08 3.885 ;
      RECT 11.75 1.565 11.92 1.735 ;
      RECT 11.75 4.285 11.92 4.455 ;
      RECT 11.51 3.7 11.68 3.87 ;
      RECT 11.49 8.605 11.66 8.775 ;
      RECT 11.47 2.185 11.64 2.355 ;
      RECT 11.42 5.945 11.59 6.115 ;
      RECT 11.29 1.565 11.46 1.735 ;
      RECT 11.29 4.285 11.46 4.455 ;
      RECT 10.83 1.565 11 1.735 ;
      RECT 10.83 4.285 11 4.455 ;
      RECT 10.57 2.685 10.74 2.855 ;
      RECT 10.57 3.145 10.74 3.315 ;
      RECT 10.57 3.66 10.74 3.83 ;
      RECT 10.455 2.22 10.625 2.39 ;
      RECT 10.37 1.565 10.54 1.735 ;
      RECT 10.37 4.285 10.54 4.455 ;
      RECT 9.99 3.73 10.16 3.9 ;
      RECT 9.91 1.565 10.08 1.735 ;
      RECT 9.91 4.285 10.08 4.455 ;
      RECT 9.51 2.26 9.68 2.43 ;
      RECT 9.45 1.565 9.62 1.735 ;
      RECT 9.45 4.285 9.62 4.455 ;
      RECT 9.295 2.635 9.465 2.805 ;
      RECT 8.99 1.565 9.16 1.735 ;
      RECT 8.99 4.285 9.16 4.455 ;
      RECT 8.795 3.235 8.965 3.405 ;
      RECT 8.68 2.685 8.85 2.855 ;
      RECT 8.53 1.565 8.7 1.735 ;
      RECT 8.53 4.285 8.7 4.455 ;
      RECT 8.51 2.135 8.68 2.305 ;
      RECT 8.135 3.165 8.305 3.335 ;
      RECT 8.07 1.565 8.24 1.735 ;
      RECT 8.07 4.285 8.24 4.455 ;
      RECT 7.65 2.765 7.82 2.935 ;
      RECT 7.61 1.565 7.78 1.735 ;
      RECT 7.61 4.285 7.78 4.455 ;
      RECT 7.6 3.54 7.77 3.71 ;
      RECT 7.15 1.565 7.32 1.735 ;
      RECT 7.15 4.285 7.32 4.455 ;
      RECT 7.11 3.165 7.28 3.335 ;
      RECT 7.075 2.27 7.245 2.44 ;
      RECT 6.715 2.67 6.885 2.84 ;
      RECT 6.69 1.565 6.86 1.735 ;
      RECT 6.69 4.285 6.86 4.455 ;
      RECT 6.51 3.48 6.68 3.65 ;
      RECT 6.23 1.565 6.4 1.735 ;
      RECT 6.23 4.285 6.4 4.455 ;
      RECT 6.205 2.91 6.375 3.08 ;
      RECT 5.77 1.565 5.94 1.735 ;
      RECT 5.77 4.285 5.94 4.455 ;
      RECT 5.505 2.7 5.675 2.87 ;
      RECT 5.31 1.565 5.48 1.735 ;
      RECT 5.31 4.285 5.48 4.455 ;
      RECT 5.185 3.145 5.355 3.315 ;
      RECT 4.85 1.565 5.02 1.735 ;
      RECT 4.85 4.285 5.02 4.455 ;
      RECT 4.77 3.18 4.94 3.35 ;
      RECT 4.6 2.165 4.77 2.335 ;
      RECT 4.425 2.62 4.595 2.79 ;
      RECT 4.39 1.565 4.56 1.735 ;
      RECT 4.39 4.285 4.56 4.455 ;
      RECT 3.93 1.565 4.1 1.735 ;
      RECT 3.93 4.285 4.1 4.455 ;
      RECT 3.505 2.27 3.675 2.44 ;
      RECT 3.5 3.585 3.67 3.755 ;
      RECT 3.47 1.565 3.64 1.735 ;
      RECT 3.47 4.285 3.64 4.455 ;
      RECT 2.5 4.545 2.67 4.715 ;
      RECT 2.5 8.605 2.67 8.775 ;
      RECT 2.19 6.685 2.36 6.855 ;
      RECT 1.82 8.605 1.99 8.775 ;
      RECT 1.76 7.055 1.93 7.225 ;
      RECT 1.76 7.795 1.93 7.965 ;
      RECT 1.385 6.315 1.555 6.485 ;
      RECT 1.14 8.605 1.31 8.775 ;
      RECT 0.46 8.605 0.63 8.775 ;
      RECT 0.39 5.945 0.56 6.115 ;
    LAYER li ;
      RECT 86.075 0 86.245 2.235 ;
      RECT 85.115 0 85.285 2.235 ;
      RECT 84.155 0 84.325 2.235 ;
      RECT 83.635 0 83.805 2.235 ;
      RECT 82.675 0 82.845 2.235 ;
      RECT 81.675 0 81.845 2.235 ;
      RECT 80.715 0 80.885 2.235 ;
      RECT 79.235 0 79.405 2.235 ;
      RECT 77.315 0 77.485 2.235 ;
      RECT 75.835 0 76.005 2.235 ;
      RECT 68.15 0 68.32 2.235 ;
      RECT 67.19 0 67.36 2.235 ;
      RECT 66.23 0 66.4 2.235 ;
      RECT 65.71 0 65.88 2.235 ;
      RECT 64.75 0 64.92 2.235 ;
      RECT 63.75 0 63.92 2.235 ;
      RECT 62.79 0 62.96 2.235 ;
      RECT 61.31 0 61.48 2.235 ;
      RECT 59.39 0 59.56 2.235 ;
      RECT 57.91 0 58.08 2.235 ;
      RECT 50.225 0 50.395 2.235 ;
      RECT 49.265 0 49.435 2.235 ;
      RECT 48.305 0 48.475 2.235 ;
      RECT 47.785 0 47.955 2.235 ;
      RECT 46.825 0 46.995 2.235 ;
      RECT 45.825 0 45.995 2.235 ;
      RECT 44.865 0 45.035 2.235 ;
      RECT 43.385 0 43.555 2.235 ;
      RECT 41.465 0 41.635 2.235 ;
      RECT 39.985 0 40.155 2.235 ;
      RECT 32.3 0 32.47 2.235 ;
      RECT 31.34 0 31.51 2.235 ;
      RECT 30.38 0 30.55 2.235 ;
      RECT 29.86 0 30.03 2.235 ;
      RECT 28.9 0 29.07 2.235 ;
      RECT 27.9 0 28.07 2.235 ;
      RECT 26.94 0 27.11 2.235 ;
      RECT 25.46 0 25.63 2.235 ;
      RECT 23.54 0 23.71 2.235 ;
      RECT 22.06 0 22.23 2.235 ;
      RECT 14.375 0 14.545 2.235 ;
      RECT 13.415 0 13.585 2.235 ;
      RECT 12.455 0 12.625 2.235 ;
      RECT 11.935 0 12.105 2.235 ;
      RECT 10.975 0 11.145 2.235 ;
      RECT 9.975 0 10.145 2.235 ;
      RECT 9.015 0 9.185 2.235 ;
      RECT 7.535 0 7.705 2.235 ;
      RECT 5.615 0 5.785 2.235 ;
      RECT 4.135 0 4.305 2.235 ;
      RECT 75.025 0 86.985 1.735 ;
      RECT 57.1 0 69.06 1.735 ;
      RECT 39.175 0 51.135 1.735 ;
      RECT 21.25 0 33.21 1.735 ;
      RECT 3.325 0 15.285 1.735 ;
      RECT 75.02 0 86.985 1.68 ;
      RECT 57.095 0 69.06 1.68 ;
      RECT 39.17 0 51.135 1.68 ;
      RECT 21.245 0 33.21 1.68 ;
      RECT 3.32 0 15.285 1.68 ;
      RECT 91.605 0 91.775 0.935 ;
      RECT 90.615 0 90.785 0.935 ;
      RECT 87.87 0 88.04 0.935 ;
      RECT 73.68 0 73.85 0.935 ;
      RECT 72.69 0 72.86 0.935 ;
      RECT 69.945 0 70.115 0.935 ;
      RECT 55.755 0 55.925 0.935 ;
      RECT 54.765 0 54.935 0.935 ;
      RECT 52.02 0 52.19 0.935 ;
      RECT 37.83 0 38 0.935 ;
      RECT 36.84 0 37.01 0.935 ;
      RECT 34.095 0 34.265 0.935 ;
      RECT 19.905 0 20.075 0.935 ;
      RECT 18.915 0 19.085 0.935 ;
      RECT 16.17 0 16.34 0.935 ;
      RECT 0 0 92.575 0.305 ;
      RECT 2.19 4.285 2.36 8.305 ;
      RECT 91.605 3.405 91.775 5.475 ;
      RECT 90.615 3.405 90.785 5.475 ;
      RECT 87.87 3.405 88.04 5.475 ;
      RECT 83.11 4.285 83.28 5.475 ;
      RECT 73.68 3.405 73.85 5.475 ;
      RECT 72.69 3.405 72.86 5.475 ;
      RECT 69.945 3.405 70.115 5.475 ;
      RECT 65.185 4.285 65.355 5.475 ;
      RECT 55.755 3.405 55.925 5.475 ;
      RECT 54.765 3.405 54.935 5.475 ;
      RECT 52.02 3.405 52.19 5.475 ;
      RECT 47.26 4.285 47.43 5.475 ;
      RECT 37.83 3.405 38 5.475 ;
      RECT 36.84 3.405 37.01 5.475 ;
      RECT 34.095 3.405 34.265 5.475 ;
      RECT 29.335 4.285 29.505 5.475 ;
      RECT 19.905 3.405 20.075 5.475 ;
      RECT 18.915 3.405 19.085 5.475 ;
      RECT 16.17 3.405 16.34 5.475 ;
      RECT 11.41 4.285 11.58 5.475 ;
      RECT 0.38 4.285 0.55 5.475 ;
      RECT 0 4.285 92.575 4.745 ;
      RECT 86.615 4.135 92.575 4.745 ;
      RECT 85.115 3.785 85.285 4.745 ;
      RECT 82.675 3.785 82.845 4.745 ;
      RECT 80.715 3.785 80.885 4.745 ;
      RECT 79.755 3.785 79.925 4.745 ;
      RECT 77.795 3.785 77.965 4.745 ;
      RECT 76.795 3.785 76.965 4.745 ;
      RECT 75.835 3.785 76.005 4.745 ;
      RECT 68.69 4.135 74.65 4.745 ;
      RECT 67.19 3.785 67.36 4.745 ;
      RECT 64.75 3.785 64.92 4.745 ;
      RECT 62.79 3.785 62.96 4.745 ;
      RECT 61.83 3.785 62 4.745 ;
      RECT 59.87 3.785 60.04 4.745 ;
      RECT 58.87 3.785 59.04 4.745 ;
      RECT 57.91 3.785 58.08 4.745 ;
      RECT 50.765 4.135 56.725 4.745 ;
      RECT 49.265 3.785 49.435 4.745 ;
      RECT 46.825 3.785 46.995 4.745 ;
      RECT 44.865 3.785 45.035 4.745 ;
      RECT 43.905 3.785 44.075 4.745 ;
      RECT 41.945 3.785 42.115 4.745 ;
      RECT 40.945 3.785 41.115 4.745 ;
      RECT 39.985 3.785 40.155 4.745 ;
      RECT 32.84 4.135 38.8 4.745 ;
      RECT 31.34 3.785 31.51 4.745 ;
      RECT 28.9 3.785 29.07 4.745 ;
      RECT 26.94 3.785 27.11 4.745 ;
      RECT 25.98 3.785 26.15 4.745 ;
      RECT 24.02 3.785 24.19 4.745 ;
      RECT 23.02 3.785 23.19 4.745 ;
      RECT 22.06 3.785 22.23 4.745 ;
      RECT 14.915 4.135 20.875 4.745 ;
      RECT 13.415 3.785 13.585 4.745 ;
      RECT 10.975 3.785 11.145 4.745 ;
      RECT 9.015 3.785 9.185 4.745 ;
      RECT 8.055 3.785 8.225 4.745 ;
      RECT 6.095 3.785 6.265 4.745 ;
      RECT 5.095 3.785 5.265 4.745 ;
      RECT 4.135 3.785 4.305 4.745 ;
      RECT 0 8.575 92.575 8.88 ;
      RECT 91.605 7.945 91.775 8.88 ;
      RECT 90.615 7.945 90.785 8.88 ;
      RECT 87.87 7.945 88.04 8.88 ;
      RECT 83.11 7.945 83.28 8.88 ;
      RECT 73.68 7.945 73.85 8.88 ;
      RECT 72.69 7.945 72.86 8.88 ;
      RECT 69.945 7.945 70.115 8.88 ;
      RECT 65.185 7.945 65.355 8.88 ;
      RECT 55.755 7.945 55.925 8.88 ;
      RECT 54.765 7.945 54.935 8.88 ;
      RECT 52.02 7.945 52.19 8.88 ;
      RECT 47.26 7.945 47.43 8.88 ;
      RECT 37.83 7.945 38 8.88 ;
      RECT 36.84 7.945 37.01 8.88 ;
      RECT 34.095 7.945 34.265 8.88 ;
      RECT 29.335 7.945 29.505 8.88 ;
      RECT 19.905 7.945 20.075 8.88 ;
      RECT 18.915 7.945 19.085 8.88 ;
      RECT 16.17 7.945 16.34 8.88 ;
      RECT 11.41 7.945 11.58 8.88 ;
      RECT 0.38 7.945 0.55 8.88 ;
      RECT 91.665 1.74 91.835 2.935 ;
      RECT 91.665 1.74 92.13 1.91 ;
      RECT 91.665 6.97 92.13 7.14 ;
      RECT 91.665 5.945 91.835 7.14 ;
      RECT 90.675 1.74 90.845 2.935 ;
      RECT 90.675 1.74 91.14 1.91 ;
      RECT 90.675 6.97 91.14 7.14 ;
      RECT 90.675 5.945 90.845 7.14 ;
      RECT 88.82 2.635 88.99 3.865 ;
      RECT 88.875 0.855 89.045 2.805 ;
      RECT 88.82 0.575 88.99 1.025 ;
      RECT 88.82 7.855 88.99 8.305 ;
      RECT 88.875 6.075 89.045 8.025 ;
      RECT 88.82 5.015 88.99 6.245 ;
      RECT 88.3 0.575 88.47 3.865 ;
      RECT 88.3 2.075 88.705 2.405 ;
      RECT 88.3 1.235 88.705 1.565 ;
      RECT 88.3 5.015 88.47 8.305 ;
      RECT 88.3 7.315 88.705 7.645 ;
      RECT 88.3 6.475 88.705 6.805 ;
      RECT 86.4 3.392 86.415 3.443 ;
      RECT 86.395 3.372 86.4 3.49 ;
      RECT 86.38 3.362 86.395 3.558 ;
      RECT 86.355 3.342 86.38 3.613 ;
      RECT 86.315 3.327 86.355 3.633 ;
      RECT 86.27 3.321 86.315 3.661 ;
      RECT 86.2 3.311 86.27 3.678 ;
      RECT 86.18 3.303 86.2 3.678 ;
      RECT 86.12 3.297 86.18 3.67 ;
      RECT 86.061 3.288 86.12 3.658 ;
      RECT 85.975 3.277 86.061 3.641 ;
      RECT 85.953 3.268 85.975 3.629 ;
      RECT 85.867 3.261 85.953 3.616 ;
      RECT 85.781 3.248 85.867 3.597 ;
      RECT 85.695 3.236 85.781 3.577 ;
      RECT 85.665 3.225 85.695 3.564 ;
      RECT 85.615 3.211 85.665 3.556 ;
      RECT 85.595 3.2 85.615 3.548 ;
      RECT 85.546 3.189 85.595 3.54 ;
      RECT 85.46 3.168 85.546 3.525 ;
      RECT 85.415 3.155 85.46 3.51 ;
      RECT 85.37 3.155 85.415 3.49 ;
      RECT 85.315 3.155 85.37 3.425 ;
      RECT 85.29 3.155 85.315 3.348 ;
      RECT 85.815 2.892 85.985 3.075 ;
      RECT 85.815 2.892 86 3.033 ;
      RECT 85.815 2.892 86.005 2.975 ;
      RECT 85.875 2.66 86.01 2.951 ;
      RECT 85.875 2.664 86.015 2.934 ;
      RECT 85.82 2.827 86.015 2.934 ;
      RECT 85.845 2.672 85.985 3.075 ;
      RECT 85.845 2.676 86.025 2.875 ;
      RECT 85.83 2.762 86.025 2.875 ;
      RECT 85.84 2.692 85.985 3.075 ;
      RECT 85.84 2.695 86.035 2.788 ;
      RECT 85.835 2.712 86.035 2.788 ;
      RECT 85.605 1.932 85.775 2.415 ;
      RECT 85.6 1.927 85.75 2.405 ;
      RECT 85.6 1.934 85.78 2.399 ;
      RECT 85.59 1.928 85.75 2.378 ;
      RECT 85.59 1.944 85.795 2.337 ;
      RECT 85.56 1.929 85.75 2.3 ;
      RECT 85.56 1.959 85.805 2.24 ;
      RECT 85.555 1.931 85.75 2.238 ;
      RECT 85.535 1.94 85.78 2.195 ;
      RECT 85.51 1.956 85.795 2.107 ;
      RECT 85.51 1.975 85.82 2.098 ;
      RECT 85.505 2.012 85.82 2.05 ;
      RECT 85.51 1.992 85.825 2.018 ;
      RECT 85.605 1.926 85.715 2.415 ;
      RECT 85.691 1.925 85.715 2.415 ;
      RECT 84.925 2.71 84.93 2.921 ;
      RECT 85.525 2.71 85.53 2.895 ;
      RECT 85.59 2.75 85.595 2.863 ;
      RECT 85.585 2.742 85.59 2.869 ;
      RECT 85.58 2.732 85.585 2.877 ;
      RECT 85.575 2.722 85.58 2.886 ;
      RECT 85.57 2.712 85.575 2.89 ;
      RECT 85.53 2.71 85.57 2.893 ;
      RECT 85.502 2.709 85.525 2.897 ;
      RECT 85.416 2.706 85.502 2.904 ;
      RECT 85.33 2.702 85.416 2.915 ;
      RECT 85.31 2.7 85.33 2.921 ;
      RECT 85.292 2.699 85.31 2.924 ;
      RECT 85.206 2.697 85.292 2.931 ;
      RECT 85.12 2.692 85.206 2.944 ;
      RECT 85.101 2.689 85.12 2.949 ;
      RECT 85.015 2.687 85.101 2.94 ;
      RECT 85.005 2.687 85.015 2.933 ;
      RECT 84.93 2.7 85.005 2.927 ;
      RECT 84.915 2.711 84.925 2.921 ;
      RECT 84.905 2.713 84.915 2.92 ;
      RECT 84.895 2.717 84.905 2.916 ;
      RECT 84.89 2.72 84.895 2.91 ;
      RECT 84.88 2.722 84.89 2.904 ;
      RECT 84.875 2.725 84.88 2.898 ;
      RECT 84.855 3.311 84.86 3.515 ;
      RECT 84.84 3.298 84.855 3.608 ;
      RECT 84.825 3.279 84.84 3.885 ;
      RECT 84.79 3.245 84.825 3.885 ;
      RECT 84.786 3.215 84.79 3.885 ;
      RECT 84.7 3.097 84.786 3.885 ;
      RECT 84.69 2.972 84.7 3.885 ;
      RECT 84.675 2.94 84.69 3.885 ;
      RECT 84.67 2.915 84.675 3.885 ;
      RECT 84.665 2.905 84.67 3.841 ;
      RECT 84.65 2.877 84.665 3.746 ;
      RECT 84.635 2.843 84.65 3.645 ;
      RECT 84.63 2.821 84.635 3.598 ;
      RECT 84.625 2.81 84.63 3.568 ;
      RECT 84.62 2.8 84.625 3.534 ;
      RECT 84.61 2.787 84.62 3.502 ;
      RECT 84.585 2.763 84.61 3.428 ;
      RECT 84.58 2.743 84.585 3.353 ;
      RECT 84.575 2.737 84.58 3.328 ;
      RECT 84.57 2.732 84.575 3.293 ;
      RECT 84.565 2.727 84.57 3.268 ;
      RECT 84.56 2.725 84.565 3.248 ;
      RECT 84.555 2.725 84.56 3.233 ;
      RECT 84.55 2.725 84.555 3.193 ;
      RECT 84.54 2.725 84.55 3.165 ;
      RECT 84.53 2.725 84.54 3.11 ;
      RECT 84.515 2.725 84.53 3.048 ;
      RECT 84.51 2.724 84.515 2.993 ;
      RECT 84.495 2.723 84.51 2.973 ;
      RECT 84.435 2.721 84.495 2.947 ;
      RECT 84.4 2.722 84.435 2.927 ;
      RECT 84.395 2.724 84.4 2.917 ;
      RECT 84.385 2.743 84.395 2.907 ;
      RECT 84.38 2.77 84.385 2.838 ;
      RECT 84.495 2.195 84.665 2.44 ;
      RECT 84.53 1.966 84.665 2.44 ;
      RECT 84.53 1.968 84.675 2.435 ;
      RECT 84.53 1.97 84.7 2.423 ;
      RECT 84.53 1.973 84.725 2.405 ;
      RECT 84.53 1.978 84.775 2.378 ;
      RECT 84.53 1.983 84.795 2.343 ;
      RECT 84.51 1.985 84.805 2.318 ;
      RECT 84.5 2.08 84.805 2.318 ;
      RECT 84.53 1.965 84.64 2.44 ;
      RECT 84.54 1.962 84.635 2.44 ;
      RECT 84.06 3.227 84.25 3.585 ;
      RECT 84.06 3.239 84.285 3.584 ;
      RECT 84.06 3.267 84.305 3.582 ;
      RECT 84.06 3.292 84.31 3.581 ;
      RECT 84.06 3.35 84.325 3.58 ;
      RECT 84.045 3.223 84.205 3.565 ;
      RECT 84.025 3.232 84.25 3.518 ;
      RECT 84 3.243 84.285 3.455 ;
      RECT 84 3.327 84.32 3.455 ;
      RECT 84 3.302 84.315 3.455 ;
      RECT 84.06 3.218 84.205 3.585 ;
      RECT 84.146 3.217 84.205 3.585 ;
      RECT 84.146 3.216 84.19 3.585 ;
      RECT 84.06 7.855 84.23 8.305 ;
      RECT 84.115 6.075 84.285 8.025 ;
      RECT 84.06 5.015 84.23 6.245 ;
      RECT 83.54 5.015 83.71 8.305 ;
      RECT 83.54 7.315 83.945 7.645 ;
      RECT 83.54 6.475 83.945 6.805 ;
      RECT 83.845 2.732 83.85 3.11 ;
      RECT 83.84 2.7 83.845 3.11 ;
      RECT 83.835 2.672 83.84 3.11 ;
      RECT 83.83 2.652 83.835 3.11 ;
      RECT 83.775 2.635 83.83 3.11 ;
      RECT 83.735 2.62 83.775 3.11 ;
      RECT 83.68 2.607 83.735 3.11 ;
      RECT 83.645 2.598 83.68 3.11 ;
      RECT 83.641 2.596 83.645 3.109 ;
      RECT 83.555 2.592 83.641 3.092 ;
      RECT 83.47 2.584 83.555 3.055 ;
      RECT 83.46 2.58 83.47 3.028 ;
      RECT 83.45 2.58 83.46 3.01 ;
      RECT 83.44 2.582 83.45 2.993 ;
      RECT 83.435 2.587 83.44 2.979 ;
      RECT 83.43 2.591 83.435 2.966 ;
      RECT 83.42 2.596 83.43 2.95 ;
      RECT 83.405 2.61 83.42 2.925 ;
      RECT 83.4 2.616 83.405 2.905 ;
      RECT 83.395 2.618 83.4 2.898 ;
      RECT 83.39 2.622 83.395 2.773 ;
      RECT 83.57 3.422 83.815 3.885 ;
      RECT 83.49 3.395 83.81 3.881 ;
      RECT 83.42 3.43 83.815 3.874 ;
      RECT 83.21 3.685 83.815 3.87 ;
      RECT 83.39 3.453 83.815 3.87 ;
      RECT 83.23 3.645 83.815 3.87 ;
      RECT 83.38 3.465 83.815 3.87 ;
      RECT 83.265 3.582 83.815 3.87 ;
      RECT 83.32 3.507 83.815 3.87 ;
      RECT 83.57 3.372 83.81 3.885 ;
      RECT 83.6 3.365 83.81 3.885 ;
      RECT 83.59 3.367 83.81 3.885 ;
      RECT 83.6 3.362 83.73 3.885 ;
      RECT 83.155 1.925 83.241 2.364 ;
      RECT 83.15 1.925 83.241 2.362 ;
      RECT 83.15 1.925 83.31 2.361 ;
      RECT 83.15 1.925 83.34 2.358 ;
      RECT 83.135 1.932 83.34 2.349 ;
      RECT 83.135 1.932 83.345 2.345 ;
      RECT 83.13 1.942 83.345 2.338 ;
      RECT 83.125 1.947 83.345 2.313 ;
      RECT 83.125 1.947 83.36 2.295 ;
      RECT 83.15 1.925 83.38 2.21 ;
      RECT 83.12 1.952 83.38 2.208 ;
      RECT 83.13 1.945 83.385 2.146 ;
      RECT 83.12 2.067 83.39 2.129 ;
      RECT 83.105 1.962 83.385 2.08 ;
      RECT 83.1 1.972 83.385 1.98 ;
      RECT 83.18 2.743 83.185 2.82 ;
      RECT 83.17 2.737 83.18 3.01 ;
      RECT 83.16 2.729 83.17 3.031 ;
      RECT 83.15 2.72 83.16 3.053 ;
      RECT 83.145 2.715 83.15 3.07 ;
      RECT 83.105 2.715 83.145 3.11 ;
      RECT 83.085 2.715 83.105 3.165 ;
      RECT 83.08 2.715 83.085 3.193 ;
      RECT 83.07 2.715 83.08 3.208 ;
      RECT 83.035 2.715 83.07 3.25 ;
      RECT 83.03 2.715 83.035 3.293 ;
      RECT 83.02 2.715 83.03 3.308 ;
      RECT 83.005 2.715 83.02 3.328 ;
      RECT 82.99 2.715 83.005 3.355 ;
      RECT 82.985 2.716 82.99 3.373 ;
      RECT 82.965 2.717 82.985 3.38 ;
      RECT 82.91 2.718 82.965 3.4 ;
      RECT 82.9 2.719 82.91 3.414 ;
      RECT 82.895 2.722 82.9 3.413 ;
      RECT 82.855 2.795 82.895 3.411 ;
      RECT 82.84 2.875 82.855 3.409 ;
      RECT 82.815 2.93 82.84 3.407 ;
      RECT 82.8 2.995 82.815 3.406 ;
      RECT 82.755 3.027 82.8 3.403 ;
      RECT 82.67 3.05 82.755 3.398 ;
      RECT 82.645 3.07 82.67 3.393 ;
      RECT 82.575 3.075 82.645 3.389 ;
      RECT 82.555 3.077 82.575 3.386 ;
      RECT 82.47 3.088 82.555 3.38 ;
      RECT 82.465 3.099 82.47 3.375 ;
      RECT 82.455 3.101 82.465 3.375 ;
      RECT 82.42 3.105 82.455 3.373 ;
      RECT 82.37 3.115 82.42 3.36 ;
      RECT 82.35 3.123 82.37 3.345 ;
      RECT 82.27 3.135 82.35 3.328 ;
      RECT 82.435 2.685 82.605 2.895 ;
      RECT 82.551 2.681 82.605 2.895 ;
      RECT 82.356 2.685 82.605 2.886 ;
      RECT 82.356 2.685 82.61 2.875 ;
      RECT 82.27 2.685 82.61 2.866 ;
      RECT 82.27 2.693 82.62 2.81 ;
      RECT 82.27 2.705 82.625 2.723 ;
      RECT 82.27 2.712 82.63 2.715 ;
      RECT 82.465 2.683 82.605 2.895 ;
      RECT 82.22 3.628 82.465 3.96 ;
      RECT 82.215 3.62 82.22 3.957 ;
      RECT 82.185 3.64 82.465 3.938 ;
      RECT 82.165 3.672 82.465 3.911 ;
      RECT 82.215 3.625 82.392 3.957 ;
      RECT 82.215 3.622 82.306 3.957 ;
      RECT 82.155 1.97 82.325 2.39 ;
      RECT 82.15 1.97 82.325 2.388 ;
      RECT 82.15 1.97 82.35 2.378 ;
      RECT 82.15 1.97 82.37 2.353 ;
      RECT 82.145 1.97 82.37 2.348 ;
      RECT 82.145 1.97 82.38 2.338 ;
      RECT 82.145 1.97 82.385 2.333 ;
      RECT 82.145 1.975 82.39 2.328 ;
      RECT 82.145 2.007 82.405 2.318 ;
      RECT 82.145 2.077 82.43 2.301 ;
      RECT 82.125 2.077 82.43 2.293 ;
      RECT 82.125 2.137 82.44 2.27 ;
      RECT 82.125 2.177 82.45 2.215 ;
      RECT 82.11 1.97 82.385 2.195 ;
      RECT 82.1 1.985 82.39 2.093 ;
      RECT 81.69 3.375 81.86 3.9 ;
      RECT 81.685 3.375 81.86 3.893 ;
      RECT 81.675 3.375 81.865 3.858 ;
      RECT 81.67 3.385 81.865 3.83 ;
      RECT 81.665 3.405 81.865 3.813 ;
      RECT 81.675 3.38 81.87 3.803 ;
      RECT 81.66 3.425 81.87 3.795 ;
      RECT 81.655 3.445 81.87 3.78 ;
      RECT 81.65 3.475 81.87 3.77 ;
      RECT 81.64 3.52 81.87 3.745 ;
      RECT 81.67 3.39 81.875 3.728 ;
      RECT 81.635 3.572 81.875 3.723 ;
      RECT 81.67 3.4 81.88 3.693 ;
      RECT 81.63 3.605 81.88 3.69 ;
      RECT 81.625 3.63 81.88 3.67 ;
      RECT 81.665 3.417 81.89 3.61 ;
      RECT 81.66 3.439 81.9 3.503 ;
      RECT 81.61 2.686 81.625 2.955 ;
      RECT 81.565 2.67 81.61 3 ;
      RECT 81.56 2.658 81.565 3.05 ;
      RECT 81.55 2.654 81.56 3.083 ;
      RECT 81.545 2.651 81.55 3.111 ;
      RECT 81.53 2.653 81.545 3.153 ;
      RECT 81.525 2.657 81.53 3.193 ;
      RECT 81.505 2.662 81.525 3.245 ;
      RECT 81.501 2.667 81.505 3.302 ;
      RECT 81.415 2.686 81.501 3.339 ;
      RECT 81.405 2.707 81.415 3.375 ;
      RECT 81.4 2.715 81.405 3.376 ;
      RECT 81.395 2.757 81.4 3.377 ;
      RECT 81.38 2.845 81.395 3.378 ;
      RECT 81.37 2.995 81.38 3.38 ;
      RECT 81.365 3.04 81.37 3.382 ;
      RECT 81.33 3.082 81.365 3.385 ;
      RECT 81.325 3.1 81.33 3.388 ;
      RECT 81.248 3.106 81.325 3.394 ;
      RECT 81.162 3.12 81.248 3.407 ;
      RECT 81.076 3.134 81.162 3.421 ;
      RECT 80.99 3.148 81.076 3.434 ;
      RECT 80.93 3.16 80.99 3.446 ;
      RECT 80.905 3.167 80.93 3.453 ;
      RECT 80.891 3.17 80.905 3.458 ;
      RECT 80.805 3.178 80.891 3.474 ;
      RECT 80.8 3.185 80.805 3.489 ;
      RECT 80.776 3.185 80.8 3.496 ;
      RECT 80.69 3.188 80.776 3.524 ;
      RECT 80.605 3.192 80.69 3.568 ;
      RECT 80.54 3.196 80.605 3.605 ;
      RECT 80.515 3.199 80.54 3.621 ;
      RECT 80.44 3.212 80.515 3.625 ;
      RECT 80.415 3.23 80.44 3.629 ;
      RECT 80.405 3.237 80.415 3.631 ;
      RECT 80.39 3.24 80.405 3.632 ;
      RECT 80.33 3.252 80.39 3.636 ;
      RECT 80.32 3.266 80.33 3.64 ;
      RECT 80.265 3.276 80.32 3.628 ;
      RECT 80.24 3.297 80.265 3.611 ;
      RECT 80.22 3.317 80.24 3.602 ;
      RECT 80.215 3.33 80.22 3.597 ;
      RECT 80.2 3.342 80.215 3.593 ;
      RECT 81.435 1.997 81.44 2.02 ;
      RECT 81.43 1.988 81.435 2.06 ;
      RECT 81.425 1.986 81.43 2.103 ;
      RECT 81.42 1.977 81.425 2.138 ;
      RECT 81.415 1.967 81.42 2.21 ;
      RECT 81.41 1.957 81.415 2.275 ;
      RECT 81.405 1.954 81.41 2.315 ;
      RECT 81.38 1.948 81.405 2.405 ;
      RECT 81.345 1.936 81.38 2.43 ;
      RECT 81.335 1.927 81.345 2.43 ;
      RECT 81.2 1.925 81.21 2.413 ;
      RECT 81.19 1.925 81.2 2.38 ;
      RECT 81.185 1.925 81.19 2.355 ;
      RECT 81.18 1.925 81.185 2.343 ;
      RECT 81.175 1.925 81.18 2.325 ;
      RECT 81.165 1.925 81.175 2.29 ;
      RECT 81.16 1.927 81.165 2.268 ;
      RECT 81.155 1.933 81.16 2.253 ;
      RECT 81.15 1.939 81.155 2.238 ;
      RECT 81.135 1.951 81.15 2.211 ;
      RECT 81.13 1.962 81.135 2.179 ;
      RECT 81.125 1.972 81.13 2.163 ;
      RECT 81.115 1.98 81.125 2.132 ;
      RECT 81.11 1.99 81.115 2.106 ;
      RECT 81.105 2.047 81.11 2.089 ;
      RECT 81.21 1.925 81.335 2.43 ;
      RECT 80.925 2.612 81.185 2.91 ;
      RECT 80.92 2.619 81.185 2.908 ;
      RECT 80.925 2.614 81.2 2.903 ;
      RECT 80.915 2.627 81.2 2.9 ;
      RECT 80.915 2.632 81.205 2.893 ;
      RECT 80.91 2.64 81.205 2.89 ;
      RECT 80.91 2.657 81.21 2.688 ;
      RECT 80.925 2.609 81.156 2.91 ;
      RECT 80.98 2.608 81.156 2.91 ;
      RECT 80.98 2.605 81.07 2.91 ;
      RECT 80.98 2.602 81.066 2.91 ;
      RECT 80.67 2.875 80.675 2.888 ;
      RECT 80.665 2.842 80.67 2.893 ;
      RECT 80.66 2.797 80.665 2.9 ;
      RECT 80.655 2.752 80.66 2.908 ;
      RECT 80.65 2.72 80.655 2.916 ;
      RECT 80.645 2.68 80.65 2.917 ;
      RECT 80.63 2.66 80.645 2.919 ;
      RECT 80.555 2.642 80.63 2.931 ;
      RECT 80.545 2.635 80.555 2.942 ;
      RECT 80.54 2.635 80.545 2.944 ;
      RECT 80.51 2.641 80.54 2.948 ;
      RECT 80.47 2.654 80.51 2.948 ;
      RECT 80.445 2.665 80.47 2.934 ;
      RECT 80.43 2.671 80.445 2.917 ;
      RECT 80.42 2.673 80.43 2.908 ;
      RECT 80.415 2.674 80.42 2.903 ;
      RECT 80.41 2.675 80.415 2.898 ;
      RECT 80.405 2.676 80.41 2.895 ;
      RECT 80.38 2.681 80.405 2.885 ;
      RECT 80.37 2.697 80.38 2.872 ;
      RECT 80.365 2.717 80.37 2.867 ;
      RECT 80.375 2.11 80.38 2.306 ;
      RECT 80.36 2.074 80.375 2.308 ;
      RECT 80.35 2.056 80.36 2.313 ;
      RECT 80.34 2.042 80.35 2.317 ;
      RECT 80.295 2.026 80.34 2.327 ;
      RECT 80.29 2.016 80.295 2.336 ;
      RECT 80.245 2.005 80.29 2.342 ;
      RECT 80.24 1.993 80.245 2.349 ;
      RECT 80.225 1.988 80.24 2.353 ;
      RECT 80.21 1.98 80.225 2.358 ;
      RECT 80.2 1.973 80.21 2.363 ;
      RECT 80.19 1.97 80.2 2.368 ;
      RECT 80.18 1.97 80.19 2.369 ;
      RECT 80.175 1.967 80.18 2.368 ;
      RECT 80.14 1.962 80.165 2.367 ;
      RECT 80.116 1.958 80.14 2.366 ;
      RECT 80.03 1.949 80.116 2.363 ;
      RECT 80.015 1.941 80.03 2.36 ;
      RECT 79.993 1.94 80.015 2.359 ;
      RECT 79.907 1.94 79.993 2.357 ;
      RECT 79.821 1.94 79.907 2.355 ;
      RECT 79.735 1.94 79.821 2.352 ;
      RECT 79.725 1.94 79.735 2.343 ;
      RECT 79.695 1.94 79.725 2.303 ;
      RECT 79.685 1.95 79.695 2.258 ;
      RECT 79.68 1.99 79.685 2.243 ;
      RECT 79.675 2.005 79.68 2.23 ;
      RECT 79.645 2.085 79.675 2.192 ;
      RECT 80.165 1.965 80.175 2.368 ;
      RECT 79.99 2.73 80.005 3.335 ;
      RECT 79.995 2.725 80.005 3.335 ;
      RECT 80.16 2.725 80.165 2.908 ;
      RECT 80.15 2.725 80.16 2.938 ;
      RECT 80.135 2.725 80.15 2.998 ;
      RECT 80.13 2.725 80.135 3.043 ;
      RECT 80.125 2.725 80.13 3.073 ;
      RECT 80.12 2.725 80.125 3.093 ;
      RECT 80.11 2.725 80.12 3.128 ;
      RECT 80.095 2.725 80.11 3.16 ;
      RECT 80.05 2.725 80.095 3.188 ;
      RECT 80.045 2.725 80.05 3.218 ;
      RECT 80.04 2.725 80.045 3.23 ;
      RECT 80.035 2.725 80.04 3.238 ;
      RECT 80.025 2.725 80.035 3.253 ;
      RECT 80.02 2.725 80.025 3.275 ;
      RECT 80.01 2.725 80.02 3.298 ;
      RECT 80.005 2.725 80.01 3.318 ;
      RECT 79.97 2.74 79.99 3.335 ;
      RECT 79.945 2.757 79.97 3.335 ;
      RECT 79.94 2.767 79.945 3.335 ;
      RECT 79.91 2.782 79.94 3.335 ;
      RECT 79.835 2.824 79.91 3.335 ;
      RECT 79.83 2.855 79.835 3.318 ;
      RECT 79.825 2.859 79.83 3.3 ;
      RECT 79.82 2.863 79.825 3.263 ;
      RECT 79.815 3.047 79.82 3.23 ;
      RECT 79.3 3.236 79.386 3.801 ;
      RECT 79.255 3.238 79.42 3.795 ;
      RECT 79.386 3.235 79.42 3.795 ;
      RECT 79.3 3.237 79.505 3.789 ;
      RECT 79.255 3.247 79.515 3.785 ;
      RECT 79.23 3.239 79.505 3.781 ;
      RECT 79.225 3.242 79.505 3.776 ;
      RECT 79.2 3.257 79.515 3.77 ;
      RECT 79.2 3.282 79.555 3.765 ;
      RECT 79.16 3.29 79.555 3.74 ;
      RECT 79.16 3.317 79.57 3.738 ;
      RECT 79.16 3.347 79.58 3.725 ;
      RECT 79.155 3.492 79.58 3.713 ;
      RECT 79.16 3.421 79.6 3.71 ;
      RECT 79.16 3.478 79.605 3.518 ;
      RECT 79.35 2.757 79.52 2.935 ;
      RECT 79.3 2.696 79.35 2.92 ;
      RECT 79.035 2.676 79.3 2.905 ;
      RECT 78.995 2.74 79.47 2.905 ;
      RECT 78.995 2.73 79.425 2.905 ;
      RECT 78.995 2.727 79.415 2.905 ;
      RECT 78.995 2.715 79.405 2.905 ;
      RECT 78.995 2.7 79.35 2.905 ;
      RECT 79.035 2.672 79.236 2.905 ;
      RECT 79.045 2.65 79.236 2.905 ;
      RECT 79.07 2.635 79.15 2.905 ;
      RECT 78.825 3.165 78.945 3.61 ;
      RECT 78.81 3.165 78.945 3.609 ;
      RECT 78.765 3.187 78.945 3.604 ;
      RECT 78.725 3.236 78.945 3.598 ;
      RECT 78.725 3.236 78.95 3.573 ;
      RECT 78.725 3.236 78.97 3.463 ;
      RECT 78.72 3.266 78.97 3.46 ;
      RECT 78.81 3.165 78.98 3.355 ;
      RECT 78.47 1.95 78.475 2.395 ;
      RECT 78.28 1.95 78.3 2.36 ;
      RECT 78.25 1.95 78.255 2.335 ;
      RECT 78.93 2.257 78.945 2.445 ;
      RECT 78.925 2.242 78.93 2.451 ;
      RECT 78.905 2.215 78.925 2.454 ;
      RECT 78.855 2.182 78.905 2.463 ;
      RECT 78.825 2.162 78.855 2.467 ;
      RECT 78.806 2.15 78.825 2.463 ;
      RECT 78.72 2.122 78.806 2.453 ;
      RECT 78.71 2.097 78.72 2.443 ;
      RECT 78.64 2.065 78.71 2.435 ;
      RECT 78.615 2.025 78.64 2.427 ;
      RECT 78.595 2.007 78.615 2.421 ;
      RECT 78.585 1.997 78.595 2.418 ;
      RECT 78.575 1.99 78.585 2.416 ;
      RECT 78.555 1.977 78.575 2.413 ;
      RECT 78.545 1.967 78.555 2.41 ;
      RECT 78.535 1.96 78.545 2.408 ;
      RECT 78.485 1.952 78.535 2.402 ;
      RECT 78.475 1.95 78.485 2.396 ;
      RECT 78.445 1.95 78.47 2.393 ;
      RECT 78.416 1.95 78.445 2.388 ;
      RECT 78.33 1.95 78.416 2.378 ;
      RECT 78.3 1.95 78.33 2.365 ;
      RECT 78.255 1.95 78.28 2.348 ;
      RECT 78.24 1.95 78.25 2.33 ;
      RECT 78.22 1.957 78.24 2.315 ;
      RECT 78.215 1.972 78.22 2.303 ;
      RECT 78.21 1.977 78.215 2.243 ;
      RECT 78.205 1.982 78.21 2.085 ;
      RECT 78.2 1.985 78.205 2.003 ;
      RECT 78.465 2.67 78.551 2.991 ;
      RECT 78.465 2.67 78.585 2.984 ;
      RECT 78.415 2.67 78.585 2.98 ;
      RECT 78.415 2.672 78.671 2.978 ;
      RECT 78.415 2.674 78.695 2.972 ;
      RECT 78.415 2.681 78.705 2.971 ;
      RECT 78.415 2.69 78.71 2.968 ;
      RECT 78.415 2.696 78.715 2.963 ;
      RECT 78.415 2.74 78.72 2.96 ;
      RECT 78.415 2.832 78.725 2.957 ;
      RECT 77.94 3.275 77.975 3.595 ;
      RECT 78.525 3.46 78.53 3.642 ;
      RECT 78.48 3.342 78.525 3.661 ;
      RECT 78.465 3.319 78.48 3.684 ;
      RECT 78.455 3.309 78.465 3.694 ;
      RECT 78.435 3.304 78.455 3.707 ;
      RECT 78.41 3.302 78.435 3.728 ;
      RECT 78.391 3.301 78.41 3.74 ;
      RECT 78.305 3.298 78.391 3.74 ;
      RECT 78.235 3.293 78.305 3.728 ;
      RECT 78.16 3.289 78.235 3.703 ;
      RECT 78.095 3.285 78.16 3.67 ;
      RECT 78.025 3.282 78.095 3.63 ;
      RECT 77.995 3.278 78.025 3.605 ;
      RECT 77.975 3.276 77.995 3.598 ;
      RECT 77.891 3.274 77.94 3.596 ;
      RECT 77.805 3.271 77.891 3.597 ;
      RECT 77.73 3.27 77.805 3.599 ;
      RECT 77.645 3.27 77.73 3.625 ;
      RECT 77.568 3.271 77.645 3.65 ;
      RECT 77.482 3.272 77.568 3.65 ;
      RECT 77.396 3.272 77.482 3.65 ;
      RECT 77.31 3.273 77.396 3.65 ;
      RECT 77.29 3.274 77.31 3.642 ;
      RECT 77.275 3.28 77.29 3.627 ;
      RECT 77.24 3.3 77.275 3.607 ;
      RECT 77.23 3.32 77.24 3.589 ;
      RECT 78.2 2.625 78.205 2.895 ;
      RECT 78.195 2.616 78.2 2.9 ;
      RECT 78.185 2.606 78.195 2.912 ;
      RECT 78.18 2.595 78.185 2.923 ;
      RECT 78.16 2.589 78.18 2.941 ;
      RECT 78.115 2.586 78.16 2.99 ;
      RECT 78.1 2.585 78.115 3.035 ;
      RECT 78.095 2.585 78.1 3.048 ;
      RECT 78.085 2.585 78.095 3.06 ;
      RECT 78.08 2.586 78.085 3.075 ;
      RECT 78.06 2.594 78.08 3.08 ;
      RECT 78.03 2.61 78.06 3.08 ;
      RECT 78.02 2.622 78.025 3.08 ;
      RECT 77.985 2.637 78.02 3.08 ;
      RECT 77.955 2.657 77.985 3.08 ;
      RECT 77.945 2.682 77.955 3.08 ;
      RECT 77.94 2.71 77.945 3.08 ;
      RECT 77.935 2.74 77.94 3.08 ;
      RECT 77.93 2.757 77.935 3.08 ;
      RECT 77.92 2.785 77.93 3.08 ;
      RECT 77.91 2.82 77.92 3.08 ;
      RECT 77.905 2.855 77.91 3.08 ;
      RECT 78.025 2.62 78.03 3.08 ;
      RECT 77.54 2.722 77.725 2.895 ;
      RECT 77.5 2.64 77.685 2.893 ;
      RECT 77.461 2.645 77.685 2.889 ;
      RECT 77.375 2.654 77.685 2.884 ;
      RECT 77.291 2.67 77.69 2.879 ;
      RECT 77.205 2.69 77.715 2.873 ;
      RECT 77.205 2.71 77.72 2.873 ;
      RECT 77.291 2.68 77.715 2.879 ;
      RECT 77.375 2.655 77.69 2.884 ;
      RECT 77.54 2.637 77.685 2.895 ;
      RECT 77.54 2.632 77.64 2.895 ;
      RECT 77.626 2.626 77.64 2.895 ;
      RECT 77.015 1.95 77.02 2.349 ;
      RECT 76.76 1.95 76.795 2.347 ;
      RECT 76.355 1.985 76.36 2.341 ;
      RECT 77.1 1.988 77.105 2.243 ;
      RECT 77.095 1.986 77.1 2.249 ;
      RECT 77.09 1.985 77.095 2.256 ;
      RECT 77.065 1.978 77.09 2.28 ;
      RECT 77.06 1.971 77.065 2.304 ;
      RECT 77.055 1.967 77.06 2.313 ;
      RECT 77.045 1.962 77.055 2.326 ;
      RECT 77.04 1.959 77.045 2.335 ;
      RECT 77.035 1.957 77.04 2.34 ;
      RECT 77.02 1.953 77.035 2.35 ;
      RECT 77.005 1.947 77.015 2.349 ;
      RECT 76.967 1.945 77.005 2.349 ;
      RECT 76.881 1.947 76.967 2.349 ;
      RECT 76.795 1.949 76.881 2.348 ;
      RECT 76.724 1.95 76.76 2.347 ;
      RECT 76.638 1.952 76.724 2.347 ;
      RECT 76.552 1.954 76.638 2.346 ;
      RECT 76.466 1.956 76.552 2.346 ;
      RECT 76.38 1.959 76.466 2.345 ;
      RECT 76.37 1.965 76.38 2.344 ;
      RECT 76.36 1.977 76.37 2.342 ;
      RECT 76.3 2.012 76.355 2.338 ;
      RECT 76.295 2.042 76.3 2.1 ;
      RECT 77.04 3.122 77.055 3.315 ;
      RECT 77.035 3.09 77.04 3.315 ;
      RECT 77.025 3.065 77.035 3.315 ;
      RECT 77.02 3.037 77.025 3.315 ;
      RECT 76.99 2.96 77.02 3.315 ;
      RECT 76.965 2.842 76.99 3.315 ;
      RECT 76.96 2.78 76.965 3.315 ;
      RECT 76.95 2.767 76.96 3.315 ;
      RECT 76.93 2.757 76.95 3.315 ;
      RECT 76.915 2.74 76.93 3.315 ;
      RECT 76.885 2.728 76.915 3.315 ;
      RECT 76.88 2.727 76.885 3.26 ;
      RECT 76.875 2.727 76.88 3.218 ;
      RECT 76.86 2.726 76.875 3.17 ;
      RECT 76.845 2.726 76.86 3.108 ;
      RECT 76.825 2.726 76.845 3.068 ;
      RECT 76.82 2.726 76.825 3.053 ;
      RECT 76.795 2.725 76.82 3.048 ;
      RECT 76.725 2.724 76.795 3.035 ;
      RECT 76.71 2.723 76.725 3.02 ;
      RECT 76.68 2.722 76.71 3.003 ;
      RECT 76.675 2.722 76.68 2.988 ;
      RECT 76.625 2.721 76.675 2.968 ;
      RECT 76.56 2.72 76.625 2.923 ;
      RECT 76.555 2.72 76.56 2.895 ;
      RECT 76.64 3.257 76.645 3.514 ;
      RECT 76.62 3.176 76.64 3.531 ;
      RECT 76.6 3.17 76.62 3.56 ;
      RECT 76.54 3.157 76.6 3.58 ;
      RECT 76.495 3.141 76.54 3.581 ;
      RECT 76.411 3.129 76.495 3.569 ;
      RECT 76.325 3.116 76.411 3.553 ;
      RECT 76.315 3.109 76.325 3.545 ;
      RECT 76.27 3.106 76.315 3.485 ;
      RECT 76.25 3.102 76.27 3.4 ;
      RECT 76.235 3.1 76.25 3.353 ;
      RECT 76.205 3.097 76.235 3.323 ;
      RECT 76.17 3.093 76.205 3.3 ;
      RECT 76.127 3.088 76.17 3.288 ;
      RECT 76.041 3.079 76.127 3.297 ;
      RECT 75.955 3.068 76.041 3.309 ;
      RECT 75.89 3.059 75.955 3.318 ;
      RECT 75.87 3.05 75.89 3.323 ;
      RECT 75.865 3.043 75.87 3.325 ;
      RECT 75.825 3.028 75.865 3.322 ;
      RECT 75.805 3.007 75.825 3.317 ;
      RECT 75.79 2.995 75.805 3.31 ;
      RECT 75.785 2.987 75.79 3.303 ;
      RECT 75.77 2.967 75.785 3.296 ;
      RECT 75.765 2.83 75.77 3.29 ;
      RECT 75.685 2.719 75.765 3.262 ;
      RECT 75.676 2.712 75.685 3.228 ;
      RECT 75.59 2.706 75.676 3.153 ;
      RECT 75.565 2.697 75.59 3.065 ;
      RECT 75.535 2.692 75.565 3.04 ;
      RECT 75.47 2.701 75.535 3.025 ;
      RECT 75.45 2.717 75.47 3 ;
      RECT 75.44 2.723 75.45 2.948 ;
      RECT 75.42 2.745 75.44 2.83 ;
      RECT 76.075 2.71 76.245 2.895 ;
      RECT 76.075 2.71 76.28 2.893 ;
      RECT 76.125 2.62 76.295 2.884 ;
      RECT 76.075 2.777 76.3 2.877 ;
      RECT 76.09 2.655 76.295 2.884 ;
      RECT 75.29 3.388 75.355 3.831 ;
      RECT 75.23 3.413 75.355 3.829 ;
      RECT 75.23 3.413 75.41 3.823 ;
      RECT 75.215 3.438 75.41 3.822 ;
      RECT 75.355 3.375 75.43 3.819 ;
      RECT 75.29 3.4 75.51 3.813 ;
      RECT 75.215 3.439 75.555 3.807 ;
      RECT 75.2 3.466 75.555 3.798 ;
      RECT 75.215 3.459 75.575 3.79 ;
      RECT 75.2 3.468 75.58 3.773 ;
      RECT 75.195 3.485 75.58 3.6 ;
      RECT 75.2 2.207 75.235 2.445 ;
      RECT 75.2 2.207 75.265 2.444 ;
      RECT 75.2 2.207 75.38 2.44 ;
      RECT 75.2 2.207 75.435 2.418 ;
      RECT 75.21 2.15 75.49 2.318 ;
      RECT 75.315 1.99 75.345 2.441 ;
      RECT 75.345 1.985 75.525 2.198 ;
      RECT 75.215 2.126 75.525 2.198 ;
      RECT 75.265 2.022 75.315 2.442 ;
      RECT 75.235 2.078 75.525 2.198 ;
      RECT 73.74 1.74 73.91 2.935 ;
      RECT 73.74 1.74 74.205 1.91 ;
      RECT 73.74 6.97 74.205 7.14 ;
      RECT 73.74 5.945 73.91 7.14 ;
      RECT 72.75 1.74 72.92 2.935 ;
      RECT 72.75 1.74 73.215 1.91 ;
      RECT 72.75 6.97 73.215 7.14 ;
      RECT 72.75 5.945 72.92 7.14 ;
      RECT 70.895 2.635 71.065 3.865 ;
      RECT 70.95 0.855 71.12 2.805 ;
      RECT 70.895 0.575 71.065 1.025 ;
      RECT 70.895 7.855 71.065 8.305 ;
      RECT 70.95 6.075 71.12 8.025 ;
      RECT 70.895 5.015 71.065 6.245 ;
      RECT 70.375 0.575 70.545 3.865 ;
      RECT 70.375 2.075 70.78 2.405 ;
      RECT 70.375 1.235 70.78 1.565 ;
      RECT 70.375 5.015 70.545 8.305 ;
      RECT 70.375 7.315 70.78 7.645 ;
      RECT 70.375 6.475 70.78 6.805 ;
      RECT 68.475 3.392 68.49 3.443 ;
      RECT 68.47 3.372 68.475 3.49 ;
      RECT 68.455 3.362 68.47 3.558 ;
      RECT 68.43 3.342 68.455 3.613 ;
      RECT 68.39 3.327 68.43 3.633 ;
      RECT 68.345 3.321 68.39 3.661 ;
      RECT 68.275 3.311 68.345 3.678 ;
      RECT 68.255 3.303 68.275 3.678 ;
      RECT 68.195 3.297 68.255 3.67 ;
      RECT 68.136 3.288 68.195 3.658 ;
      RECT 68.05 3.277 68.136 3.641 ;
      RECT 68.028 3.268 68.05 3.629 ;
      RECT 67.942 3.261 68.028 3.616 ;
      RECT 67.856 3.248 67.942 3.597 ;
      RECT 67.77 3.236 67.856 3.577 ;
      RECT 67.74 3.225 67.77 3.564 ;
      RECT 67.69 3.211 67.74 3.556 ;
      RECT 67.67 3.2 67.69 3.548 ;
      RECT 67.621 3.189 67.67 3.54 ;
      RECT 67.535 3.168 67.621 3.525 ;
      RECT 67.49 3.155 67.535 3.51 ;
      RECT 67.445 3.155 67.49 3.49 ;
      RECT 67.39 3.155 67.445 3.425 ;
      RECT 67.365 3.155 67.39 3.348 ;
      RECT 67.89 2.892 68.06 3.075 ;
      RECT 67.89 2.892 68.075 3.033 ;
      RECT 67.89 2.892 68.08 2.975 ;
      RECT 67.95 2.66 68.085 2.951 ;
      RECT 67.95 2.664 68.09 2.934 ;
      RECT 67.895 2.827 68.09 2.934 ;
      RECT 67.92 2.672 68.06 3.075 ;
      RECT 67.92 2.676 68.1 2.875 ;
      RECT 67.905 2.762 68.1 2.875 ;
      RECT 67.915 2.692 68.06 3.075 ;
      RECT 67.915 2.695 68.11 2.788 ;
      RECT 67.91 2.712 68.11 2.788 ;
      RECT 67.68 1.932 67.85 2.415 ;
      RECT 67.675 1.927 67.825 2.405 ;
      RECT 67.675 1.934 67.855 2.399 ;
      RECT 67.665 1.928 67.825 2.378 ;
      RECT 67.665 1.944 67.87 2.337 ;
      RECT 67.635 1.929 67.825 2.3 ;
      RECT 67.635 1.959 67.88 2.24 ;
      RECT 67.63 1.931 67.825 2.238 ;
      RECT 67.61 1.94 67.855 2.195 ;
      RECT 67.585 1.956 67.87 2.107 ;
      RECT 67.585 1.975 67.895 2.098 ;
      RECT 67.58 2.012 67.895 2.05 ;
      RECT 67.585 1.992 67.9 2.018 ;
      RECT 67.68 1.926 67.79 2.415 ;
      RECT 67.766 1.925 67.79 2.415 ;
      RECT 67 2.71 67.005 2.921 ;
      RECT 67.6 2.71 67.605 2.895 ;
      RECT 67.665 2.75 67.67 2.863 ;
      RECT 67.66 2.742 67.665 2.869 ;
      RECT 67.655 2.732 67.66 2.877 ;
      RECT 67.65 2.722 67.655 2.886 ;
      RECT 67.645 2.712 67.65 2.89 ;
      RECT 67.605 2.71 67.645 2.893 ;
      RECT 67.577 2.709 67.6 2.897 ;
      RECT 67.491 2.706 67.577 2.904 ;
      RECT 67.405 2.702 67.491 2.915 ;
      RECT 67.385 2.7 67.405 2.921 ;
      RECT 67.367 2.699 67.385 2.924 ;
      RECT 67.281 2.697 67.367 2.931 ;
      RECT 67.195 2.692 67.281 2.944 ;
      RECT 67.176 2.689 67.195 2.949 ;
      RECT 67.09 2.687 67.176 2.94 ;
      RECT 67.08 2.687 67.09 2.933 ;
      RECT 67.005 2.7 67.08 2.927 ;
      RECT 66.99 2.711 67 2.921 ;
      RECT 66.98 2.713 66.99 2.92 ;
      RECT 66.97 2.717 66.98 2.916 ;
      RECT 66.965 2.72 66.97 2.91 ;
      RECT 66.955 2.722 66.965 2.904 ;
      RECT 66.95 2.725 66.955 2.898 ;
      RECT 66.93 3.311 66.935 3.515 ;
      RECT 66.915 3.298 66.93 3.608 ;
      RECT 66.9 3.279 66.915 3.885 ;
      RECT 66.865 3.245 66.9 3.885 ;
      RECT 66.861 3.215 66.865 3.885 ;
      RECT 66.775 3.097 66.861 3.885 ;
      RECT 66.765 2.972 66.775 3.885 ;
      RECT 66.75 2.94 66.765 3.885 ;
      RECT 66.745 2.915 66.75 3.885 ;
      RECT 66.74 2.905 66.745 3.841 ;
      RECT 66.725 2.877 66.74 3.746 ;
      RECT 66.71 2.843 66.725 3.645 ;
      RECT 66.705 2.821 66.71 3.598 ;
      RECT 66.7 2.81 66.705 3.568 ;
      RECT 66.695 2.8 66.7 3.534 ;
      RECT 66.685 2.787 66.695 3.502 ;
      RECT 66.66 2.763 66.685 3.428 ;
      RECT 66.655 2.743 66.66 3.353 ;
      RECT 66.65 2.737 66.655 3.328 ;
      RECT 66.645 2.732 66.65 3.293 ;
      RECT 66.64 2.727 66.645 3.268 ;
      RECT 66.635 2.725 66.64 3.248 ;
      RECT 66.63 2.725 66.635 3.233 ;
      RECT 66.625 2.725 66.63 3.193 ;
      RECT 66.615 2.725 66.625 3.165 ;
      RECT 66.605 2.725 66.615 3.11 ;
      RECT 66.59 2.725 66.605 3.048 ;
      RECT 66.585 2.724 66.59 2.993 ;
      RECT 66.57 2.723 66.585 2.973 ;
      RECT 66.51 2.721 66.57 2.947 ;
      RECT 66.475 2.722 66.51 2.927 ;
      RECT 66.47 2.724 66.475 2.917 ;
      RECT 66.46 2.743 66.47 2.907 ;
      RECT 66.455 2.77 66.46 2.838 ;
      RECT 66.57 2.195 66.74 2.44 ;
      RECT 66.605 1.966 66.74 2.44 ;
      RECT 66.605 1.968 66.75 2.435 ;
      RECT 66.605 1.97 66.775 2.423 ;
      RECT 66.605 1.973 66.8 2.405 ;
      RECT 66.605 1.978 66.85 2.378 ;
      RECT 66.605 1.983 66.87 2.343 ;
      RECT 66.585 1.985 66.88 2.318 ;
      RECT 66.575 2.08 66.88 2.318 ;
      RECT 66.605 1.965 66.715 2.44 ;
      RECT 66.615 1.962 66.71 2.44 ;
      RECT 66.135 3.227 66.325 3.585 ;
      RECT 66.135 3.239 66.36 3.584 ;
      RECT 66.135 3.267 66.38 3.582 ;
      RECT 66.135 3.292 66.385 3.581 ;
      RECT 66.135 3.35 66.4 3.58 ;
      RECT 66.12 3.223 66.28 3.565 ;
      RECT 66.1 3.232 66.325 3.518 ;
      RECT 66.075 3.243 66.36 3.455 ;
      RECT 66.075 3.327 66.395 3.455 ;
      RECT 66.075 3.302 66.39 3.455 ;
      RECT 66.135 3.218 66.28 3.585 ;
      RECT 66.221 3.217 66.28 3.585 ;
      RECT 66.221 3.216 66.265 3.585 ;
      RECT 66.135 7.855 66.305 8.305 ;
      RECT 66.19 6.075 66.36 8.025 ;
      RECT 66.135 5.015 66.305 6.245 ;
      RECT 65.615 5.015 65.785 8.305 ;
      RECT 65.615 7.315 66.02 7.645 ;
      RECT 65.615 6.475 66.02 6.805 ;
      RECT 65.92 2.732 65.925 3.11 ;
      RECT 65.915 2.7 65.92 3.11 ;
      RECT 65.91 2.672 65.915 3.11 ;
      RECT 65.905 2.652 65.91 3.11 ;
      RECT 65.85 2.635 65.905 3.11 ;
      RECT 65.81 2.62 65.85 3.11 ;
      RECT 65.755 2.607 65.81 3.11 ;
      RECT 65.72 2.598 65.755 3.11 ;
      RECT 65.716 2.596 65.72 3.109 ;
      RECT 65.63 2.592 65.716 3.092 ;
      RECT 65.545 2.584 65.63 3.055 ;
      RECT 65.535 2.58 65.545 3.028 ;
      RECT 65.525 2.58 65.535 3.01 ;
      RECT 65.515 2.582 65.525 2.993 ;
      RECT 65.51 2.587 65.515 2.979 ;
      RECT 65.505 2.591 65.51 2.966 ;
      RECT 65.495 2.596 65.505 2.95 ;
      RECT 65.48 2.61 65.495 2.925 ;
      RECT 65.475 2.616 65.48 2.905 ;
      RECT 65.47 2.618 65.475 2.898 ;
      RECT 65.465 2.622 65.47 2.773 ;
      RECT 65.645 3.422 65.89 3.885 ;
      RECT 65.565 3.395 65.885 3.881 ;
      RECT 65.495 3.43 65.89 3.874 ;
      RECT 65.285 3.685 65.89 3.87 ;
      RECT 65.465 3.453 65.89 3.87 ;
      RECT 65.305 3.645 65.89 3.87 ;
      RECT 65.455 3.465 65.89 3.87 ;
      RECT 65.34 3.582 65.89 3.87 ;
      RECT 65.395 3.507 65.89 3.87 ;
      RECT 65.645 3.372 65.885 3.885 ;
      RECT 65.675 3.365 65.885 3.885 ;
      RECT 65.665 3.367 65.885 3.885 ;
      RECT 65.675 3.362 65.805 3.885 ;
      RECT 65.23 1.925 65.316 2.364 ;
      RECT 65.225 1.925 65.316 2.362 ;
      RECT 65.225 1.925 65.385 2.361 ;
      RECT 65.225 1.925 65.415 2.358 ;
      RECT 65.21 1.932 65.415 2.349 ;
      RECT 65.21 1.932 65.42 2.345 ;
      RECT 65.205 1.942 65.42 2.338 ;
      RECT 65.2 1.947 65.42 2.313 ;
      RECT 65.2 1.947 65.435 2.295 ;
      RECT 65.225 1.925 65.455 2.21 ;
      RECT 65.195 1.952 65.455 2.208 ;
      RECT 65.205 1.945 65.46 2.146 ;
      RECT 65.195 2.067 65.465 2.129 ;
      RECT 65.18 1.962 65.46 2.08 ;
      RECT 65.175 1.972 65.46 1.98 ;
      RECT 65.255 2.743 65.26 2.82 ;
      RECT 65.245 2.737 65.255 3.01 ;
      RECT 65.235 2.729 65.245 3.031 ;
      RECT 65.225 2.72 65.235 3.053 ;
      RECT 65.22 2.715 65.225 3.07 ;
      RECT 65.18 2.715 65.22 3.11 ;
      RECT 65.16 2.715 65.18 3.165 ;
      RECT 65.155 2.715 65.16 3.193 ;
      RECT 65.145 2.715 65.155 3.208 ;
      RECT 65.11 2.715 65.145 3.25 ;
      RECT 65.105 2.715 65.11 3.293 ;
      RECT 65.095 2.715 65.105 3.308 ;
      RECT 65.08 2.715 65.095 3.328 ;
      RECT 65.065 2.715 65.08 3.355 ;
      RECT 65.06 2.716 65.065 3.373 ;
      RECT 65.04 2.717 65.06 3.38 ;
      RECT 64.985 2.718 65.04 3.4 ;
      RECT 64.975 2.719 64.985 3.414 ;
      RECT 64.97 2.722 64.975 3.413 ;
      RECT 64.93 2.795 64.97 3.411 ;
      RECT 64.915 2.875 64.93 3.409 ;
      RECT 64.89 2.93 64.915 3.407 ;
      RECT 64.875 2.995 64.89 3.406 ;
      RECT 64.83 3.027 64.875 3.403 ;
      RECT 64.745 3.05 64.83 3.398 ;
      RECT 64.72 3.07 64.745 3.393 ;
      RECT 64.65 3.075 64.72 3.389 ;
      RECT 64.63 3.077 64.65 3.386 ;
      RECT 64.545 3.088 64.63 3.38 ;
      RECT 64.54 3.099 64.545 3.375 ;
      RECT 64.53 3.101 64.54 3.375 ;
      RECT 64.495 3.105 64.53 3.373 ;
      RECT 64.445 3.115 64.495 3.36 ;
      RECT 64.425 3.123 64.445 3.345 ;
      RECT 64.345 3.135 64.425 3.328 ;
      RECT 64.51 2.685 64.68 2.895 ;
      RECT 64.626 2.681 64.68 2.895 ;
      RECT 64.431 2.685 64.68 2.886 ;
      RECT 64.431 2.685 64.685 2.875 ;
      RECT 64.345 2.685 64.685 2.866 ;
      RECT 64.345 2.693 64.695 2.81 ;
      RECT 64.345 2.705 64.7 2.723 ;
      RECT 64.345 2.712 64.705 2.715 ;
      RECT 64.54 2.683 64.68 2.895 ;
      RECT 64.295 3.628 64.54 3.96 ;
      RECT 64.29 3.62 64.295 3.957 ;
      RECT 64.26 3.64 64.54 3.938 ;
      RECT 64.24 3.672 64.54 3.911 ;
      RECT 64.29 3.625 64.467 3.957 ;
      RECT 64.29 3.622 64.381 3.957 ;
      RECT 64.23 1.97 64.4 2.39 ;
      RECT 64.225 1.97 64.4 2.388 ;
      RECT 64.225 1.97 64.425 2.378 ;
      RECT 64.225 1.97 64.445 2.353 ;
      RECT 64.22 1.97 64.445 2.348 ;
      RECT 64.22 1.97 64.455 2.338 ;
      RECT 64.22 1.97 64.46 2.333 ;
      RECT 64.22 1.975 64.465 2.328 ;
      RECT 64.22 2.007 64.48 2.318 ;
      RECT 64.22 2.077 64.505 2.301 ;
      RECT 64.2 2.077 64.505 2.293 ;
      RECT 64.2 2.137 64.515 2.27 ;
      RECT 64.2 2.177 64.525 2.215 ;
      RECT 64.185 1.97 64.46 2.195 ;
      RECT 64.175 1.985 64.465 2.093 ;
      RECT 63.765 3.375 63.935 3.9 ;
      RECT 63.76 3.375 63.935 3.893 ;
      RECT 63.75 3.375 63.94 3.858 ;
      RECT 63.745 3.385 63.94 3.83 ;
      RECT 63.74 3.405 63.94 3.813 ;
      RECT 63.75 3.38 63.945 3.803 ;
      RECT 63.735 3.425 63.945 3.795 ;
      RECT 63.73 3.445 63.945 3.78 ;
      RECT 63.725 3.475 63.945 3.77 ;
      RECT 63.715 3.52 63.945 3.745 ;
      RECT 63.745 3.39 63.95 3.728 ;
      RECT 63.71 3.572 63.95 3.723 ;
      RECT 63.745 3.4 63.955 3.693 ;
      RECT 63.705 3.605 63.955 3.69 ;
      RECT 63.7 3.63 63.955 3.67 ;
      RECT 63.74 3.417 63.965 3.61 ;
      RECT 63.735 3.439 63.975 3.503 ;
      RECT 63.685 2.686 63.7 2.955 ;
      RECT 63.64 2.67 63.685 3 ;
      RECT 63.635 2.658 63.64 3.05 ;
      RECT 63.625 2.654 63.635 3.083 ;
      RECT 63.62 2.651 63.625 3.111 ;
      RECT 63.605 2.653 63.62 3.153 ;
      RECT 63.6 2.657 63.605 3.193 ;
      RECT 63.58 2.662 63.6 3.245 ;
      RECT 63.576 2.667 63.58 3.302 ;
      RECT 63.49 2.686 63.576 3.339 ;
      RECT 63.48 2.707 63.49 3.375 ;
      RECT 63.475 2.715 63.48 3.376 ;
      RECT 63.47 2.757 63.475 3.377 ;
      RECT 63.455 2.845 63.47 3.378 ;
      RECT 63.445 2.995 63.455 3.38 ;
      RECT 63.44 3.04 63.445 3.382 ;
      RECT 63.405 3.082 63.44 3.385 ;
      RECT 63.4 3.1 63.405 3.388 ;
      RECT 63.323 3.106 63.4 3.394 ;
      RECT 63.237 3.12 63.323 3.407 ;
      RECT 63.151 3.134 63.237 3.421 ;
      RECT 63.065 3.148 63.151 3.434 ;
      RECT 63.005 3.16 63.065 3.446 ;
      RECT 62.98 3.167 63.005 3.453 ;
      RECT 62.966 3.17 62.98 3.458 ;
      RECT 62.88 3.178 62.966 3.474 ;
      RECT 62.875 3.185 62.88 3.489 ;
      RECT 62.851 3.185 62.875 3.496 ;
      RECT 62.765 3.188 62.851 3.524 ;
      RECT 62.68 3.192 62.765 3.568 ;
      RECT 62.615 3.196 62.68 3.605 ;
      RECT 62.59 3.199 62.615 3.621 ;
      RECT 62.515 3.212 62.59 3.625 ;
      RECT 62.49 3.23 62.515 3.629 ;
      RECT 62.48 3.237 62.49 3.631 ;
      RECT 62.465 3.24 62.48 3.632 ;
      RECT 62.405 3.252 62.465 3.636 ;
      RECT 62.395 3.266 62.405 3.64 ;
      RECT 62.34 3.276 62.395 3.628 ;
      RECT 62.315 3.297 62.34 3.611 ;
      RECT 62.295 3.317 62.315 3.602 ;
      RECT 62.29 3.33 62.295 3.597 ;
      RECT 62.275 3.342 62.29 3.593 ;
      RECT 63.51 1.997 63.515 2.02 ;
      RECT 63.505 1.988 63.51 2.06 ;
      RECT 63.5 1.986 63.505 2.103 ;
      RECT 63.495 1.977 63.5 2.138 ;
      RECT 63.49 1.967 63.495 2.21 ;
      RECT 63.485 1.957 63.49 2.275 ;
      RECT 63.48 1.954 63.485 2.315 ;
      RECT 63.455 1.948 63.48 2.405 ;
      RECT 63.42 1.936 63.455 2.43 ;
      RECT 63.41 1.927 63.42 2.43 ;
      RECT 63.275 1.925 63.285 2.413 ;
      RECT 63.265 1.925 63.275 2.38 ;
      RECT 63.26 1.925 63.265 2.355 ;
      RECT 63.255 1.925 63.26 2.343 ;
      RECT 63.25 1.925 63.255 2.325 ;
      RECT 63.24 1.925 63.25 2.29 ;
      RECT 63.235 1.927 63.24 2.268 ;
      RECT 63.23 1.933 63.235 2.253 ;
      RECT 63.225 1.939 63.23 2.238 ;
      RECT 63.21 1.951 63.225 2.211 ;
      RECT 63.205 1.962 63.21 2.179 ;
      RECT 63.2 1.972 63.205 2.163 ;
      RECT 63.19 1.98 63.2 2.132 ;
      RECT 63.185 1.99 63.19 2.106 ;
      RECT 63.18 2.047 63.185 2.089 ;
      RECT 63.285 1.925 63.41 2.43 ;
      RECT 63 2.612 63.26 2.91 ;
      RECT 62.995 2.619 63.26 2.908 ;
      RECT 63 2.614 63.275 2.903 ;
      RECT 62.99 2.627 63.275 2.9 ;
      RECT 62.99 2.632 63.28 2.893 ;
      RECT 62.985 2.64 63.28 2.89 ;
      RECT 62.985 2.657 63.285 2.688 ;
      RECT 63 2.609 63.231 2.91 ;
      RECT 63.055 2.608 63.231 2.91 ;
      RECT 63.055 2.605 63.145 2.91 ;
      RECT 63.055 2.602 63.141 2.91 ;
      RECT 62.745 2.875 62.75 2.888 ;
      RECT 62.74 2.842 62.745 2.893 ;
      RECT 62.735 2.797 62.74 2.9 ;
      RECT 62.73 2.752 62.735 2.908 ;
      RECT 62.725 2.72 62.73 2.916 ;
      RECT 62.72 2.68 62.725 2.917 ;
      RECT 62.705 2.66 62.72 2.919 ;
      RECT 62.63 2.642 62.705 2.931 ;
      RECT 62.62 2.635 62.63 2.942 ;
      RECT 62.615 2.635 62.62 2.944 ;
      RECT 62.585 2.641 62.615 2.948 ;
      RECT 62.545 2.654 62.585 2.948 ;
      RECT 62.52 2.665 62.545 2.934 ;
      RECT 62.505 2.671 62.52 2.917 ;
      RECT 62.495 2.673 62.505 2.908 ;
      RECT 62.49 2.674 62.495 2.903 ;
      RECT 62.485 2.675 62.49 2.898 ;
      RECT 62.48 2.676 62.485 2.895 ;
      RECT 62.455 2.681 62.48 2.885 ;
      RECT 62.445 2.697 62.455 2.872 ;
      RECT 62.44 2.717 62.445 2.867 ;
      RECT 62.45 2.11 62.455 2.306 ;
      RECT 62.435 2.074 62.45 2.308 ;
      RECT 62.425 2.056 62.435 2.313 ;
      RECT 62.415 2.042 62.425 2.317 ;
      RECT 62.37 2.026 62.415 2.327 ;
      RECT 62.365 2.016 62.37 2.336 ;
      RECT 62.32 2.005 62.365 2.342 ;
      RECT 62.315 1.993 62.32 2.349 ;
      RECT 62.3 1.988 62.315 2.353 ;
      RECT 62.285 1.98 62.3 2.358 ;
      RECT 62.275 1.973 62.285 2.363 ;
      RECT 62.265 1.97 62.275 2.368 ;
      RECT 62.255 1.97 62.265 2.369 ;
      RECT 62.25 1.967 62.255 2.368 ;
      RECT 62.215 1.962 62.24 2.367 ;
      RECT 62.191 1.958 62.215 2.366 ;
      RECT 62.105 1.949 62.191 2.363 ;
      RECT 62.09 1.941 62.105 2.36 ;
      RECT 62.068 1.94 62.09 2.359 ;
      RECT 61.982 1.94 62.068 2.357 ;
      RECT 61.896 1.94 61.982 2.355 ;
      RECT 61.81 1.94 61.896 2.352 ;
      RECT 61.8 1.94 61.81 2.343 ;
      RECT 61.77 1.94 61.8 2.303 ;
      RECT 61.76 1.95 61.77 2.258 ;
      RECT 61.755 1.99 61.76 2.243 ;
      RECT 61.75 2.005 61.755 2.23 ;
      RECT 61.72 2.085 61.75 2.192 ;
      RECT 62.24 1.965 62.25 2.368 ;
      RECT 62.065 2.73 62.08 3.335 ;
      RECT 62.07 2.725 62.08 3.335 ;
      RECT 62.235 2.725 62.24 2.908 ;
      RECT 62.225 2.725 62.235 2.938 ;
      RECT 62.21 2.725 62.225 2.998 ;
      RECT 62.205 2.725 62.21 3.043 ;
      RECT 62.2 2.725 62.205 3.073 ;
      RECT 62.195 2.725 62.2 3.093 ;
      RECT 62.185 2.725 62.195 3.128 ;
      RECT 62.17 2.725 62.185 3.16 ;
      RECT 62.125 2.725 62.17 3.188 ;
      RECT 62.12 2.725 62.125 3.218 ;
      RECT 62.115 2.725 62.12 3.23 ;
      RECT 62.11 2.725 62.115 3.238 ;
      RECT 62.1 2.725 62.11 3.253 ;
      RECT 62.095 2.725 62.1 3.275 ;
      RECT 62.085 2.725 62.095 3.298 ;
      RECT 62.08 2.725 62.085 3.318 ;
      RECT 62.045 2.74 62.065 3.335 ;
      RECT 62.02 2.757 62.045 3.335 ;
      RECT 62.015 2.767 62.02 3.335 ;
      RECT 61.985 2.782 62.015 3.335 ;
      RECT 61.91 2.824 61.985 3.335 ;
      RECT 61.905 2.855 61.91 3.318 ;
      RECT 61.9 2.859 61.905 3.3 ;
      RECT 61.895 2.863 61.9 3.263 ;
      RECT 61.89 3.047 61.895 3.23 ;
      RECT 61.375 3.236 61.461 3.801 ;
      RECT 61.33 3.238 61.495 3.795 ;
      RECT 61.461 3.235 61.495 3.795 ;
      RECT 61.375 3.237 61.58 3.789 ;
      RECT 61.33 3.247 61.59 3.785 ;
      RECT 61.305 3.239 61.58 3.781 ;
      RECT 61.3 3.242 61.58 3.776 ;
      RECT 61.275 3.257 61.59 3.77 ;
      RECT 61.275 3.282 61.63 3.765 ;
      RECT 61.235 3.29 61.63 3.74 ;
      RECT 61.235 3.317 61.645 3.738 ;
      RECT 61.235 3.347 61.655 3.725 ;
      RECT 61.23 3.492 61.655 3.713 ;
      RECT 61.235 3.421 61.675 3.71 ;
      RECT 61.235 3.478 61.68 3.518 ;
      RECT 61.425 2.757 61.595 2.935 ;
      RECT 61.375 2.696 61.425 2.92 ;
      RECT 61.11 2.676 61.375 2.905 ;
      RECT 61.07 2.74 61.545 2.905 ;
      RECT 61.07 2.73 61.5 2.905 ;
      RECT 61.07 2.727 61.49 2.905 ;
      RECT 61.07 2.715 61.48 2.905 ;
      RECT 61.07 2.7 61.425 2.905 ;
      RECT 61.11 2.672 61.311 2.905 ;
      RECT 61.12 2.65 61.311 2.905 ;
      RECT 61.145 2.635 61.225 2.905 ;
      RECT 60.9 3.165 61.02 3.61 ;
      RECT 60.885 3.165 61.02 3.609 ;
      RECT 60.84 3.187 61.02 3.604 ;
      RECT 60.8 3.236 61.02 3.598 ;
      RECT 60.8 3.236 61.025 3.573 ;
      RECT 60.8 3.236 61.045 3.463 ;
      RECT 60.795 3.266 61.045 3.46 ;
      RECT 60.885 3.165 61.055 3.355 ;
      RECT 60.545 1.95 60.55 2.395 ;
      RECT 60.355 1.95 60.375 2.36 ;
      RECT 60.325 1.95 60.33 2.335 ;
      RECT 61.005 2.257 61.02 2.445 ;
      RECT 61 2.242 61.005 2.451 ;
      RECT 60.98 2.215 61 2.454 ;
      RECT 60.93 2.182 60.98 2.463 ;
      RECT 60.9 2.162 60.93 2.467 ;
      RECT 60.881 2.15 60.9 2.463 ;
      RECT 60.795 2.122 60.881 2.453 ;
      RECT 60.785 2.097 60.795 2.443 ;
      RECT 60.715 2.065 60.785 2.435 ;
      RECT 60.69 2.025 60.715 2.427 ;
      RECT 60.67 2.007 60.69 2.421 ;
      RECT 60.66 1.997 60.67 2.418 ;
      RECT 60.65 1.99 60.66 2.416 ;
      RECT 60.63 1.977 60.65 2.413 ;
      RECT 60.62 1.967 60.63 2.41 ;
      RECT 60.61 1.96 60.62 2.408 ;
      RECT 60.56 1.952 60.61 2.402 ;
      RECT 60.55 1.95 60.56 2.396 ;
      RECT 60.52 1.95 60.545 2.393 ;
      RECT 60.491 1.95 60.52 2.388 ;
      RECT 60.405 1.95 60.491 2.378 ;
      RECT 60.375 1.95 60.405 2.365 ;
      RECT 60.33 1.95 60.355 2.348 ;
      RECT 60.315 1.95 60.325 2.33 ;
      RECT 60.295 1.957 60.315 2.315 ;
      RECT 60.29 1.972 60.295 2.303 ;
      RECT 60.285 1.977 60.29 2.243 ;
      RECT 60.28 1.982 60.285 2.085 ;
      RECT 60.275 1.985 60.28 2.003 ;
      RECT 60.54 2.67 60.626 2.991 ;
      RECT 60.54 2.67 60.66 2.984 ;
      RECT 60.49 2.67 60.66 2.98 ;
      RECT 60.49 2.672 60.746 2.978 ;
      RECT 60.49 2.674 60.77 2.972 ;
      RECT 60.49 2.681 60.78 2.971 ;
      RECT 60.49 2.69 60.785 2.968 ;
      RECT 60.49 2.696 60.79 2.963 ;
      RECT 60.49 2.74 60.795 2.96 ;
      RECT 60.49 2.832 60.8 2.957 ;
      RECT 60.015 3.275 60.05 3.595 ;
      RECT 60.6 3.46 60.605 3.642 ;
      RECT 60.555 3.342 60.6 3.661 ;
      RECT 60.54 3.319 60.555 3.684 ;
      RECT 60.53 3.309 60.54 3.694 ;
      RECT 60.51 3.304 60.53 3.707 ;
      RECT 60.485 3.302 60.51 3.728 ;
      RECT 60.466 3.301 60.485 3.74 ;
      RECT 60.38 3.298 60.466 3.74 ;
      RECT 60.31 3.293 60.38 3.728 ;
      RECT 60.235 3.289 60.31 3.703 ;
      RECT 60.17 3.285 60.235 3.67 ;
      RECT 60.1 3.282 60.17 3.63 ;
      RECT 60.07 3.278 60.1 3.605 ;
      RECT 60.05 3.276 60.07 3.598 ;
      RECT 59.966 3.274 60.015 3.596 ;
      RECT 59.88 3.271 59.966 3.597 ;
      RECT 59.805 3.27 59.88 3.599 ;
      RECT 59.72 3.27 59.805 3.625 ;
      RECT 59.643 3.271 59.72 3.65 ;
      RECT 59.557 3.272 59.643 3.65 ;
      RECT 59.471 3.272 59.557 3.65 ;
      RECT 59.385 3.273 59.471 3.65 ;
      RECT 59.365 3.274 59.385 3.642 ;
      RECT 59.35 3.28 59.365 3.627 ;
      RECT 59.315 3.3 59.35 3.607 ;
      RECT 59.305 3.32 59.315 3.589 ;
      RECT 60.275 2.625 60.28 2.895 ;
      RECT 60.27 2.616 60.275 2.9 ;
      RECT 60.26 2.606 60.27 2.912 ;
      RECT 60.255 2.595 60.26 2.923 ;
      RECT 60.235 2.589 60.255 2.941 ;
      RECT 60.19 2.586 60.235 2.99 ;
      RECT 60.175 2.585 60.19 3.035 ;
      RECT 60.17 2.585 60.175 3.048 ;
      RECT 60.16 2.585 60.17 3.06 ;
      RECT 60.155 2.586 60.16 3.075 ;
      RECT 60.135 2.594 60.155 3.08 ;
      RECT 60.105 2.61 60.135 3.08 ;
      RECT 60.095 2.622 60.1 3.08 ;
      RECT 60.06 2.637 60.095 3.08 ;
      RECT 60.03 2.657 60.06 3.08 ;
      RECT 60.02 2.682 60.03 3.08 ;
      RECT 60.015 2.71 60.02 3.08 ;
      RECT 60.01 2.74 60.015 3.08 ;
      RECT 60.005 2.757 60.01 3.08 ;
      RECT 59.995 2.785 60.005 3.08 ;
      RECT 59.985 2.82 59.995 3.08 ;
      RECT 59.98 2.855 59.985 3.08 ;
      RECT 60.1 2.62 60.105 3.08 ;
      RECT 59.615 2.722 59.8 2.895 ;
      RECT 59.575 2.64 59.76 2.893 ;
      RECT 59.536 2.645 59.76 2.889 ;
      RECT 59.45 2.654 59.76 2.884 ;
      RECT 59.366 2.67 59.765 2.879 ;
      RECT 59.28 2.69 59.79 2.873 ;
      RECT 59.28 2.71 59.795 2.873 ;
      RECT 59.366 2.68 59.79 2.879 ;
      RECT 59.45 2.655 59.765 2.884 ;
      RECT 59.615 2.637 59.76 2.895 ;
      RECT 59.615 2.632 59.715 2.895 ;
      RECT 59.701 2.626 59.715 2.895 ;
      RECT 59.09 1.95 59.095 2.349 ;
      RECT 58.835 1.95 58.87 2.347 ;
      RECT 58.43 1.985 58.435 2.341 ;
      RECT 59.175 1.988 59.18 2.243 ;
      RECT 59.17 1.986 59.175 2.249 ;
      RECT 59.165 1.985 59.17 2.256 ;
      RECT 59.14 1.978 59.165 2.28 ;
      RECT 59.135 1.971 59.14 2.304 ;
      RECT 59.13 1.967 59.135 2.313 ;
      RECT 59.12 1.962 59.13 2.326 ;
      RECT 59.115 1.959 59.12 2.335 ;
      RECT 59.11 1.957 59.115 2.34 ;
      RECT 59.095 1.953 59.11 2.35 ;
      RECT 59.08 1.947 59.09 2.349 ;
      RECT 59.042 1.945 59.08 2.349 ;
      RECT 58.956 1.947 59.042 2.349 ;
      RECT 58.87 1.949 58.956 2.348 ;
      RECT 58.799 1.95 58.835 2.347 ;
      RECT 58.713 1.952 58.799 2.347 ;
      RECT 58.627 1.954 58.713 2.346 ;
      RECT 58.541 1.956 58.627 2.346 ;
      RECT 58.455 1.959 58.541 2.345 ;
      RECT 58.445 1.965 58.455 2.344 ;
      RECT 58.435 1.977 58.445 2.342 ;
      RECT 58.375 2.012 58.43 2.338 ;
      RECT 58.37 2.042 58.375 2.1 ;
      RECT 59.115 3.122 59.13 3.315 ;
      RECT 59.11 3.09 59.115 3.315 ;
      RECT 59.1 3.065 59.11 3.315 ;
      RECT 59.095 3.037 59.1 3.315 ;
      RECT 59.065 2.96 59.095 3.315 ;
      RECT 59.04 2.842 59.065 3.315 ;
      RECT 59.035 2.78 59.04 3.315 ;
      RECT 59.025 2.767 59.035 3.315 ;
      RECT 59.005 2.757 59.025 3.315 ;
      RECT 58.99 2.74 59.005 3.315 ;
      RECT 58.96 2.728 58.99 3.315 ;
      RECT 58.955 2.727 58.96 3.26 ;
      RECT 58.95 2.727 58.955 3.218 ;
      RECT 58.935 2.726 58.95 3.17 ;
      RECT 58.92 2.726 58.935 3.108 ;
      RECT 58.9 2.726 58.92 3.068 ;
      RECT 58.895 2.726 58.9 3.053 ;
      RECT 58.87 2.725 58.895 3.048 ;
      RECT 58.8 2.724 58.87 3.035 ;
      RECT 58.785 2.723 58.8 3.02 ;
      RECT 58.755 2.722 58.785 3.003 ;
      RECT 58.75 2.722 58.755 2.988 ;
      RECT 58.7 2.721 58.75 2.968 ;
      RECT 58.635 2.72 58.7 2.923 ;
      RECT 58.63 2.72 58.635 2.895 ;
      RECT 58.715 3.257 58.72 3.514 ;
      RECT 58.695 3.176 58.715 3.531 ;
      RECT 58.675 3.17 58.695 3.56 ;
      RECT 58.615 3.157 58.675 3.58 ;
      RECT 58.57 3.141 58.615 3.581 ;
      RECT 58.486 3.129 58.57 3.569 ;
      RECT 58.4 3.116 58.486 3.553 ;
      RECT 58.39 3.109 58.4 3.545 ;
      RECT 58.345 3.106 58.39 3.485 ;
      RECT 58.325 3.102 58.345 3.4 ;
      RECT 58.31 3.1 58.325 3.353 ;
      RECT 58.28 3.097 58.31 3.323 ;
      RECT 58.245 3.093 58.28 3.3 ;
      RECT 58.202 3.088 58.245 3.288 ;
      RECT 58.116 3.079 58.202 3.297 ;
      RECT 58.03 3.068 58.116 3.309 ;
      RECT 57.965 3.059 58.03 3.318 ;
      RECT 57.945 3.05 57.965 3.323 ;
      RECT 57.94 3.043 57.945 3.325 ;
      RECT 57.9 3.028 57.94 3.322 ;
      RECT 57.88 3.007 57.9 3.317 ;
      RECT 57.865 2.995 57.88 3.31 ;
      RECT 57.86 2.987 57.865 3.303 ;
      RECT 57.845 2.967 57.86 3.296 ;
      RECT 57.84 2.83 57.845 3.29 ;
      RECT 57.76 2.719 57.84 3.262 ;
      RECT 57.751 2.712 57.76 3.228 ;
      RECT 57.665 2.706 57.751 3.153 ;
      RECT 57.64 2.697 57.665 3.065 ;
      RECT 57.61 2.692 57.64 3.04 ;
      RECT 57.545 2.701 57.61 3.025 ;
      RECT 57.525 2.717 57.545 3 ;
      RECT 57.515 2.723 57.525 2.948 ;
      RECT 57.495 2.745 57.515 2.83 ;
      RECT 58.15 2.71 58.32 2.895 ;
      RECT 58.15 2.71 58.355 2.893 ;
      RECT 58.2 2.62 58.37 2.884 ;
      RECT 58.15 2.777 58.375 2.877 ;
      RECT 58.165 2.655 58.37 2.884 ;
      RECT 57.365 3.388 57.43 3.831 ;
      RECT 57.305 3.413 57.43 3.829 ;
      RECT 57.305 3.413 57.485 3.823 ;
      RECT 57.29 3.438 57.485 3.822 ;
      RECT 57.43 3.375 57.505 3.819 ;
      RECT 57.365 3.4 57.585 3.813 ;
      RECT 57.29 3.439 57.63 3.807 ;
      RECT 57.275 3.466 57.63 3.798 ;
      RECT 57.29 3.459 57.65 3.79 ;
      RECT 57.275 3.468 57.655 3.773 ;
      RECT 57.27 3.485 57.655 3.6 ;
      RECT 57.275 2.207 57.31 2.445 ;
      RECT 57.275 2.207 57.34 2.444 ;
      RECT 57.275 2.207 57.455 2.44 ;
      RECT 57.275 2.207 57.51 2.418 ;
      RECT 57.285 2.15 57.565 2.318 ;
      RECT 57.39 1.99 57.42 2.441 ;
      RECT 57.42 1.985 57.6 2.198 ;
      RECT 57.29 2.126 57.6 2.198 ;
      RECT 57.34 2.022 57.39 2.442 ;
      RECT 57.31 2.078 57.6 2.198 ;
      RECT 55.815 1.74 55.985 2.935 ;
      RECT 55.815 1.74 56.28 1.91 ;
      RECT 55.815 6.97 56.28 7.14 ;
      RECT 55.815 5.945 55.985 7.14 ;
      RECT 54.825 1.74 54.995 2.935 ;
      RECT 54.825 1.74 55.29 1.91 ;
      RECT 54.825 6.97 55.29 7.14 ;
      RECT 54.825 5.945 54.995 7.14 ;
      RECT 52.97 2.635 53.14 3.865 ;
      RECT 53.025 0.855 53.195 2.805 ;
      RECT 52.97 0.575 53.14 1.025 ;
      RECT 52.97 7.855 53.14 8.305 ;
      RECT 53.025 6.075 53.195 8.025 ;
      RECT 52.97 5.015 53.14 6.245 ;
      RECT 52.45 0.575 52.62 3.865 ;
      RECT 52.45 2.075 52.855 2.405 ;
      RECT 52.45 1.235 52.855 1.565 ;
      RECT 52.45 5.015 52.62 8.305 ;
      RECT 52.45 7.315 52.855 7.645 ;
      RECT 52.45 6.475 52.855 6.805 ;
      RECT 50.55 3.392 50.565 3.443 ;
      RECT 50.545 3.372 50.55 3.49 ;
      RECT 50.53 3.362 50.545 3.558 ;
      RECT 50.505 3.342 50.53 3.613 ;
      RECT 50.465 3.327 50.505 3.633 ;
      RECT 50.42 3.321 50.465 3.661 ;
      RECT 50.35 3.311 50.42 3.678 ;
      RECT 50.33 3.303 50.35 3.678 ;
      RECT 50.27 3.297 50.33 3.67 ;
      RECT 50.211 3.288 50.27 3.658 ;
      RECT 50.125 3.277 50.211 3.641 ;
      RECT 50.103 3.268 50.125 3.629 ;
      RECT 50.017 3.261 50.103 3.616 ;
      RECT 49.931 3.248 50.017 3.597 ;
      RECT 49.845 3.236 49.931 3.577 ;
      RECT 49.815 3.225 49.845 3.564 ;
      RECT 49.765 3.211 49.815 3.556 ;
      RECT 49.745 3.2 49.765 3.548 ;
      RECT 49.696 3.189 49.745 3.54 ;
      RECT 49.61 3.168 49.696 3.525 ;
      RECT 49.565 3.155 49.61 3.51 ;
      RECT 49.52 3.155 49.565 3.49 ;
      RECT 49.465 3.155 49.52 3.425 ;
      RECT 49.44 3.155 49.465 3.348 ;
      RECT 49.965 2.892 50.135 3.075 ;
      RECT 49.965 2.892 50.15 3.033 ;
      RECT 49.965 2.892 50.155 2.975 ;
      RECT 50.025 2.66 50.16 2.951 ;
      RECT 50.025 2.664 50.165 2.934 ;
      RECT 49.97 2.827 50.165 2.934 ;
      RECT 49.995 2.672 50.135 3.075 ;
      RECT 49.995 2.676 50.175 2.875 ;
      RECT 49.98 2.762 50.175 2.875 ;
      RECT 49.99 2.692 50.135 3.075 ;
      RECT 49.99 2.695 50.185 2.788 ;
      RECT 49.985 2.712 50.185 2.788 ;
      RECT 49.755 1.932 49.925 2.415 ;
      RECT 49.75 1.927 49.9 2.405 ;
      RECT 49.75 1.934 49.93 2.399 ;
      RECT 49.74 1.928 49.9 2.378 ;
      RECT 49.74 1.944 49.945 2.337 ;
      RECT 49.71 1.929 49.9 2.3 ;
      RECT 49.71 1.959 49.955 2.24 ;
      RECT 49.705 1.931 49.9 2.238 ;
      RECT 49.685 1.94 49.93 2.195 ;
      RECT 49.66 1.956 49.945 2.107 ;
      RECT 49.66 1.975 49.97 2.098 ;
      RECT 49.655 2.012 49.97 2.05 ;
      RECT 49.66 1.992 49.975 2.018 ;
      RECT 49.755 1.926 49.865 2.415 ;
      RECT 49.841 1.925 49.865 2.415 ;
      RECT 49.075 2.71 49.08 2.921 ;
      RECT 49.675 2.71 49.68 2.895 ;
      RECT 49.74 2.75 49.745 2.863 ;
      RECT 49.735 2.742 49.74 2.869 ;
      RECT 49.73 2.732 49.735 2.877 ;
      RECT 49.725 2.722 49.73 2.886 ;
      RECT 49.72 2.712 49.725 2.89 ;
      RECT 49.68 2.71 49.72 2.893 ;
      RECT 49.652 2.709 49.675 2.897 ;
      RECT 49.566 2.706 49.652 2.904 ;
      RECT 49.48 2.702 49.566 2.915 ;
      RECT 49.46 2.7 49.48 2.921 ;
      RECT 49.442 2.699 49.46 2.924 ;
      RECT 49.356 2.697 49.442 2.931 ;
      RECT 49.27 2.692 49.356 2.944 ;
      RECT 49.251 2.689 49.27 2.949 ;
      RECT 49.165 2.687 49.251 2.94 ;
      RECT 49.155 2.687 49.165 2.933 ;
      RECT 49.08 2.7 49.155 2.927 ;
      RECT 49.065 2.711 49.075 2.921 ;
      RECT 49.055 2.713 49.065 2.92 ;
      RECT 49.045 2.717 49.055 2.916 ;
      RECT 49.04 2.72 49.045 2.91 ;
      RECT 49.03 2.722 49.04 2.904 ;
      RECT 49.025 2.725 49.03 2.898 ;
      RECT 49.005 3.311 49.01 3.515 ;
      RECT 48.99 3.298 49.005 3.608 ;
      RECT 48.975 3.279 48.99 3.885 ;
      RECT 48.94 3.245 48.975 3.885 ;
      RECT 48.936 3.215 48.94 3.885 ;
      RECT 48.85 3.097 48.936 3.885 ;
      RECT 48.84 2.972 48.85 3.885 ;
      RECT 48.825 2.94 48.84 3.885 ;
      RECT 48.82 2.915 48.825 3.885 ;
      RECT 48.815 2.905 48.82 3.841 ;
      RECT 48.8 2.877 48.815 3.746 ;
      RECT 48.785 2.843 48.8 3.645 ;
      RECT 48.78 2.821 48.785 3.598 ;
      RECT 48.775 2.81 48.78 3.568 ;
      RECT 48.77 2.8 48.775 3.534 ;
      RECT 48.76 2.787 48.77 3.502 ;
      RECT 48.735 2.763 48.76 3.428 ;
      RECT 48.73 2.743 48.735 3.353 ;
      RECT 48.725 2.737 48.73 3.328 ;
      RECT 48.72 2.732 48.725 3.293 ;
      RECT 48.715 2.727 48.72 3.268 ;
      RECT 48.71 2.725 48.715 3.248 ;
      RECT 48.705 2.725 48.71 3.233 ;
      RECT 48.7 2.725 48.705 3.193 ;
      RECT 48.69 2.725 48.7 3.165 ;
      RECT 48.68 2.725 48.69 3.11 ;
      RECT 48.665 2.725 48.68 3.048 ;
      RECT 48.66 2.724 48.665 2.993 ;
      RECT 48.645 2.723 48.66 2.973 ;
      RECT 48.585 2.721 48.645 2.947 ;
      RECT 48.55 2.722 48.585 2.927 ;
      RECT 48.545 2.724 48.55 2.917 ;
      RECT 48.535 2.743 48.545 2.907 ;
      RECT 48.53 2.77 48.535 2.838 ;
      RECT 48.645 2.195 48.815 2.44 ;
      RECT 48.68 1.966 48.815 2.44 ;
      RECT 48.68 1.968 48.825 2.435 ;
      RECT 48.68 1.97 48.85 2.423 ;
      RECT 48.68 1.973 48.875 2.405 ;
      RECT 48.68 1.978 48.925 2.378 ;
      RECT 48.68 1.983 48.945 2.343 ;
      RECT 48.66 1.985 48.955 2.318 ;
      RECT 48.65 2.08 48.955 2.318 ;
      RECT 48.68 1.965 48.79 2.44 ;
      RECT 48.69 1.962 48.785 2.44 ;
      RECT 48.21 3.227 48.4 3.585 ;
      RECT 48.21 3.239 48.435 3.584 ;
      RECT 48.21 3.267 48.455 3.582 ;
      RECT 48.21 3.292 48.46 3.581 ;
      RECT 48.21 3.35 48.475 3.58 ;
      RECT 48.195 3.223 48.355 3.565 ;
      RECT 48.175 3.232 48.4 3.518 ;
      RECT 48.15 3.243 48.435 3.455 ;
      RECT 48.15 3.327 48.47 3.455 ;
      RECT 48.15 3.302 48.465 3.455 ;
      RECT 48.21 3.218 48.355 3.585 ;
      RECT 48.296 3.217 48.355 3.585 ;
      RECT 48.296 3.216 48.34 3.585 ;
      RECT 48.21 7.855 48.38 8.305 ;
      RECT 48.265 6.075 48.435 8.025 ;
      RECT 48.21 5.015 48.38 6.245 ;
      RECT 47.69 5.015 47.86 8.305 ;
      RECT 47.69 7.315 48.095 7.645 ;
      RECT 47.69 6.475 48.095 6.805 ;
      RECT 47.995 2.732 48 3.11 ;
      RECT 47.99 2.7 47.995 3.11 ;
      RECT 47.985 2.672 47.99 3.11 ;
      RECT 47.98 2.652 47.985 3.11 ;
      RECT 47.925 2.635 47.98 3.11 ;
      RECT 47.885 2.62 47.925 3.11 ;
      RECT 47.83 2.607 47.885 3.11 ;
      RECT 47.795 2.598 47.83 3.11 ;
      RECT 47.791 2.596 47.795 3.109 ;
      RECT 47.705 2.592 47.791 3.092 ;
      RECT 47.62 2.584 47.705 3.055 ;
      RECT 47.61 2.58 47.62 3.028 ;
      RECT 47.6 2.58 47.61 3.01 ;
      RECT 47.59 2.582 47.6 2.993 ;
      RECT 47.585 2.587 47.59 2.979 ;
      RECT 47.58 2.591 47.585 2.966 ;
      RECT 47.57 2.596 47.58 2.95 ;
      RECT 47.555 2.61 47.57 2.925 ;
      RECT 47.55 2.616 47.555 2.905 ;
      RECT 47.545 2.618 47.55 2.898 ;
      RECT 47.54 2.622 47.545 2.773 ;
      RECT 47.72 3.422 47.965 3.885 ;
      RECT 47.64 3.395 47.96 3.881 ;
      RECT 47.57 3.43 47.965 3.874 ;
      RECT 47.36 3.685 47.965 3.87 ;
      RECT 47.54 3.453 47.965 3.87 ;
      RECT 47.38 3.645 47.965 3.87 ;
      RECT 47.53 3.465 47.965 3.87 ;
      RECT 47.415 3.582 47.965 3.87 ;
      RECT 47.47 3.507 47.965 3.87 ;
      RECT 47.72 3.372 47.96 3.885 ;
      RECT 47.75 3.365 47.96 3.885 ;
      RECT 47.74 3.367 47.96 3.885 ;
      RECT 47.75 3.362 47.88 3.885 ;
      RECT 47.305 1.925 47.391 2.364 ;
      RECT 47.3 1.925 47.391 2.362 ;
      RECT 47.3 1.925 47.46 2.361 ;
      RECT 47.3 1.925 47.49 2.358 ;
      RECT 47.285 1.932 47.49 2.349 ;
      RECT 47.285 1.932 47.495 2.345 ;
      RECT 47.28 1.942 47.495 2.338 ;
      RECT 47.275 1.947 47.495 2.313 ;
      RECT 47.275 1.947 47.51 2.295 ;
      RECT 47.3 1.925 47.53 2.21 ;
      RECT 47.27 1.952 47.53 2.208 ;
      RECT 47.28 1.945 47.535 2.146 ;
      RECT 47.27 2.067 47.54 2.129 ;
      RECT 47.255 1.962 47.535 2.08 ;
      RECT 47.25 1.972 47.535 1.98 ;
      RECT 47.33 2.743 47.335 2.82 ;
      RECT 47.32 2.737 47.33 3.01 ;
      RECT 47.31 2.729 47.32 3.031 ;
      RECT 47.3 2.72 47.31 3.053 ;
      RECT 47.295 2.715 47.3 3.07 ;
      RECT 47.255 2.715 47.295 3.11 ;
      RECT 47.235 2.715 47.255 3.165 ;
      RECT 47.23 2.715 47.235 3.193 ;
      RECT 47.22 2.715 47.23 3.208 ;
      RECT 47.185 2.715 47.22 3.25 ;
      RECT 47.18 2.715 47.185 3.293 ;
      RECT 47.17 2.715 47.18 3.308 ;
      RECT 47.155 2.715 47.17 3.328 ;
      RECT 47.14 2.715 47.155 3.355 ;
      RECT 47.135 2.716 47.14 3.373 ;
      RECT 47.115 2.717 47.135 3.38 ;
      RECT 47.06 2.718 47.115 3.4 ;
      RECT 47.05 2.719 47.06 3.414 ;
      RECT 47.045 2.722 47.05 3.413 ;
      RECT 47.005 2.795 47.045 3.411 ;
      RECT 46.99 2.875 47.005 3.409 ;
      RECT 46.965 2.93 46.99 3.407 ;
      RECT 46.95 2.995 46.965 3.406 ;
      RECT 46.905 3.027 46.95 3.403 ;
      RECT 46.82 3.05 46.905 3.398 ;
      RECT 46.795 3.07 46.82 3.393 ;
      RECT 46.725 3.075 46.795 3.389 ;
      RECT 46.705 3.077 46.725 3.386 ;
      RECT 46.62 3.088 46.705 3.38 ;
      RECT 46.615 3.099 46.62 3.375 ;
      RECT 46.605 3.101 46.615 3.375 ;
      RECT 46.57 3.105 46.605 3.373 ;
      RECT 46.52 3.115 46.57 3.36 ;
      RECT 46.5 3.123 46.52 3.345 ;
      RECT 46.42 3.135 46.5 3.328 ;
      RECT 46.585 2.685 46.755 2.895 ;
      RECT 46.701 2.681 46.755 2.895 ;
      RECT 46.506 2.685 46.755 2.886 ;
      RECT 46.506 2.685 46.76 2.875 ;
      RECT 46.42 2.685 46.76 2.866 ;
      RECT 46.42 2.693 46.77 2.81 ;
      RECT 46.42 2.705 46.775 2.723 ;
      RECT 46.42 2.712 46.78 2.715 ;
      RECT 46.615 2.683 46.755 2.895 ;
      RECT 46.37 3.628 46.615 3.96 ;
      RECT 46.365 3.62 46.37 3.957 ;
      RECT 46.335 3.64 46.615 3.938 ;
      RECT 46.315 3.672 46.615 3.911 ;
      RECT 46.365 3.625 46.542 3.957 ;
      RECT 46.365 3.622 46.456 3.957 ;
      RECT 46.305 1.97 46.475 2.39 ;
      RECT 46.3 1.97 46.475 2.388 ;
      RECT 46.3 1.97 46.5 2.378 ;
      RECT 46.3 1.97 46.52 2.353 ;
      RECT 46.295 1.97 46.52 2.348 ;
      RECT 46.295 1.97 46.53 2.338 ;
      RECT 46.295 1.97 46.535 2.333 ;
      RECT 46.295 1.975 46.54 2.328 ;
      RECT 46.295 2.007 46.555 2.318 ;
      RECT 46.295 2.077 46.58 2.301 ;
      RECT 46.275 2.077 46.58 2.293 ;
      RECT 46.275 2.137 46.59 2.27 ;
      RECT 46.275 2.177 46.6 2.215 ;
      RECT 46.26 1.97 46.535 2.195 ;
      RECT 46.25 1.985 46.54 2.093 ;
      RECT 45.84 3.375 46.01 3.9 ;
      RECT 45.835 3.375 46.01 3.893 ;
      RECT 45.825 3.375 46.015 3.858 ;
      RECT 45.82 3.385 46.015 3.83 ;
      RECT 45.815 3.405 46.015 3.813 ;
      RECT 45.825 3.38 46.02 3.803 ;
      RECT 45.81 3.425 46.02 3.795 ;
      RECT 45.805 3.445 46.02 3.78 ;
      RECT 45.8 3.475 46.02 3.77 ;
      RECT 45.79 3.52 46.02 3.745 ;
      RECT 45.82 3.39 46.025 3.728 ;
      RECT 45.785 3.572 46.025 3.723 ;
      RECT 45.82 3.4 46.03 3.693 ;
      RECT 45.78 3.605 46.03 3.69 ;
      RECT 45.775 3.63 46.03 3.67 ;
      RECT 45.815 3.417 46.04 3.61 ;
      RECT 45.81 3.439 46.05 3.503 ;
      RECT 45.76 2.686 45.775 2.955 ;
      RECT 45.715 2.67 45.76 3 ;
      RECT 45.71 2.658 45.715 3.05 ;
      RECT 45.7 2.654 45.71 3.083 ;
      RECT 45.695 2.651 45.7 3.111 ;
      RECT 45.68 2.653 45.695 3.153 ;
      RECT 45.675 2.657 45.68 3.193 ;
      RECT 45.655 2.662 45.675 3.245 ;
      RECT 45.651 2.667 45.655 3.302 ;
      RECT 45.565 2.686 45.651 3.339 ;
      RECT 45.555 2.707 45.565 3.375 ;
      RECT 45.55 2.715 45.555 3.376 ;
      RECT 45.545 2.757 45.55 3.377 ;
      RECT 45.53 2.845 45.545 3.378 ;
      RECT 45.52 2.995 45.53 3.38 ;
      RECT 45.515 3.04 45.52 3.382 ;
      RECT 45.48 3.082 45.515 3.385 ;
      RECT 45.475 3.1 45.48 3.388 ;
      RECT 45.398 3.106 45.475 3.394 ;
      RECT 45.312 3.12 45.398 3.407 ;
      RECT 45.226 3.134 45.312 3.421 ;
      RECT 45.14 3.148 45.226 3.434 ;
      RECT 45.08 3.16 45.14 3.446 ;
      RECT 45.055 3.167 45.08 3.453 ;
      RECT 45.041 3.17 45.055 3.458 ;
      RECT 44.955 3.178 45.041 3.474 ;
      RECT 44.95 3.185 44.955 3.489 ;
      RECT 44.926 3.185 44.95 3.496 ;
      RECT 44.84 3.188 44.926 3.524 ;
      RECT 44.755 3.192 44.84 3.568 ;
      RECT 44.69 3.196 44.755 3.605 ;
      RECT 44.665 3.199 44.69 3.621 ;
      RECT 44.59 3.212 44.665 3.625 ;
      RECT 44.565 3.23 44.59 3.629 ;
      RECT 44.555 3.237 44.565 3.631 ;
      RECT 44.54 3.24 44.555 3.632 ;
      RECT 44.48 3.252 44.54 3.636 ;
      RECT 44.47 3.266 44.48 3.64 ;
      RECT 44.415 3.276 44.47 3.628 ;
      RECT 44.39 3.297 44.415 3.611 ;
      RECT 44.37 3.317 44.39 3.602 ;
      RECT 44.365 3.33 44.37 3.597 ;
      RECT 44.35 3.342 44.365 3.593 ;
      RECT 45.585 1.997 45.59 2.02 ;
      RECT 45.58 1.988 45.585 2.06 ;
      RECT 45.575 1.986 45.58 2.103 ;
      RECT 45.57 1.977 45.575 2.138 ;
      RECT 45.565 1.967 45.57 2.21 ;
      RECT 45.56 1.957 45.565 2.275 ;
      RECT 45.555 1.954 45.56 2.315 ;
      RECT 45.53 1.948 45.555 2.405 ;
      RECT 45.495 1.936 45.53 2.43 ;
      RECT 45.485 1.927 45.495 2.43 ;
      RECT 45.35 1.925 45.36 2.413 ;
      RECT 45.34 1.925 45.35 2.38 ;
      RECT 45.335 1.925 45.34 2.355 ;
      RECT 45.33 1.925 45.335 2.343 ;
      RECT 45.325 1.925 45.33 2.325 ;
      RECT 45.315 1.925 45.325 2.29 ;
      RECT 45.31 1.927 45.315 2.268 ;
      RECT 45.305 1.933 45.31 2.253 ;
      RECT 45.3 1.939 45.305 2.238 ;
      RECT 45.285 1.951 45.3 2.211 ;
      RECT 45.28 1.962 45.285 2.179 ;
      RECT 45.275 1.972 45.28 2.163 ;
      RECT 45.265 1.98 45.275 2.132 ;
      RECT 45.26 1.99 45.265 2.106 ;
      RECT 45.255 2.047 45.26 2.089 ;
      RECT 45.36 1.925 45.485 2.43 ;
      RECT 45.075 2.612 45.335 2.91 ;
      RECT 45.07 2.619 45.335 2.908 ;
      RECT 45.075 2.614 45.35 2.903 ;
      RECT 45.065 2.627 45.35 2.9 ;
      RECT 45.065 2.632 45.355 2.893 ;
      RECT 45.06 2.64 45.355 2.89 ;
      RECT 45.06 2.657 45.36 2.688 ;
      RECT 45.075 2.609 45.306 2.91 ;
      RECT 45.13 2.608 45.306 2.91 ;
      RECT 45.13 2.605 45.22 2.91 ;
      RECT 45.13 2.602 45.216 2.91 ;
      RECT 44.82 2.875 44.825 2.888 ;
      RECT 44.815 2.842 44.82 2.893 ;
      RECT 44.81 2.797 44.815 2.9 ;
      RECT 44.805 2.752 44.81 2.908 ;
      RECT 44.8 2.72 44.805 2.916 ;
      RECT 44.795 2.68 44.8 2.917 ;
      RECT 44.78 2.66 44.795 2.919 ;
      RECT 44.705 2.642 44.78 2.931 ;
      RECT 44.695 2.635 44.705 2.942 ;
      RECT 44.69 2.635 44.695 2.944 ;
      RECT 44.66 2.641 44.69 2.948 ;
      RECT 44.62 2.654 44.66 2.948 ;
      RECT 44.595 2.665 44.62 2.934 ;
      RECT 44.58 2.671 44.595 2.917 ;
      RECT 44.57 2.673 44.58 2.908 ;
      RECT 44.565 2.674 44.57 2.903 ;
      RECT 44.56 2.675 44.565 2.898 ;
      RECT 44.555 2.676 44.56 2.895 ;
      RECT 44.53 2.681 44.555 2.885 ;
      RECT 44.52 2.697 44.53 2.872 ;
      RECT 44.515 2.717 44.52 2.867 ;
      RECT 44.525 2.11 44.53 2.306 ;
      RECT 44.51 2.074 44.525 2.308 ;
      RECT 44.5 2.056 44.51 2.313 ;
      RECT 44.49 2.042 44.5 2.317 ;
      RECT 44.445 2.026 44.49 2.327 ;
      RECT 44.44 2.016 44.445 2.336 ;
      RECT 44.395 2.005 44.44 2.342 ;
      RECT 44.39 1.993 44.395 2.349 ;
      RECT 44.375 1.988 44.39 2.353 ;
      RECT 44.36 1.98 44.375 2.358 ;
      RECT 44.35 1.973 44.36 2.363 ;
      RECT 44.34 1.97 44.35 2.368 ;
      RECT 44.33 1.97 44.34 2.369 ;
      RECT 44.325 1.967 44.33 2.368 ;
      RECT 44.29 1.962 44.315 2.367 ;
      RECT 44.266 1.958 44.29 2.366 ;
      RECT 44.18 1.949 44.266 2.363 ;
      RECT 44.165 1.941 44.18 2.36 ;
      RECT 44.143 1.94 44.165 2.359 ;
      RECT 44.057 1.94 44.143 2.357 ;
      RECT 43.971 1.94 44.057 2.355 ;
      RECT 43.885 1.94 43.971 2.352 ;
      RECT 43.875 1.94 43.885 2.343 ;
      RECT 43.845 1.94 43.875 2.303 ;
      RECT 43.835 1.95 43.845 2.258 ;
      RECT 43.83 1.99 43.835 2.243 ;
      RECT 43.825 2.005 43.83 2.23 ;
      RECT 43.795 2.085 43.825 2.192 ;
      RECT 44.315 1.965 44.325 2.368 ;
      RECT 44.14 2.73 44.155 3.335 ;
      RECT 44.145 2.725 44.155 3.335 ;
      RECT 44.31 2.725 44.315 2.908 ;
      RECT 44.3 2.725 44.31 2.938 ;
      RECT 44.285 2.725 44.3 2.998 ;
      RECT 44.28 2.725 44.285 3.043 ;
      RECT 44.275 2.725 44.28 3.073 ;
      RECT 44.27 2.725 44.275 3.093 ;
      RECT 44.26 2.725 44.27 3.128 ;
      RECT 44.245 2.725 44.26 3.16 ;
      RECT 44.2 2.725 44.245 3.188 ;
      RECT 44.195 2.725 44.2 3.218 ;
      RECT 44.19 2.725 44.195 3.23 ;
      RECT 44.185 2.725 44.19 3.238 ;
      RECT 44.175 2.725 44.185 3.253 ;
      RECT 44.17 2.725 44.175 3.275 ;
      RECT 44.16 2.725 44.17 3.298 ;
      RECT 44.155 2.725 44.16 3.318 ;
      RECT 44.12 2.74 44.14 3.335 ;
      RECT 44.095 2.757 44.12 3.335 ;
      RECT 44.09 2.767 44.095 3.335 ;
      RECT 44.06 2.782 44.09 3.335 ;
      RECT 43.985 2.824 44.06 3.335 ;
      RECT 43.98 2.855 43.985 3.318 ;
      RECT 43.975 2.859 43.98 3.3 ;
      RECT 43.97 2.863 43.975 3.263 ;
      RECT 43.965 3.047 43.97 3.23 ;
      RECT 43.45 3.236 43.536 3.801 ;
      RECT 43.405 3.238 43.57 3.795 ;
      RECT 43.536 3.235 43.57 3.795 ;
      RECT 43.45 3.237 43.655 3.789 ;
      RECT 43.405 3.247 43.665 3.785 ;
      RECT 43.38 3.239 43.655 3.781 ;
      RECT 43.375 3.242 43.655 3.776 ;
      RECT 43.35 3.257 43.665 3.77 ;
      RECT 43.35 3.282 43.705 3.765 ;
      RECT 43.31 3.29 43.705 3.74 ;
      RECT 43.31 3.317 43.72 3.738 ;
      RECT 43.31 3.347 43.73 3.725 ;
      RECT 43.305 3.492 43.73 3.713 ;
      RECT 43.31 3.421 43.75 3.71 ;
      RECT 43.31 3.478 43.755 3.518 ;
      RECT 43.5 2.757 43.67 2.935 ;
      RECT 43.45 2.696 43.5 2.92 ;
      RECT 43.185 2.676 43.45 2.905 ;
      RECT 43.145 2.74 43.62 2.905 ;
      RECT 43.145 2.73 43.575 2.905 ;
      RECT 43.145 2.727 43.565 2.905 ;
      RECT 43.145 2.715 43.555 2.905 ;
      RECT 43.145 2.7 43.5 2.905 ;
      RECT 43.185 2.672 43.386 2.905 ;
      RECT 43.195 2.65 43.386 2.905 ;
      RECT 43.22 2.635 43.3 2.905 ;
      RECT 42.975 3.165 43.095 3.61 ;
      RECT 42.96 3.165 43.095 3.609 ;
      RECT 42.915 3.187 43.095 3.604 ;
      RECT 42.875 3.236 43.095 3.598 ;
      RECT 42.875 3.236 43.1 3.573 ;
      RECT 42.875 3.236 43.12 3.463 ;
      RECT 42.87 3.266 43.12 3.46 ;
      RECT 42.96 3.165 43.13 3.355 ;
      RECT 42.62 1.95 42.625 2.395 ;
      RECT 42.43 1.95 42.45 2.36 ;
      RECT 42.4 1.95 42.405 2.335 ;
      RECT 43.08 2.257 43.095 2.445 ;
      RECT 43.075 2.242 43.08 2.451 ;
      RECT 43.055 2.215 43.075 2.454 ;
      RECT 43.005 2.182 43.055 2.463 ;
      RECT 42.975 2.162 43.005 2.467 ;
      RECT 42.956 2.15 42.975 2.463 ;
      RECT 42.87 2.122 42.956 2.453 ;
      RECT 42.86 2.097 42.87 2.443 ;
      RECT 42.79 2.065 42.86 2.435 ;
      RECT 42.765 2.025 42.79 2.427 ;
      RECT 42.745 2.007 42.765 2.421 ;
      RECT 42.735 1.997 42.745 2.418 ;
      RECT 42.725 1.99 42.735 2.416 ;
      RECT 42.705 1.977 42.725 2.413 ;
      RECT 42.695 1.967 42.705 2.41 ;
      RECT 42.685 1.96 42.695 2.408 ;
      RECT 42.635 1.952 42.685 2.402 ;
      RECT 42.625 1.95 42.635 2.396 ;
      RECT 42.595 1.95 42.62 2.393 ;
      RECT 42.566 1.95 42.595 2.388 ;
      RECT 42.48 1.95 42.566 2.378 ;
      RECT 42.45 1.95 42.48 2.365 ;
      RECT 42.405 1.95 42.43 2.348 ;
      RECT 42.39 1.95 42.4 2.33 ;
      RECT 42.37 1.957 42.39 2.315 ;
      RECT 42.365 1.972 42.37 2.303 ;
      RECT 42.36 1.977 42.365 2.243 ;
      RECT 42.355 1.982 42.36 2.085 ;
      RECT 42.35 1.985 42.355 2.003 ;
      RECT 42.615 2.67 42.701 2.991 ;
      RECT 42.615 2.67 42.735 2.984 ;
      RECT 42.565 2.67 42.735 2.98 ;
      RECT 42.565 2.672 42.821 2.978 ;
      RECT 42.565 2.674 42.845 2.972 ;
      RECT 42.565 2.681 42.855 2.971 ;
      RECT 42.565 2.69 42.86 2.968 ;
      RECT 42.565 2.696 42.865 2.963 ;
      RECT 42.565 2.74 42.87 2.96 ;
      RECT 42.565 2.832 42.875 2.957 ;
      RECT 42.09 3.275 42.125 3.595 ;
      RECT 42.675 3.46 42.68 3.642 ;
      RECT 42.63 3.342 42.675 3.661 ;
      RECT 42.615 3.319 42.63 3.684 ;
      RECT 42.605 3.309 42.615 3.694 ;
      RECT 42.585 3.304 42.605 3.707 ;
      RECT 42.56 3.302 42.585 3.728 ;
      RECT 42.541 3.301 42.56 3.74 ;
      RECT 42.455 3.298 42.541 3.74 ;
      RECT 42.385 3.293 42.455 3.728 ;
      RECT 42.31 3.289 42.385 3.703 ;
      RECT 42.245 3.285 42.31 3.67 ;
      RECT 42.175 3.282 42.245 3.63 ;
      RECT 42.145 3.278 42.175 3.605 ;
      RECT 42.125 3.276 42.145 3.598 ;
      RECT 42.041 3.274 42.09 3.596 ;
      RECT 41.955 3.271 42.041 3.597 ;
      RECT 41.88 3.27 41.955 3.599 ;
      RECT 41.795 3.27 41.88 3.625 ;
      RECT 41.718 3.271 41.795 3.65 ;
      RECT 41.632 3.272 41.718 3.65 ;
      RECT 41.546 3.272 41.632 3.65 ;
      RECT 41.46 3.273 41.546 3.65 ;
      RECT 41.44 3.274 41.46 3.642 ;
      RECT 41.425 3.28 41.44 3.627 ;
      RECT 41.39 3.3 41.425 3.607 ;
      RECT 41.38 3.32 41.39 3.589 ;
      RECT 42.35 2.625 42.355 2.895 ;
      RECT 42.345 2.616 42.35 2.9 ;
      RECT 42.335 2.606 42.345 2.912 ;
      RECT 42.33 2.595 42.335 2.923 ;
      RECT 42.31 2.589 42.33 2.941 ;
      RECT 42.265 2.586 42.31 2.99 ;
      RECT 42.25 2.585 42.265 3.035 ;
      RECT 42.245 2.585 42.25 3.048 ;
      RECT 42.235 2.585 42.245 3.06 ;
      RECT 42.23 2.586 42.235 3.075 ;
      RECT 42.21 2.594 42.23 3.08 ;
      RECT 42.18 2.61 42.21 3.08 ;
      RECT 42.17 2.622 42.175 3.08 ;
      RECT 42.135 2.637 42.17 3.08 ;
      RECT 42.105 2.657 42.135 3.08 ;
      RECT 42.095 2.682 42.105 3.08 ;
      RECT 42.09 2.71 42.095 3.08 ;
      RECT 42.085 2.74 42.09 3.08 ;
      RECT 42.08 2.757 42.085 3.08 ;
      RECT 42.07 2.785 42.08 3.08 ;
      RECT 42.06 2.82 42.07 3.08 ;
      RECT 42.055 2.855 42.06 3.08 ;
      RECT 42.175 2.62 42.18 3.08 ;
      RECT 41.69 2.722 41.875 2.895 ;
      RECT 41.65 2.64 41.835 2.893 ;
      RECT 41.611 2.645 41.835 2.889 ;
      RECT 41.525 2.654 41.835 2.884 ;
      RECT 41.441 2.67 41.84 2.879 ;
      RECT 41.355 2.69 41.865 2.873 ;
      RECT 41.355 2.71 41.87 2.873 ;
      RECT 41.441 2.68 41.865 2.879 ;
      RECT 41.525 2.655 41.84 2.884 ;
      RECT 41.69 2.637 41.835 2.895 ;
      RECT 41.69 2.632 41.79 2.895 ;
      RECT 41.776 2.626 41.79 2.895 ;
      RECT 41.165 1.95 41.17 2.349 ;
      RECT 40.91 1.95 40.945 2.347 ;
      RECT 40.505 1.985 40.51 2.341 ;
      RECT 41.25 1.988 41.255 2.243 ;
      RECT 41.245 1.986 41.25 2.249 ;
      RECT 41.24 1.985 41.245 2.256 ;
      RECT 41.215 1.978 41.24 2.28 ;
      RECT 41.21 1.971 41.215 2.304 ;
      RECT 41.205 1.967 41.21 2.313 ;
      RECT 41.195 1.962 41.205 2.326 ;
      RECT 41.19 1.959 41.195 2.335 ;
      RECT 41.185 1.957 41.19 2.34 ;
      RECT 41.17 1.953 41.185 2.35 ;
      RECT 41.155 1.947 41.165 2.349 ;
      RECT 41.117 1.945 41.155 2.349 ;
      RECT 41.031 1.947 41.117 2.349 ;
      RECT 40.945 1.949 41.031 2.348 ;
      RECT 40.874 1.95 40.91 2.347 ;
      RECT 40.788 1.952 40.874 2.347 ;
      RECT 40.702 1.954 40.788 2.346 ;
      RECT 40.616 1.956 40.702 2.346 ;
      RECT 40.53 1.959 40.616 2.345 ;
      RECT 40.52 1.965 40.53 2.344 ;
      RECT 40.51 1.977 40.52 2.342 ;
      RECT 40.45 2.012 40.505 2.338 ;
      RECT 40.445 2.042 40.45 2.1 ;
      RECT 41.19 3.122 41.205 3.315 ;
      RECT 41.185 3.09 41.19 3.315 ;
      RECT 41.175 3.065 41.185 3.315 ;
      RECT 41.17 3.037 41.175 3.315 ;
      RECT 41.14 2.96 41.17 3.315 ;
      RECT 41.115 2.842 41.14 3.315 ;
      RECT 41.11 2.78 41.115 3.315 ;
      RECT 41.1 2.767 41.11 3.315 ;
      RECT 41.08 2.757 41.1 3.315 ;
      RECT 41.065 2.74 41.08 3.315 ;
      RECT 41.035 2.728 41.065 3.315 ;
      RECT 41.03 2.727 41.035 3.26 ;
      RECT 41.025 2.727 41.03 3.218 ;
      RECT 41.01 2.726 41.025 3.17 ;
      RECT 40.995 2.726 41.01 3.108 ;
      RECT 40.975 2.726 40.995 3.068 ;
      RECT 40.97 2.726 40.975 3.053 ;
      RECT 40.945 2.725 40.97 3.048 ;
      RECT 40.875 2.724 40.945 3.035 ;
      RECT 40.86 2.723 40.875 3.02 ;
      RECT 40.83 2.722 40.86 3.003 ;
      RECT 40.825 2.722 40.83 2.988 ;
      RECT 40.775 2.721 40.825 2.968 ;
      RECT 40.71 2.72 40.775 2.923 ;
      RECT 40.705 2.72 40.71 2.895 ;
      RECT 40.79 3.257 40.795 3.514 ;
      RECT 40.77 3.176 40.79 3.531 ;
      RECT 40.75 3.17 40.77 3.56 ;
      RECT 40.69 3.157 40.75 3.58 ;
      RECT 40.645 3.141 40.69 3.581 ;
      RECT 40.561 3.129 40.645 3.569 ;
      RECT 40.475 3.116 40.561 3.553 ;
      RECT 40.465 3.109 40.475 3.545 ;
      RECT 40.42 3.106 40.465 3.485 ;
      RECT 40.4 3.102 40.42 3.4 ;
      RECT 40.385 3.1 40.4 3.353 ;
      RECT 40.355 3.097 40.385 3.323 ;
      RECT 40.32 3.093 40.355 3.3 ;
      RECT 40.277 3.088 40.32 3.288 ;
      RECT 40.191 3.079 40.277 3.297 ;
      RECT 40.105 3.068 40.191 3.309 ;
      RECT 40.04 3.059 40.105 3.318 ;
      RECT 40.02 3.05 40.04 3.323 ;
      RECT 40.015 3.043 40.02 3.325 ;
      RECT 39.975 3.028 40.015 3.322 ;
      RECT 39.955 3.007 39.975 3.317 ;
      RECT 39.94 2.995 39.955 3.31 ;
      RECT 39.935 2.987 39.94 3.303 ;
      RECT 39.92 2.967 39.935 3.296 ;
      RECT 39.915 2.83 39.92 3.29 ;
      RECT 39.835 2.719 39.915 3.262 ;
      RECT 39.826 2.712 39.835 3.228 ;
      RECT 39.74 2.706 39.826 3.153 ;
      RECT 39.715 2.697 39.74 3.065 ;
      RECT 39.685 2.692 39.715 3.04 ;
      RECT 39.62 2.701 39.685 3.025 ;
      RECT 39.6 2.717 39.62 3 ;
      RECT 39.59 2.723 39.6 2.948 ;
      RECT 39.57 2.745 39.59 2.83 ;
      RECT 40.225 2.71 40.395 2.895 ;
      RECT 40.225 2.71 40.43 2.893 ;
      RECT 40.275 2.62 40.445 2.884 ;
      RECT 40.225 2.777 40.45 2.877 ;
      RECT 40.24 2.655 40.445 2.884 ;
      RECT 39.44 3.388 39.505 3.831 ;
      RECT 39.38 3.413 39.505 3.829 ;
      RECT 39.38 3.413 39.56 3.823 ;
      RECT 39.365 3.438 39.56 3.822 ;
      RECT 39.505 3.375 39.58 3.819 ;
      RECT 39.44 3.4 39.66 3.813 ;
      RECT 39.365 3.439 39.705 3.807 ;
      RECT 39.35 3.466 39.705 3.798 ;
      RECT 39.365 3.459 39.725 3.79 ;
      RECT 39.35 3.468 39.73 3.773 ;
      RECT 39.345 3.485 39.73 3.6 ;
      RECT 39.35 2.207 39.385 2.445 ;
      RECT 39.35 2.207 39.415 2.444 ;
      RECT 39.35 2.207 39.53 2.44 ;
      RECT 39.35 2.207 39.585 2.418 ;
      RECT 39.36 2.15 39.64 2.318 ;
      RECT 39.465 1.99 39.495 2.441 ;
      RECT 39.495 1.985 39.675 2.198 ;
      RECT 39.365 2.126 39.675 2.198 ;
      RECT 39.415 2.022 39.465 2.442 ;
      RECT 39.385 2.078 39.675 2.198 ;
      RECT 37.89 1.74 38.06 2.935 ;
      RECT 37.89 1.74 38.355 1.91 ;
      RECT 37.89 6.97 38.355 7.14 ;
      RECT 37.89 5.945 38.06 7.14 ;
      RECT 36.9 1.74 37.07 2.935 ;
      RECT 36.9 1.74 37.365 1.91 ;
      RECT 36.9 6.97 37.365 7.14 ;
      RECT 36.9 5.945 37.07 7.14 ;
      RECT 35.045 2.635 35.215 3.865 ;
      RECT 35.1 0.855 35.27 2.805 ;
      RECT 35.045 0.575 35.215 1.025 ;
      RECT 35.045 7.855 35.215 8.305 ;
      RECT 35.1 6.075 35.27 8.025 ;
      RECT 35.045 5.015 35.215 6.245 ;
      RECT 34.525 0.575 34.695 3.865 ;
      RECT 34.525 2.075 34.93 2.405 ;
      RECT 34.525 1.235 34.93 1.565 ;
      RECT 34.525 5.015 34.695 8.305 ;
      RECT 34.525 7.315 34.93 7.645 ;
      RECT 34.525 6.475 34.93 6.805 ;
      RECT 32.625 3.392 32.64 3.443 ;
      RECT 32.62 3.372 32.625 3.49 ;
      RECT 32.605 3.362 32.62 3.558 ;
      RECT 32.58 3.342 32.605 3.613 ;
      RECT 32.54 3.327 32.58 3.633 ;
      RECT 32.495 3.321 32.54 3.661 ;
      RECT 32.425 3.311 32.495 3.678 ;
      RECT 32.405 3.303 32.425 3.678 ;
      RECT 32.345 3.297 32.405 3.67 ;
      RECT 32.286 3.288 32.345 3.658 ;
      RECT 32.2 3.277 32.286 3.641 ;
      RECT 32.178 3.268 32.2 3.629 ;
      RECT 32.092 3.261 32.178 3.616 ;
      RECT 32.006 3.248 32.092 3.597 ;
      RECT 31.92 3.236 32.006 3.577 ;
      RECT 31.89 3.225 31.92 3.564 ;
      RECT 31.84 3.211 31.89 3.556 ;
      RECT 31.82 3.2 31.84 3.548 ;
      RECT 31.771 3.189 31.82 3.54 ;
      RECT 31.685 3.168 31.771 3.525 ;
      RECT 31.64 3.155 31.685 3.51 ;
      RECT 31.595 3.155 31.64 3.49 ;
      RECT 31.54 3.155 31.595 3.425 ;
      RECT 31.515 3.155 31.54 3.348 ;
      RECT 32.04 2.892 32.21 3.075 ;
      RECT 32.04 2.892 32.225 3.033 ;
      RECT 32.04 2.892 32.23 2.975 ;
      RECT 32.1 2.66 32.235 2.951 ;
      RECT 32.1 2.664 32.24 2.934 ;
      RECT 32.045 2.827 32.24 2.934 ;
      RECT 32.07 2.672 32.21 3.075 ;
      RECT 32.07 2.676 32.25 2.875 ;
      RECT 32.055 2.762 32.25 2.875 ;
      RECT 32.065 2.692 32.21 3.075 ;
      RECT 32.065 2.695 32.26 2.788 ;
      RECT 32.06 2.712 32.26 2.788 ;
      RECT 31.83 1.932 32 2.415 ;
      RECT 31.825 1.927 31.975 2.405 ;
      RECT 31.825 1.934 32.005 2.399 ;
      RECT 31.815 1.928 31.975 2.378 ;
      RECT 31.815 1.944 32.02 2.337 ;
      RECT 31.785 1.929 31.975 2.3 ;
      RECT 31.785 1.959 32.03 2.24 ;
      RECT 31.78 1.931 31.975 2.238 ;
      RECT 31.76 1.94 32.005 2.195 ;
      RECT 31.735 1.956 32.02 2.107 ;
      RECT 31.735 1.975 32.045 2.098 ;
      RECT 31.73 2.012 32.045 2.05 ;
      RECT 31.735 1.992 32.05 2.018 ;
      RECT 31.83 1.926 31.94 2.415 ;
      RECT 31.916 1.925 31.94 2.415 ;
      RECT 31.15 2.71 31.155 2.921 ;
      RECT 31.75 2.71 31.755 2.895 ;
      RECT 31.815 2.75 31.82 2.863 ;
      RECT 31.81 2.742 31.815 2.869 ;
      RECT 31.805 2.732 31.81 2.877 ;
      RECT 31.8 2.722 31.805 2.886 ;
      RECT 31.795 2.712 31.8 2.89 ;
      RECT 31.755 2.71 31.795 2.893 ;
      RECT 31.727 2.709 31.75 2.897 ;
      RECT 31.641 2.706 31.727 2.904 ;
      RECT 31.555 2.702 31.641 2.915 ;
      RECT 31.535 2.7 31.555 2.921 ;
      RECT 31.517 2.699 31.535 2.924 ;
      RECT 31.431 2.697 31.517 2.931 ;
      RECT 31.345 2.692 31.431 2.944 ;
      RECT 31.326 2.689 31.345 2.949 ;
      RECT 31.24 2.687 31.326 2.94 ;
      RECT 31.23 2.687 31.24 2.933 ;
      RECT 31.155 2.7 31.23 2.927 ;
      RECT 31.14 2.711 31.15 2.921 ;
      RECT 31.13 2.713 31.14 2.92 ;
      RECT 31.12 2.717 31.13 2.916 ;
      RECT 31.115 2.72 31.12 2.91 ;
      RECT 31.105 2.722 31.115 2.904 ;
      RECT 31.1 2.725 31.105 2.898 ;
      RECT 31.08 3.311 31.085 3.515 ;
      RECT 31.065 3.298 31.08 3.608 ;
      RECT 31.05 3.279 31.065 3.885 ;
      RECT 31.015 3.245 31.05 3.885 ;
      RECT 31.011 3.215 31.015 3.885 ;
      RECT 30.925 3.097 31.011 3.885 ;
      RECT 30.915 2.972 30.925 3.885 ;
      RECT 30.9 2.94 30.915 3.885 ;
      RECT 30.895 2.915 30.9 3.885 ;
      RECT 30.89 2.905 30.895 3.841 ;
      RECT 30.875 2.877 30.89 3.746 ;
      RECT 30.86 2.843 30.875 3.645 ;
      RECT 30.855 2.821 30.86 3.598 ;
      RECT 30.85 2.81 30.855 3.568 ;
      RECT 30.845 2.8 30.85 3.534 ;
      RECT 30.835 2.787 30.845 3.502 ;
      RECT 30.81 2.763 30.835 3.428 ;
      RECT 30.805 2.743 30.81 3.353 ;
      RECT 30.8 2.737 30.805 3.328 ;
      RECT 30.795 2.732 30.8 3.293 ;
      RECT 30.79 2.727 30.795 3.268 ;
      RECT 30.785 2.725 30.79 3.248 ;
      RECT 30.78 2.725 30.785 3.233 ;
      RECT 30.775 2.725 30.78 3.193 ;
      RECT 30.765 2.725 30.775 3.165 ;
      RECT 30.755 2.725 30.765 3.11 ;
      RECT 30.74 2.725 30.755 3.048 ;
      RECT 30.735 2.724 30.74 2.993 ;
      RECT 30.72 2.723 30.735 2.973 ;
      RECT 30.66 2.721 30.72 2.947 ;
      RECT 30.625 2.722 30.66 2.927 ;
      RECT 30.62 2.724 30.625 2.917 ;
      RECT 30.61 2.743 30.62 2.907 ;
      RECT 30.605 2.77 30.61 2.838 ;
      RECT 30.72 2.195 30.89 2.44 ;
      RECT 30.755 1.966 30.89 2.44 ;
      RECT 30.755 1.968 30.9 2.435 ;
      RECT 30.755 1.97 30.925 2.423 ;
      RECT 30.755 1.973 30.95 2.405 ;
      RECT 30.755 1.978 31 2.378 ;
      RECT 30.755 1.983 31.02 2.343 ;
      RECT 30.735 1.985 31.03 2.318 ;
      RECT 30.725 2.08 31.03 2.318 ;
      RECT 30.755 1.965 30.865 2.44 ;
      RECT 30.765 1.962 30.86 2.44 ;
      RECT 30.285 3.227 30.475 3.585 ;
      RECT 30.285 3.239 30.51 3.584 ;
      RECT 30.285 3.267 30.53 3.582 ;
      RECT 30.285 3.292 30.535 3.581 ;
      RECT 30.285 3.35 30.55 3.58 ;
      RECT 30.27 3.223 30.43 3.565 ;
      RECT 30.25 3.232 30.475 3.518 ;
      RECT 30.225 3.243 30.51 3.455 ;
      RECT 30.225 3.327 30.545 3.455 ;
      RECT 30.225 3.302 30.54 3.455 ;
      RECT 30.285 3.218 30.43 3.585 ;
      RECT 30.371 3.217 30.43 3.585 ;
      RECT 30.371 3.216 30.415 3.585 ;
      RECT 30.285 7.855 30.455 8.305 ;
      RECT 30.34 6.075 30.51 8.025 ;
      RECT 30.285 5.015 30.455 6.245 ;
      RECT 29.765 5.015 29.935 8.305 ;
      RECT 29.765 7.315 30.17 7.645 ;
      RECT 29.765 6.475 30.17 6.805 ;
      RECT 30.07 2.732 30.075 3.11 ;
      RECT 30.065 2.7 30.07 3.11 ;
      RECT 30.06 2.672 30.065 3.11 ;
      RECT 30.055 2.652 30.06 3.11 ;
      RECT 30 2.635 30.055 3.11 ;
      RECT 29.96 2.62 30 3.11 ;
      RECT 29.905 2.607 29.96 3.11 ;
      RECT 29.87 2.598 29.905 3.11 ;
      RECT 29.866 2.596 29.87 3.109 ;
      RECT 29.78 2.592 29.866 3.092 ;
      RECT 29.695 2.584 29.78 3.055 ;
      RECT 29.685 2.58 29.695 3.028 ;
      RECT 29.675 2.58 29.685 3.01 ;
      RECT 29.665 2.582 29.675 2.993 ;
      RECT 29.66 2.587 29.665 2.979 ;
      RECT 29.655 2.591 29.66 2.966 ;
      RECT 29.645 2.596 29.655 2.95 ;
      RECT 29.63 2.61 29.645 2.925 ;
      RECT 29.625 2.616 29.63 2.905 ;
      RECT 29.62 2.618 29.625 2.898 ;
      RECT 29.615 2.622 29.62 2.773 ;
      RECT 29.795 3.422 30.04 3.885 ;
      RECT 29.715 3.395 30.035 3.881 ;
      RECT 29.645 3.43 30.04 3.874 ;
      RECT 29.435 3.685 30.04 3.87 ;
      RECT 29.615 3.453 30.04 3.87 ;
      RECT 29.455 3.645 30.04 3.87 ;
      RECT 29.605 3.465 30.04 3.87 ;
      RECT 29.49 3.582 30.04 3.87 ;
      RECT 29.545 3.507 30.04 3.87 ;
      RECT 29.795 3.372 30.035 3.885 ;
      RECT 29.825 3.365 30.035 3.885 ;
      RECT 29.815 3.367 30.035 3.885 ;
      RECT 29.825 3.362 29.955 3.885 ;
      RECT 29.38 1.925 29.466 2.364 ;
      RECT 29.375 1.925 29.466 2.362 ;
      RECT 29.375 1.925 29.535 2.361 ;
      RECT 29.375 1.925 29.565 2.358 ;
      RECT 29.36 1.932 29.565 2.349 ;
      RECT 29.36 1.932 29.57 2.345 ;
      RECT 29.355 1.942 29.57 2.338 ;
      RECT 29.35 1.947 29.57 2.313 ;
      RECT 29.35 1.947 29.585 2.295 ;
      RECT 29.375 1.925 29.605 2.21 ;
      RECT 29.345 1.952 29.605 2.208 ;
      RECT 29.355 1.945 29.61 2.146 ;
      RECT 29.345 2.067 29.615 2.129 ;
      RECT 29.33 1.962 29.61 2.08 ;
      RECT 29.325 1.972 29.61 1.98 ;
      RECT 29.405 2.743 29.41 2.82 ;
      RECT 29.395 2.737 29.405 3.01 ;
      RECT 29.385 2.729 29.395 3.031 ;
      RECT 29.375 2.72 29.385 3.053 ;
      RECT 29.37 2.715 29.375 3.07 ;
      RECT 29.33 2.715 29.37 3.11 ;
      RECT 29.31 2.715 29.33 3.165 ;
      RECT 29.305 2.715 29.31 3.193 ;
      RECT 29.295 2.715 29.305 3.208 ;
      RECT 29.26 2.715 29.295 3.25 ;
      RECT 29.255 2.715 29.26 3.293 ;
      RECT 29.245 2.715 29.255 3.308 ;
      RECT 29.23 2.715 29.245 3.328 ;
      RECT 29.215 2.715 29.23 3.355 ;
      RECT 29.21 2.716 29.215 3.373 ;
      RECT 29.19 2.717 29.21 3.38 ;
      RECT 29.135 2.718 29.19 3.4 ;
      RECT 29.125 2.719 29.135 3.414 ;
      RECT 29.12 2.722 29.125 3.413 ;
      RECT 29.08 2.795 29.12 3.411 ;
      RECT 29.065 2.875 29.08 3.409 ;
      RECT 29.04 2.93 29.065 3.407 ;
      RECT 29.025 2.995 29.04 3.406 ;
      RECT 28.98 3.027 29.025 3.403 ;
      RECT 28.895 3.05 28.98 3.398 ;
      RECT 28.87 3.07 28.895 3.393 ;
      RECT 28.8 3.075 28.87 3.389 ;
      RECT 28.78 3.077 28.8 3.386 ;
      RECT 28.695 3.088 28.78 3.38 ;
      RECT 28.69 3.099 28.695 3.375 ;
      RECT 28.68 3.101 28.69 3.375 ;
      RECT 28.645 3.105 28.68 3.373 ;
      RECT 28.595 3.115 28.645 3.36 ;
      RECT 28.575 3.123 28.595 3.345 ;
      RECT 28.495 3.135 28.575 3.328 ;
      RECT 28.66 2.685 28.83 2.895 ;
      RECT 28.776 2.681 28.83 2.895 ;
      RECT 28.581 2.685 28.83 2.886 ;
      RECT 28.581 2.685 28.835 2.875 ;
      RECT 28.495 2.685 28.835 2.866 ;
      RECT 28.495 2.693 28.845 2.81 ;
      RECT 28.495 2.705 28.85 2.723 ;
      RECT 28.495 2.712 28.855 2.715 ;
      RECT 28.69 2.683 28.83 2.895 ;
      RECT 28.445 3.628 28.69 3.96 ;
      RECT 28.44 3.62 28.445 3.957 ;
      RECT 28.41 3.64 28.69 3.938 ;
      RECT 28.39 3.672 28.69 3.911 ;
      RECT 28.44 3.625 28.617 3.957 ;
      RECT 28.44 3.622 28.531 3.957 ;
      RECT 28.38 1.97 28.55 2.39 ;
      RECT 28.375 1.97 28.55 2.388 ;
      RECT 28.375 1.97 28.575 2.378 ;
      RECT 28.375 1.97 28.595 2.353 ;
      RECT 28.37 1.97 28.595 2.348 ;
      RECT 28.37 1.97 28.605 2.338 ;
      RECT 28.37 1.97 28.61 2.333 ;
      RECT 28.37 1.975 28.615 2.328 ;
      RECT 28.37 2.007 28.63 2.318 ;
      RECT 28.37 2.077 28.655 2.301 ;
      RECT 28.35 2.077 28.655 2.293 ;
      RECT 28.35 2.137 28.665 2.27 ;
      RECT 28.35 2.177 28.675 2.215 ;
      RECT 28.335 1.97 28.61 2.195 ;
      RECT 28.325 1.985 28.615 2.093 ;
      RECT 27.915 3.375 28.085 3.9 ;
      RECT 27.91 3.375 28.085 3.893 ;
      RECT 27.9 3.375 28.09 3.858 ;
      RECT 27.895 3.385 28.09 3.83 ;
      RECT 27.89 3.405 28.09 3.813 ;
      RECT 27.9 3.38 28.095 3.803 ;
      RECT 27.885 3.425 28.095 3.795 ;
      RECT 27.88 3.445 28.095 3.78 ;
      RECT 27.875 3.475 28.095 3.77 ;
      RECT 27.865 3.52 28.095 3.745 ;
      RECT 27.895 3.39 28.1 3.728 ;
      RECT 27.86 3.572 28.1 3.723 ;
      RECT 27.895 3.4 28.105 3.693 ;
      RECT 27.855 3.605 28.105 3.69 ;
      RECT 27.85 3.63 28.105 3.67 ;
      RECT 27.89 3.417 28.115 3.61 ;
      RECT 27.885 3.439 28.125 3.503 ;
      RECT 27.835 2.686 27.85 2.955 ;
      RECT 27.79 2.67 27.835 3 ;
      RECT 27.785 2.658 27.79 3.05 ;
      RECT 27.775 2.654 27.785 3.083 ;
      RECT 27.77 2.651 27.775 3.111 ;
      RECT 27.755 2.653 27.77 3.153 ;
      RECT 27.75 2.657 27.755 3.193 ;
      RECT 27.73 2.662 27.75 3.245 ;
      RECT 27.726 2.667 27.73 3.302 ;
      RECT 27.64 2.686 27.726 3.339 ;
      RECT 27.63 2.707 27.64 3.375 ;
      RECT 27.625 2.715 27.63 3.376 ;
      RECT 27.62 2.757 27.625 3.377 ;
      RECT 27.605 2.845 27.62 3.378 ;
      RECT 27.595 2.995 27.605 3.38 ;
      RECT 27.59 3.04 27.595 3.382 ;
      RECT 27.555 3.082 27.59 3.385 ;
      RECT 27.55 3.1 27.555 3.388 ;
      RECT 27.473 3.106 27.55 3.394 ;
      RECT 27.387 3.12 27.473 3.407 ;
      RECT 27.301 3.134 27.387 3.421 ;
      RECT 27.215 3.148 27.301 3.434 ;
      RECT 27.155 3.16 27.215 3.446 ;
      RECT 27.13 3.167 27.155 3.453 ;
      RECT 27.116 3.17 27.13 3.458 ;
      RECT 27.03 3.178 27.116 3.474 ;
      RECT 27.025 3.185 27.03 3.489 ;
      RECT 27.001 3.185 27.025 3.496 ;
      RECT 26.915 3.188 27.001 3.524 ;
      RECT 26.83 3.192 26.915 3.568 ;
      RECT 26.765 3.196 26.83 3.605 ;
      RECT 26.74 3.199 26.765 3.621 ;
      RECT 26.665 3.212 26.74 3.625 ;
      RECT 26.64 3.23 26.665 3.629 ;
      RECT 26.63 3.237 26.64 3.631 ;
      RECT 26.615 3.24 26.63 3.632 ;
      RECT 26.555 3.252 26.615 3.636 ;
      RECT 26.545 3.266 26.555 3.64 ;
      RECT 26.49 3.276 26.545 3.628 ;
      RECT 26.465 3.297 26.49 3.611 ;
      RECT 26.445 3.317 26.465 3.602 ;
      RECT 26.44 3.33 26.445 3.597 ;
      RECT 26.425 3.342 26.44 3.593 ;
      RECT 27.66 1.997 27.665 2.02 ;
      RECT 27.655 1.988 27.66 2.06 ;
      RECT 27.65 1.986 27.655 2.103 ;
      RECT 27.645 1.977 27.65 2.138 ;
      RECT 27.64 1.967 27.645 2.21 ;
      RECT 27.635 1.957 27.64 2.275 ;
      RECT 27.63 1.954 27.635 2.315 ;
      RECT 27.605 1.948 27.63 2.405 ;
      RECT 27.57 1.936 27.605 2.43 ;
      RECT 27.56 1.927 27.57 2.43 ;
      RECT 27.425 1.925 27.435 2.413 ;
      RECT 27.415 1.925 27.425 2.38 ;
      RECT 27.41 1.925 27.415 2.355 ;
      RECT 27.405 1.925 27.41 2.343 ;
      RECT 27.4 1.925 27.405 2.325 ;
      RECT 27.39 1.925 27.4 2.29 ;
      RECT 27.385 1.927 27.39 2.268 ;
      RECT 27.38 1.933 27.385 2.253 ;
      RECT 27.375 1.939 27.38 2.238 ;
      RECT 27.36 1.951 27.375 2.211 ;
      RECT 27.355 1.962 27.36 2.179 ;
      RECT 27.35 1.972 27.355 2.163 ;
      RECT 27.34 1.98 27.35 2.132 ;
      RECT 27.335 1.99 27.34 2.106 ;
      RECT 27.33 2.047 27.335 2.089 ;
      RECT 27.435 1.925 27.56 2.43 ;
      RECT 27.15 2.612 27.41 2.91 ;
      RECT 27.145 2.619 27.41 2.908 ;
      RECT 27.15 2.614 27.425 2.903 ;
      RECT 27.14 2.627 27.425 2.9 ;
      RECT 27.14 2.632 27.43 2.893 ;
      RECT 27.135 2.64 27.43 2.89 ;
      RECT 27.135 2.657 27.435 2.688 ;
      RECT 27.15 2.609 27.381 2.91 ;
      RECT 27.205 2.608 27.381 2.91 ;
      RECT 27.205 2.605 27.295 2.91 ;
      RECT 27.205 2.602 27.291 2.91 ;
      RECT 26.895 2.875 26.9 2.888 ;
      RECT 26.89 2.842 26.895 2.893 ;
      RECT 26.885 2.797 26.89 2.9 ;
      RECT 26.88 2.752 26.885 2.908 ;
      RECT 26.875 2.72 26.88 2.916 ;
      RECT 26.87 2.68 26.875 2.917 ;
      RECT 26.855 2.66 26.87 2.919 ;
      RECT 26.78 2.642 26.855 2.931 ;
      RECT 26.77 2.635 26.78 2.942 ;
      RECT 26.765 2.635 26.77 2.944 ;
      RECT 26.735 2.641 26.765 2.948 ;
      RECT 26.695 2.654 26.735 2.948 ;
      RECT 26.67 2.665 26.695 2.934 ;
      RECT 26.655 2.671 26.67 2.917 ;
      RECT 26.645 2.673 26.655 2.908 ;
      RECT 26.64 2.674 26.645 2.903 ;
      RECT 26.635 2.675 26.64 2.898 ;
      RECT 26.63 2.676 26.635 2.895 ;
      RECT 26.605 2.681 26.63 2.885 ;
      RECT 26.595 2.697 26.605 2.872 ;
      RECT 26.59 2.717 26.595 2.867 ;
      RECT 26.6 2.11 26.605 2.306 ;
      RECT 26.585 2.074 26.6 2.308 ;
      RECT 26.575 2.056 26.585 2.313 ;
      RECT 26.565 2.042 26.575 2.317 ;
      RECT 26.52 2.026 26.565 2.327 ;
      RECT 26.515 2.016 26.52 2.336 ;
      RECT 26.47 2.005 26.515 2.342 ;
      RECT 26.465 1.993 26.47 2.349 ;
      RECT 26.45 1.988 26.465 2.353 ;
      RECT 26.435 1.98 26.45 2.358 ;
      RECT 26.425 1.973 26.435 2.363 ;
      RECT 26.415 1.97 26.425 2.368 ;
      RECT 26.405 1.97 26.415 2.369 ;
      RECT 26.4 1.967 26.405 2.368 ;
      RECT 26.365 1.962 26.39 2.367 ;
      RECT 26.341 1.958 26.365 2.366 ;
      RECT 26.255 1.949 26.341 2.363 ;
      RECT 26.24 1.941 26.255 2.36 ;
      RECT 26.218 1.94 26.24 2.359 ;
      RECT 26.132 1.94 26.218 2.357 ;
      RECT 26.046 1.94 26.132 2.355 ;
      RECT 25.96 1.94 26.046 2.352 ;
      RECT 25.95 1.94 25.96 2.343 ;
      RECT 25.92 1.94 25.95 2.303 ;
      RECT 25.91 1.95 25.92 2.258 ;
      RECT 25.905 1.99 25.91 2.243 ;
      RECT 25.9 2.005 25.905 2.23 ;
      RECT 25.87 2.085 25.9 2.192 ;
      RECT 26.39 1.965 26.4 2.368 ;
      RECT 26.215 2.73 26.23 3.335 ;
      RECT 26.22 2.725 26.23 3.335 ;
      RECT 26.385 2.725 26.39 2.908 ;
      RECT 26.375 2.725 26.385 2.938 ;
      RECT 26.36 2.725 26.375 2.998 ;
      RECT 26.355 2.725 26.36 3.043 ;
      RECT 26.35 2.725 26.355 3.073 ;
      RECT 26.345 2.725 26.35 3.093 ;
      RECT 26.335 2.725 26.345 3.128 ;
      RECT 26.32 2.725 26.335 3.16 ;
      RECT 26.275 2.725 26.32 3.188 ;
      RECT 26.27 2.725 26.275 3.218 ;
      RECT 26.265 2.725 26.27 3.23 ;
      RECT 26.26 2.725 26.265 3.238 ;
      RECT 26.25 2.725 26.26 3.253 ;
      RECT 26.245 2.725 26.25 3.275 ;
      RECT 26.235 2.725 26.245 3.298 ;
      RECT 26.23 2.725 26.235 3.318 ;
      RECT 26.195 2.74 26.215 3.335 ;
      RECT 26.17 2.757 26.195 3.335 ;
      RECT 26.165 2.767 26.17 3.335 ;
      RECT 26.135 2.782 26.165 3.335 ;
      RECT 26.06 2.824 26.135 3.335 ;
      RECT 26.055 2.855 26.06 3.318 ;
      RECT 26.05 2.859 26.055 3.3 ;
      RECT 26.045 2.863 26.05 3.263 ;
      RECT 26.04 3.047 26.045 3.23 ;
      RECT 25.525 3.236 25.611 3.801 ;
      RECT 25.48 3.238 25.645 3.795 ;
      RECT 25.611 3.235 25.645 3.795 ;
      RECT 25.525 3.237 25.73 3.789 ;
      RECT 25.48 3.247 25.74 3.785 ;
      RECT 25.455 3.239 25.73 3.781 ;
      RECT 25.45 3.242 25.73 3.776 ;
      RECT 25.425 3.257 25.74 3.77 ;
      RECT 25.425 3.282 25.78 3.765 ;
      RECT 25.385 3.29 25.78 3.74 ;
      RECT 25.385 3.317 25.795 3.738 ;
      RECT 25.385 3.347 25.805 3.725 ;
      RECT 25.38 3.492 25.805 3.713 ;
      RECT 25.385 3.421 25.825 3.71 ;
      RECT 25.385 3.478 25.83 3.518 ;
      RECT 25.575 2.757 25.745 2.935 ;
      RECT 25.525 2.696 25.575 2.92 ;
      RECT 25.26 2.676 25.525 2.905 ;
      RECT 25.22 2.74 25.695 2.905 ;
      RECT 25.22 2.73 25.65 2.905 ;
      RECT 25.22 2.727 25.64 2.905 ;
      RECT 25.22 2.715 25.63 2.905 ;
      RECT 25.22 2.7 25.575 2.905 ;
      RECT 25.26 2.672 25.461 2.905 ;
      RECT 25.27 2.65 25.461 2.905 ;
      RECT 25.295 2.635 25.375 2.905 ;
      RECT 25.05 3.165 25.17 3.61 ;
      RECT 25.035 3.165 25.17 3.609 ;
      RECT 24.99 3.187 25.17 3.604 ;
      RECT 24.95 3.236 25.17 3.598 ;
      RECT 24.95 3.236 25.175 3.573 ;
      RECT 24.95 3.236 25.195 3.463 ;
      RECT 24.945 3.266 25.195 3.46 ;
      RECT 25.035 3.165 25.205 3.355 ;
      RECT 24.695 1.95 24.7 2.395 ;
      RECT 24.505 1.95 24.525 2.36 ;
      RECT 24.475 1.95 24.48 2.335 ;
      RECT 25.155 2.257 25.17 2.445 ;
      RECT 25.15 2.242 25.155 2.451 ;
      RECT 25.13 2.215 25.15 2.454 ;
      RECT 25.08 2.182 25.13 2.463 ;
      RECT 25.05 2.162 25.08 2.467 ;
      RECT 25.031 2.15 25.05 2.463 ;
      RECT 24.945 2.122 25.031 2.453 ;
      RECT 24.935 2.097 24.945 2.443 ;
      RECT 24.865 2.065 24.935 2.435 ;
      RECT 24.84 2.025 24.865 2.427 ;
      RECT 24.82 2.007 24.84 2.421 ;
      RECT 24.81 1.997 24.82 2.418 ;
      RECT 24.8 1.99 24.81 2.416 ;
      RECT 24.78 1.977 24.8 2.413 ;
      RECT 24.77 1.967 24.78 2.41 ;
      RECT 24.76 1.96 24.77 2.408 ;
      RECT 24.71 1.952 24.76 2.402 ;
      RECT 24.7 1.95 24.71 2.396 ;
      RECT 24.67 1.95 24.695 2.393 ;
      RECT 24.641 1.95 24.67 2.388 ;
      RECT 24.555 1.95 24.641 2.378 ;
      RECT 24.525 1.95 24.555 2.365 ;
      RECT 24.48 1.95 24.505 2.348 ;
      RECT 24.465 1.95 24.475 2.33 ;
      RECT 24.445 1.957 24.465 2.315 ;
      RECT 24.44 1.972 24.445 2.303 ;
      RECT 24.435 1.977 24.44 2.243 ;
      RECT 24.43 1.982 24.435 2.085 ;
      RECT 24.425 1.985 24.43 2.003 ;
      RECT 24.69 2.67 24.776 2.991 ;
      RECT 24.69 2.67 24.81 2.984 ;
      RECT 24.64 2.67 24.81 2.98 ;
      RECT 24.64 2.672 24.896 2.978 ;
      RECT 24.64 2.674 24.92 2.972 ;
      RECT 24.64 2.681 24.93 2.971 ;
      RECT 24.64 2.69 24.935 2.968 ;
      RECT 24.64 2.696 24.94 2.963 ;
      RECT 24.64 2.74 24.945 2.96 ;
      RECT 24.64 2.832 24.95 2.957 ;
      RECT 24.165 3.275 24.2 3.595 ;
      RECT 24.75 3.46 24.755 3.642 ;
      RECT 24.705 3.342 24.75 3.661 ;
      RECT 24.69 3.319 24.705 3.684 ;
      RECT 24.68 3.309 24.69 3.694 ;
      RECT 24.66 3.304 24.68 3.707 ;
      RECT 24.635 3.302 24.66 3.728 ;
      RECT 24.616 3.301 24.635 3.74 ;
      RECT 24.53 3.298 24.616 3.74 ;
      RECT 24.46 3.293 24.53 3.728 ;
      RECT 24.385 3.289 24.46 3.703 ;
      RECT 24.32 3.285 24.385 3.67 ;
      RECT 24.25 3.282 24.32 3.63 ;
      RECT 24.22 3.278 24.25 3.605 ;
      RECT 24.2 3.276 24.22 3.598 ;
      RECT 24.116 3.274 24.165 3.596 ;
      RECT 24.03 3.271 24.116 3.597 ;
      RECT 23.955 3.27 24.03 3.599 ;
      RECT 23.87 3.27 23.955 3.625 ;
      RECT 23.793 3.271 23.87 3.65 ;
      RECT 23.707 3.272 23.793 3.65 ;
      RECT 23.621 3.272 23.707 3.65 ;
      RECT 23.535 3.273 23.621 3.65 ;
      RECT 23.515 3.274 23.535 3.642 ;
      RECT 23.5 3.28 23.515 3.627 ;
      RECT 23.465 3.3 23.5 3.607 ;
      RECT 23.455 3.32 23.465 3.589 ;
      RECT 24.425 2.625 24.43 2.895 ;
      RECT 24.42 2.616 24.425 2.9 ;
      RECT 24.41 2.606 24.42 2.912 ;
      RECT 24.405 2.595 24.41 2.923 ;
      RECT 24.385 2.589 24.405 2.941 ;
      RECT 24.34 2.586 24.385 2.99 ;
      RECT 24.325 2.585 24.34 3.035 ;
      RECT 24.32 2.585 24.325 3.048 ;
      RECT 24.31 2.585 24.32 3.06 ;
      RECT 24.305 2.586 24.31 3.075 ;
      RECT 24.285 2.594 24.305 3.08 ;
      RECT 24.255 2.61 24.285 3.08 ;
      RECT 24.245 2.622 24.25 3.08 ;
      RECT 24.21 2.637 24.245 3.08 ;
      RECT 24.18 2.657 24.21 3.08 ;
      RECT 24.17 2.682 24.18 3.08 ;
      RECT 24.165 2.71 24.17 3.08 ;
      RECT 24.16 2.74 24.165 3.08 ;
      RECT 24.155 2.757 24.16 3.08 ;
      RECT 24.145 2.785 24.155 3.08 ;
      RECT 24.135 2.82 24.145 3.08 ;
      RECT 24.13 2.855 24.135 3.08 ;
      RECT 24.25 2.62 24.255 3.08 ;
      RECT 23.765 2.722 23.95 2.895 ;
      RECT 23.725 2.64 23.91 2.893 ;
      RECT 23.686 2.645 23.91 2.889 ;
      RECT 23.6 2.654 23.91 2.884 ;
      RECT 23.516 2.67 23.915 2.879 ;
      RECT 23.43 2.69 23.94 2.873 ;
      RECT 23.43 2.71 23.945 2.873 ;
      RECT 23.516 2.68 23.94 2.879 ;
      RECT 23.6 2.655 23.915 2.884 ;
      RECT 23.765 2.637 23.91 2.895 ;
      RECT 23.765 2.632 23.865 2.895 ;
      RECT 23.851 2.626 23.865 2.895 ;
      RECT 23.24 1.95 23.245 2.349 ;
      RECT 22.985 1.95 23.02 2.347 ;
      RECT 22.58 1.985 22.585 2.341 ;
      RECT 23.325 1.988 23.33 2.243 ;
      RECT 23.32 1.986 23.325 2.249 ;
      RECT 23.315 1.985 23.32 2.256 ;
      RECT 23.29 1.978 23.315 2.28 ;
      RECT 23.285 1.971 23.29 2.304 ;
      RECT 23.28 1.967 23.285 2.313 ;
      RECT 23.27 1.962 23.28 2.326 ;
      RECT 23.265 1.959 23.27 2.335 ;
      RECT 23.26 1.957 23.265 2.34 ;
      RECT 23.245 1.953 23.26 2.35 ;
      RECT 23.23 1.947 23.24 2.349 ;
      RECT 23.192 1.945 23.23 2.349 ;
      RECT 23.106 1.947 23.192 2.349 ;
      RECT 23.02 1.949 23.106 2.348 ;
      RECT 22.949 1.95 22.985 2.347 ;
      RECT 22.863 1.952 22.949 2.347 ;
      RECT 22.777 1.954 22.863 2.346 ;
      RECT 22.691 1.956 22.777 2.346 ;
      RECT 22.605 1.959 22.691 2.345 ;
      RECT 22.595 1.965 22.605 2.344 ;
      RECT 22.585 1.977 22.595 2.342 ;
      RECT 22.525 2.012 22.58 2.338 ;
      RECT 22.52 2.042 22.525 2.1 ;
      RECT 23.265 3.122 23.28 3.315 ;
      RECT 23.26 3.09 23.265 3.315 ;
      RECT 23.25 3.065 23.26 3.315 ;
      RECT 23.245 3.037 23.25 3.315 ;
      RECT 23.215 2.96 23.245 3.315 ;
      RECT 23.19 2.842 23.215 3.315 ;
      RECT 23.185 2.78 23.19 3.315 ;
      RECT 23.175 2.767 23.185 3.315 ;
      RECT 23.155 2.757 23.175 3.315 ;
      RECT 23.14 2.74 23.155 3.315 ;
      RECT 23.11 2.728 23.14 3.315 ;
      RECT 23.105 2.727 23.11 3.26 ;
      RECT 23.1 2.727 23.105 3.218 ;
      RECT 23.085 2.726 23.1 3.17 ;
      RECT 23.07 2.726 23.085 3.108 ;
      RECT 23.05 2.726 23.07 3.068 ;
      RECT 23.045 2.726 23.05 3.053 ;
      RECT 23.02 2.725 23.045 3.048 ;
      RECT 22.95 2.724 23.02 3.035 ;
      RECT 22.935 2.723 22.95 3.02 ;
      RECT 22.905 2.722 22.935 3.003 ;
      RECT 22.9 2.722 22.905 2.988 ;
      RECT 22.85 2.721 22.9 2.968 ;
      RECT 22.785 2.72 22.85 2.923 ;
      RECT 22.78 2.72 22.785 2.895 ;
      RECT 22.865 3.257 22.87 3.514 ;
      RECT 22.845 3.176 22.865 3.531 ;
      RECT 22.825 3.17 22.845 3.56 ;
      RECT 22.765 3.157 22.825 3.58 ;
      RECT 22.72 3.141 22.765 3.581 ;
      RECT 22.636 3.129 22.72 3.569 ;
      RECT 22.55 3.116 22.636 3.553 ;
      RECT 22.54 3.109 22.55 3.545 ;
      RECT 22.495 3.106 22.54 3.485 ;
      RECT 22.475 3.102 22.495 3.4 ;
      RECT 22.46 3.1 22.475 3.353 ;
      RECT 22.43 3.097 22.46 3.323 ;
      RECT 22.395 3.093 22.43 3.3 ;
      RECT 22.352 3.088 22.395 3.288 ;
      RECT 22.266 3.079 22.352 3.297 ;
      RECT 22.18 3.068 22.266 3.309 ;
      RECT 22.115 3.059 22.18 3.318 ;
      RECT 22.095 3.05 22.115 3.323 ;
      RECT 22.09 3.043 22.095 3.325 ;
      RECT 22.05 3.028 22.09 3.322 ;
      RECT 22.03 3.007 22.05 3.317 ;
      RECT 22.015 2.995 22.03 3.31 ;
      RECT 22.01 2.987 22.015 3.303 ;
      RECT 21.995 2.967 22.01 3.296 ;
      RECT 21.99 2.83 21.995 3.29 ;
      RECT 21.91 2.719 21.99 3.262 ;
      RECT 21.901 2.712 21.91 3.228 ;
      RECT 21.815 2.706 21.901 3.153 ;
      RECT 21.79 2.697 21.815 3.065 ;
      RECT 21.76 2.692 21.79 3.04 ;
      RECT 21.695 2.701 21.76 3.025 ;
      RECT 21.675 2.717 21.695 3 ;
      RECT 21.665 2.723 21.675 2.948 ;
      RECT 21.645 2.745 21.665 2.83 ;
      RECT 22.3 2.71 22.47 2.895 ;
      RECT 22.3 2.71 22.505 2.893 ;
      RECT 22.35 2.62 22.52 2.884 ;
      RECT 22.3 2.777 22.525 2.877 ;
      RECT 22.315 2.655 22.52 2.884 ;
      RECT 21.515 3.388 21.58 3.831 ;
      RECT 21.455 3.413 21.58 3.829 ;
      RECT 21.455 3.413 21.635 3.823 ;
      RECT 21.44 3.438 21.635 3.822 ;
      RECT 21.58 3.375 21.655 3.819 ;
      RECT 21.515 3.4 21.735 3.813 ;
      RECT 21.44 3.439 21.78 3.807 ;
      RECT 21.425 3.466 21.78 3.798 ;
      RECT 21.44 3.459 21.8 3.79 ;
      RECT 21.425 3.468 21.805 3.773 ;
      RECT 21.42 3.485 21.805 3.6 ;
      RECT 21.425 2.207 21.46 2.445 ;
      RECT 21.425 2.207 21.49 2.444 ;
      RECT 21.425 2.207 21.605 2.44 ;
      RECT 21.425 2.207 21.66 2.418 ;
      RECT 21.435 2.15 21.715 2.318 ;
      RECT 21.54 1.99 21.57 2.441 ;
      RECT 21.57 1.985 21.75 2.198 ;
      RECT 21.44 2.126 21.75 2.198 ;
      RECT 21.49 2.022 21.54 2.442 ;
      RECT 21.46 2.078 21.75 2.198 ;
      RECT 19.965 1.74 20.135 2.935 ;
      RECT 19.965 1.74 20.43 1.91 ;
      RECT 19.965 6.97 20.43 7.14 ;
      RECT 19.965 5.945 20.135 7.14 ;
      RECT 18.975 1.74 19.145 2.935 ;
      RECT 18.975 1.74 19.44 1.91 ;
      RECT 18.975 6.97 19.44 7.14 ;
      RECT 18.975 5.945 19.145 7.14 ;
      RECT 17.12 2.635 17.29 3.865 ;
      RECT 17.175 0.855 17.345 2.805 ;
      RECT 17.12 0.575 17.29 1.025 ;
      RECT 17.12 7.855 17.29 8.305 ;
      RECT 17.175 6.075 17.345 8.025 ;
      RECT 17.12 5.015 17.29 6.245 ;
      RECT 16.6 0.575 16.77 3.865 ;
      RECT 16.6 2.075 17.005 2.405 ;
      RECT 16.6 1.235 17.005 1.565 ;
      RECT 16.6 5.015 16.77 8.305 ;
      RECT 16.6 7.315 17.005 7.645 ;
      RECT 16.6 6.475 17.005 6.805 ;
      RECT 14.7 3.392 14.715 3.443 ;
      RECT 14.695 3.372 14.7 3.49 ;
      RECT 14.68 3.362 14.695 3.558 ;
      RECT 14.655 3.342 14.68 3.613 ;
      RECT 14.615 3.327 14.655 3.633 ;
      RECT 14.57 3.321 14.615 3.661 ;
      RECT 14.5 3.311 14.57 3.678 ;
      RECT 14.48 3.303 14.5 3.678 ;
      RECT 14.42 3.297 14.48 3.67 ;
      RECT 14.361 3.288 14.42 3.658 ;
      RECT 14.275 3.277 14.361 3.641 ;
      RECT 14.253 3.268 14.275 3.629 ;
      RECT 14.167 3.261 14.253 3.616 ;
      RECT 14.081 3.248 14.167 3.597 ;
      RECT 13.995 3.236 14.081 3.577 ;
      RECT 13.965 3.225 13.995 3.564 ;
      RECT 13.915 3.211 13.965 3.556 ;
      RECT 13.895 3.2 13.915 3.548 ;
      RECT 13.846 3.189 13.895 3.54 ;
      RECT 13.76 3.168 13.846 3.525 ;
      RECT 13.715 3.155 13.76 3.51 ;
      RECT 13.67 3.155 13.715 3.49 ;
      RECT 13.615 3.155 13.67 3.425 ;
      RECT 13.59 3.155 13.615 3.348 ;
      RECT 14.115 2.892 14.285 3.075 ;
      RECT 14.115 2.892 14.3 3.033 ;
      RECT 14.115 2.892 14.305 2.975 ;
      RECT 14.175 2.66 14.31 2.951 ;
      RECT 14.175 2.664 14.315 2.934 ;
      RECT 14.12 2.827 14.315 2.934 ;
      RECT 14.145 2.672 14.285 3.075 ;
      RECT 14.145 2.676 14.325 2.875 ;
      RECT 14.13 2.762 14.325 2.875 ;
      RECT 14.14 2.692 14.285 3.075 ;
      RECT 14.14 2.695 14.335 2.788 ;
      RECT 14.135 2.712 14.335 2.788 ;
      RECT 13.905 1.932 14.075 2.415 ;
      RECT 13.9 1.927 14.05 2.405 ;
      RECT 13.9 1.934 14.08 2.399 ;
      RECT 13.89 1.928 14.05 2.378 ;
      RECT 13.89 1.944 14.095 2.337 ;
      RECT 13.86 1.929 14.05 2.3 ;
      RECT 13.86 1.959 14.105 2.24 ;
      RECT 13.855 1.931 14.05 2.238 ;
      RECT 13.835 1.94 14.08 2.195 ;
      RECT 13.81 1.956 14.095 2.107 ;
      RECT 13.81 1.975 14.12 2.098 ;
      RECT 13.805 2.012 14.12 2.05 ;
      RECT 13.81 1.992 14.125 2.018 ;
      RECT 13.905 1.926 14.015 2.415 ;
      RECT 13.991 1.925 14.015 2.415 ;
      RECT 13.225 2.71 13.23 2.921 ;
      RECT 13.825 2.71 13.83 2.895 ;
      RECT 13.89 2.75 13.895 2.863 ;
      RECT 13.885 2.742 13.89 2.869 ;
      RECT 13.88 2.732 13.885 2.877 ;
      RECT 13.875 2.722 13.88 2.886 ;
      RECT 13.87 2.712 13.875 2.89 ;
      RECT 13.83 2.71 13.87 2.893 ;
      RECT 13.802 2.709 13.825 2.897 ;
      RECT 13.716 2.706 13.802 2.904 ;
      RECT 13.63 2.702 13.716 2.915 ;
      RECT 13.61 2.7 13.63 2.921 ;
      RECT 13.592 2.699 13.61 2.924 ;
      RECT 13.506 2.697 13.592 2.931 ;
      RECT 13.42 2.692 13.506 2.944 ;
      RECT 13.401 2.689 13.42 2.949 ;
      RECT 13.315 2.687 13.401 2.94 ;
      RECT 13.305 2.687 13.315 2.933 ;
      RECT 13.23 2.7 13.305 2.927 ;
      RECT 13.215 2.711 13.225 2.921 ;
      RECT 13.205 2.713 13.215 2.92 ;
      RECT 13.195 2.717 13.205 2.916 ;
      RECT 13.19 2.72 13.195 2.91 ;
      RECT 13.18 2.722 13.19 2.904 ;
      RECT 13.175 2.725 13.18 2.898 ;
      RECT 13.155 3.311 13.16 3.515 ;
      RECT 13.14 3.298 13.155 3.608 ;
      RECT 13.125 3.279 13.14 3.885 ;
      RECT 13.09 3.245 13.125 3.885 ;
      RECT 13.086 3.215 13.09 3.885 ;
      RECT 13 3.097 13.086 3.885 ;
      RECT 12.99 2.972 13 3.885 ;
      RECT 12.975 2.94 12.99 3.885 ;
      RECT 12.97 2.915 12.975 3.885 ;
      RECT 12.965 2.905 12.97 3.841 ;
      RECT 12.95 2.877 12.965 3.746 ;
      RECT 12.935 2.843 12.95 3.645 ;
      RECT 12.93 2.821 12.935 3.598 ;
      RECT 12.925 2.81 12.93 3.568 ;
      RECT 12.92 2.8 12.925 3.534 ;
      RECT 12.91 2.787 12.92 3.502 ;
      RECT 12.885 2.763 12.91 3.428 ;
      RECT 12.88 2.743 12.885 3.353 ;
      RECT 12.875 2.737 12.88 3.328 ;
      RECT 12.87 2.732 12.875 3.293 ;
      RECT 12.865 2.727 12.87 3.268 ;
      RECT 12.86 2.725 12.865 3.248 ;
      RECT 12.855 2.725 12.86 3.233 ;
      RECT 12.85 2.725 12.855 3.193 ;
      RECT 12.84 2.725 12.85 3.165 ;
      RECT 12.83 2.725 12.84 3.11 ;
      RECT 12.815 2.725 12.83 3.048 ;
      RECT 12.81 2.724 12.815 2.993 ;
      RECT 12.795 2.723 12.81 2.973 ;
      RECT 12.735 2.721 12.795 2.947 ;
      RECT 12.7 2.722 12.735 2.927 ;
      RECT 12.695 2.724 12.7 2.917 ;
      RECT 12.685 2.743 12.695 2.907 ;
      RECT 12.68 2.77 12.685 2.838 ;
      RECT 12.795 2.195 12.965 2.44 ;
      RECT 12.83 1.966 12.965 2.44 ;
      RECT 12.83 1.968 12.975 2.435 ;
      RECT 12.83 1.97 13 2.423 ;
      RECT 12.83 1.973 13.025 2.405 ;
      RECT 12.83 1.978 13.075 2.378 ;
      RECT 12.83 1.983 13.095 2.343 ;
      RECT 12.81 1.985 13.105 2.318 ;
      RECT 12.8 2.08 13.105 2.318 ;
      RECT 12.83 1.965 12.94 2.44 ;
      RECT 12.84 1.962 12.935 2.44 ;
      RECT 12.36 3.227 12.55 3.585 ;
      RECT 12.36 3.239 12.585 3.584 ;
      RECT 12.36 3.267 12.605 3.582 ;
      RECT 12.36 3.292 12.61 3.581 ;
      RECT 12.36 3.35 12.625 3.58 ;
      RECT 12.345 3.223 12.505 3.565 ;
      RECT 12.325 3.232 12.55 3.518 ;
      RECT 12.3 3.243 12.585 3.455 ;
      RECT 12.3 3.327 12.62 3.455 ;
      RECT 12.3 3.302 12.615 3.455 ;
      RECT 12.36 3.218 12.505 3.585 ;
      RECT 12.446 3.217 12.505 3.585 ;
      RECT 12.446 3.216 12.49 3.585 ;
      RECT 12.36 7.855 12.53 8.305 ;
      RECT 12.415 6.075 12.585 8.025 ;
      RECT 12.36 5.015 12.53 6.245 ;
      RECT 11.84 5.015 12.01 8.305 ;
      RECT 11.84 7.315 12.245 7.645 ;
      RECT 11.84 6.475 12.245 6.805 ;
      RECT 12.145 2.732 12.15 3.11 ;
      RECT 12.14 2.7 12.145 3.11 ;
      RECT 12.135 2.672 12.14 3.11 ;
      RECT 12.13 2.652 12.135 3.11 ;
      RECT 12.075 2.635 12.13 3.11 ;
      RECT 12.035 2.62 12.075 3.11 ;
      RECT 11.98 2.607 12.035 3.11 ;
      RECT 11.945 2.598 11.98 3.11 ;
      RECT 11.941 2.596 11.945 3.109 ;
      RECT 11.855 2.592 11.941 3.092 ;
      RECT 11.77 2.584 11.855 3.055 ;
      RECT 11.76 2.58 11.77 3.028 ;
      RECT 11.75 2.58 11.76 3.01 ;
      RECT 11.74 2.582 11.75 2.993 ;
      RECT 11.735 2.587 11.74 2.979 ;
      RECT 11.73 2.591 11.735 2.966 ;
      RECT 11.72 2.596 11.73 2.95 ;
      RECT 11.705 2.61 11.72 2.925 ;
      RECT 11.7 2.616 11.705 2.905 ;
      RECT 11.695 2.618 11.7 2.898 ;
      RECT 11.69 2.622 11.695 2.773 ;
      RECT 11.87 3.422 12.115 3.885 ;
      RECT 11.79 3.395 12.11 3.881 ;
      RECT 11.72 3.43 12.115 3.874 ;
      RECT 11.51 3.685 12.115 3.87 ;
      RECT 11.69 3.453 12.115 3.87 ;
      RECT 11.53 3.645 12.115 3.87 ;
      RECT 11.68 3.465 12.115 3.87 ;
      RECT 11.565 3.582 12.115 3.87 ;
      RECT 11.62 3.507 12.115 3.87 ;
      RECT 11.87 3.372 12.11 3.885 ;
      RECT 11.9 3.365 12.11 3.885 ;
      RECT 11.89 3.367 12.11 3.885 ;
      RECT 11.9 3.362 12.03 3.885 ;
      RECT 11.455 1.925 11.541 2.364 ;
      RECT 11.45 1.925 11.541 2.362 ;
      RECT 11.45 1.925 11.61 2.361 ;
      RECT 11.45 1.925 11.64 2.358 ;
      RECT 11.435 1.932 11.64 2.349 ;
      RECT 11.435 1.932 11.645 2.345 ;
      RECT 11.43 1.942 11.645 2.338 ;
      RECT 11.425 1.947 11.645 2.313 ;
      RECT 11.425 1.947 11.66 2.295 ;
      RECT 11.45 1.925 11.68 2.21 ;
      RECT 11.42 1.952 11.68 2.208 ;
      RECT 11.43 1.945 11.685 2.146 ;
      RECT 11.42 2.067 11.69 2.129 ;
      RECT 11.405 1.962 11.685 2.08 ;
      RECT 11.4 1.972 11.685 1.98 ;
      RECT 11.48 2.743 11.485 2.82 ;
      RECT 11.47 2.737 11.48 3.01 ;
      RECT 11.46 2.729 11.47 3.031 ;
      RECT 11.45 2.72 11.46 3.053 ;
      RECT 11.445 2.715 11.45 3.07 ;
      RECT 11.405 2.715 11.445 3.11 ;
      RECT 11.385 2.715 11.405 3.165 ;
      RECT 11.38 2.715 11.385 3.193 ;
      RECT 11.37 2.715 11.38 3.208 ;
      RECT 11.335 2.715 11.37 3.25 ;
      RECT 11.33 2.715 11.335 3.293 ;
      RECT 11.32 2.715 11.33 3.308 ;
      RECT 11.305 2.715 11.32 3.328 ;
      RECT 11.29 2.715 11.305 3.355 ;
      RECT 11.285 2.716 11.29 3.373 ;
      RECT 11.265 2.717 11.285 3.38 ;
      RECT 11.21 2.718 11.265 3.4 ;
      RECT 11.2 2.719 11.21 3.414 ;
      RECT 11.195 2.722 11.2 3.413 ;
      RECT 11.155 2.795 11.195 3.411 ;
      RECT 11.14 2.875 11.155 3.409 ;
      RECT 11.115 2.93 11.14 3.407 ;
      RECT 11.1 2.995 11.115 3.406 ;
      RECT 11.055 3.027 11.1 3.403 ;
      RECT 10.97 3.05 11.055 3.398 ;
      RECT 10.945 3.07 10.97 3.393 ;
      RECT 10.875 3.075 10.945 3.389 ;
      RECT 10.855 3.077 10.875 3.386 ;
      RECT 10.77 3.088 10.855 3.38 ;
      RECT 10.765 3.099 10.77 3.375 ;
      RECT 10.755 3.101 10.765 3.375 ;
      RECT 10.72 3.105 10.755 3.373 ;
      RECT 10.67 3.115 10.72 3.36 ;
      RECT 10.65 3.123 10.67 3.345 ;
      RECT 10.57 3.135 10.65 3.328 ;
      RECT 10.735 2.685 10.905 2.895 ;
      RECT 10.851 2.681 10.905 2.895 ;
      RECT 10.656 2.685 10.905 2.886 ;
      RECT 10.656 2.685 10.91 2.875 ;
      RECT 10.57 2.685 10.91 2.866 ;
      RECT 10.57 2.693 10.92 2.81 ;
      RECT 10.57 2.705 10.925 2.723 ;
      RECT 10.57 2.712 10.93 2.715 ;
      RECT 10.765 2.683 10.905 2.895 ;
      RECT 10.52 3.628 10.765 3.96 ;
      RECT 10.515 3.62 10.52 3.957 ;
      RECT 10.485 3.64 10.765 3.938 ;
      RECT 10.465 3.672 10.765 3.911 ;
      RECT 10.515 3.625 10.692 3.957 ;
      RECT 10.515 3.622 10.606 3.957 ;
      RECT 10.455 1.97 10.625 2.39 ;
      RECT 10.45 1.97 10.625 2.388 ;
      RECT 10.45 1.97 10.65 2.378 ;
      RECT 10.45 1.97 10.67 2.353 ;
      RECT 10.445 1.97 10.67 2.348 ;
      RECT 10.445 1.97 10.68 2.338 ;
      RECT 10.445 1.97 10.685 2.333 ;
      RECT 10.445 1.975 10.69 2.328 ;
      RECT 10.445 2.007 10.705 2.318 ;
      RECT 10.445 2.077 10.73 2.301 ;
      RECT 10.425 2.077 10.73 2.293 ;
      RECT 10.425 2.137 10.74 2.27 ;
      RECT 10.425 2.177 10.75 2.215 ;
      RECT 10.41 1.97 10.685 2.195 ;
      RECT 10.4 1.985 10.69 2.093 ;
      RECT 9.99 3.375 10.16 3.9 ;
      RECT 9.985 3.375 10.16 3.893 ;
      RECT 9.975 3.375 10.165 3.858 ;
      RECT 9.97 3.385 10.165 3.83 ;
      RECT 9.965 3.405 10.165 3.813 ;
      RECT 9.975 3.38 10.17 3.803 ;
      RECT 9.96 3.425 10.17 3.795 ;
      RECT 9.955 3.445 10.17 3.78 ;
      RECT 9.95 3.475 10.17 3.77 ;
      RECT 9.94 3.52 10.17 3.745 ;
      RECT 9.97 3.39 10.175 3.728 ;
      RECT 9.935 3.572 10.175 3.723 ;
      RECT 9.97 3.4 10.18 3.693 ;
      RECT 9.93 3.605 10.18 3.69 ;
      RECT 9.925 3.63 10.18 3.67 ;
      RECT 9.965 3.417 10.19 3.61 ;
      RECT 9.96 3.439 10.2 3.503 ;
      RECT 9.91 2.686 9.925 2.955 ;
      RECT 9.865 2.67 9.91 3 ;
      RECT 9.86 2.658 9.865 3.05 ;
      RECT 9.85 2.654 9.86 3.083 ;
      RECT 9.845 2.651 9.85 3.111 ;
      RECT 9.83 2.653 9.845 3.153 ;
      RECT 9.825 2.657 9.83 3.193 ;
      RECT 9.805 2.662 9.825 3.245 ;
      RECT 9.801 2.667 9.805 3.302 ;
      RECT 9.715 2.686 9.801 3.339 ;
      RECT 9.705 2.707 9.715 3.375 ;
      RECT 9.7 2.715 9.705 3.376 ;
      RECT 9.695 2.757 9.7 3.377 ;
      RECT 9.68 2.845 9.695 3.378 ;
      RECT 9.67 2.995 9.68 3.38 ;
      RECT 9.665 3.04 9.67 3.382 ;
      RECT 9.63 3.082 9.665 3.385 ;
      RECT 9.625 3.1 9.63 3.388 ;
      RECT 9.548 3.106 9.625 3.394 ;
      RECT 9.462 3.12 9.548 3.407 ;
      RECT 9.376 3.134 9.462 3.421 ;
      RECT 9.29 3.148 9.376 3.434 ;
      RECT 9.23 3.16 9.29 3.446 ;
      RECT 9.205 3.167 9.23 3.453 ;
      RECT 9.191 3.17 9.205 3.458 ;
      RECT 9.105 3.178 9.191 3.474 ;
      RECT 9.1 3.185 9.105 3.489 ;
      RECT 9.076 3.185 9.1 3.496 ;
      RECT 8.99 3.188 9.076 3.524 ;
      RECT 8.905 3.192 8.99 3.568 ;
      RECT 8.84 3.196 8.905 3.605 ;
      RECT 8.815 3.199 8.84 3.621 ;
      RECT 8.74 3.212 8.815 3.625 ;
      RECT 8.715 3.23 8.74 3.629 ;
      RECT 8.705 3.237 8.715 3.631 ;
      RECT 8.69 3.24 8.705 3.632 ;
      RECT 8.63 3.252 8.69 3.636 ;
      RECT 8.62 3.266 8.63 3.64 ;
      RECT 8.565 3.276 8.62 3.628 ;
      RECT 8.54 3.297 8.565 3.611 ;
      RECT 8.52 3.317 8.54 3.602 ;
      RECT 8.515 3.33 8.52 3.597 ;
      RECT 8.5 3.342 8.515 3.593 ;
      RECT 9.735 1.997 9.74 2.02 ;
      RECT 9.73 1.988 9.735 2.06 ;
      RECT 9.725 1.986 9.73 2.103 ;
      RECT 9.72 1.977 9.725 2.138 ;
      RECT 9.715 1.967 9.72 2.21 ;
      RECT 9.71 1.957 9.715 2.275 ;
      RECT 9.705 1.954 9.71 2.315 ;
      RECT 9.68 1.948 9.705 2.405 ;
      RECT 9.645 1.936 9.68 2.43 ;
      RECT 9.635 1.927 9.645 2.43 ;
      RECT 9.5 1.925 9.51 2.413 ;
      RECT 9.49 1.925 9.5 2.38 ;
      RECT 9.485 1.925 9.49 2.355 ;
      RECT 9.48 1.925 9.485 2.343 ;
      RECT 9.475 1.925 9.48 2.325 ;
      RECT 9.465 1.925 9.475 2.29 ;
      RECT 9.46 1.927 9.465 2.268 ;
      RECT 9.455 1.933 9.46 2.253 ;
      RECT 9.45 1.939 9.455 2.238 ;
      RECT 9.435 1.951 9.45 2.211 ;
      RECT 9.43 1.962 9.435 2.179 ;
      RECT 9.425 1.972 9.43 2.163 ;
      RECT 9.415 1.98 9.425 2.132 ;
      RECT 9.41 1.99 9.415 2.106 ;
      RECT 9.405 2.047 9.41 2.089 ;
      RECT 9.51 1.925 9.635 2.43 ;
      RECT 9.225 2.612 9.485 2.91 ;
      RECT 9.22 2.619 9.485 2.908 ;
      RECT 9.225 2.614 9.5 2.903 ;
      RECT 9.215 2.627 9.5 2.9 ;
      RECT 9.215 2.632 9.505 2.893 ;
      RECT 9.21 2.64 9.505 2.89 ;
      RECT 9.21 2.657 9.51 2.688 ;
      RECT 9.225 2.609 9.456 2.91 ;
      RECT 9.28 2.608 9.456 2.91 ;
      RECT 9.28 2.605 9.37 2.91 ;
      RECT 9.28 2.602 9.366 2.91 ;
      RECT 8.97 2.875 8.975 2.888 ;
      RECT 8.965 2.842 8.97 2.893 ;
      RECT 8.96 2.797 8.965 2.9 ;
      RECT 8.955 2.752 8.96 2.908 ;
      RECT 8.95 2.72 8.955 2.916 ;
      RECT 8.945 2.68 8.95 2.917 ;
      RECT 8.93 2.66 8.945 2.919 ;
      RECT 8.855 2.642 8.93 2.931 ;
      RECT 8.845 2.635 8.855 2.942 ;
      RECT 8.84 2.635 8.845 2.944 ;
      RECT 8.81 2.641 8.84 2.948 ;
      RECT 8.77 2.654 8.81 2.948 ;
      RECT 8.745 2.665 8.77 2.934 ;
      RECT 8.73 2.671 8.745 2.917 ;
      RECT 8.72 2.673 8.73 2.908 ;
      RECT 8.715 2.674 8.72 2.903 ;
      RECT 8.71 2.675 8.715 2.898 ;
      RECT 8.705 2.676 8.71 2.895 ;
      RECT 8.68 2.681 8.705 2.885 ;
      RECT 8.67 2.697 8.68 2.872 ;
      RECT 8.665 2.717 8.67 2.867 ;
      RECT 8.675 2.11 8.68 2.306 ;
      RECT 8.66 2.074 8.675 2.308 ;
      RECT 8.65 2.056 8.66 2.313 ;
      RECT 8.64 2.042 8.65 2.317 ;
      RECT 8.595 2.026 8.64 2.327 ;
      RECT 8.59 2.016 8.595 2.336 ;
      RECT 8.545 2.005 8.59 2.342 ;
      RECT 8.54 1.993 8.545 2.349 ;
      RECT 8.525 1.988 8.54 2.353 ;
      RECT 8.51 1.98 8.525 2.358 ;
      RECT 8.5 1.973 8.51 2.363 ;
      RECT 8.49 1.97 8.5 2.368 ;
      RECT 8.48 1.97 8.49 2.369 ;
      RECT 8.475 1.967 8.48 2.368 ;
      RECT 8.44 1.962 8.465 2.367 ;
      RECT 8.416 1.958 8.44 2.366 ;
      RECT 8.33 1.949 8.416 2.363 ;
      RECT 8.315 1.941 8.33 2.36 ;
      RECT 8.293 1.94 8.315 2.359 ;
      RECT 8.207 1.94 8.293 2.357 ;
      RECT 8.121 1.94 8.207 2.355 ;
      RECT 8.035 1.94 8.121 2.352 ;
      RECT 8.025 1.94 8.035 2.343 ;
      RECT 7.995 1.94 8.025 2.303 ;
      RECT 7.985 1.95 7.995 2.258 ;
      RECT 7.98 1.99 7.985 2.243 ;
      RECT 7.975 2.005 7.98 2.23 ;
      RECT 7.945 2.085 7.975 2.192 ;
      RECT 8.465 1.965 8.475 2.368 ;
      RECT 8.29 2.73 8.305 3.335 ;
      RECT 8.295 2.725 8.305 3.335 ;
      RECT 8.46 2.725 8.465 2.908 ;
      RECT 8.45 2.725 8.46 2.938 ;
      RECT 8.435 2.725 8.45 2.998 ;
      RECT 8.43 2.725 8.435 3.043 ;
      RECT 8.425 2.725 8.43 3.073 ;
      RECT 8.42 2.725 8.425 3.093 ;
      RECT 8.41 2.725 8.42 3.128 ;
      RECT 8.395 2.725 8.41 3.16 ;
      RECT 8.35 2.725 8.395 3.188 ;
      RECT 8.345 2.725 8.35 3.218 ;
      RECT 8.34 2.725 8.345 3.23 ;
      RECT 8.335 2.725 8.34 3.238 ;
      RECT 8.325 2.725 8.335 3.253 ;
      RECT 8.32 2.725 8.325 3.275 ;
      RECT 8.31 2.725 8.32 3.298 ;
      RECT 8.305 2.725 8.31 3.318 ;
      RECT 8.27 2.74 8.29 3.335 ;
      RECT 8.245 2.757 8.27 3.335 ;
      RECT 8.24 2.767 8.245 3.335 ;
      RECT 8.21 2.782 8.24 3.335 ;
      RECT 8.135 2.824 8.21 3.335 ;
      RECT 8.13 2.855 8.135 3.318 ;
      RECT 8.125 2.859 8.13 3.3 ;
      RECT 8.12 2.863 8.125 3.263 ;
      RECT 8.115 3.047 8.12 3.23 ;
      RECT 7.6 3.236 7.686 3.801 ;
      RECT 7.555 3.238 7.72 3.795 ;
      RECT 7.686 3.235 7.72 3.795 ;
      RECT 7.6 3.237 7.805 3.789 ;
      RECT 7.555 3.247 7.815 3.785 ;
      RECT 7.53 3.239 7.805 3.781 ;
      RECT 7.525 3.242 7.805 3.776 ;
      RECT 7.5 3.257 7.815 3.77 ;
      RECT 7.5 3.282 7.855 3.765 ;
      RECT 7.46 3.29 7.855 3.74 ;
      RECT 7.46 3.317 7.87 3.738 ;
      RECT 7.46 3.347 7.88 3.725 ;
      RECT 7.455 3.492 7.88 3.713 ;
      RECT 7.46 3.421 7.9 3.71 ;
      RECT 7.46 3.478 7.905 3.518 ;
      RECT 7.65 2.757 7.82 2.935 ;
      RECT 7.6 2.696 7.65 2.92 ;
      RECT 7.335 2.676 7.6 2.905 ;
      RECT 7.295 2.74 7.77 2.905 ;
      RECT 7.295 2.73 7.725 2.905 ;
      RECT 7.295 2.727 7.715 2.905 ;
      RECT 7.295 2.715 7.705 2.905 ;
      RECT 7.295 2.7 7.65 2.905 ;
      RECT 7.335 2.672 7.536 2.905 ;
      RECT 7.345 2.65 7.536 2.905 ;
      RECT 7.37 2.635 7.45 2.905 ;
      RECT 7.125 3.165 7.245 3.61 ;
      RECT 7.11 3.165 7.245 3.609 ;
      RECT 7.065 3.187 7.245 3.604 ;
      RECT 7.025 3.236 7.245 3.598 ;
      RECT 7.025 3.236 7.25 3.573 ;
      RECT 7.025 3.236 7.27 3.463 ;
      RECT 7.02 3.266 7.27 3.46 ;
      RECT 7.11 3.165 7.28 3.355 ;
      RECT 6.77 1.95 6.775 2.395 ;
      RECT 6.58 1.95 6.6 2.36 ;
      RECT 6.55 1.95 6.555 2.335 ;
      RECT 7.23 2.257 7.245 2.445 ;
      RECT 7.225 2.242 7.23 2.451 ;
      RECT 7.205 2.215 7.225 2.454 ;
      RECT 7.155 2.182 7.205 2.463 ;
      RECT 7.125 2.162 7.155 2.467 ;
      RECT 7.106 2.15 7.125 2.463 ;
      RECT 7.02 2.122 7.106 2.453 ;
      RECT 7.01 2.097 7.02 2.443 ;
      RECT 6.94 2.065 7.01 2.435 ;
      RECT 6.915 2.025 6.94 2.427 ;
      RECT 6.895 2.007 6.915 2.421 ;
      RECT 6.885 1.997 6.895 2.418 ;
      RECT 6.875 1.99 6.885 2.416 ;
      RECT 6.855 1.977 6.875 2.413 ;
      RECT 6.845 1.967 6.855 2.41 ;
      RECT 6.835 1.96 6.845 2.408 ;
      RECT 6.785 1.952 6.835 2.402 ;
      RECT 6.775 1.95 6.785 2.396 ;
      RECT 6.745 1.95 6.77 2.393 ;
      RECT 6.716 1.95 6.745 2.388 ;
      RECT 6.63 1.95 6.716 2.378 ;
      RECT 6.6 1.95 6.63 2.365 ;
      RECT 6.555 1.95 6.58 2.348 ;
      RECT 6.54 1.95 6.55 2.33 ;
      RECT 6.52 1.957 6.54 2.315 ;
      RECT 6.515 1.972 6.52 2.303 ;
      RECT 6.51 1.977 6.515 2.243 ;
      RECT 6.505 1.982 6.51 2.085 ;
      RECT 6.5 1.985 6.505 2.003 ;
      RECT 6.765 2.67 6.851 2.991 ;
      RECT 6.765 2.67 6.885 2.984 ;
      RECT 6.715 2.67 6.885 2.98 ;
      RECT 6.715 2.672 6.971 2.978 ;
      RECT 6.715 2.674 6.995 2.972 ;
      RECT 6.715 2.681 7.005 2.971 ;
      RECT 6.715 2.69 7.01 2.968 ;
      RECT 6.715 2.696 7.015 2.963 ;
      RECT 6.715 2.74 7.02 2.96 ;
      RECT 6.715 2.832 7.025 2.957 ;
      RECT 6.24 3.275 6.275 3.595 ;
      RECT 6.825 3.46 6.83 3.642 ;
      RECT 6.78 3.342 6.825 3.661 ;
      RECT 6.765 3.319 6.78 3.684 ;
      RECT 6.755 3.309 6.765 3.694 ;
      RECT 6.735 3.304 6.755 3.707 ;
      RECT 6.71 3.302 6.735 3.728 ;
      RECT 6.691 3.301 6.71 3.74 ;
      RECT 6.605 3.298 6.691 3.74 ;
      RECT 6.535 3.293 6.605 3.728 ;
      RECT 6.46 3.289 6.535 3.703 ;
      RECT 6.395 3.285 6.46 3.67 ;
      RECT 6.325 3.282 6.395 3.63 ;
      RECT 6.295 3.278 6.325 3.605 ;
      RECT 6.275 3.276 6.295 3.598 ;
      RECT 6.191 3.274 6.24 3.596 ;
      RECT 6.105 3.271 6.191 3.597 ;
      RECT 6.03 3.27 6.105 3.599 ;
      RECT 5.945 3.27 6.03 3.625 ;
      RECT 5.868 3.271 5.945 3.65 ;
      RECT 5.782 3.272 5.868 3.65 ;
      RECT 5.696 3.272 5.782 3.65 ;
      RECT 5.61 3.273 5.696 3.65 ;
      RECT 5.59 3.274 5.61 3.642 ;
      RECT 5.575 3.28 5.59 3.627 ;
      RECT 5.54 3.3 5.575 3.607 ;
      RECT 5.53 3.32 5.54 3.589 ;
      RECT 6.5 2.625 6.505 2.895 ;
      RECT 6.495 2.616 6.5 2.9 ;
      RECT 6.485 2.606 6.495 2.912 ;
      RECT 6.48 2.595 6.485 2.923 ;
      RECT 6.46 2.589 6.48 2.941 ;
      RECT 6.415 2.586 6.46 2.99 ;
      RECT 6.4 2.585 6.415 3.035 ;
      RECT 6.395 2.585 6.4 3.048 ;
      RECT 6.385 2.585 6.395 3.06 ;
      RECT 6.38 2.586 6.385 3.075 ;
      RECT 6.36 2.594 6.38 3.08 ;
      RECT 6.33 2.61 6.36 3.08 ;
      RECT 6.32 2.622 6.325 3.08 ;
      RECT 6.285 2.637 6.32 3.08 ;
      RECT 6.255 2.657 6.285 3.08 ;
      RECT 6.245 2.682 6.255 3.08 ;
      RECT 6.24 2.71 6.245 3.08 ;
      RECT 6.235 2.74 6.24 3.08 ;
      RECT 6.23 2.757 6.235 3.08 ;
      RECT 6.22 2.785 6.23 3.08 ;
      RECT 6.21 2.82 6.22 3.08 ;
      RECT 6.205 2.855 6.21 3.08 ;
      RECT 6.325 2.62 6.33 3.08 ;
      RECT 5.84 2.722 6.025 2.895 ;
      RECT 5.8 2.64 5.985 2.893 ;
      RECT 5.761 2.645 5.985 2.889 ;
      RECT 5.675 2.654 5.985 2.884 ;
      RECT 5.591 2.67 5.99 2.879 ;
      RECT 5.505 2.69 6.015 2.873 ;
      RECT 5.505 2.71 6.02 2.873 ;
      RECT 5.591 2.68 6.015 2.879 ;
      RECT 5.675 2.655 5.99 2.884 ;
      RECT 5.84 2.637 5.985 2.895 ;
      RECT 5.84 2.632 5.94 2.895 ;
      RECT 5.926 2.626 5.94 2.895 ;
      RECT 5.315 1.95 5.32 2.349 ;
      RECT 5.06 1.95 5.095 2.347 ;
      RECT 4.655 1.985 4.66 2.341 ;
      RECT 5.4 1.988 5.405 2.243 ;
      RECT 5.395 1.986 5.4 2.249 ;
      RECT 5.39 1.985 5.395 2.256 ;
      RECT 5.365 1.978 5.39 2.28 ;
      RECT 5.36 1.971 5.365 2.304 ;
      RECT 5.355 1.967 5.36 2.313 ;
      RECT 5.345 1.962 5.355 2.326 ;
      RECT 5.34 1.959 5.345 2.335 ;
      RECT 5.335 1.957 5.34 2.34 ;
      RECT 5.32 1.953 5.335 2.35 ;
      RECT 5.305 1.947 5.315 2.349 ;
      RECT 5.267 1.945 5.305 2.349 ;
      RECT 5.181 1.947 5.267 2.349 ;
      RECT 5.095 1.949 5.181 2.348 ;
      RECT 5.024 1.95 5.06 2.347 ;
      RECT 4.938 1.952 5.024 2.347 ;
      RECT 4.852 1.954 4.938 2.346 ;
      RECT 4.766 1.956 4.852 2.346 ;
      RECT 4.68 1.959 4.766 2.345 ;
      RECT 4.67 1.965 4.68 2.344 ;
      RECT 4.66 1.977 4.67 2.342 ;
      RECT 4.6 2.012 4.655 2.338 ;
      RECT 4.595 2.042 4.6 2.1 ;
      RECT 5.34 3.122 5.355 3.315 ;
      RECT 5.335 3.09 5.34 3.315 ;
      RECT 5.325 3.065 5.335 3.315 ;
      RECT 5.32 3.037 5.325 3.315 ;
      RECT 5.29 2.96 5.32 3.315 ;
      RECT 5.265 2.842 5.29 3.315 ;
      RECT 5.26 2.78 5.265 3.315 ;
      RECT 5.25 2.767 5.26 3.315 ;
      RECT 5.23 2.757 5.25 3.315 ;
      RECT 5.215 2.74 5.23 3.315 ;
      RECT 5.185 2.728 5.215 3.315 ;
      RECT 5.18 2.727 5.185 3.26 ;
      RECT 5.175 2.727 5.18 3.218 ;
      RECT 5.16 2.726 5.175 3.17 ;
      RECT 5.145 2.726 5.16 3.108 ;
      RECT 5.125 2.726 5.145 3.068 ;
      RECT 5.12 2.726 5.125 3.053 ;
      RECT 5.095 2.725 5.12 3.048 ;
      RECT 5.025 2.724 5.095 3.035 ;
      RECT 5.01 2.723 5.025 3.02 ;
      RECT 4.98 2.722 5.01 3.003 ;
      RECT 4.975 2.722 4.98 2.988 ;
      RECT 4.925 2.721 4.975 2.968 ;
      RECT 4.86 2.72 4.925 2.923 ;
      RECT 4.855 2.72 4.86 2.895 ;
      RECT 4.94 3.257 4.945 3.514 ;
      RECT 4.92 3.176 4.94 3.531 ;
      RECT 4.9 3.17 4.92 3.56 ;
      RECT 4.84 3.157 4.9 3.58 ;
      RECT 4.795 3.141 4.84 3.581 ;
      RECT 4.711 3.129 4.795 3.569 ;
      RECT 4.625 3.116 4.711 3.553 ;
      RECT 4.615 3.109 4.625 3.545 ;
      RECT 4.57 3.106 4.615 3.485 ;
      RECT 4.55 3.102 4.57 3.4 ;
      RECT 4.535 3.1 4.55 3.353 ;
      RECT 4.505 3.097 4.535 3.323 ;
      RECT 4.47 3.093 4.505 3.3 ;
      RECT 4.427 3.088 4.47 3.288 ;
      RECT 4.341 3.079 4.427 3.297 ;
      RECT 4.255 3.068 4.341 3.309 ;
      RECT 4.19 3.059 4.255 3.318 ;
      RECT 4.17 3.05 4.19 3.323 ;
      RECT 4.165 3.043 4.17 3.325 ;
      RECT 4.125 3.028 4.165 3.322 ;
      RECT 4.105 3.007 4.125 3.317 ;
      RECT 4.09 2.995 4.105 3.31 ;
      RECT 4.085 2.987 4.09 3.303 ;
      RECT 4.07 2.967 4.085 3.296 ;
      RECT 4.065 2.83 4.07 3.29 ;
      RECT 3.985 2.719 4.065 3.262 ;
      RECT 3.976 2.712 3.985 3.228 ;
      RECT 3.89 2.706 3.976 3.153 ;
      RECT 3.865 2.697 3.89 3.065 ;
      RECT 3.835 2.692 3.865 3.04 ;
      RECT 3.77 2.701 3.835 3.025 ;
      RECT 3.75 2.717 3.77 3 ;
      RECT 3.74 2.723 3.75 2.948 ;
      RECT 3.72 2.745 3.74 2.83 ;
      RECT 4.375 2.71 4.545 2.895 ;
      RECT 4.375 2.71 4.58 2.893 ;
      RECT 4.425 2.62 4.595 2.884 ;
      RECT 4.375 2.777 4.6 2.877 ;
      RECT 4.39 2.655 4.595 2.884 ;
      RECT 3.59 3.388 3.655 3.831 ;
      RECT 3.53 3.413 3.655 3.829 ;
      RECT 3.53 3.413 3.71 3.823 ;
      RECT 3.515 3.438 3.71 3.822 ;
      RECT 3.655 3.375 3.73 3.819 ;
      RECT 3.59 3.4 3.81 3.813 ;
      RECT 3.515 3.439 3.855 3.807 ;
      RECT 3.5 3.466 3.855 3.798 ;
      RECT 3.515 3.459 3.875 3.79 ;
      RECT 3.5 3.468 3.88 3.773 ;
      RECT 3.495 3.485 3.88 3.6 ;
      RECT 3.5 2.207 3.535 2.445 ;
      RECT 3.5 2.207 3.565 2.444 ;
      RECT 3.5 2.207 3.68 2.44 ;
      RECT 3.5 2.207 3.735 2.418 ;
      RECT 3.51 2.15 3.79 2.318 ;
      RECT 3.615 1.99 3.645 2.441 ;
      RECT 3.645 1.985 3.825 2.198 ;
      RECT 3.515 2.126 3.825 2.198 ;
      RECT 3.565 2.022 3.615 2.442 ;
      RECT 3.535 2.078 3.825 2.198 ;
      RECT 1.33 7.855 1.5 8.305 ;
      RECT 1.385 6.075 1.555 8.025 ;
      RECT 1.33 5.015 1.5 6.245 ;
      RECT 0.81 5.015 0.98 8.305 ;
      RECT 0.81 7.315 1.215 7.645 ;
      RECT 0.81 6.475 1.215 6.805 ;
      RECT 92.035 0.575 92.205 1.085 ;
      RECT 92.035 2.395 92.205 3.865 ;
      RECT 92.035 5.015 92.205 6.485 ;
      RECT 92.035 7.795 92.205 8.305 ;
      RECT 91.045 0.575 91.215 1.085 ;
      RECT 91.045 2.395 91.215 3.865 ;
      RECT 91.045 5.015 91.215 6.485 ;
      RECT 91.045 7.795 91.215 8.305 ;
      RECT 89.68 0.575 89.85 3.865 ;
      RECT 89.68 5.015 89.85 8.305 ;
      RECT 89.25 0.575 89.42 1.085 ;
      RECT 89.25 1.655 89.42 3.865 ;
      RECT 89.25 5.015 89.42 7.225 ;
      RECT 89.25 7.795 89.42 8.305 ;
      RECT 87.88 1.66 88.05 2.935 ;
      RECT 87.88 5.945 88.05 7.22 ;
      RECT 84.92 5.015 85.09 8.305 ;
      RECT 84.49 5.015 84.66 7.225 ;
      RECT 84.49 7.795 84.66 8.305 ;
      RECT 83.12 5.945 83.29 7.22 ;
      RECT 74.11 0.575 74.28 1.085 ;
      RECT 74.11 2.395 74.28 3.865 ;
      RECT 74.11 5.015 74.28 6.485 ;
      RECT 74.11 7.795 74.28 8.305 ;
      RECT 73.12 0.575 73.29 1.085 ;
      RECT 73.12 2.395 73.29 3.865 ;
      RECT 73.12 5.015 73.29 6.485 ;
      RECT 73.12 7.795 73.29 8.305 ;
      RECT 71.755 0.575 71.925 3.865 ;
      RECT 71.755 5.015 71.925 8.305 ;
      RECT 71.325 0.575 71.495 1.085 ;
      RECT 71.325 1.655 71.495 3.865 ;
      RECT 71.325 5.015 71.495 7.225 ;
      RECT 71.325 7.795 71.495 8.305 ;
      RECT 69.955 1.66 70.125 2.935 ;
      RECT 69.955 5.945 70.125 7.22 ;
      RECT 66.995 5.015 67.165 8.305 ;
      RECT 66.565 5.015 66.735 7.225 ;
      RECT 66.565 7.795 66.735 8.305 ;
      RECT 65.195 5.945 65.365 7.22 ;
      RECT 56.185 0.575 56.355 1.085 ;
      RECT 56.185 2.395 56.355 3.865 ;
      RECT 56.185 5.015 56.355 6.485 ;
      RECT 56.185 7.795 56.355 8.305 ;
      RECT 55.195 0.575 55.365 1.085 ;
      RECT 55.195 2.395 55.365 3.865 ;
      RECT 55.195 5.015 55.365 6.485 ;
      RECT 55.195 7.795 55.365 8.305 ;
      RECT 53.83 0.575 54 3.865 ;
      RECT 53.83 5.015 54 8.305 ;
      RECT 53.4 0.575 53.57 1.085 ;
      RECT 53.4 1.655 53.57 3.865 ;
      RECT 53.4 5.015 53.57 7.225 ;
      RECT 53.4 7.795 53.57 8.305 ;
      RECT 52.03 1.66 52.2 2.935 ;
      RECT 52.03 5.945 52.2 7.22 ;
      RECT 49.07 5.015 49.24 8.305 ;
      RECT 48.64 5.015 48.81 7.225 ;
      RECT 48.64 7.795 48.81 8.305 ;
      RECT 47.27 5.945 47.44 7.22 ;
      RECT 38.26 0.575 38.43 1.085 ;
      RECT 38.26 2.395 38.43 3.865 ;
      RECT 38.26 5.015 38.43 6.485 ;
      RECT 38.26 7.795 38.43 8.305 ;
      RECT 37.27 0.575 37.44 1.085 ;
      RECT 37.27 2.395 37.44 3.865 ;
      RECT 37.27 5.015 37.44 6.485 ;
      RECT 37.27 7.795 37.44 8.305 ;
      RECT 35.905 0.575 36.075 3.865 ;
      RECT 35.905 5.015 36.075 8.305 ;
      RECT 35.475 0.575 35.645 1.085 ;
      RECT 35.475 1.655 35.645 3.865 ;
      RECT 35.475 5.015 35.645 7.225 ;
      RECT 35.475 7.795 35.645 8.305 ;
      RECT 34.105 1.66 34.275 2.935 ;
      RECT 34.105 5.945 34.275 7.22 ;
      RECT 31.145 5.015 31.315 8.305 ;
      RECT 30.715 5.015 30.885 7.225 ;
      RECT 30.715 7.795 30.885 8.305 ;
      RECT 29.345 5.945 29.515 7.22 ;
      RECT 20.335 0.575 20.505 1.085 ;
      RECT 20.335 2.395 20.505 3.865 ;
      RECT 20.335 5.015 20.505 6.485 ;
      RECT 20.335 7.795 20.505 8.305 ;
      RECT 19.345 0.575 19.515 1.085 ;
      RECT 19.345 2.395 19.515 3.865 ;
      RECT 19.345 5.015 19.515 6.485 ;
      RECT 19.345 7.795 19.515 8.305 ;
      RECT 17.98 0.575 18.15 3.865 ;
      RECT 17.98 5.015 18.15 8.305 ;
      RECT 17.55 0.575 17.72 1.085 ;
      RECT 17.55 1.655 17.72 3.865 ;
      RECT 17.55 5.015 17.72 7.225 ;
      RECT 17.55 7.795 17.72 8.305 ;
      RECT 16.18 1.66 16.35 2.935 ;
      RECT 16.18 5.945 16.35 7.22 ;
      RECT 13.22 5.015 13.39 8.305 ;
      RECT 12.79 5.015 12.96 7.225 ;
      RECT 12.79 7.795 12.96 8.305 ;
      RECT 11.42 5.945 11.59 7.22 ;
      RECT 1.76 5.015 1.93 7.225 ;
      RECT 1.76 7.795 1.93 8.305 ;
      RECT 0.39 5.945 0.56 7.22 ;
  END
END sky130_osu_ring_oscillator_mpr2at_8_b0r2

MACRO sky130_osu_ring_oscillator_mpr2ca_8_b0r1
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 0.025 0 ;
  SIZE 85.755 BY 8.88 ;
  SYMMETRY X Y R90 ;
  SITE CoreSite ;
  OBS
    LAYER met3 ;
      RECT 77.605 2.735 77.935 3.065 ;
      RECT 77.605 2.75 78.405 3.05 ;
      RECT 77.605 2.73 77.925 3.065 ;
      RECT 71.925 7.97 76.205 8.27 ;
      RECT 75.9 5.795 76.2 8.27 ;
      RECT 71.925 7.03 72.225 8.27 ;
      RECT 71.05 6.995 71.42 7.365 ;
      RECT 71.05 7.03 72.225 7.33 ;
      RECT 76.925 5.795 77.255 6.125 ;
      RECT 75.275 5.795 76.21 6.125 ;
      RECT 75.275 5.81 77.725 6.11 ;
      RECT 75.275 5.795 77.255 6.11 ;
      RECT 76.93 5.79 77.23 6.125 ;
      RECT 75.275 3.765 75.605 6.125 ;
      RECT 75.275 3.765 77.57 4.095 ;
      RECT 75.275 3.765 77.935 4.085 ;
      RECT 77.605 3.755 77.935 4.085 ;
      RECT 75.275 3.77 78.405 4.07 ;
      RECT 77.61 3.705 77.91 4.085 ;
      RECT 76.905 3.075 77.235 3.405 ;
      RECT 76.435 3.09 77.235 3.39 ;
      RECT 76.93 3.06 77.23 3.405 ;
      RECT 76.245 4.775 76.575 5.105 ;
      RECT 76.245 4.79 77.045 5.09 ;
      RECT 75.565 2.39 75.895 2.72 ;
      RECT 75.095 2.41 75.455 2.71 ;
      RECT 75.455 2.405 75.895 2.705 ;
      RECT 75.175 6.49 75.475 6.905 ;
      RECT 75.205 6.475 75.535 6.805 ;
      RECT 74.735 6.49 75.535 6.79 ;
      RECT 61.025 2.735 61.355 3.065 ;
      RECT 61.025 2.75 61.825 3.05 ;
      RECT 61.025 2.73 61.345 3.065 ;
      RECT 55.345 7.97 59.625 8.27 ;
      RECT 59.32 5.795 59.62 8.27 ;
      RECT 55.345 7.03 55.645 8.27 ;
      RECT 54.47 6.995 54.84 7.365 ;
      RECT 54.47 7.03 55.645 7.33 ;
      RECT 60.345 5.795 60.675 6.125 ;
      RECT 58.695 5.795 59.63 6.125 ;
      RECT 58.695 5.81 61.145 6.11 ;
      RECT 58.695 5.795 60.675 6.11 ;
      RECT 60.35 5.79 60.65 6.125 ;
      RECT 58.695 3.765 59.025 6.125 ;
      RECT 58.695 3.765 60.99 4.095 ;
      RECT 58.695 3.765 61.355 4.085 ;
      RECT 61.025 3.755 61.355 4.085 ;
      RECT 58.695 3.77 61.825 4.07 ;
      RECT 61.03 3.705 61.33 4.085 ;
      RECT 60.325 3.075 60.655 3.405 ;
      RECT 59.855 3.09 60.655 3.39 ;
      RECT 60.35 3.06 60.65 3.405 ;
      RECT 59.665 4.775 59.995 5.105 ;
      RECT 59.665 4.79 60.465 5.09 ;
      RECT 58.985 2.39 59.315 2.72 ;
      RECT 58.515 2.41 58.875 2.71 ;
      RECT 58.875 2.405 59.315 2.705 ;
      RECT 58.595 6.49 58.895 6.905 ;
      RECT 58.625 6.475 58.955 6.805 ;
      RECT 58.155 6.49 58.955 6.79 ;
      RECT 44.44 2.735 44.77 3.065 ;
      RECT 44.44 2.75 45.24 3.05 ;
      RECT 44.44 2.73 44.76 3.065 ;
      RECT 38.76 7.97 43.04 8.27 ;
      RECT 42.735 5.795 43.035 8.27 ;
      RECT 38.76 7.03 39.06 8.27 ;
      RECT 37.885 6.995 38.255 7.365 ;
      RECT 37.885 7.03 39.06 7.33 ;
      RECT 43.76 5.795 44.09 6.125 ;
      RECT 42.11 5.795 43.045 6.125 ;
      RECT 42.11 5.81 44.56 6.11 ;
      RECT 42.11 5.795 44.09 6.11 ;
      RECT 43.765 5.79 44.065 6.125 ;
      RECT 42.11 3.765 42.44 6.125 ;
      RECT 42.11 3.765 44.405 4.095 ;
      RECT 42.11 3.765 44.77 4.085 ;
      RECT 44.44 3.755 44.77 4.085 ;
      RECT 42.11 3.77 45.24 4.07 ;
      RECT 44.445 3.705 44.745 4.085 ;
      RECT 43.74 3.075 44.07 3.405 ;
      RECT 43.27 3.09 44.07 3.39 ;
      RECT 43.765 3.06 44.065 3.405 ;
      RECT 43.08 4.775 43.41 5.105 ;
      RECT 43.08 4.79 43.88 5.09 ;
      RECT 42.4 2.39 42.73 2.72 ;
      RECT 41.93 2.41 42.29 2.71 ;
      RECT 42.29 2.405 42.73 2.705 ;
      RECT 42.01 6.49 42.31 6.905 ;
      RECT 42.04 6.475 42.37 6.805 ;
      RECT 41.57 6.49 42.37 6.79 ;
      RECT 27.855 2.735 28.185 3.065 ;
      RECT 27.855 2.75 28.655 3.05 ;
      RECT 27.855 2.73 28.175 3.065 ;
      RECT 22.175 7.97 26.455 8.27 ;
      RECT 26.15 5.795 26.45 8.27 ;
      RECT 22.175 7.03 22.475 8.27 ;
      RECT 21.3 6.995 21.67 7.365 ;
      RECT 21.3 7.03 22.475 7.33 ;
      RECT 27.175 5.795 27.505 6.125 ;
      RECT 25.525 5.795 26.46 6.125 ;
      RECT 25.525 5.81 27.975 6.11 ;
      RECT 25.525 5.795 27.505 6.11 ;
      RECT 27.18 5.79 27.48 6.125 ;
      RECT 25.525 3.765 25.855 6.125 ;
      RECT 25.525 3.765 27.82 4.095 ;
      RECT 25.525 3.765 28.185 4.085 ;
      RECT 27.855 3.755 28.185 4.085 ;
      RECT 25.525 3.77 28.655 4.07 ;
      RECT 27.86 3.705 28.16 4.085 ;
      RECT 27.155 3.075 27.485 3.405 ;
      RECT 26.685 3.09 27.485 3.39 ;
      RECT 27.18 3.06 27.48 3.405 ;
      RECT 26.495 4.775 26.825 5.105 ;
      RECT 26.495 4.79 27.295 5.09 ;
      RECT 25.815 2.39 26.145 2.72 ;
      RECT 25.345 2.41 25.705 2.71 ;
      RECT 25.705 2.405 26.145 2.705 ;
      RECT 25.425 6.49 25.725 6.905 ;
      RECT 25.455 6.475 25.785 6.805 ;
      RECT 24.985 6.49 25.785 6.79 ;
      RECT 11.27 2.735 11.6 3.065 ;
      RECT 11.27 2.75 12.07 3.05 ;
      RECT 11.27 2.73 11.59 3.065 ;
      RECT 5.59 7.97 9.87 8.27 ;
      RECT 9.565 5.795 9.865 8.27 ;
      RECT 5.59 7.03 5.89 8.27 ;
      RECT 4.715 6.995 5.085 7.365 ;
      RECT 4.715 7.03 5.89 7.33 ;
      RECT 10.59 5.795 10.92 6.125 ;
      RECT 8.94 5.795 9.875 6.125 ;
      RECT 8.94 5.81 11.39 6.11 ;
      RECT 8.94 5.795 10.92 6.11 ;
      RECT 10.595 5.79 10.895 6.125 ;
      RECT 8.94 3.765 9.27 6.125 ;
      RECT 8.94 3.765 11.235 4.095 ;
      RECT 8.94 3.765 11.6 4.085 ;
      RECT 11.27 3.755 11.6 4.085 ;
      RECT 8.94 3.77 12.07 4.07 ;
      RECT 11.275 3.705 11.575 4.085 ;
      RECT 10.57 3.075 10.9 3.405 ;
      RECT 10.1 3.09 10.9 3.39 ;
      RECT 10.595 3.06 10.895 3.405 ;
      RECT 9.91 4.775 10.24 5.105 ;
      RECT 9.91 4.79 10.71 5.09 ;
      RECT 9.23 2.39 9.56 2.72 ;
      RECT 8.76 2.41 9.12 2.71 ;
      RECT 9.12 2.405 9.56 2.705 ;
      RECT 8.84 6.49 9.14 6.905 ;
      RECT 8.87 6.475 9.2 6.805 ;
      RECT 8.4 6.49 9.2 6.79 ;
    LAYER via2 ;
      RECT 77.67 2.8 77.87 3 ;
      RECT 77.67 3.82 77.87 4.02 ;
      RECT 76.99 5.86 77.19 6.06 ;
      RECT 76.97 3.14 77.17 3.34 ;
      RECT 76.31 4.84 76.51 5.04 ;
      RECT 75.945 5.86 76.145 6.06 ;
      RECT 75.63 2.455 75.83 2.655 ;
      RECT 75.27 6.54 75.47 6.74 ;
      RECT 71.135 7.08 71.335 7.28 ;
      RECT 61.09 2.8 61.29 3 ;
      RECT 61.09 3.82 61.29 4.02 ;
      RECT 60.41 5.86 60.61 6.06 ;
      RECT 60.39 3.14 60.59 3.34 ;
      RECT 59.73 4.84 59.93 5.04 ;
      RECT 59.365 5.86 59.565 6.06 ;
      RECT 59.05 2.455 59.25 2.655 ;
      RECT 58.69 6.54 58.89 6.74 ;
      RECT 54.555 7.08 54.755 7.28 ;
      RECT 44.505 2.8 44.705 3 ;
      RECT 44.505 3.82 44.705 4.02 ;
      RECT 43.825 5.86 44.025 6.06 ;
      RECT 43.805 3.14 44.005 3.34 ;
      RECT 43.145 4.84 43.345 5.04 ;
      RECT 42.78 5.86 42.98 6.06 ;
      RECT 42.465 2.455 42.665 2.655 ;
      RECT 42.105 6.54 42.305 6.74 ;
      RECT 37.97 7.08 38.17 7.28 ;
      RECT 27.92 2.8 28.12 3 ;
      RECT 27.92 3.82 28.12 4.02 ;
      RECT 27.24 5.86 27.44 6.06 ;
      RECT 27.22 3.14 27.42 3.34 ;
      RECT 26.56 4.84 26.76 5.04 ;
      RECT 26.195 5.86 26.395 6.06 ;
      RECT 25.88 2.455 26.08 2.655 ;
      RECT 25.52 6.54 25.72 6.74 ;
      RECT 21.385 7.08 21.585 7.28 ;
      RECT 11.335 2.8 11.535 3 ;
      RECT 11.335 3.82 11.535 4.02 ;
      RECT 10.655 5.86 10.855 6.06 ;
      RECT 10.635 3.14 10.835 3.34 ;
      RECT 9.975 4.84 10.175 5.04 ;
      RECT 9.61 5.86 9.81 6.06 ;
      RECT 9.295 2.455 9.495 2.655 ;
      RECT 8.935 6.54 9.135 6.74 ;
      RECT 4.8 7.08 5 7.28 ;
    LAYER met2 ;
      RECT 1.205 8.6 85.33 8.77 ;
      RECT 85.16 7.3 85.33 8.77 ;
      RECT 1.205 6.255 1.375 8.77 ;
      RECT 85.125 7.3 85.45 7.625 ;
      RECT 1.15 6.255 1.43 6.595 ;
      RECT 81.97 6.28 82.29 6.605 ;
      RECT 82 5.695 82.17 6.605 ;
      RECT 82 5.695 82.175 6.045 ;
      RECT 82 5.695 82.975 5.87 ;
      RECT 82.8 1.965 82.975 5.87 ;
      RECT 82.745 1.965 83.095 2.315 ;
      RECT 71.635 8.29 81.815 8.46 ;
      RECT 81.655 2.395 81.815 8.46 ;
      RECT 71.635 6.6 71.805 8.46 ;
      RECT 82.77 6.655 83.095 6.98 ;
      RECT 68.58 6.655 68.905 6.98 ;
      RECT 71.58 6.6 71.86 6.94 ;
      RECT 81.655 6.745 83.095 6.915 ;
      RECT 68.58 6.685 71.86 6.855 ;
      RECT 81.97 2.365 82.29 2.685 ;
      RECT 81.655 2.395 82.29 2.565 ;
      RECT 72.085 7.885 81.17 8.055 ;
      RECT 80.995 3.635 81.17 8.055 ;
      RECT 72.085 5.86 72.255 8.055 ;
      RECT 72.03 5.86 72.31 6.2 ;
      RECT 80.93 5.865 81.255 6.19 ;
      RECT 80.925 3.635 81.25 3.96 ;
      RECT 79.715 3.185 80.04 3.51 ;
      RECT 79.715 3.215 80.545 3.4 ;
      RECT 80.375 1.995 80.545 3.4 ;
      RECT 80.3 1.995 80.625 2.32 ;
      RECT 79.33 4.78 79.59 5.1 ;
      RECT 79.39 2.74 79.53 5.1 ;
      RECT 79.33 2.74 79.59 3.06 ;
      RECT 78.31 5.8 78.57 6.12 ;
      RECT 77.69 5.89 78.57 6.03 ;
      RECT 77.69 3.735 77.83 6.03 ;
      RECT 77.63 3.735 77.91 4.105 ;
      RECT 76.95 5.775 77.23 6.145 ;
      RECT 77.01 3.85 77.15 6.145 ;
      RECT 77.01 3.85 77.49 3.99 ;
      RECT 77.35 2.06 77.49 3.99 ;
      RECT 77.29 2.06 77.55 2.38 ;
      RECT 76.27 4.755 76.55 5.125 ;
      RECT 76.33 2.4 76.47 5.125 ;
      RECT 76.27 2.4 76.53 2.72 ;
      RECT 75.905 5.775 76.185 6.145 ;
      RECT 75.905 5.8 76.19 6.12 ;
      RECT 71.05 6.995 71.42 7.365 ;
      RECT 71.05 6.995 71.425 7.005 ;
      RECT 65.39 6.28 65.71 6.605 ;
      RECT 65.42 5.695 65.59 6.605 ;
      RECT 65.42 5.695 65.595 6.045 ;
      RECT 65.42 5.695 66.395 5.87 ;
      RECT 66.22 1.965 66.395 5.87 ;
      RECT 66.165 1.965 66.515 2.315 ;
      RECT 55.055 8.29 65.235 8.46 ;
      RECT 65.075 2.395 65.235 8.46 ;
      RECT 55.055 6.6 55.225 8.46 ;
      RECT 66.19 6.655 66.515 6.98 ;
      RECT 51.995 6.655 52.32 6.98 ;
      RECT 55 6.6 55.28 6.94 ;
      RECT 65.075 6.745 66.515 6.915 ;
      RECT 51.995 6.685 55.28 6.855 ;
      RECT 65.39 2.365 65.71 2.685 ;
      RECT 65.075 2.395 65.71 2.565 ;
      RECT 55.505 7.885 64.59 8.055 ;
      RECT 64.415 3.635 64.59 8.055 ;
      RECT 55.505 5.86 55.675 8.055 ;
      RECT 55.45 5.86 55.73 6.2 ;
      RECT 64.35 5.865 64.675 6.19 ;
      RECT 64.345 3.635 64.67 3.96 ;
      RECT 63.135 3.185 63.46 3.51 ;
      RECT 63.135 3.215 63.965 3.4 ;
      RECT 63.795 1.995 63.965 3.4 ;
      RECT 63.72 1.995 64.045 2.32 ;
      RECT 62.75 4.78 63.01 5.1 ;
      RECT 62.81 2.74 62.95 5.1 ;
      RECT 62.75 2.74 63.01 3.06 ;
      RECT 61.73 5.8 61.99 6.12 ;
      RECT 61.11 5.89 61.99 6.03 ;
      RECT 61.11 3.735 61.25 6.03 ;
      RECT 61.05 3.735 61.33 4.105 ;
      RECT 60.37 5.775 60.65 6.145 ;
      RECT 60.43 3.85 60.57 6.145 ;
      RECT 60.43 3.85 60.91 3.99 ;
      RECT 60.77 2.06 60.91 3.99 ;
      RECT 60.71 2.06 60.97 2.38 ;
      RECT 59.69 4.755 59.97 5.125 ;
      RECT 59.75 2.4 59.89 5.125 ;
      RECT 59.69 2.4 59.95 2.72 ;
      RECT 59.325 5.775 59.605 6.145 ;
      RECT 59.325 5.8 59.61 6.12 ;
      RECT 48.805 6.28 49.125 6.605 ;
      RECT 48.835 5.695 49.005 6.605 ;
      RECT 48.835 5.695 49.01 6.045 ;
      RECT 48.835 5.695 49.81 5.87 ;
      RECT 49.635 1.965 49.81 5.87 ;
      RECT 49.58 1.965 49.93 2.315 ;
      RECT 38.47 8.29 48.65 8.46 ;
      RECT 48.49 2.395 48.65 8.46 ;
      RECT 38.47 6.6 38.64 8.46 ;
      RECT 49.605 6.655 49.93 6.98 ;
      RECT 35.41 6.655 35.735 6.98 ;
      RECT 38.415 6.6 38.695 6.94 ;
      RECT 48.49 6.745 49.93 6.915 ;
      RECT 35.41 6.685 38.695 6.855 ;
      RECT 48.805 2.365 49.125 2.685 ;
      RECT 48.49 2.395 49.125 2.565 ;
      RECT 38.92 7.885 48.005 8.055 ;
      RECT 47.83 3.635 48.005 8.055 ;
      RECT 38.92 5.86 39.09 8.055 ;
      RECT 38.865 5.86 39.145 6.2 ;
      RECT 47.765 5.865 48.09 6.19 ;
      RECT 47.76 3.635 48.085 3.96 ;
      RECT 46.55 3.185 46.875 3.51 ;
      RECT 46.55 3.215 47.38 3.4 ;
      RECT 47.21 1.995 47.38 3.4 ;
      RECT 47.135 1.995 47.46 2.32 ;
      RECT 46.165 4.78 46.425 5.1 ;
      RECT 46.225 2.74 46.365 5.1 ;
      RECT 46.165 2.74 46.425 3.06 ;
      RECT 45.145 5.8 45.405 6.12 ;
      RECT 44.525 5.89 45.405 6.03 ;
      RECT 44.525 3.735 44.665 6.03 ;
      RECT 44.465 3.735 44.745 4.105 ;
      RECT 43.785 5.775 44.065 6.145 ;
      RECT 43.845 3.85 43.985 6.145 ;
      RECT 43.845 3.85 44.325 3.99 ;
      RECT 44.185 2.06 44.325 3.99 ;
      RECT 44.125 2.06 44.385 2.38 ;
      RECT 43.105 4.755 43.385 5.125 ;
      RECT 43.165 2.4 43.305 5.125 ;
      RECT 43.105 2.4 43.365 2.72 ;
      RECT 42.74 5.775 43.02 6.145 ;
      RECT 42.74 5.8 43.025 6.12 ;
      RECT 32.22 6.28 32.54 6.605 ;
      RECT 32.25 5.695 32.42 6.605 ;
      RECT 32.25 5.695 32.425 6.045 ;
      RECT 32.25 5.695 33.225 5.87 ;
      RECT 33.05 1.965 33.225 5.87 ;
      RECT 32.995 1.965 33.345 2.315 ;
      RECT 21.885 8.29 32.065 8.46 ;
      RECT 31.905 2.395 32.065 8.46 ;
      RECT 21.885 6.6 22.055 8.46 ;
      RECT 33.02 6.655 33.345 6.98 ;
      RECT 18.825 6.655 19.15 6.98 ;
      RECT 21.83 6.6 22.11 6.94 ;
      RECT 31.905 6.745 33.345 6.915 ;
      RECT 18.825 6.685 22.11 6.855 ;
      RECT 32.22 2.365 32.54 2.685 ;
      RECT 31.905 2.395 32.54 2.565 ;
      RECT 22.335 7.885 31.42 8.055 ;
      RECT 31.245 3.635 31.42 8.055 ;
      RECT 22.335 5.86 22.505 8.055 ;
      RECT 22.28 5.86 22.56 6.2 ;
      RECT 31.18 5.865 31.505 6.19 ;
      RECT 31.175 3.635 31.5 3.96 ;
      RECT 29.965 3.185 30.29 3.51 ;
      RECT 29.965 3.215 30.795 3.4 ;
      RECT 30.625 1.995 30.795 3.4 ;
      RECT 30.55 1.995 30.875 2.32 ;
      RECT 29.58 4.78 29.84 5.1 ;
      RECT 29.64 2.74 29.78 5.1 ;
      RECT 29.58 2.74 29.84 3.06 ;
      RECT 28.56 5.8 28.82 6.12 ;
      RECT 27.94 5.89 28.82 6.03 ;
      RECT 27.94 3.735 28.08 6.03 ;
      RECT 27.88 3.735 28.16 4.105 ;
      RECT 27.2 5.775 27.48 6.145 ;
      RECT 27.26 3.85 27.4 6.145 ;
      RECT 27.26 3.85 27.74 3.99 ;
      RECT 27.6 2.06 27.74 3.99 ;
      RECT 27.54 2.06 27.8 2.38 ;
      RECT 26.52 4.755 26.8 5.125 ;
      RECT 26.58 2.4 26.72 5.125 ;
      RECT 26.52 2.4 26.78 2.72 ;
      RECT 26.155 5.775 26.435 6.145 ;
      RECT 26.155 5.8 26.44 6.12 ;
      RECT 15.635 6.28 15.955 6.605 ;
      RECT 15.665 5.695 15.835 6.605 ;
      RECT 15.665 5.695 15.84 6.045 ;
      RECT 15.665 5.695 16.64 5.87 ;
      RECT 16.465 1.965 16.64 5.87 ;
      RECT 16.41 1.965 16.76 2.315 ;
      RECT 5.3 8.29 15.48 8.46 ;
      RECT 15.32 2.395 15.48 8.46 ;
      RECT 5.3 6.6 5.47 8.46 ;
      RECT 1.525 6.995 1.805 7.335 ;
      RECT 1.525 7.06 2.69 7.23 ;
      RECT 2.52 6.685 2.69 7.23 ;
      RECT 16.435 6.655 16.76 6.98 ;
      RECT 5.245 6.6 5.525 6.94 ;
      RECT 15.32 6.745 16.76 6.915 ;
      RECT 2.52 6.685 5.525 6.855 ;
      RECT 15.635 2.365 15.955 2.685 ;
      RECT 15.32 2.395 15.955 2.565 ;
      RECT 5.75 7.885 14.835 8.055 ;
      RECT 14.66 3.635 14.835 8.055 ;
      RECT 5.75 5.86 5.92 8.055 ;
      RECT 5.695 5.86 5.975 6.2 ;
      RECT 14.595 5.865 14.92 6.19 ;
      RECT 14.59 3.635 14.915 3.96 ;
      RECT 13.38 3.185 13.705 3.51 ;
      RECT 13.38 3.215 14.21 3.4 ;
      RECT 14.04 1.995 14.21 3.4 ;
      RECT 13.965 1.995 14.29 2.32 ;
      RECT 12.995 4.78 13.255 5.1 ;
      RECT 13.055 2.74 13.195 5.1 ;
      RECT 12.995 2.74 13.255 3.06 ;
      RECT 11.975 5.8 12.235 6.12 ;
      RECT 11.355 5.89 12.235 6.03 ;
      RECT 11.355 3.735 11.495 6.03 ;
      RECT 11.295 3.735 11.575 4.105 ;
      RECT 10.615 5.775 10.895 6.145 ;
      RECT 10.675 3.85 10.815 6.145 ;
      RECT 10.675 3.85 11.155 3.99 ;
      RECT 11.015 2.06 11.155 3.99 ;
      RECT 10.955 2.06 11.215 2.38 ;
      RECT 9.935 4.755 10.215 5.125 ;
      RECT 9.995 2.4 10.135 5.125 ;
      RECT 9.935 2.4 10.195 2.72 ;
      RECT 9.57 5.775 9.85 6.145 ;
      RECT 9.57 5.8 9.855 6.12 ;
      RECT 77.63 2.715 77.91 3.085 ;
      RECT 76.93 3.055 77.21 3.425 ;
      RECT 75.59 2.37 75.87 2.74 ;
      RECT 75.23 6.455 75.51 6.825 ;
      RECT 61.05 2.715 61.33 3.085 ;
      RECT 60.35 3.055 60.63 3.425 ;
      RECT 59.01 2.37 59.29 2.74 ;
      RECT 58.65 6.455 58.93 6.825 ;
      RECT 54.47 6.995 54.84 7.365 ;
      RECT 44.465 2.715 44.745 3.085 ;
      RECT 43.765 3.055 44.045 3.425 ;
      RECT 42.425 2.37 42.705 2.74 ;
      RECT 42.065 6.455 42.345 6.825 ;
      RECT 37.885 6.995 38.255 7.365 ;
      RECT 27.88 2.715 28.16 3.085 ;
      RECT 27.18 3.055 27.46 3.425 ;
      RECT 25.84 2.37 26.12 2.74 ;
      RECT 25.48 6.455 25.76 6.825 ;
      RECT 21.3 6.995 21.67 7.365 ;
      RECT 11.295 2.715 11.575 3.085 ;
      RECT 10.595 3.055 10.875 3.425 ;
      RECT 9.255 2.37 9.535 2.74 ;
      RECT 8.895 6.455 9.175 6.825 ;
      RECT 4.715 6.995 5.085 7.365 ;
    LAYER via1 ;
      RECT 85.215 7.385 85.365 7.535 ;
      RECT 82.86 6.74 83.01 6.89 ;
      RECT 82.845 2.065 82.995 2.215 ;
      RECT 82.055 2.45 82.205 2.6 ;
      RECT 82.055 6.37 82.205 6.52 ;
      RECT 81.02 5.95 81.17 6.1 ;
      RECT 81.015 3.72 81.165 3.87 ;
      RECT 80.39 2.08 80.54 2.23 ;
      RECT 79.805 3.27 79.955 3.42 ;
      RECT 79.385 2.825 79.535 2.975 ;
      RECT 79.385 4.865 79.535 5.015 ;
      RECT 78.365 5.885 78.515 6.035 ;
      RECT 77.685 2.825 77.835 2.975 ;
      RECT 77.685 3.845 77.835 3.995 ;
      RECT 77.345 2.145 77.495 2.295 ;
      RECT 77.005 3.165 77.155 3.315 ;
      RECT 77.005 5.885 77.155 6.035 ;
      RECT 76.325 2.485 76.475 2.635 ;
      RECT 76.325 4.865 76.475 5.015 ;
      RECT 75.985 5.885 76.135 6.035 ;
      RECT 75.645 2.48 75.795 2.63 ;
      RECT 75.305 6.565 75.455 6.715 ;
      RECT 72.095 5.955 72.245 6.105 ;
      RECT 71.645 6.695 71.795 6.845 ;
      RECT 71.16 7.105 71.31 7.255 ;
      RECT 68.67 6.74 68.82 6.89 ;
      RECT 66.28 6.74 66.43 6.89 ;
      RECT 66.265 2.065 66.415 2.215 ;
      RECT 65.475 2.45 65.625 2.6 ;
      RECT 65.475 6.37 65.625 6.52 ;
      RECT 64.44 5.95 64.59 6.1 ;
      RECT 64.435 3.72 64.585 3.87 ;
      RECT 63.81 2.08 63.96 2.23 ;
      RECT 63.225 3.27 63.375 3.42 ;
      RECT 62.805 2.825 62.955 2.975 ;
      RECT 62.805 4.865 62.955 5.015 ;
      RECT 61.785 5.885 61.935 6.035 ;
      RECT 61.105 2.825 61.255 2.975 ;
      RECT 61.105 3.845 61.255 3.995 ;
      RECT 60.765 2.145 60.915 2.295 ;
      RECT 60.425 3.165 60.575 3.315 ;
      RECT 60.425 5.885 60.575 6.035 ;
      RECT 59.745 2.485 59.895 2.635 ;
      RECT 59.745 4.865 59.895 5.015 ;
      RECT 59.405 5.885 59.555 6.035 ;
      RECT 59.065 2.48 59.215 2.63 ;
      RECT 58.725 6.565 58.875 6.715 ;
      RECT 55.515 5.955 55.665 6.105 ;
      RECT 55.065 6.695 55.215 6.845 ;
      RECT 54.58 7.105 54.73 7.255 ;
      RECT 52.085 6.74 52.235 6.89 ;
      RECT 49.695 6.74 49.845 6.89 ;
      RECT 49.68 2.065 49.83 2.215 ;
      RECT 48.89 2.45 49.04 2.6 ;
      RECT 48.89 6.37 49.04 6.52 ;
      RECT 47.855 5.95 48.005 6.1 ;
      RECT 47.85 3.72 48 3.87 ;
      RECT 47.225 2.08 47.375 2.23 ;
      RECT 46.64 3.27 46.79 3.42 ;
      RECT 46.22 2.825 46.37 2.975 ;
      RECT 46.22 4.865 46.37 5.015 ;
      RECT 45.2 5.885 45.35 6.035 ;
      RECT 44.52 2.825 44.67 2.975 ;
      RECT 44.52 3.845 44.67 3.995 ;
      RECT 44.18 2.145 44.33 2.295 ;
      RECT 43.84 3.165 43.99 3.315 ;
      RECT 43.84 5.885 43.99 6.035 ;
      RECT 43.16 2.485 43.31 2.635 ;
      RECT 43.16 4.865 43.31 5.015 ;
      RECT 42.82 5.885 42.97 6.035 ;
      RECT 42.48 2.48 42.63 2.63 ;
      RECT 42.14 6.565 42.29 6.715 ;
      RECT 38.93 5.955 39.08 6.105 ;
      RECT 38.48 6.695 38.63 6.845 ;
      RECT 37.995 7.105 38.145 7.255 ;
      RECT 35.5 6.74 35.65 6.89 ;
      RECT 33.11 6.74 33.26 6.89 ;
      RECT 33.095 2.065 33.245 2.215 ;
      RECT 32.305 2.45 32.455 2.6 ;
      RECT 32.305 6.37 32.455 6.52 ;
      RECT 31.27 5.95 31.42 6.1 ;
      RECT 31.265 3.72 31.415 3.87 ;
      RECT 30.64 2.08 30.79 2.23 ;
      RECT 30.055 3.27 30.205 3.42 ;
      RECT 29.635 2.825 29.785 2.975 ;
      RECT 29.635 4.865 29.785 5.015 ;
      RECT 28.615 5.885 28.765 6.035 ;
      RECT 27.935 2.825 28.085 2.975 ;
      RECT 27.935 3.845 28.085 3.995 ;
      RECT 27.595 2.145 27.745 2.295 ;
      RECT 27.255 3.165 27.405 3.315 ;
      RECT 27.255 5.885 27.405 6.035 ;
      RECT 26.575 2.485 26.725 2.635 ;
      RECT 26.575 4.865 26.725 5.015 ;
      RECT 26.235 5.885 26.385 6.035 ;
      RECT 25.895 2.48 26.045 2.63 ;
      RECT 25.555 6.565 25.705 6.715 ;
      RECT 22.345 5.955 22.495 6.105 ;
      RECT 21.895 6.695 22.045 6.845 ;
      RECT 21.41 7.105 21.56 7.255 ;
      RECT 18.915 6.74 19.065 6.89 ;
      RECT 16.525 6.74 16.675 6.89 ;
      RECT 16.51 2.065 16.66 2.215 ;
      RECT 15.72 2.45 15.87 2.6 ;
      RECT 15.72 6.37 15.87 6.52 ;
      RECT 14.685 5.95 14.835 6.1 ;
      RECT 14.68 3.72 14.83 3.87 ;
      RECT 14.055 2.08 14.205 2.23 ;
      RECT 13.47 3.27 13.62 3.42 ;
      RECT 13.05 2.825 13.2 2.975 ;
      RECT 13.05 4.865 13.2 5.015 ;
      RECT 12.03 5.885 12.18 6.035 ;
      RECT 11.35 2.825 11.5 2.975 ;
      RECT 11.35 3.845 11.5 3.995 ;
      RECT 11.01 2.145 11.16 2.295 ;
      RECT 10.67 3.165 10.82 3.315 ;
      RECT 10.67 5.885 10.82 6.035 ;
      RECT 9.99 2.485 10.14 2.635 ;
      RECT 9.99 4.865 10.14 5.015 ;
      RECT 9.65 5.885 9.8 6.035 ;
      RECT 9.31 2.48 9.46 2.63 ;
      RECT 8.97 6.565 9.12 6.715 ;
      RECT 5.76 5.955 5.91 6.105 ;
      RECT 5.31 6.695 5.46 6.845 ;
      RECT 4.825 7.105 4.975 7.255 ;
      RECT 1.59 7.09 1.74 7.24 ;
      RECT 1.215 6.35 1.365 6.5 ;
    LAYER met1 ;
      RECT 0.025 8.57 85.73 8.88 ;
      RECT 72.535 7.18 79.735 8.88 ;
      RECT 70.555 6.315 70.725 8.88 ;
      RECT 55.955 7.18 63.155 8.88 ;
      RECT 53.975 6.315 54.145 8.88 ;
      RECT 39.37 7.18 46.57 8.88 ;
      RECT 37.39 6.315 37.56 8.88 ;
      RECT 22.785 7.18 29.985 8.88 ;
      RECT 20.805 6.315 20.975 8.88 ;
      RECT 6.2 7.18 13.4 8.88 ;
      RECT 4.22 6.315 4.39 8.88 ;
      RECT 72.83 6.91 79.73 8.88 ;
      RECT 56.25 6.91 63.15 8.88 ;
      RECT 39.665 6.91 46.565 8.88 ;
      RECT 23.08 6.91 29.98 8.88 ;
      RECT 6.495 6.91 13.395 8.88 ;
      RECT 75.255 6.51 75.51 8.88 ;
      RECT 58.675 6.51 58.93 8.88 ;
      RECT 42.09 6.51 42.345 8.88 ;
      RECT 25.505 6.51 25.76 8.88 ;
      RECT 8.92 6.51 9.175 8.88 ;
      RECT 75.22 6.51 75.54 6.77 ;
      RECT 58.64 6.51 58.96 6.77 ;
      RECT 42.055 6.51 42.375 6.77 ;
      RECT 25.47 6.51 25.79 6.77 ;
      RECT 8.885 6.51 9.205 6.77 ;
      RECT 74.29 6.57 76.64 6.71 ;
      RECT 76.5 5.845 76.64 6.71 ;
      RECT 57.71 6.57 60.06 6.71 ;
      RECT 59.92 5.845 60.06 6.71 ;
      RECT 41.125 6.57 43.475 6.71 ;
      RECT 43.335 5.845 43.475 6.71 ;
      RECT 24.54 6.57 26.89 6.71 ;
      RECT 26.75 5.845 26.89 6.71 ;
      RECT 7.955 6.57 10.305 6.71 ;
      RECT 10.165 5.845 10.305 6.71 ;
      RECT 74.29 5.845 74.43 6.71 ;
      RECT 57.71 5.845 57.85 6.71 ;
      RECT 41.125 5.845 41.265 6.71 ;
      RECT 24.54 5.845 24.68 6.71 ;
      RECT 7.955 5.845 8.095 6.71 ;
      RECT 70.715 6.285 71.005 6.515 ;
      RECT 54.135 6.285 54.425 6.515 ;
      RECT 37.55 6.285 37.84 6.515 ;
      RECT 20.965 6.285 21.255 6.515 ;
      RECT 4.38 6.285 4.67 6.515 ;
      RECT 70.545 6.315 71.005 6.485 ;
      RECT 53.965 6.315 54.425 6.485 ;
      RECT 37.38 6.315 37.84 6.485 ;
      RECT 20.795 6.315 21.255 6.485 ;
      RECT 4.21 6.315 4.67 6.485 ;
      RECT 76.425 5.845 76.715 6.075 ;
      RECT 74.215 5.845 74.505 6.075 ;
      RECT 59.845 5.845 60.135 6.075 ;
      RECT 57.635 5.845 57.925 6.075 ;
      RECT 43.26 5.845 43.55 6.075 ;
      RECT 41.05 5.845 41.34 6.075 ;
      RECT 26.675 5.845 26.965 6.075 ;
      RECT 24.465 5.845 24.755 6.075 ;
      RECT 10.09 5.845 10.38 6.075 ;
      RECT 7.88 5.845 8.17 6.075 ;
      RECT 72.83 0 79.73 1.95 ;
      RECT 56.25 0 63.15 1.95 ;
      RECT 39.665 0 46.565 1.95 ;
      RECT 23.08 0 29.98 1.95 ;
      RECT 6.495 0 13.395 1.95 ;
      RECT 72.83 0 79.92 1.795 ;
      RECT 56.25 0 63.34 1.795 ;
      RECT 39.665 0 46.755 1.795 ;
      RECT 23.08 0 30.17 1.795 ;
      RECT 6.495 0 13.585 1.795 ;
      RECT 72.575 0 79.92 1.655 ;
      RECT 55.995 0 63.34 1.655 ;
      RECT 39.41 0 46.755 1.655 ;
      RECT 22.825 0 30.17 1.655 ;
      RECT 6.24 0 13.585 1.655 ;
      RECT 0 0 85.705 0.31 ;
      RECT 79.76 4.15 85.7 4.745 ;
      RECT 80.22 4.135 85.7 4.745 ;
      RECT 69.595 4.13 72.345 4.745 ;
      RECT 63.18 4.15 69.12 4.745 ;
      RECT 53.015 4.13 55.765 4.745 ;
      RECT 46.595 4.15 52.535 4.745 ;
      RECT 36.43 4.13 39.18 4.745 ;
      RECT 30.01 4.15 35.95 4.745 ;
      RECT 19.845 4.13 22.595 4.745 ;
      RECT 13.425 4.15 19.365 4.745 ;
      RECT 3.26 4.13 6.01 4.745 ;
      RECT 0.03 4.13 2.78 4.745 ;
      RECT 69.115 4.13 72.69 4.74 ;
      RECT 52.535 4.13 56.11 4.74 ;
      RECT 35.95 4.13 39.525 4.74 ;
      RECT 19.365 4.13 22.94 4.74 ;
      RECT 0.03 4.13 6.355 4.74 ;
      RECT 0.03 4.19 85.7 4.67 ;
      RECT 79.63 4.15 85.7 4.67 ;
      RECT 63.05 4.15 72.69 4.67 ;
      RECT 46.465 4.15 56.11 4.67 ;
      RECT 29.88 4.15 39.525 4.67 ;
      RECT 13.295 4.15 22.94 4.67 ;
      RECT 63.64 4.135 72.69 4.74 ;
      RECT 47.055 4.135 56.11 4.74 ;
      RECT 30.47 4.135 39.525 4.74 ;
      RECT 13.885 4.135 22.94 4.74 ;
      RECT 85.1 7.765 85.39 7.995 ;
      RECT 85.16 6.285 85.33 7.995 ;
      RECT 85.125 7.3 85.45 7.625 ;
      RECT 85.1 6.285 85.39 6.515 ;
      RECT 85.1 2.365 85.39 2.595 ;
      RECT 85.16 0.885 85.33 2.595 ;
      RECT 85.1 0.885 85.39 1.115 ;
      RECT 84.69 2.735 85.02 2.965 ;
      RECT 84.69 2.765 85.19 2.935 ;
      RECT 84.69 2.395 84.88 2.965 ;
      RECT 84.11 2.365 84.4 2.595 ;
      RECT 84.11 2.395 84.88 2.565 ;
      RECT 84.17 0.885 84.34 2.595 ;
      RECT 84.11 0.885 84.4 1.115 ;
      RECT 84.11 7.765 84.4 7.995 ;
      RECT 84.17 6.285 84.34 7.995 ;
      RECT 84.11 6.285 84.4 6.515 ;
      RECT 84.11 6.325 84.96 6.485 ;
      RECT 84.79 5.915 84.96 6.485 ;
      RECT 84.11 6.32 84.5 6.485 ;
      RECT 84.73 5.915 85.02 6.145 ;
      RECT 84.73 5.945 85.19 6.115 ;
      RECT 83.74 2.735 84.03 2.965 ;
      RECT 83.74 2.765 84.2 2.935 ;
      RECT 83.8 1.655 83.965 2.965 ;
      RECT 82.315 1.625 82.605 1.855 ;
      RECT 82.315 1.655 83.965 1.825 ;
      RECT 82.375 0.885 82.545 1.855 ;
      RECT 82.315 0.885 82.605 1.115 ;
      RECT 82.315 7.765 82.605 7.995 ;
      RECT 82.375 7.025 82.545 7.995 ;
      RECT 82.375 7.12 83.965 7.29 ;
      RECT 83.795 5.915 83.965 7.29 ;
      RECT 82.315 7.025 82.605 7.255 ;
      RECT 83.74 5.915 84.03 6.145 ;
      RECT 83.74 5.945 84.2 6.115 ;
      RECT 80.3 1.995 80.625 2.32 ;
      RECT 82.745 1.965 83.095 2.315 ;
      RECT 80.3 2.025 83.095 2.195 ;
      RECT 82.77 6.655 83.095 6.98 ;
      RECT 82.745 6.655 83.095 6.885 ;
      RECT 82.575 6.685 83.095 6.855 ;
      RECT 81.97 2.365 82.29 2.685 ;
      RECT 81.94 2.365 82.29 2.595 ;
      RECT 81.655 2.395 82.29 2.565 ;
      RECT 81.97 6.28 82.29 6.605 ;
      RECT 81.94 6.285 82.29 6.515 ;
      RECT 81.77 6.315 82.29 6.485 ;
      RECT 80.925 3.635 81.25 3.96 ;
      RECT 81 2.735 81.18 3.96 ;
      RECT 80.945 2.735 81.235 2.965 ;
      RECT 80.945 2.765 81.405 2.935 ;
      RECT 80.93 5.865 81.255 6.19 ;
      RECT 80.93 5.945 81.405 6.115 ;
      RECT 79.715 3.185 80.04 3.51 ;
      RECT 76.92 3.11 77.24 3.37 ;
      RECT 78.895 3.125 79.185 3.355 ;
      RECT 79.615 3.185 80.04 3.325 ;
      RECT 76.92 3.17 79.755 3.31 ;
      RECT 79.3 2.77 79.62 3.03 ;
      RECT 79.025 2.83 79.62 2.97 ;
      RECT 78.28 5.83 78.6 6.09 ;
      RECT 78.28 5.89 78.875 6.03 ;
      RECT 77.6 2.77 77.92 3.03 ;
      RECT 72.86 2.785 73.15 3.015 ;
      RECT 72.86 2.83 77.92 2.97 ;
      RECT 77.69 2.49 77.83 3.03 ;
      RECT 77.69 2.49 78.17 2.63 ;
      RECT 78.03 2.105 78.17 2.63 ;
      RECT 77.955 2.105 78.245 2.335 ;
      RECT 77.6 3.79 77.92 4.05 ;
      RECT 76.935 3.805 77.225 4.035 ;
      RECT 74.725 3.805 75.015 4.035 ;
      RECT 74.725 3.85 77.92 3.99 ;
      RECT 75.9 5.83 76.22 6.09 ;
      RECT 77.615 5.845 77.905 6.075 ;
      RECT 75.235 5.845 75.525 6.075 ;
      RECT 75.235 5.89 76.22 6.03 ;
      RECT 77.69 5.55 77.83 6.075 ;
      RECT 75.99 5.55 76.13 6.09 ;
      RECT 75.99 5.55 77.83 5.69 ;
      RECT 74.895 2.445 75.185 2.675 ;
      RECT 74.97 2.15 75.11 2.675 ;
      RECT 77.26 2.09 77.58 2.35 ;
      RECT 77.16 2.105 77.58 2.335 ;
      RECT 74.97 2.15 77.58 2.29 ;
      RECT 76.24 2.43 76.56 2.69 ;
      RECT 76.24 2.49 76.835 2.63 ;
      RECT 76.24 4.81 76.56 5.07 ;
      RECT 73.535 4.825 73.825 5.055 ;
      RECT 73.535 4.87 76.56 5.01 ;
      RECT 75.565 2.39 75.895 2.72 ;
      RECT 75.56 2.425 75.895 2.685 ;
      RECT 75.91 2.445 76.025 2.675 ;
      RECT 75.56 2.44 75.91 2.67 ;
      RECT 75.56 2.49 76.04 2.63 ;
      RECT 75.445 2.49 75.455 2.63 ;
      RECT 75.455 2.485 76.025 2.625 ;
      RECT 72 5.89 72.34 6.17 ;
      RECT 69.72 5.915 70.01 6.145 ;
      RECT 69.72 5.945 72.34 6.115 ;
      RECT 71.55 6.63 71.89 6.91 ;
      RECT 71.52 6.655 71.89 6.885 ;
      RECT 71.35 6.685 71.89 6.855 ;
      RECT 71.09 7.765 71.38 7.995 ;
      RECT 71.15 6.995 71.32 7.995 ;
      RECT 71.05 6.995 71.42 7.365 ;
      RECT 68.52 7.765 68.81 7.995 ;
      RECT 68.58 6.285 68.75 7.995 ;
      RECT 68.58 6.655 68.905 6.98 ;
      RECT 68.52 6.285 68.81 6.515 ;
      RECT 68.52 2.365 68.81 2.595 ;
      RECT 68.58 0.885 68.75 2.595 ;
      RECT 68.52 0.885 68.81 1.115 ;
      RECT 68.11 2.735 68.44 2.965 ;
      RECT 68.11 2.765 68.61 2.935 ;
      RECT 68.11 2.395 68.3 2.965 ;
      RECT 67.53 2.365 67.82 2.595 ;
      RECT 67.53 2.395 68.3 2.565 ;
      RECT 67.59 0.885 67.76 2.595 ;
      RECT 67.53 0.885 67.82 1.115 ;
      RECT 67.53 7.765 67.82 7.995 ;
      RECT 67.59 6.285 67.76 7.995 ;
      RECT 67.53 6.285 67.82 6.515 ;
      RECT 67.53 6.325 68.38 6.485 ;
      RECT 68.21 5.915 68.38 6.485 ;
      RECT 67.53 6.32 67.92 6.485 ;
      RECT 68.15 5.915 68.44 6.145 ;
      RECT 68.15 5.945 68.61 6.115 ;
      RECT 67.16 2.735 67.45 2.965 ;
      RECT 67.16 2.765 67.62 2.935 ;
      RECT 67.22 1.655 67.385 2.965 ;
      RECT 65.735 1.625 66.025 1.855 ;
      RECT 65.735 1.655 67.385 1.825 ;
      RECT 65.795 0.885 65.965 1.855 ;
      RECT 65.735 0.885 66.025 1.115 ;
      RECT 65.735 7.765 66.025 7.995 ;
      RECT 65.795 7.025 65.965 7.995 ;
      RECT 65.795 7.12 67.385 7.29 ;
      RECT 67.215 5.915 67.385 7.29 ;
      RECT 65.735 7.025 66.025 7.255 ;
      RECT 67.16 5.915 67.45 6.145 ;
      RECT 67.16 5.945 67.62 6.115 ;
      RECT 63.72 1.995 64.045 2.32 ;
      RECT 66.165 1.965 66.515 2.315 ;
      RECT 63.72 2.025 66.515 2.195 ;
      RECT 66.19 6.655 66.515 6.98 ;
      RECT 66.165 6.655 66.515 6.885 ;
      RECT 65.995 6.685 66.515 6.855 ;
      RECT 65.39 2.365 65.71 2.685 ;
      RECT 65.36 2.365 65.71 2.595 ;
      RECT 65.075 2.395 65.71 2.565 ;
      RECT 65.39 6.28 65.71 6.605 ;
      RECT 65.36 6.285 65.71 6.515 ;
      RECT 65.19 6.315 65.71 6.485 ;
      RECT 64.345 3.635 64.67 3.96 ;
      RECT 64.42 2.735 64.6 3.96 ;
      RECT 64.365 2.735 64.655 2.965 ;
      RECT 64.365 2.765 64.825 2.935 ;
      RECT 64.35 5.865 64.675 6.19 ;
      RECT 64.35 5.945 64.825 6.115 ;
      RECT 63.135 3.185 63.46 3.51 ;
      RECT 60.34 3.11 60.66 3.37 ;
      RECT 62.315 3.125 62.605 3.355 ;
      RECT 63.035 3.185 63.46 3.325 ;
      RECT 60.34 3.17 63.175 3.31 ;
      RECT 62.72 2.77 63.04 3.03 ;
      RECT 62.445 2.83 63.04 2.97 ;
      RECT 61.7 5.83 62.02 6.09 ;
      RECT 61.7 5.89 62.295 6.03 ;
      RECT 61.02 2.77 61.34 3.03 ;
      RECT 56.28 2.785 56.57 3.015 ;
      RECT 56.28 2.83 61.34 2.97 ;
      RECT 61.11 2.49 61.25 3.03 ;
      RECT 61.11 2.49 61.59 2.63 ;
      RECT 61.45 2.105 61.59 2.63 ;
      RECT 61.375 2.105 61.665 2.335 ;
      RECT 61.02 3.79 61.34 4.05 ;
      RECT 60.355 3.805 60.645 4.035 ;
      RECT 58.145 3.805 58.435 4.035 ;
      RECT 58.145 3.85 61.34 3.99 ;
      RECT 59.32 5.83 59.64 6.09 ;
      RECT 61.035 5.845 61.325 6.075 ;
      RECT 58.655 5.845 58.945 6.075 ;
      RECT 58.655 5.89 59.64 6.03 ;
      RECT 61.11 5.55 61.25 6.075 ;
      RECT 59.41 5.55 59.55 6.09 ;
      RECT 59.41 5.55 61.25 5.69 ;
      RECT 58.315 2.445 58.605 2.675 ;
      RECT 58.39 2.15 58.53 2.675 ;
      RECT 60.68 2.09 61 2.35 ;
      RECT 60.58 2.105 61 2.335 ;
      RECT 58.39 2.15 61 2.29 ;
      RECT 59.66 2.43 59.98 2.69 ;
      RECT 59.66 2.49 60.255 2.63 ;
      RECT 59.66 4.81 59.98 5.07 ;
      RECT 56.955 4.825 57.245 5.055 ;
      RECT 56.955 4.87 59.98 5.01 ;
      RECT 58.985 2.39 59.315 2.72 ;
      RECT 58.98 2.425 59.315 2.685 ;
      RECT 59.33 2.445 59.445 2.675 ;
      RECT 58.98 2.44 59.33 2.67 ;
      RECT 58.98 2.49 59.46 2.63 ;
      RECT 58.865 2.49 58.875 2.63 ;
      RECT 58.875 2.485 59.445 2.625 ;
      RECT 55.42 5.89 55.76 6.17 ;
      RECT 53.14 5.915 53.43 6.145 ;
      RECT 53.14 5.945 55.76 6.115 ;
      RECT 54.97 6.63 55.31 6.91 ;
      RECT 54.94 6.655 55.31 6.885 ;
      RECT 54.77 6.685 55.31 6.855 ;
      RECT 54.51 7.765 54.8 7.995 ;
      RECT 54.57 6.995 54.74 7.995 ;
      RECT 54.47 6.995 54.84 7.365 ;
      RECT 51.935 7.765 52.225 7.995 ;
      RECT 51.995 6.285 52.165 7.995 ;
      RECT 51.995 6.655 52.32 6.98 ;
      RECT 51.935 6.285 52.225 6.515 ;
      RECT 51.935 2.365 52.225 2.595 ;
      RECT 51.995 0.885 52.165 2.595 ;
      RECT 51.935 0.885 52.225 1.115 ;
      RECT 51.525 2.735 51.855 2.965 ;
      RECT 51.525 2.765 52.025 2.935 ;
      RECT 51.525 2.395 51.715 2.965 ;
      RECT 50.945 2.365 51.235 2.595 ;
      RECT 50.945 2.395 51.715 2.565 ;
      RECT 51.005 0.885 51.175 2.595 ;
      RECT 50.945 0.885 51.235 1.115 ;
      RECT 50.945 7.765 51.235 7.995 ;
      RECT 51.005 6.285 51.175 7.995 ;
      RECT 50.945 6.285 51.235 6.515 ;
      RECT 50.945 6.325 51.795 6.485 ;
      RECT 51.625 5.915 51.795 6.485 ;
      RECT 50.945 6.32 51.335 6.485 ;
      RECT 51.565 5.915 51.855 6.145 ;
      RECT 51.565 5.945 52.025 6.115 ;
      RECT 50.575 2.735 50.865 2.965 ;
      RECT 50.575 2.765 51.035 2.935 ;
      RECT 50.635 1.655 50.8 2.965 ;
      RECT 49.15 1.625 49.44 1.855 ;
      RECT 49.15 1.655 50.8 1.825 ;
      RECT 49.21 0.885 49.38 1.855 ;
      RECT 49.15 0.885 49.44 1.115 ;
      RECT 49.15 7.765 49.44 7.995 ;
      RECT 49.21 7.025 49.38 7.995 ;
      RECT 49.21 7.12 50.8 7.29 ;
      RECT 50.63 5.915 50.8 7.29 ;
      RECT 49.15 7.025 49.44 7.255 ;
      RECT 50.575 5.915 50.865 6.145 ;
      RECT 50.575 5.945 51.035 6.115 ;
      RECT 47.135 1.995 47.46 2.32 ;
      RECT 49.58 1.965 49.93 2.315 ;
      RECT 47.135 2.025 49.93 2.195 ;
      RECT 49.605 6.655 49.93 6.98 ;
      RECT 49.58 6.655 49.93 6.885 ;
      RECT 49.41 6.685 49.93 6.855 ;
      RECT 48.805 2.365 49.125 2.685 ;
      RECT 48.775 2.365 49.125 2.595 ;
      RECT 48.49 2.395 49.125 2.565 ;
      RECT 48.805 6.28 49.125 6.605 ;
      RECT 48.775 6.285 49.125 6.515 ;
      RECT 48.605 6.315 49.125 6.485 ;
      RECT 47.76 3.635 48.085 3.96 ;
      RECT 47.835 2.735 48.015 3.96 ;
      RECT 47.78 2.735 48.07 2.965 ;
      RECT 47.78 2.765 48.24 2.935 ;
      RECT 47.765 5.865 48.09 6.19 ;
      RECT 47.765 5.945 48.24 6.115 ;
      RECT 46.55 3.185 46.875 3.51 ;
      RECT 43.755 3.11 44.075 3.37 ;
      RECT 45.73 3.125 46.02 3.355 ;
      RECT 46.45 3.185 46.875 3.325 ;
      RECT 43.755 3.17 46.59 3.31 ;
      RECT 46.135 2.77 46.455 3.03 ;
      RECT 45.86 2.83 46.455 2.97 ;
      RECT 45.115 5.83 45.435 6.09 ;
      RECT 45.115 5.89 45.71 6.03 ;
      RECT 44.435 2.77 44.755 3.03 ;
      RECT 39.695 2.785 39.985 3.015 ;
      RECT 39.695 2.83 44.755 2.97 ;
      RECT 44.525 2.49 44.665 3.03 ;
      RECT 44.525 2.49 45.005 2.63 ;
      RECT 44.865 2.105 45.005 2.63 ;
      RECT 44.79 2.105 45.08 2.335 ;
      RECT 44.435 3.79 44.755 4.05 ;
      RECT 43.77 3.805 44.06 4.035 ;
      RECT 41.56 3.805 41.85 4.035 ;
      RECT 41.56 3.85 44.755 3.99 ;
      RECT 42.735 5.83 43.055 6.09 ;
      RECT 44.45 5.845 44.74 6.075 ;
      RECT 42.07 5.845 42.36 6.075 ;
      RECT 42.07 5.89 43.055 6.03 ;
      RECT 44.525 5.55 44.665 6.075 ;
      RECT 42.825 5.55 42.965 6.09 ;
      RECT 42.825 5.55 44.665 5.69 ;
      RECT 41.73 2.445 42.02 2.675 ;
      RECT 41.805 2.15 41.945 2.675 ;
      RECT 44.095 2.09 44.415 2.35 ;
      RECT 43.995 2.105 44.415 2.335 ;
      RECT 41.805 2.15 44.415 2.29 ;
      RECT 43.075 2.43 43.395 2.69 ;
      RECT 43.075 2.49 43.67 2.63 ;
      RECT 43.075 4.81 43.395 5.07 ;
      RECT 40.37 4.825 40.66 5.055 ;
      RECT 40.37 4.87 43.395 5.01 ;
      RECT 42.4 2.39 42.73 2.72 ;
      RECT 42.395 2.425 42.73 2.685 ;
      RECT 42.745 2.445 42.86 2.675 ;
      RECT 42.395 2.44 42.745 2.67 ;
      RECT 42.395 2.49 42.875 2.63 ;
      RECT 42.28 2.49 42.29 2.63 ;
      RECT 42.29 2.485 42.86 2.625 ;
      RECT 38.835 5.89 39.175 6.17 ;
      RECT 36.555 5.915 36.845 6.145 ;
      RECT 36.555 5.945 39.175 6.115 ;
      RECT 38.385 6.63 38.725 6.91 ;
      RECT 38.355 6.655 38.725 6.885 ;
      RECT 38.185 6.685 38.725 6.855 ;
      RECT 37.925 7.765 38.215 7.995 ;
      RECT 37.985 6.995 38.155 7.995 ;
      RECT 37.885 6.995 38.255 7.365 ;
      RECT 35.35 7.765 35.64 7.995 ;
      RECT 35.41 6.285 35.58 7.995 ;
      RECT 35.41 6.655 35.735 6.98 ;
      RECT 35.35 6.285 35.64 6.515 ;
      RECT 35.35 2.365 35.64 2.595 ;
      RECT 35.41 0.885 35.58 2.595 ;
      RECT 35.35 0.885 35.64 1.115 ;
      RECT 34.94 2.735 35.27 2.965 ;
      RECT 34.94 2.765 35.44 2.935 ;
      RECT 34.94 2.395 35.13 2.965 ;
      RECT 34.36 2.365 34.65 2.595 ;
      RECT 34.36 2.395 35.13 2.565 ;
      RECT 34.42 0.885 34.59 2.595 ;
      RECT 34.36 0.885 34.65 1.115 ;
      RECT 34.36 7.765 34.65 7.995 ;
      RECT 34.42 6.285 34.59 7.995 ;
      RECT 34.36 6.285 34.65 6.515 ;
      RECT 34.36 6.325 35.21 6.485 ;
      RECT 35.04 5.915 35.21 6.485 ;
      RECT 34.36 6.32 34.75 6.485 ;
      RECT 34.98 5.915 35.27 6.145 ;
      RECT 34.98 5.945 35.44 6.115 ;
      RECT 33.99 2.735 34.28 2.965 ;
      RECT 33.99 2.765 34.45 2.935 ;
      RECT 34.05 1.655 34.215 2.965 ;
      RECT 32.565 1.625 32.855 1.855 ;
      RECT 32.565 1.655 34.215 1.825 ;
      RECT 32.625 0.885 32.795 1.855 ;
      RECT 32.565 0.885 32.855 1.115 ;
      RECT 32.565 7.765 32.855 7.995 ;
      RECT 32.625 7.025 32.795 7.995 ;
      RECT 32.625 7.12 34.215 7.29 ;
      RECT 34.045 5.915 34.215 7.29 ;
      RECT 32.565 7.025 32.855 7.255 ;
      RECT 33.99 5.915 34.28 6.145 ;
      RECT 33.99 5.945 34.45 6.115 ;
      RECT 30.55 1.995 30.875 2.32 ;
      RECT 32.995 1.965 33.345 2.315 ;
      RECT 30.55 2.025 33.345 2.195 ;
      RECT 33.02 6.655 33.345 6.98 ;
      RECT 32.995 6.655 33.345 6.885 ;
      RECT 32.825 6.685 33.345 6.855 ;
      RECT 32.22 2.365 32.54 2.685 ;
      RECT 32.19 2.365 32.54 2.595 ;
      RECT 31.905 2.395 32.54 2.565 ;
      RECT 32.22 6.28 32.54 6.605 ;
      RECT 32.19 6.285 32.54 6.515 ;
      RECT 32.02 6.315 32.54 6.485 ;
      RECT 31.175 3.635 31.5 3.96 ;
      RECT 31.25 2.735 31.43 3.96 ;
      RECT 31.195 2.735 31.485 2.965 ;
      RECT 31.195 2.765 31.655 2.935 ;
      RECT 31.18 5.865 31.505 6.19 ;
      RECT 31.18 5.945 31.655 6.115 ;
      RECT 29.965 3.185 30.29 3.51 ;
      RECT 27.17 3.11 27.49 3.37 ;
      RECT 29.145 3.125 29.435 3.355 ;
      RECT 29.865 3.185 30.29 3.325 ;
      RECT 27.17 3.17 30.005 3.31 ;
      RECT 29.55 2.77 29.87 3.03 ;
      RECT 29.275 2.83 29.87 2.97 ;
      RECT 28.53 5.83 28.85 6.09 ;
      RECT 28.53 5.89 29.125 6.03 ;
      RECT 27.85 2.77 28.17 3.03 ;
      RECT 23.11 2.785 23.4 3.015 ;
      RECT 23.11 2.83 28.17 2.97 ;
      RECT 27.94 2.49 28.08 3.03 ;
      RECT 27.94 2.49 28.42 2.63 ;
      RECT 28.28 2.105 28.42 2.63 ;
      RECT 28.205 2.105 28.495 2.335 ;
      RECT 27.85 3.79 28.17 4.05 ;
      RECT 27.185 3.805 27.475 4.035 ;
      RECT 24.975 3.805 25.265 4.035 ;
      RECT 24.975 3.85 28.17 3.99 ;
      RECT 26.15 5.83 26.47 6.09 ;
      RECT 27.865 5.845 28.155 6.075 ;
      RECT 25.485 5.845 25.775 6.075 ;
      RECT 25.485 5.89 26.47 6.03 ;
      RECT 27.94 5.55 28.08 6.075 ;
      RECT 26.24 5.55 26.38 6.09 ;
      RECT 26.24 5.55 28.08 5.69 ;
      RECT 25.145 2.445 25.435 2.675 ;
      RECT 25.22 2.15 25.36 2.675 ;
      RECT 27.51 2.09 27.83 2.35 ;
      RECT 27.41 2.105 27.83 2.335 ;
      RECT 25.22 2.15 27.83 2.29 ;
      RECT 26.49 2.43 26.81 2.69 ;
      RECT 26.49 2.49 27.085 2.63 ;
      RECT 26.49 4.81 26.81 5.07 ;
      RECT 23.785 4.825 24.075 5.055 ;
      RECT 23.785 4.87 26.81 5.01 ;
      RECT 25.815 2.39 26.145 2.72 ;
      RECT 25.81 2.425 26.145 2.685 ;
      RECT 26.16 2.445 26.275 2.675 ;
      RECT 25.81 2.44 26.16 2.67 ;
      RECT 25.81 2.49 26.29 2.63 ;
      RECT 25.695 2.49 25.705 2.63 ;
      RECT 25.705 2.485 26.275 2.625 ;
      RECT 22.25 5.89 22.59 6.17 ;
      RECT 19.97 5.915 20.26 6.145 ;
      RECT 19.97 5.945 22.59 6.115 ;
      RECT 21.8 6.63 22.14 6.91 ;
      RECT 21.77 6.655 22.14 6.885 ;
      RECT 21.6 6.685 22.14 6.855 ;
      RECT 21.34 7.765 21.63 7.995 ;
      RECT 21.4 6.995 21.57 7.995 ;
      RECT 21.3 6.995 21.67 7.365 ;
      RECT 18.765 7.765 19.055 7.995 ;
      RECT 18.825 6.285 18.995 7.995 ;
      RECT 18.825 6.655 19.15 6.98 ;
      RECT 18.765 6.285 19.055 6.515 ;
      RECT 18.765 2.365 19.055 2.595 ;
      RECT 18.825 0.885 18.995 2.595 ;
      RECT 18.765 0.885 19.055 1.115 ;
      RECT 18.355 2.735 18.685 2.965 ;
      RECT 18.355 2.765 18.855 2.935 ;
      RECT 18.355 2.395 18.545 2.965 ;
      RECT 17.775 2.365 18.065 2.595 ;
      RECT 17.775 2.395 18.545 2.565 ;
      RECT 17.835 0.885 18.005 2.595 ;
      RECT 17.775 0.885 18.065 1.115 ;
      RECT 17.775 7.765 18.065 7.995 ;
      RECT 17.835 6.285 18.005 7.995 ;
      RECT 17.775 6.285 18.065 6.515 ;
      RECT 17.775 6.325 18.625 6.485 ;
      RECT 18.455 5.915 18.625 6.485 ;
      RECT 17.775 6.32 18.165 6.485 ;
      RECT 18.395 5.915 18.685 6.145 ;
      RECT 18.395 5.945 18.855 6.115 ;
      RECT 17.405 2.735 17.695 2.965 ;
      RECT 17.405 2.765 17.865 2.935 ;
      RECT 17.465 1.655 17.63 2.965 ;
      RECT 15.98 1.625 16.27 1.855 ;
      RECT 15.98 1.655 17.63 1.825 ;
      RECT 16.04 0.885 16.21 1.855 ;
      RECT 15.98 0.885 16.27 1.115 ;
      RECT 15.98 7.765 16.27 7.995 ;
      RECT 16.04 7.025 16.21 7.995 ;
      RECT 16.04 7.12 17.63 7.29 ;
      RECT 17.46 5.915 17.63 7.29 ;
      RECT 15.98 7.025 16.27 7.255 ;
      RECT 17.405 5.915 17.695 6.145 ;
      RECT 17.405 5.945 17.865 6.115 ;
      RECT 13.965 1.995 14.29 2.32 ;
      RECT 16.41 1.965 16.76 2.315 ;
      RECT 13.965 2.025 16.76 2.195 ;
      RECT 16.435 6.655 16.76 6.98 ;
      RECT 16.41 6.655 16.76 6.885 ;
      RECT 16.24 6.685 16.76 6.855 ;
      RECT 15.635 2.365 15.955 2.685 ;
      RECT 15.605 2.365 15.955 2.595 ;
      RECT 15.32 2.395 15.955 2.565 ;
      RECT 15.635 6.28 15.955 6.605 ;
      RECT 15.605 6.285 15.955 6.515 ;
      RECT 15.435 6.315 15.955 6.485 ;
      RECT 14.59 3.635 14.915 3.96 ;
      RECT 14.665 2.735 14.845 3.96 ;
      RECT 14.61 2.735 14.9 2.965 ;
      RECT 14.61 2.765 15.07 2.935 ;
      RECT 14.595 5.865 14.92 6.19 ;
      RECT 14.595 5.945 15.07 6.115 ;
      RECT 13.38 3.185 13.705 3.51 ;
      RECT 10.585 3.11 10.905 3.37 ;
      RECT 12.56 3.125 12.85 3.355 ;
      RECT 13.28 3.185 13.705 3.325 ;
      RECT 10.585 3.17 13.42 3.31 ;
      RECT 12.965 2.77 13.285 3.03 ;
      RECT 12.69 2.83 13.285 2.97 ;
      RECT 11.945 5.83 12.265 6.09 ;
      RECT 11.945 5.89 12.54 6.03 ;
      RECT 11.265 2.77 11.585 3.03 ;
      RECT 6.525 2.785 6.815 3.015 ;
      RECT 6.525 2.83 11.585 2.97 ;
      RECT 11.355 2.49 11.495 3.03 ;
      RECT 11.355 2.49 11.835 2.63 ;
      RECT 11.695 2.105 11.835 2.63 ;
      RECT 11.62 2.105 11.91 2.335 ;
      RECT 11.265 3.79 11.585 4.05 ;
      RECT 10.6 3.805 10.89 4.035 ;
      RECT 8.39 3.805 8.68 4.035 ;
      RECT 8.39 3.85 11.585 3.99 ;
      RECT 9.565 5.83 9.885 6.09 ;
      RECT 11.28 5.845 11.57 6.075 ;
      RECT 8.9 5.845 9.19 6.075 ;
      RECT 8.9 5.89 9.885 6.03 ;
      RECT 11.355 5.55 11.495 6.075 ;
      RECT 9.655 5.55 9.795 6.09 ;
      RECT 9.655 5.55 11.495 5.69 ;
      RECT 8.56 2.445 8.85 2.675 ;
      RECT 8.635 2.15 8.775 2.675 ;
      RECT 10.925 2.09 11.245 2.35 ;
      RECT 10.825 2.105 11.245 2.335 ;
      RECT 8.635 2.15 11.245 2.29 ;
      RECT 9.905 2.43 10.225 2.69 ;
      RECT 9.905 2.49 10.5 2.63 ;
      RECT 9.905 4.81 10.225 5.07 ;
      RECT 7.2 4.825 7.49 5.055 ;
      RECT 7.2 4.87 10.225 5.01 ;
      RECT 9.23 2.39 9.56 2.72 ;
      RECT 9.225 2.425 9.56 2.685 ;
      RECT 9.575 2.445 9.69 2.675 ;
      RECT 9.225 2.44 9.575 2.67 ;
      RECT 9.225 2.49 9.705 2.63 ;
      RECT 9.11 2.49 9.12 2.63 ;
      RECT 9.12 2.485 9.69 2.625 ;
      RECT 5.665 5.89 6.005 6.17 ;
      RECT 3.385 5.915 3.675 6.145 ;
      RECT 3.385 5.945 6.005 6.115 ;
      RECT 5.215 6.63 5.555 6.91 ;
      RECT 5.185 6.655 5.555 6.885 ;
      RECT 5.015 6.685 5.555 6.855 ;
      RECT 4.755 7.765 5.045 7.995 ;
      RECT 4.815 6.995 4.985 7.995 ;
      RECT 4.715 6.995 5.085 7.365 ;
      RECT 1.955 6.655 2.245 6.885 ;
      RECT 1.785 6.685 2.245 6.855 ;
      RECT 1.525 7.765 1.815 7.995 ;
      RECT 1.585 7.025 1.755 7.995 ;
      RECT 1.495 7.025 1.835 7.305 ;
      RECT 1.12 6.285 1.46 6.565 ;
      RECT 0.98 6.315 1.46 6.485 ;
      RECT 0.155 5.915 0.445 6.145 ;
      RECT 0.155 5.945 0.615 6.115 ;
      RECT 78.975 4.81 79.62 5.07 ;
      RECT 76.92 5.83 77.24 6.09 ;
      RECT 62.395 4.81 63.04 5.07 ;
      RECT 60.34 5.83 60.66 6.09 ;
      RECT 45.81 4.81 46.455 5.07 ;
      RECT 43.755 5.83 44.075 6.09 ;
      RECT 29.225 4.81 29.87 5.07 ;
      RECT 27.17 5.83 27.49 6.09 ;
      RECT 12.64 4.81 13.285 5.07 ;
      RECT 10.585 5.83 10.905 6.09 ;
    LAYER mcon ;
      RECT 85.16 0.915 85.33 1.085 ;
      RECT 85.16 2.395 85.33 2.565 ;
      RECT 85.16 6.315 85.33 6.485 ;
      RECT 85.16 7.795 85.33 7.965 ;
      RECT 84.81 0.105 84.98 0.275 ;
      RECT 84.81 4.165 84.98 4.335 ;
      RECT 84.81 4.545 84.98 4.715 ;
      RECT 84.81 8.605 84.98 8.775 ;
      RECT 84.79 2.765 84.96 2.935 ;
      RECT 84.79 5.945 84.96 6.115 ;
      RECT 84.17 0.915 84.34 1.085 ;
      RECT 84.17 2.395 84.34 2.565 ;
      RECT 84.17 6.315 84.34 6.485 ;
      RECT 84.17 7.795 84.34 7.965 ;
      RECT 83.82 0.105 83.99 0.275 ;
      RECT 83.82 4.165 83.99 4.335 ;
      RECT 83.82 4.545 83.99 4.715 ;
      RECT 83.82 8.605 83.99 8.775 ;
      RECT 83.8 2.765 83.97 2.935 ;
      RECT 83.8 5.945 83.97 6.115 ;
      RECT 83.115 0.105 83.285 0.275 ;
      RECT 83.115 4.165 83.285 4.335 ;
      RECT 83.115 4.545 83.285 4.715 ;
      RECT 83.115 8.605 83.285 8.775 ;
      RECT 82.805 2.025 82.975 2.195 ;
      RECT 82.805 6.685 82.975 6.855 ;
      RECT 82.435 0.105 82.605 0.275 ;
      RECT 82.435 8.605 82.605 8.775 ;
      RECT 82.375 0.915 82.545 1.085 ;
      RECT 82.375 1.655 82.545 1.825 ;
      RECT 82.375 7.055 82.545 7.225 ;
      RECT 82.375 7.795 82.545 7.965 ;
      RECT 82 2.395 82.17 2.565 ;
      RECT 82 6.315 82.17 6.485 ;
      RECT 81.755 0.105 81.925 0.275 ;
      RECT 81.755 8.605 81.925 8.775 ;
      RECT 81.075 0.105 81.245 0.275 ;
      RECT 81.075 8.605 81.245 8.775 ;
      RECT 81.005 2.765 81.175 2.935 ;
      RECT 81.005 5.945 81.175 6.115 ;
      RECT 79.415 1.625 79.585 1.795 ;
      RECT 79.415 4.345 79.585 4.515 ;
      RECT 79.415 7.065 79.585 7.235 ;
      RECT 79.375 2.815 79.545 2.985 ;
      RECT 79.035 4.855 79.205 5.025 ;
      RECT 78.955 1.625 79.125 1.795 ;
      RECT 78.955 3.155 79.125 3.325 ;
      RECT 78.955 4.345 79.125 4.515 ;
      RECT 78.955 7.065 79.125 7.235 ;
      RECT 78.495 1.625 78.665 1.795 ;
      RECT 78.495 4.345 78.665 4.515 ;
      RECT 78.495 7.065 78.665 7.235 ;
      RECT 78.355 5.875 78.525 6.045 ;
      RECT 78.035 1.625 78.205 1.795 ;
      RECT 78.035 4.345 78.205 4.515 ;
      RECT 78.035 7.065 78.205 7.235 ;
      RECT 78.015 2.135 78.185 2.305 ;
      RECT 77.675 5.875 77.845 6.045 ;
      RECT 77.575 1.625 77.745 1.795 ;
      RECT 77.575 4.345 77.745 4.515 ;
      RECT 77.575 7.065 77.745 7.235 ;
      RECT 77.22 2.135 77.39 2.305 ;
      RECT 77.115 1.625 77.285 1.795 ;
      RECT 77.115 4.345 77.285 4.515 ;
      RECT 77.115 7.065 77.285 7.235 ;
      RECT 76.995 3.835 77.165 4.005 ;
      RECT 76.995 5.875 77.165 6.045 ;
      RECT 76.655 1.625 76.825 1.795 ;
      RECT 76.655 4.345 76.825 4.515 ;
      RECT 76.655 7.065 76.825 7.235 ;
      RECT 76.485 5.875 76.655 6.045 ;
      RECT 76.315 2.475 76.485 2.645 ;
      RECT 76.195 1.625 76.365 1.795 ;
      RECT 76.195 4.345 76.365 4.515 ;
      RECT 76.195 7.065 76.365 7.235 ;
      RECT 75.735 1.625 75.905 1.795 ;
      RECT 75.735 4.345 75.905 4.515 ;
      RECT 75.735 7.065 75.905 7.235 ;
      RECT 75.295 5.875 75.465 6.045 ;
      RECT 75.275 1.625 75.445 1.795 ;
      RECT 75.275 4.345 75.445 4.515 ;
      RECT 75.275 7.065 75.445 7.235 ;
      RECT 74.955 2.475 75.125 2.645 ;
      RECT 74.815 1.625 74.985 1.795 ;
      RECT 74.815 4.345 74.985 4.515 ;
      RECT 74.815 7.065 74.985 7.235 ;
      RECT 74.785 3.835 74.955 4.005 ;
      RECT 74.355 1.625 74.525 1.795 ;
      RECT 74.355 4.345 74.525 4.515 ;
      RECT 74.355 7.065 74.525 7.235 ;
      RECT 74.275 5.875 74.445 6.045 ;
      RECT 73.895 1.625 74.065 1.795 ;
      RECT 73.895 4.345 74.065 4.515 ;
      RECT 73.895 7.065 74.065 7.235 ;
      RECT 73.595 4.855 73.765 5.025 ;
      RECT 73.435 1.625 73.605 1.795 ;
      RECT 73.435 4.345 73.605 4.515 ;
      RECT 73.435 7.065 73.605 7.235 ;
      RECT 72.975 1.625 73.145 1.795 ;
      RECT 72.975 4.345 73.145 4.515 ;
      RECT 72.975 7.065 73.145 7.235 ;
      RECT 72.92 2.815 73.09 2.985 ;
      RECT 71.89 4.545 72.06 4.715 ;
      RECT 71.89 8.605 72.06 8.775 ;
      RECT 71.58 6.685 71.75 6.855 ;
      RECT 71.21 8.605 71.38 8.775 ;
      RECT 71.15 7.055 71.32 7.225 ;
      RECT 71.15 7.795 71.32 7.965 ;
      RECT 70.775 6.315 70.945 6.485 ;
      RECT 70.53 8.605 70.7 8.775 ;
      RECT 69.85 8.605 70.02 8.775 ;
      RECT 69.78 5.945 69.95 6.115 ;
      RECT 68.58 0.915 68.75 1.085 ;
      RECT 68.58 2.395 68.75 2.565 ;
      RECT 68.58 6.315 68.75 6.485 ;
      RECT 68.58 7.795 68.75 7.965 ;
      RECT 68.23 0.105 68.4 0.275 ;
      RECT 68.23 4.165 68.4 4.335 ;
      RECT 68.23 4.545 68.4 4.715 ;
      RECT 68.23 8.605 68.4 8.775 ;
      RECT 68.21 2.765 68.38 2.935 ;
      RECT 68.21 5.945 68.38 6.115 ;
      RECT 67.59 0.915 67.76 1.085 ;
      RECT 67.59 2.395 67.76 2.565 ;
      RECT 67.59 6.315 67.76 6.485 ;
      RECT 67.59 7.795 67.76 7.965 ;
      RECT 67.24 0.105 67.41 0.275 ;
      RECT 67.24 4.165 67.41 4.335 ;
      RECT 67.24 4.545 67.41 4.715 ;
      RECT 67.24 8.605 67.41 8.775 ;
      RECT 67.22 2.765 67.39 2.935 ;
      RECT 67.22 5.945 67.39 6.115 ;
      RECT 66.535 0.105 66.705 0.275 ;
      RECT 66.535 4.165 66.705 4.335 ;
      RECT 66.535 4.545 66.705 4.715 ;
      RECT 66.535 8.605 66.705 8.775 ;
      RECT 66.225 2.025 66.395 2.195 ;
      RECT 66.225 6.685 66.395 6.855 ;
      RECT 65.855 0.105 66.025 0.275 ;
      RECT 65.855 8.605 66.025 8.775 ;
      RECT 65.795 0.915 65.965 1.085 ;
      RECT 65.795 1.655 65.965 1.825 ;
      RECT 65.795 7.055 65.965 7.225 ;
      RECT 65.795 7.795 65.965 7.965 ;
      RECT 65.42 2.395 65.59 2.565 ;
      RECT 65.42 6.315 65.59 6.485 ;
      RECT 65.175 0.105 65.345 0.275 ;
      RECT 65.175 8.605 65.345 8.775 ;
      RECT 64.495 0.105 64.665 0.275 ;
      RECT 64.495 8.605 64.665 8.775 ;
      RECT 64.425 2.765 64.595 2.935 ;
      RECT 64.425 5.945 64.595 6.115 ;
      RECT 62.835 1.625 63.005 1.795 ;
      RECT 62.835 4.345 63.005 4.515 ;
      RECT 62.835 7.065 63.005 7.235 ;
      RECT 62.795 2.815 62.965 2.985 ;
      RECT 62.455 4.855 62.625 5.025 ;
      RECT 62.375 1.625 62.545 1.795 ;
      RECT 62.375 3.155 62.545 3.325 ;
      RECT 62.375 4.345 62.545 4.515 ;
      RECT 62.375 7.065 62.545 7.235 ;
      RECT 61.915 1.625 62.085 1.795 ;
      RECT 61.915 4.345 62.085 4.515 ;
      RECT 61.915 7.065 62.085 7.235 ;
      RECT 61.775 5.875 61.945 6.045 ;
      RECT 61.455 1.625 61.625 1.795 ;
      RECT 61.455 4.345 61.625 4.515 ;
      RECT 61.455 7.065 61.625 7.235 ;
      RECT 61.435 2.135 61.605 2.305 ;
      RECT 61.095 5.875 61.265 6.045 ;
      RECT 60.995 1.625 61.165 1.795 ;
      RECT 60.995 4.345 61.165 4.515 ;
      RECT 60.995 7.065 61.165 7.235 ;
      RECT 60.64 2.135 60.81 2.305 ;
      RECT 60.535 1.625 60.705 1.795 ;
      RECT 60.535 4.345 60.705 4.515 ;
      RECT 60.535 7.065 60.705 7.235 ;
      RECT 60.415 3.835 60.585 4.005 ;
      RECT 60.415 5.875 60.585 6.045 ;
      RECT 60.075 1.625 60.245 1.795 ;
      RECT 60.075 4.345 60.245 4.515 ;
      RECT 60.075 7.065 60.245 7.235 ;
      RECT 59.905 5.875 60.075 6.045 ;
      RECT 59.735 2.475 59.905 2.645 ;
      RECT 59.615 1.625 59.785 1.795 ;
      RECT 59.615 4.345 59.785 4.515 ;
      RECT 59.615 7.065 59.785 7.235 ;
      RECT 59.155 1.625 59.325 1.795 ;
      RECT 59.155 4.345 59.325 4.515 ;
      RECT 59.155 7.065 59.325 7.235 ;
      RECT 58.715 5.875 58.885 6.045 ;
      RECT 58.695 1.625 58.865 1.795 ;
      RECT 58.695 4.345 58.865 4.515 ;
      RECT 58.695 7.065 58.865 7.235 ;
      RECT 58.375 2.475 58.545 2.645 ;
      RECT 58.235 1.625 58.405 1.795 ;
      RECT 58.235 4.345 58.405 4.515 ;
      RECT 58.235 7.065 58.405 7.235 ;
      RECT 58.205 3.835 58.375 4.005 ;
      RECT 57.775 1.625 57.945 1.795 ;
      RECT 57.775 4.345 57.945 4.515 ;
      RECT 57.775 7.065 57.945 7.235 ;
      RECT 57.695 5.875 57.865 6.045 ;
      RECT 57.315 1.625 57.485 1.795 ;
      RECT 57.315 4.345 57.485 4.515 ;
      RECT 57.315 7.065 57.485 7.235 ;
      RECT 57.015 4.855 57.185 5.025 ;
      RECT 56.855 1.625 57.025 1.795 ;
      RECT 56.855 4.345 57.025 4.515 ;
      RECT 56.855 7.065 57.025 7.235 ;
      RECT 56.395 1.625 56.565 1.795 ;
      RECT 56.395 4.345 56.565 4.515 ;
      RECT 56.395 7.065 56.565 7.235 ;
      RECT 56.34 2.815 56.51 2.985 ;
      RECT 55.31 4.545 55.48 4.715 ;
      RECT 55.31 8.605 55.48 8.775 ;
      RECT 55 6.685 55.17 6.855 ;
      RECT 54.63 8.605 54.8 8.775 ;
      RECT 54.57 7.055 54.74 7.225 ;
      RECT 54.57 7.795 54.74 7.965 ;
      RECT 54.195 6.315 54.365 6.485 ;
      RECT 53.95 8.605 54.12 8.775 ;
      RECT 53.27 8.605 53.44 8.775 ;
      RECT 53.2 5.945 53.37 6.115 ;
      RECT 51.995 0.915 52.165 1.085 ;
      RECT 51.995 2.395 52.165 2.565 ;
      RECT 51.995 6.315 52.165 6.485 ;
      RECT 51.995 7.795 52.165 7.965 ;
      RECT 51.645 0.105 51.815 0.275 ;
      RECT 51.645 4.165 51.815 4.335 ;
      RECT 51.645 4.545 51.815 4.715 ;
      RECT 51.645 8.605 51.815 8.775 ;
      RECT 51.625 2.765 51.795 2.935 ;
      RECT 51.625 5.945 51.795 6.115 ;
      RECT 51.005 0.915 51.175 1.085 ;
      RECT 51.005 2.395 51.175 2.565 ;
      RECT 51.005 6.315 51.175 6.485 ;
      RECT 51.005 7.795 51.175 7.965 ;
      RECT 50.655 0.105 50.825 0.275 ;
      RECT 50.655 4.165 50.825 4.335 ;
      RECT 50.655 4.545 50.825 4.715 ;
      RECT 50.655 8.605 50.825 8.775 ;
      RECT 50.635 2.765 50.805 2.935 ;
      RECT 50.635 5.945 50.805 6.115 ;
      RECT 49.95 0.105 50.12 0.275 ;
      RECT 49.95 4.165 50.12 4.335 ;
      RECT 49.95 4.545 50.12 4.715 ;
      RECT 49.95 8.605 50.12 8.775 ;
      RECT 49.64 2.025 49.81 2.195 ;
      RECT 49.64 6.685 49.81 6.855 ;
      RECT 49.27 0.105 49.44 0.275 ;
      RECT 49.27 8.605 49.44 8.775 ;
      RECT 49.21 0.915 49.38 1.085 ;
      RECT 49.21 1.655 49.38 1.825 ;
      RECT 49.21 7.055 49.38 7.225 ;
      RECT 49.21 7.795 49.38 7.965 ;
      RECT 48.835 2.395 49.005 2.565 ;
      RECT 48.835 6.315 49.005 6.485 ;
      RECT 48.59 0.105 48.76 0.275 ;
      RECT 48.59 8.605 48.76 8.775 ;
      RECT 47.91 0.105 48.08 0.275 ;
      RECT 47.91 8.605 48.08 8.775 ;
      RECT 47.84 2.765 48.01 2.935 ;
      RECT 47.84 5.945 48.01 6.115 ;
      RECT 46.25 1.625 46.42 1.795 ;
      RECT 46.25 4.345 46.42 4.515 ;
      RECT 46.25 7.065 46.42 7.235 ;
      RECT 46.21 2.815 46.38 2.985 ;
      RECT 45.87 4.855 46.04 5.025 ;
      RECT 45.79 1.625 45.96 1.795 ;
      RECT 45.79 3.155 45.96 3.325 ;
      RECT 45.79 4.345 45.96 4.515 ;
      RECT 45.79 7.065 45.96 7.235 ;
      RECT 45.33 1.625 45.5 1.795 ;
      RECT 45.33 4.345 45.5 4.515 ;
      RECT 45.33 7.065 45.5 7.235 ;
      RECT 45.19 5.875 45.36 6.045 ;
      RECT 44.87 1.625 45.04 1.795 ;
      RECT 44.87 4.345 45.04 4.515 ;
      RECT 44.87 7.065 45.04 7.235 ;
      RECT 44.85 2.135 45.02 2.305 ;
      RECT 44.51 5.875 44.68 6.045 ;
      RECT 44.41 1.625 44.58 1.795 ;
      RECT 44.41 4.345 44.58 4.515 ;
      RECT 44.41 7.065 44.58 7.235 ;
      RECT 44.055 2.135 44.225 2.305 ;
      RECT 43.95 1.625 44.12 1.795 ;
      RECT 43.95 4.345 44.12 4.515 ;
      RECT 43.95 7.065 44.12 7.235 ;
      RECT 43.83 3.835 44 4.005 ;
      RECT 43.83 5.875 44 6.045 ;
      RECT 43.49 1.625 43.66 1.795 ;
      RECT 43.49 4.345 43.66 4.515 ;
      RECT 43.49 7.065 43.66 7.235 ;
      RECT 43.32 5.875 43.49 6.045 ;
      RECT 43.15 2.475 43.32 2.645 ;
      RECT 43.03 1.625 43.2 1.795 ;
      RECT 43.03 4.345 43.2 4.515 ;
      RECT 43.03 7.065 43.2 7.235 ;
      RECT 42.57 1.625 42.74 1.795 ;
      RECT 42.57 4.345 42.74 4.515 ;
      RECT 42.57 7.065 42.74 7.235 ;
      RECT 42.13 5.875 42.3 6.045 ;
      RECT 42.11 1.625 42.28 1.795 ;
      RECT 42.11 4.345 42.28 4.515 ;
      RECT 42.11 7.065 42.28 7.235 ;
      RECT 41.79 2.475 41.96 2.645 ;
      RECT 41.65 1.625 41.82 1.795 ;
      RECT 41.65 4.345 41.82 4.515 ;
      RECT 41.65 7.065 41.82 7.235 ;
      RECT 41.62 3.835 41.79 4.005 ;
      RECT 41.19 1.625 41.36 1.795 ;
      RECT 41.19 4.345 41.36 4.515 ;
      RECT 41.19 7.065 41.36 7.235 ;
      RECT 41.11 5.875 41.28 6.045 ;
      RECT 40.73 1.625 40.9 1.795 ;
      RECT 40.73 4.345 40.9 4.515 ;
      RECT 40.73 7.065 40.9 7.235 ;
      RECT 40.43 4.855 40.6 5.025 ;
      RECT 40.27 1.625 40.44 1.795 ;
      RECT 40.27 4.345 40.44 4.515 ;
      RECT 40.27 7.065 40.44 7.235 ;
      RECT 39.81 1.625 39.98 1.795 ;
      RECT 39.81 4.345 39.98 4.515 ;
      RECT 39.81 7.065 39.98 7.235 ;
      RECT 39.755 2.815 39.925 2.985 ;
      RECT 38.725 4.545 38.895 4.715 ;
      RECT 38.725 8.605 38.895 8.775 ;
      RECT 38.415 6.685 38.585 6.855 ;
      RECT 38.045 8.605 38.215 8.775 ;
      RECT 37.985 7.055 38.155 7.225 ;
      RECT 37.985 7.795 38.155 7.965 ;
      RECT 37.61 6.315 37.78 6.485 ;
      RECT 37.365 8.605 37.535 8.775 ;
      RECT 36.685 8.605 36.855 8.775 ;
      RECT 36.615 5.945 36.785 6.115 ;
      RECT 35.41 0.915 35.58 1.085 ;
      RECT 35.41 2.395 35.58 2.565 ;
      RECT 35.41 6.315 35.58 6.485 ;
      RECT 35.41 7.795 35.58 7.965 ;
      RECT 35.06 0.105 35.23 0.275 ;
      RECT 35.06 4.165 35.23 4.335 ;
      RECT 35.06 4.545 35.23 4.715 ;
      RECT 35.06 8.605 35.23 8.775 ;
      RECT 35.04 2.765 35.21 2.935 ;
      RECT 35.04 5.945 35.21 6.115 ;
      RECT 34.42 0.915 34.59 1.085 ;
      RECT 34.42 2.395 34.59 2.565 ;
      RECT 34.42 6.315 34.59 6.485 ;
      RECT 34.42 7.795 34.59 7.965 ;
      RECT 34.07 0.105 34.24 0.275 ;
      RECT 34.07 4.165 34.24 4.335 ;
      RECT 34.07 4.545 34.24 4.715 ;
      RECT 34.07 8.605 34.24 8.775 ;
      RECT 34.05 2.765 34.22 2.935 ;
      RECT 34.05 5.945 34.22 6.115 ;
      RECT 33.365 0.105 33.535 0.275 ;
      RECT 33.365 4.165 33.535 4.335 ;
      RECT 33.365 4.545 33.535 4.715 ;
      RECT 33.365 8.605 33.535 8.775 ;
      RECT 33.055 2.025 33.225 2.195 ;
      RECT 33.055 6.685 33.225 6.855 ;
      RECT 32.685 0.105 32.855 0.275 ;
      RECT 32.685 8.605 32.855 8.775 ;
      RECT 32.625 0.915 32.795 1.085 ;
      RECT 32.625 1.655 32.795 1.825 ;
      RECT 32.625 7.055 32.795 7.225 ;
      RECT 32.625 7.795 32.795 7.965 ;
      RECT 32.25 2.395 32.42 2.565 ;
      RECT 32.25 6.315 32.42 6.485 ;
      RECT 32.005 0.105 32.175 0.275 ;
      RECT 32.005 8.605 32.175 8.775 ;
      RECT 31.325 0.105 31.495 0.275 ;
      RECT 31.325 8.605 31.495 8.775 ;
      RECT 31.255 2.765 31.425 2.935 ;
      RECT 31.255 5.945 31.425 6.115 ;
      RECT 29.665 1.625 29.835 1.795 ;
      RECT 29.665 4.345 29.835 4.515 ;
      RECT 29.665 7.065 29.835 7.235 ;
      RECT 29.625 2.815 29.795 2.985 ;
      RECT 29.285 4.855 29.455 5.025 ;
      RECT 29.205 1.625 29.375 1.795 ;
      RECT 29.205 3.155 29.375 3.325 ;
      RECT 29.205 4.345 29.375 4.515 ;
      RECT 29.205 7.065 29.375 7.235 ;
      RECT 28.745 1.625 28.915 1.795 ;
      RECT 28.745 4.345 28.915 4.515 ;
      RECT 28.745 7.065 28.915 7.235 ;
      RECT 28.605 5.875 28.775 6.045 ;
      RECT 28.285 1.625 28.455 1.795 ;
      RECT 28.285 4.345 28.455 4.515 ;
      RECT 28.285 7.065 28.455 7.235 ;
      RECT 28.265 2.135 28.435 2.305 ;
      RECT 27.925 5.875 28.095 6.045 ;
      RECT 27.825 1.625 27.995 1.795 ;
      RECT 27.825 4.345 27.995 4.515 ;
      RECT 27.825 7.065 27.995 7.235 ;
      RECT 27.47 2.135 27.64 2.305 ;
      RECT 27.365 1.625 27.535 1.795 ;
      RECT 27.365 4.345 27.535 4.515 ;
      RECT 27.365 7.065 27.535 7.235 ;
      RECT 27.245 3.835 27.415 4.005 ;
      RECT 27.245 5.875 27.415 6.045 ;
      RECT 26.905 1.625 27.075 1.795 ;
      RECT 26.905 4.345 27.075 4.515 ;
      RECT 26.905 7.065 27.075 7.235 ;
      RECT 26.735 5.875 26.905 6.045 ;
      RECT 26.565 2.475 26.735 2.645 ;
      RECT 26.445 1.625 26.615 1.795 ;
      RECT 26.445 4.345 26.615 4.515 ;
      RECT 26.445 7.065 26.615 7.235 ;
      RECT 25.985 1.625 26.155 1.795 ;
      RECT 25.985 4.345 26.155 4.515 ;
      RECT 25.985 7.065 26.155 7.235 ;
      RECT 25.545 5.875 25.715 6.045 ;
      RECT 25.525 1.625 25.695 1.795 ;
      RECT 25.525 4.345 25.695 4.515 ;
      RECT 25.525 7.065 25.695 7.235 ;
      RECT 25.205 2.475 25.375 2.645 ;
      RECT 25.065 1.625 25.235 1.795 ;
      RECT 25.065 4.345 25.235 4.515 ;
      RECT 25.065 7.065 25.235 7.235 ;
      RECT 25.035 3.835 25.205 4.005 ;
      RECT 24.605 1.625 24.775 1.795 ;
      RECT 24.605 4.345 24.775 4.515 ;
      RECT 24.605 7.065 24.775 7.235 ;
      RECT 24.525 5.875 24.695 6.045 ;
      RECT 24.145 1.625 24.315 1.795 ;
      RECT 24.145 4.345 24.315 4.515 ;
      RECT 24.145 7.065 24.315 7.235 ;
      RECT 23.845 4.855 24.015 5.025 ;
      RECT 23.685 1.625 23.855 1.795 ;
      RECT 23.685 4.345 23.855 4.515 ;
      RECT 23.685 7.065 23.855 7.235 ;
      RECT 23.225 1.625 23.395 1.795 ;
      RECT 23.225 4.345 23.395 4.515 ;
      RECT 23.225 7.065 23.395 7.235 ;
      RECT 23.17 2.815 23.34 2.985 ;
      RECT 22.14 4.545 22.31 4.715 ;
      RECT 22.14 8.605 22.31 8.775 ;
      RECT 21.83 6.685 22 6.855 ;
      RECT 21.46 8.605 21.63 8.775 ;
      RECT 21.4 7.055 21.57 7.225 ;
      RECT 21.4 7.795 21.57 7.965 ;
      RECT 21.025 6.315 21.195 6.485 ;
      RECT 20.78 8.605 20.95 8.775 ;
      RECT 20.1 8.605 20.27 8.775 ;
      RECT 20.03 5.945 20.2 6.115 ;
      RECT 18.825 0.915 18.995 1.085 ;
      RECT 18.825 2.395 18.995 2.565 ;
      RECT 18.825 6.315 18.995 6.485 ;
      RECT 18.825 7.795 18.995 7.965 ;
      RECT 18.475 0.105 18.645 0.275 ;
      RECT 18.475 4.165 18.645 4.335 ;
      RECT 18.475 4.545 18.645 4.715 ;
      RECT 18.475 8.605 18.645 8.775 ;
      RECT 18.455 2.765 18.625 2.935 ;
      RECT 18.455 5.945 18.625 6.115 ;
      RECT 17.835 0.915 18.005 1.085 ;
      RECT 17.835 2.395 18.005 2.565 ;
      RECT 17.835 6.315 18.005 6.485 ;
      RECT 17.835 7.795 18.005 7.965 ;
      RECT 17.485 0.105 17.655 0.275 ;
      RECT 17.485 4.165 17.655 4.335 ;
      RECT 17.485 4.545 17.655 4.715 ;
      RECT 17.485 8.605 17.655 8.775 ;
      RECT 17.465 2.765 17.635 2.935 ;
      RECT 17.465 5.945 17.635 6.115 ;
      RECT 16.78 0.105 16.95 0.275 ;
      RECT 16.78 4.165 16.95 4.335 ;
      RECT 16.78 4.545 16.95 4.715 ;
      RECT 16.78 8.605 16.95 8.775 ;
      RECT 16.47 2.025 16.64 2.195 ;
      RECT 16.47 6.685 16.64 6.855 ;
      RECT 16.1 0.105 16.27 0.275 ;
      RECT 16.1 8.605 16.27 8.775 ;
      RECT 16.04 0.915 16.21 1.085 ;
      RECT 16.04 1.655 16.21 1.825 ;
      RECT 16.04 7.055 16.21 7.225 ;
      RECT 16.04 7.795 16.21 7.965 ;
      RECT 15.665 2.395 15.835 2.565 ;
      RECT 15.665 6.315 15.835 6.485 ;
      RECT 15.42 0.105 15.59 0.275 ;
      RECT 15.42 8.605 15.59 8.775 ;
      RECT 14.74 0.105 14.91 0.275 ;
      RECT 14.74 8.605 14.91 8.775 ;
      RECT 14.67 2.765 14.84 2.935 ;
      RECT 14.67 5.945 14.84 6.115 ;
      RECT 13.08 1.625 13.25 1.795 ;
      RECT 13.08 4.345 13.25 4.515 ;
      RECT 13.08 7.065 13.25 7.235 ;
      RECT 13.04 2.815 13.21 2.985 ;
      RECT 12.7 4.855 12.87 5.025 ;
      RECT 12.62 1.625 12.79 1.795 ;
      RECT 12.62 3.155 12.79 3.325 ;
      RECT 12.62 4.345 12.79 4.515 ;
      RECT 12.62 7.065 12.79 7.235 ;
      RECT 12.16 1.625 12.33 1.795 ;
      RECT 12.16 4.345 12.33 4.515 ;
      RECT 12.16 7.065 12.33 7.235 ;
      RECT 12.02 5.875 12.19 6.045 ;
      RECT 11.7 1.625 11.87 1.795 ;
      RECT 11.7 4.345 11.87 4.515 ;
      RECT 11.7 7.065 11.87 7.235 ;
      RECT 11.68 2.135 11.85 2.305 ;
      RECT 11.34 5.875 11.51 6.045 ;
      RECT 11.24 1.625 11.41 1.795 ;
      RECT 11.24 4.345 11.41 4.515 ;
      RECT 11.24 7.065 11.41 7.235 ;
      RECT 10.885 2.135 11.055 2.305 ;
      RECT 10.78 1.625 10.95 1.795 ;
      RECT 10.78 4.345 10.95 4.515 ;
      RECT 10.78 7.065 10.95 7.235 ;
      RECT 10.66 3.835 10.83 4.005 ;
      RECT 10.66 5.875 10.83 6.045 ;
      RECT 10.32 1.625 10.49 1.795 ;
      RECT 10.32 4.345 10.49 4.515 ;
      RECT 10.32 7.065 10.49 7.235 ;
      RECT 10.15 5.875 10.32 6.045 ;
      RECT 9.98 2.475 10.15 2.645 ;
      RECT 9.86 1.625 10.03 1.795 ;
      RECT 9.86 4.345 10.03 4.515 ;
      RECT 9.86 7.065 10.03 7.235 ;
      RECT 9.4 1.625 9.57 1.795 ;
      RECT 9.4 4.345 9.57 4.515 ;
      RECT 9.4 7.065 9.57 7.235 ;
      RECT 8.96 5.875 9.13 6.045 ;
      RECT 8.94 1.625 9.11 1.795 ;
      RECT 8.94 4.345 9.11 4.515 ;
      RECT 8.94 7.065 9.11 7.235 ;
      RECT 8.62 2.475 8.79 2.645 ;
      RECT 8.48 1.625 8.65 1.795 ;
      RECT 8.48 4.345 8.65 4.515 ;
      RECT 8.48 7.065 8.65 7.235 ;
      RECT 8.45 3.835 8.62 4.005 ;
      RECT 8.02 1.625 8.19 1.795 ;
      RECT 8.02 4.345 8.19 4.515 ;
      RECT 8.02 7.065 8.19 7.235 ;
      RECT 7.94 5.875 8.11 6.045 ;
      RECT 7.56 1.625 7.73 1.795 ;
      RECT 7.56 4.345 7.73 4.515 ;
      RECT 7.56 7.065 7.73 7.235 ;
      RECT 7.26 4.855 7.43 5.025 ;
      RECT 7.1 1.625 7.27 1.795 ;
      RECT 7.1 4.345 7.27 4.515 ;
      RECT 7.1 7.065 7.27 7.235 ;
      RECT 6.64 1.625 6.81 1.795 ;
      RECT 6.64 4.345 6.81 4.515 ;
      RECT 6.64 7.065 6.81 7.235 ;
      RECT 6.585 2.815 6.755 2.985 ;
      RECT 5.555 4.545 5.725 4.715 ;
      RECT 5.555 8.605 5.725 8.775 ;
      RECT 5.245 6.685 5.415 6.855 ;
      RECT 4.875 8.605 5.045 8.775 ;
      RECT 4.815 7.055 4.985 7.225 ;
      RECT 4.815 7.795 4.985 7.965 ;
      RECT 4.44 6.315 4.61 6.485 ;
      RECT 4.195 8.605 4.365 8.775 ;
      RECT 3.515 8.605 3.685 8.775 ;
      RECT 3.445 5.945 3.615 6.115 ;
      RECT 2.325 4.545 2.495 4.715 ;
      RECT 2.325 8.605 2.495 8.775 ;
      RECT 2.015 6.685 2.185 6.855 ;
      RECT 1.645 8.605 1.815 8.775 ;
      RECT 1.585 7.055 1.755 7.225 ;
      RECT 1.585 7.795 1.755 7.965 ;
      RECT 1.21 6.315 1.38 6.485 ;
      RECT 0.965 8.605 1.135 8.775 ;
      RECT 0.285 8.605 0.455 8.775 ;
      RECT 0.215 5.945 0.385 6.115 ;
    LAYER li ;
      RECT 0.025 8.57 85.73 8.88 ;
      RECT 84.73 7.945 84.9 8.88 ;
      RECT 83.74 7.945 83.91 8.88 ;
      RECT 80.995 7.945 81.165 8.88 ;
      RECT 72.535 7.18 79.735 8.88 ;
      RECT 69.77 7.945 69.94 8.88 ;
      RECT 68.15 7.945 68.32 8.88 ;
      RECT 67.16 7.945 67.33 8.88 ;
      RECT 64.415 7.945 64.585 8.88 ;
      RECT 55.955 7.18 63.155 8.88 ;
      RECT 53.19 7.945 53.36 8.88 ;
      RECT 51.565 7.945 51.735 8.88 ;
      RECT 50.575 7.945 50.745 8.88 ;
      RECT 47.83 7.945 48 8.88 ;
      RECT 39.37 7.18 46.57 8.88 ;
      RECT 36.605 7.945 36.775 8.88 ;
      RECT 34.98 7.945 35.15 8.88 ;
      RECT 33.99 7.945 34.16 8.88 ;
      RECT 31.245 7.945 31.415 8.88 ;
      RECT 22.785 7.18 29.985 8.88 ;
      RECT 20.02 7.945 20.19 8.88 ;
      RECT 18.395 7.945 18.565 8.88 ;
      RECT 17.405 7.945 17.575 8.88 ;
      RECT 14.66 7.945 14.83 8.88 ;
      RECT 6.2 7.18 13.4 8.88 ;
      RECT 3.435 7.945 3.605 8.88 ;
      RECT 0.205 7.945 0.375 8.88 ;
      RECT 72.83 7.065 79.73 8.88 ;
      RECT 56.25 7.065 63.15 8.88 ;
      RECT 39.665 7.065 46.565 8.88 ;
      RECT 23.08 7.065 29.98 8.88 ;
      RECT 6.495 7.065 13.395 8.88 ;
      RECT 78.265 6.555 78.715 8.88 ;
      RECT 76.175 6.665 76.505 8.88 ;
      RECT 74.105 6.605 74.355 8.88 ;
      RECT 61.685 6.555 62.135 8.88 ;
      RECT 59.595 6.665 59.925 8.88 ;
      RECT 57.525 6.605 57.775 8.88 ;
      RECT 45.1 6.555 45.55 8.88 ;
      RECT 43.01 6.665 43.34 8.88 ;
      RECT 40.94 6.605 41.19 8.88 ;
      RECT 28.515 6.555 28.965 8.88 ;
      RECT 26.425 6.665 26.755 8.88 ;
      RECT 24.355 6.605 24.605 8.88 ;
      RECT 11.93 6.555 12.38 8.88 ;
      RECT 9.84 6.665 10.17 8.88 ;
      RECT 7.77 6.605 8.02 8.88 ;
      RECT 72.915 0 73.175 2.615 ;
      RECT 56.335 0 56.595 2.615 ;
      RECT 39.75 0 40.01 2.615 ;
      RECT 23.165 0 23.425 2.615 ;
      RECT 6.58 0 6.84 2.615 ;
      RECT 79.365 0 79.635 2.605 ;
      RECT 78.455 0 78.695 2.605 ;
      RECT 62.785 0 63.055 2.605 ;
      RECT 61.875 0 62.115 2.605 ;
      RECT 46.2 0 46.47 2.605 ;
      RECT 45.29 0 45.53 2.605 ;
      RECT 29.615 0 29.885 2.605 ;
      RECT 28.705 0 28.945 2.605 ;
      RECT 13.03 0 13.3 2.605 ;
      RECT 12.12 0 12.36 2.605 ;
      RECT 77.585 0 77.835 2.335 ;
      RECT 61.005 0 61.255 2.335 ;
      RECT 44.42 0 44.67 2.335 ;
      RECT 27.835 0 28.085 2.335 ;
      RECT 11.25 0 11.5 2.335 ;
      RECT 75.205 0 75.535 2.255 ;
      RECT 58.625 0 58.955 2.255 ;
      RECT 42.04 0 42.37 2.255 ;
      RECT 25.455 0 25.785 2.255 ;
      RECT 8.87 0 9.2 2.255 ;
      RECT 72.83 0 79.92 1.795 ;
      RECT 56.25 0 63.34 1.795 ;
      RECT 39.665 0 46.755 1.795 ;
      RECT 23.08 0 30.17 1.795 ;
      RECT 6.495 0 13.585 1.795 ;
      RECT 72.575 0 79.92 1.655 ;
      RECT 55.995 0 63.34 1.655 ;
      RECT 39.41 0 46.755 1.655 ;
      RECT 22.825 0 30.17 1.655 ;
      RECT 6.24 0 13.585 1.655 ;
      RECT 84.73 0 84.9 0.935 ;
      RECT 83.74 0 83.91 0.935 ;
      RECT 80.995 0 81.165 0.935 ;
      RECT 68.15 0 68.32 0.935 ;
      RECT 67.16 0 67.33 0.935 ;
      RECT 64.415 0 64.585 0.935 ;
      RECT 51.565 0 51.735 0.935 ;
      RECT 50.575 0 50.745 0.935 ;
      RECT 47.83 0 48 0.935 ;
      RECT 34.98 0 35.15 0.935 ;
      RECT 33.99 0 34.16 0.935 ;
      RECT 31.245 0 31.415 0.935 ;
      RECT 18.395 0 18.565 0.935 ;
      RECT 17.405 0 17.575 0.935 ;
      RECT 14.66 0 14.83 0.935 ;
      RECT 0 0 85.705 0.31 ;
      RECT 2.015 4.13 2.185 8.305 ;
      RECT 84.73 3.405 84.9 5.475 ;
      RECT 83.74 3.405 83.91 5.475 ;
      RECT 80.995 3.405 81.165 5.475 ;
      RECT 69.77 4.13 69.94 5.475 ;
      RECT 68.15 3.405 68.32 5.475 ;
      RECT 67.16 3.405 67.33 5.475 ;
      RECT 64.415 3.405 64.585 5.475 ;
      RECT 53.19 4.13 53.36 5.475 ;
      RECT 51.565 3.405 51.735 5.475 ;
      RECT 50.575 3.405 50.745 5.475 ;
      RECT 47.83 3.405 48 5.475 ;
      RECT 36.605 4.13 36.775 5.475 ;
      RECT 34.98 3.405 35.15 5.475 ;
      RECT 33.99 3.405 34.16 5.475 ;
      RECT 31.245 3.405 31.415 5.475 ;
      RECT 20.02 4.13 20.19 5.475 ;
      RECT 18.395 3.405 18.565 5.475 ;
      RECT 17.405 3.405 17.575 5.475 ;
      RECT 14.66 3.405 14.83 5.475 ;
      RECT 3.435 4.13 3.605 5.475 ;
      RECT 0.205 4.13 0.375 5.475 ;
      RECT 76.185 3.69 76.45 5.295 ;
      RECT 59.605 3.69 59.87 5.295 ;
      RECT 43.02 3.69 43.285 5.295 ;
      RECT 26.435 3.69 26.7 5.295 ;
      RECT 9.85 3.69 10.115 5.295 ;
      RECT 74.025 3.84 74.355 5.235 ;
      RECT 57.445 3.84 57.775 5.235 ;
      RECT 40.86 3.84 41.19 5.235 ;
      RECT 24.275 3.84 24.605 5.235 ;
      RECT 7.69 3.84 8.02 5.235 ;
      RECT 75.025 4.345 75.305 5.185 ;
      RECT 58.445 4.345 58.725 5.185 ;
      RECT 41.86 4.345 42.14 5.185 ;
      RECT 25.275 4.345 25.555 5.185 ;
      RECT 8.69 4.345 8.97 5.185 ;
      RECT 77 4.345 77.375 4.895 ;
      RECT 60.42 4.345 60.795 4.895 ;
      RECT 43.835 4.345 44.21 4.895 ;
      RECT 27.25 4.345 27.625 4.895 ;
      RECT 10.665 4.345 11.04 4.895 ;
      RECT 79.76 4.135 85.7 4.745 ;
      RECT 69.595 4.13 72.345 4.745 ;
      RECT 63.18 4.135 69.12 4.745 ;
      RECT 53.015 4.13 55.765 4.745 ;
      RECT 46.595 4.135 52.535 4.745 ;
      RECT 36.43 4.13 39.18 4.745 ;
      RECT 30.01 4.135 35.95 4.745 ;
      RECT 19.845 4.13 22.595 4.745 ;
      RECT 13.425 4.135 19.365 4.745 ;
      RECT 3.26 4.13 6.01 4.745 ;
      RECT 0.03 4.13 2.78 4.745 ;
      RECT 69.115 4.13 72.69 4.74 ;
      RECT 52.535 4.13 56.11 4.74 ;
      RECT 35.95 4.13 39.525 4.74 ;
      RECT 19.365 4.13 22.94 4.74 ;
      RECT 0.03 4.13 6.355 4.74 ;
      RECT 79.63 4.135 85.7 4.67 ;
      RECT 63.05 4.135 72.69 4.67 ;
      RECT 46.465 4.135 56.11 4.67 ;
      RECT 29.88 4.135 39.525 4.67 ;
      RECT 13.295 4.135 22.94 4.67 ;
      RECT 0.03 4.345 85.7 4.515 ;
      RECT 79.305 3.205 79.635 4.515 ;
      RECT 77.565 3.8 77.82 4.515 ;
      RECT 76.135 3.69 76.74 4.515 ;
      RECT 75.265 3.8 75.48 4.515 ;
      RECT 73.835 3.84 74.45 4.515 ;
      RECT 74.255 3.475 74.45 4.515 ;
      RECT 72.915 3.835 73.175 4.515 ;
      RECT 62.725 3.205 63.055 4.515 ;
      RECT 60.985 3.8 61.24 4.515 ;
      RECT 59.555 3.69 60.16 4.515 ;
      RECT 58.685 3.8 58.9 4.515 ;
      RECT 57.255 3.84 57.87 4.515 ;
      RECT 57.675 3.475 57.87 4.515 ;
      RECT 56.335 3.835 56.595 4.515 ;
      RECT 46.14 3.205 46.47 4.515 ;
      RECT 44.4 3.8 44.655 4.515 ;
      RECT 42.97 3.69 43.575 4.515 ;
      RECT 42.1 3.8 42.315 4.515 ;
      RECT 40.67 3.84 41.285 4.515 ;
      RECT 41.09 3.475 41.285 4.515 ;
      RECT 39.75 3.835 40.01 4.515 ;
      RECT 29.555 3.205 29.885 4.515 ;
      RECT 27.815 3.8 28.07 4.515 ;
      RECT 26.385 3.69 26.99 4.515 ;
      RECT 25.515 3.8 25.73 4.515 ;
      RECT 24.085 3.84 24.7 4.515 ;
      RECT 24.505 3.475 24.7 4.515 ;
      RECT 23.165 3.835 23.425 4.515 ;
      RECT 12.97 3.205 13.3 4.515 ;
      RECT 11.23 3.8 11.485 4.515 ;
      RECT 9.8 3.69 10.405 4.515 ;
      RECT 8.93 3.8 9.145 4.515 ;
      RECT 7.5 3.84 8.115 4.515 ;
      RECT 7.92 3.475 8.115 4.515 ;
      RECT 6.58 3.835 6.84 4.515 ;
      RECT 76.565 3.42 76.75 3.79 ;
      RECT 59.985 3.42 60.17 3.79 ;
      RECT 43.4 3.42 43.585 3.79 ;
      RECT 26.815 3.42 27 3.79 ;
      RECT 10.23 3.42 10.415 3.79 ;
      RECT 76.565 3.42 76.895 3.665 ;
      RECT 74.255 3.475 74.585 3.665 ;
      RECT 59.985 3.42 60.315 3.665 ;
      RECT 57.675 3.475 58.005 3.665 ;
      RECT 43.4 3.42 43.73 3.665 ;
      RECT 41.09 3.475 41.42 3.665 ;
      RECT 26.815 3.42 27.145 3.665 ;
      RECT 24.505 3.475 24.835 3.665 ;
      RECT 10.23 3.42 10.56 3.665 ;
      RECT 7.92 3.475 8.25 3.665 ;
      RECT 84.79 1.74 84.96 2.935 ;
      RECT 84.79 1.74 85.255 1.91 ;
      RECT 84.79 6.97 85.255 7.14 ;
      RECT 84.79 5.945 84.96 7.14 ;
      RECT 83.8 1.74 83.97 2.935 ;
      RECT 83.8 1.74 84.265 1.91 ;
      RECT 83.8 6.97 84.265 7.14 ;
      RECT 83.8 5.945 83.97 7.14 ;
      RECT 81.945 2.635 82.115 3.865 ;
      RECT 82 0.855 82.17 2.805 ;
      RECT 81.945 0.575 82.115 1.025 ;
      RECT 81.945 7.855 82.115 8.305 ;
      RECT 82 6.075 82.17 8.025 ;
      RECT 81.945 5.015 82.115 6.245 ;
      RECT 81.425 0.575 81.595 3.865 ;
      RECT 81.425 2.075 81.83 2.405 ;
      RECT 81.425 1.235 81.83 1.565 ;
      RECT 81.425 5.015 81.595 8.305 ;
      RECT 81.425 7.315 81.83 7.645 ;
      RECT 81.425 6.475 81.83 6.805 ;
      RECT 76.685 6.645 77.99 6.895 ;
      RECT 76.685 6.325 76.865 6.895 ;
      RECT 76.135 6.325 76.865 6.495 ;
      RECT 76.135 5.485 76.305 6.495 ;
      RECT 76.97 5.525 78.715 5.705 ;
      RECT 78.385 4.685 78.715 5.705 ;
      RECT 76.135 5.485 77.195 5.655 ;
      RECT 78.385 4.855 79.205 5.025 ;
      RECT 77.545 4.685 77.875 4.895 ;
      RECT 77.545 4.685 78.715 4.855 ;
      RECT 78.445 3.205 78.775 4.16 ;
      RECT 78.445 3.205 79.125 3.375 ;
      RECT 78.955 1.965 79.125 3.375 ;
      RECT 78.865 1.965 79.195 2.605 ;
      RECT 77.99 3.475 78.265 4.175 ;
      RECT 78.095 1.965 78.265 4.175 ;
      RECT 78.435 2.785 78.785 3.035 ;
      RECT 78.095 2.815 78.785 2.985 ;
      RECT 78.005 1.965 78.265 2.445 ;
      RECT 77.335 5.115 78.215 5.355 ;
      RECT 77.985 5.025 78.215 5.355 ;
      RECT 76.685 5.115 78.215 5.315 ;
      RECT 77.6 5.065 78.215 5.355 ;
      RECT 76.685 4.985 76.855 5.315 ;
      RECT 77.57 5.875 77.82 6.475 ;
      RECT 77.57 5.875 78.045 6.075 ;
      RECT 77.065 3.095 77.82 3.595 ;
      RECT 76.135 2.9 76.395 3.52 ;
      RECT 77.05 3.04 77.065 3.345 ;
      RECT 77.035 3.025 77.055 3.31 ;
      RECT 77.695 2.7 77.925 3.3 ;
      RECT 77.01 2.97 77.03 3.285 ;
      RECT 76.99 3.095 77.925 3.27 ;
      RECT 76.965 3.095 77.925 3.26 ;
      RECT 76.895 3.095 77.925 3.25 ;
      RECT 76.875 3.095 77.925 3.22 ;
      RECT 76.855 2.005 77.025 3.19 ;
      RECT 76.825 3.095 77.925 3.16 ;
      RECT 76.79 3.095 77.925 3.135 ;
      RECT 76.76 3.09 77.15 3.1 ;
      RECT 76.76 3.08 77.125 3.1 ;
      RECT 76.76 3.075 77.11 3.1 ;
      RECT 76.76 3.065 77.095 3.1 ;
      RECT 76.135 2.9 77.025 3.07 ;
      RECT 76.135 3.055 77.085 3.07 ;
      RECT 76.135 3.05 77.075 3.07 ;
      RECT 77.03 2.995 77.04 3.3 ;
      RECT 76.135 3.03 77.06 3.07 ;
      RECT 76.135 3.01 77.045 3.07 ;
      RECT 76.135 2.005 77.025 2.175 ;
      RECT 77.195 2.5 77.525 2.925 ;
      RECT 77.195 2.015 77.415 2.925 ;
      RECT 77.11 5.875 77.32 6.475 ;
      RECT 76.97 5.875 77.32 6.075 ;
      RECT 75.69 3.475 75.965 4.175 ;
      RECT 75.91 1.965 75.965 4.175 ;
      RECT 75.795 2.77 75.965 4.175 ;
      RECT 75.795 1.965 75.965 2.765 ;
      RECT 75.705 1.965 75.965 2.44 ;
      RECT 73.835 3.135 74.085 3.67 ;
      RECT 74.805 3.135 75.52 3.6 ;
      RECT 73.835 3.135 75.625 3.305 ;
      RECT 75.395 2.77 75.625 3.305 ;
      RECT 74.39 2.015 74.645 3.305 ;
      RECT 75.395 2.705 75.455 3.6 ;
      RECT 75.455 2.7 75.625 2.765 ;
      RECT 73.855 2.015 74.645 2.28 ;
      RECT 74.815 5.825 75.49 6.075 ;
      RECT 75.225 5.465 75.49 6.075 ;
      RECT 74.975 6.245 75.305 6.795 ;
      RECT 73.915 6.245 75.305 6.435 ;
      RECT 73.915 5.405 74.085 6.435 ;
      RECT 73.795 5.825 74.085 6.155 ;
      RECT 73.915 5.405 74.855 5.575 ;
      RECT 74.555 4.855 74.855 5.575 ;
      RECT 74.815 2.435 75.225 2.955 ;
      RECT 74.815 2.015 75.015 2.955 ;
      RECT 73.425 2.195 73.595 4.175 ;
      RECT 73.425 2.705 74.22 2.955 ;
      RECT 73.425 2.195 73.675 2.955 ;
      RECT 73.345 2.195 73.675 2.615 ;
      RECT 73.375 6.605 73.935 6.895 ;
      RECT 73.375 4.685 73.625 6.895 ;
      RECT 73.375 4.685 73.835 5.235 ;
      RECT 70.72 7.855 70.89 8.305 ;
      RECT 70.775 6.075 70.945 8.025 ;
      RECT 70.72 5.015 70.89 6.245 ;
      RECT 70.2 5.015 70.37 8.305 ;
      RECT 70.2 7.315 70.605 7.645 ;
      RECT 70.2 6.475 70.605 6.805 ;
      RECT 68.21 1.74 68.38 2.935 ;
      RECT 68.21 1.74 68.675 1.91 ;
      RECT 68.21 6.97 68.675 7.14 ;
      RECT 68.21 5.945 68.38 7.14 ;
      RECT 67.22 1.74 67.39 2.935 ;
      RECT 67.22 1.74 67.685 1.91 ;
      RECT 67.22 6.97 67.685 7.14 ;
      RECT 67.22 5.945 67.39 7.14 ;
      RECT 65.365 2.635 65.535 3.865 ;
      RECT 65.42 0.855 65.59 2.805 ;
      RECT 65.365 0.575 65.535 1.025 ;
      RECT 65.365 7.855 65.535 8.305 ;
      RECT 65.42 6.075 65.59 8.025 ;
      RECT 65.365 5.015 65.535 6.245 ;
      RECT 64.845 0.575 65.015 3.865 ;
      RECT 64.845 2.075 65.25 2.405 ;
      RECT 64.845 1.235 65.25 1.565 ;
      RECT 64.845 5.015 65.015 8.305 ;
      RECT 64.845 7.315 65.25 7.645 ;
      RECT 64.845 6.475 65.25 6.805 ;
      RECT 60.105 6.645 61.41 6.895 ;
      RECT 60.105 6.325 60.285 6.895 ;
      RECT 59.555 6.325 60.285 6.495 ;
      RECT 59.555 5.485 59.725 6.495 ;
      RECT 60.39 5.525 62.135 5.705 ;
      RECT 61.805 4.685 62.135 5.705 ;
      RECT 59.555 5.485 60.615 5.655 ;
      RECT 61.805 4.855 62.625 5.025 ;
      RECT 60.965 4.685 61.295 4.895 ;
      RECT 60.965 4.685 62.135 4.855 ;
      RECT 61.865 3.205 62.195 4.16 ;
      RECT 61.865 3.205 62.545 3.375 ;
      RECT 62.375 1.965 62.545 3.375 ;
      RECT 62.285 1.965 62.615 2.605 ;
      RECT 61.41 3.475 61.685 4.175 ;
      RECT 61.515 1.965 61.685 4.175 ;
      RECT 61.855 2.785 62.205 3.035 ;
      RECT 61.515 2.815 62.205 2.985 ;
      RECT 61.425 1.965 61.685 2.445 ;
      RECT 60.755 5.115 61.635 5.355 ;
      RECT 61.405 5.025 61.635 5.355 ;
      RECT 60.105 5.115 61.635 5.315 ;
      RECT 61.02 5.065 61.635 5.355 ;
      RECT 60.105 4.985 60.275 5.315 ;
      RECT 60.99 5.875 61.24 6.475 ;
      RECT 60.99 5.875 61.465 6.075 ;
      RECT 60.485 3.095 61.24 3.595 ;
      RECT 59.555 2.9 59.815 3.52 ;
      RECT 60.47 3.04 60.485 3.345 ;
      RECT 60.455 3.025 60.475 3.31 ;
      RECT 61.115 2.7 61.345 3.3 ;
      RECT 60.43 2.97 60.45 3.285 ;
      RECT 60.41 3.095 61.345 3.27 ;
      RECT 60.385 3.095 61.345 3.26 ;
      RECT 60.315 3.095 61.345 3.25 ;
      RECT 60.295 3.095 61.345 3.22 ;
      RECT 60.275 2.005 60.445 3.19 ;
      RECT 60.245 3.095 61.345 3.16 ;
      RECT 60.21 3.095 61.345 3.135 ;
      RECT 60.18 3.09 60.57 3.1 ;
      RECT 60.18 3.08 60.545 3.1 ;
      RECT 60.18 3.075 60.53 3.1 ;
      RECT 60.18 3.065 60.515 3.1 ;
      RECT 59.555 2.9 60.445 3.07 ;
      RECT 59.555 3.055 60.505 3.07 ;
      RECT 59.555 3.05 60.495 3.07 ;
      RECT 60.45 2.995 60.46 3.3 ;
      RECT 59.555 3.03 60.48 3.07 ;
      RECT 59.555 3.01 60.465 3.07 ;
      RECT 59.555 2.005 60.445 2.175 ;
      RECT 60.615 2.5 60.945 2.925 ;
      RECT 60.615 2.015 60.835 2.925 ;
      RECT 60.53 5.875 60.74 6.475 ;
      RECT 60.39 5.875 60.74 6.075 ;
      RECT 59.11 3.475 59.385 4.175 ;
      RECT 59.33 1.965 59.385 4.175 ;
      RECT 59.215 2.77 59.385 4.175 ;
      RECT 59.215 1.965 59.385 2.765 ;
      RECT 59.125 1.965 59.385 2.44 ;
      RECT 57.255 3.135 57.505 3.67 ;
      RECT 58.225 3.135 58.94 3.6 ;
      RECT 57.255 3.135 59.045 3.305 ;
      RECT 58.815 2.77 59.045 3.305 ;
      RECT 57.81 2.015 58.065 3.305 ;
      RECT 58.815 2.705 58.875 3.6 ;
      RECT 58.875 2.7 59.045 2.765 ;
      RECT 57.275 2.015 58.065 2.28 ;
      RECT 58.235 5.825 58.91 6.075 ;
      RECT 58.645 5.465 58.91 6.075 ;
      RECT 58.395 6.245 58.725 6.795 ;
      RECT 57.335 6.245 58.725 6.435 ;
      RECT 57.335 5.405 57.505 6.435 ;
      RECT 57.215 5.825 57.505 6.155 ;
      RECT 57.335 5.405 58.275 5.575 ;
      RECT 57.975 4.855 58.275 5.575 ;
      RECT 58.235 2.435 58.645 2.955 ;
      RECT 58.235 2.015 58.435 2.955 ;
      RECT 56.845 2.195 57.015 4.175 ;
      RECT 56.845 2.705 57.64 2.955 ;
      RECT 56.845 2.195 57.095 2.955 ;
      RECT 56.765 2.195 57.095 2.615 ;
      RECT 56.795 6.605 57.355 6.895 ;
      RECT 56.795 4.685 57.045 6.895 ;
      RECT 56.795 4.685 57.255 5.235 ;
      RECT 54.14 7.855 54.31 8.305 ;
      RECT 54.195 6.075 54.365 8.025 ;
      RECT 54.14 5.015 54.31 6.245 ;
      RECT 53.62 5.015 53.79 8.305 ;
      RECT 53.62 7.315 54.025 7.645 ;
      RECT 53.62 6.475 54.025 6.805 ;
      RECT 51.625 1.74 51.795 2.935 ;
      RECT 51.625 1.74 52.09 1.91 ;
      RECT 51.625 6.97 52.09 7.14 ;
      RECT 51.625 5.945 51.795 7.14 ;
      RECT 50.635 1.74 50.805 2.935 ;
      RECT 50.635 1.74 51.1 1.91 ;
      RECT 50.635 6.97 51.1 7.14 ;
      RECT 50.635 5.945 50.805 7.14 ;
      RECT 48.78 2.635 48.95 3.865 ;
      RECT 48.835 0.855 49.005 2.805 ;
      RECT 48.78 0.575 48.95 1.025 ;
      RECT 48.78 7.855 48.95 8.305 ;
      RECT 48.835 6.075 49.005 8.025 ;
      RECT 48.78 5.015 48.95 6.245 ;
      RECT 48.26 0.575 48.43 3.865 ;
      RECT 48.26 2.075 48.665 2.405 ;
      RECT 48.26 1.235 48.665 1.565 ;
      RECT 48.26 5.015 48.43 8.305 ;
      RECT 48.26 7.315 48.665 7.645 ;
      RECT 48.26 6.475 48.665 6.805 ;
      RECT 43.52 6.645 44.825 6.895 ;
      RECT 43.52 6.325 43.7 6.895 ;
      RECT 42.97 6.325 43.7 6.495 ;
      RECT 42.97 5.485 43.14 6.495 ;
      RECT 43.805 5.525 45.55 5.705 ;
      RECT 45.22 4.685 45.55 5.705 ;
      RECT 42.97 5.485 44.03 5.655 ;
      RECT 45.22 4.855 46.04 5.025 ;
      RECT 44.38 4.685 44.71 4.895 ;
      RECT 44.38 4.685 45.55 4.855 ;
      RECT 45.28 3.205 45.61 4.16 ;
      RECT 45.28 3.205 45.96 3.375 ;
      RECT 45.79 1.965 45.96 3.375 ;
      RECT 45.7 1.965 46.03 2.605 ;
      RECT 44.825 3.475 45.1 4.175 ;
      RECT 44.93 1.965 45.1 4.175 ;
      RECT 45.27 2.785 45.62 3.035 ;
      RECT 44.93 2.815 45.62 2.985 ;
      RECT 44.84 1.965 45.1 2.445 ;
      RECT 44.17 5.115 45.05 5.355 ;
      RECT 44.82 5.025 45.05 5.355 ;
      RECT 43.52 5.115 45.05 5.315 ;
      RECT 44.435 5.065 45.05 5.355 ;
      RECT 43.52 4.985 43.69 5.315 ;
      RECT 44.405 5.875 44.655 6.475 ;
      RECT 44.405 5.875 44.88 6.075 ;
      RECT 43.9 3.095 44.655 3.595 ;
      RECT 42.97 2.9 43.23 3.52 ;
      RECT 43.885 3.04 43.9 3.345 ;
      RECT 43.87 3.025 43.89 3.31 ;
      RECT 44.53 2.7 44.76 3.3 ;
      RECT 43.845 2.97 43.865 3.285 ;
      RECT 43.825 3.095 44.76 3.27 ;
      RECT 43.8 3.095 44.76 3.26 ;
      RECT 43.73 3.095 44.76 3.25 ;
      RECT 43.71 3.095 44.76 3.22 ;
      RECT 43.69 2.005 43.86 3.19 ;
      RECT 43.66 3.095 44.76 3.16 ;
      RECT 43.625 3.095 44.76 3.135 ;
      RECT 43.595 3.09 43.985 3.1 ;
      RECT 43.595 3.08 43.96 3.1 ;
      RECT 43.595 3.075 43.945 3.1 ;
      RECT 43.595 3.065 43.93 3.1 ;
      RECT 42.97 2.9 43.86 3.07 ;
      RECT 42.97 3.055 43.92 3.07 ;
      RECT 42.97 3.05 43.91 3.07 ;
      RECT 43.865 2.995 43.875 3.3 ;
      RECT 42.97 3.03 43.895 3.07 ;
      RECT 42.97 3.01 43.88 3.07 ;
      RECT 42.97 2.005 43.86 2.175 ;
      RECT 44.03 2.5 44.36 2.925 ;
      RECT 44.03 2.015 44.25 2.925 ;
      RECT 43.945 5.875 44.155 6.475 ;
      RECT 43.805 5.875 44.155 6.075 ;
      RECT 42.525 3.475 42.8 4.175 ;
      RECT 42.745 1.965 42.8 4.175 ;
      RECT 42.63 2.77 42.8 4.175 ;
      RECT 42.63 1.965 42.8 2.765 ;
      RECT 42.54 1.965 42.8 2.44 ;
      RECT 40.67 3.135 40.92 3.67 ;
      RECT 41.64 3.135 42.355 3.6 ;
      RECT 40.67 3.135 42.46 3.305 ;
      RECT 42.23 2.77 42.46 3.305 ;
      RECT 41.225 2.015 41.48 3.305 ;
      RECT 42.23 2.705 42.29 3.6 ;
      RECT 42.29 2.7 42.46 2.765 ;
      RECT 40.69 2.015 41.48 2.28 ;
      RECT 41.65 5.825 42.325 6.075 ;
      RECT 42.06 5.465 42.325 6.075 ;
      RECT 41.81 6.245 42.14 6.795 ;
      RECT 40.75 6.245 42.14 6.435 ;
      RECT 40.75 5.405 40.92 6.435 ;
      RECT 40.63 5.825 40.92 6.155 ;
      RECT 40.75 5.405 41.69 5.575 ;
      RECT 41.39 4.855 41.69 5.575 ;
      RECT 41.65 2.435 42.06 2.955 ;
      RECT 41.65 2.015 41.85 2.955 ;
      RECT 40.26 2.195 40.43 4.175 ;
      RECT 40.26 2.705 41.055 2.955 ;
      RECT 40.26 2.195 40.51 2.955 ;
      RECT 40.18 2.195 40.51 2.615 ;
      RECT 40.21 6.605 40.77 6.895 ;
      RECT 40.21 4.685 40.46 6.895 ;
      RECT 40.21 4.685 40.67 5.235 ;
      RECT 37.555 7.855 37.725 8.305 ;
      RECT 37.61 6.075 37.78 8.025 ;
      RECT 37.555 5.015 37.725 6.245 ;
      RECT 37.035 5.015 37.205 8.305 ;
      RECT 37.035 7.315 37.44 7.645 ;
      RECT 37.035 6.475 37.44 6.805 ;
      RECT 35.04 1.74 35.21 2.935 ;
      RECT 35.04 1.74 35.505 1.91 ;
      RECT 35.04 6.97 35.505 7.14 ;
      RECT 35.04 5.945 35.21 7.14 ;
      RECT 34.05 1.74 34.22 2.935 ;
      RECT 34.05 1.74 34.515 1.91 ;
      RECT 34.05 6.97 34.515 7.14 ;
      RECT 34.05 5.945 34.22 7.14 ;
      RECT 32.195 2.635 32.365 3.865 ;
      RECT 32.25 0.855 32.42 2.805 ;
      RECT 32.195 0.575 32.365 1.025 ;
      RECT 32.195 7.855 32.365 8.305 ;
      RECT 32.25 6.075 32.42 8.025 ;
      RECT 32.195 5.015 32.365 6.245 ;
      RECT 31.675 0.575 31.845 3.865 ;
      RECT 31.675 2.075 32.08 2.405 ;
      RECT 31.675 1.235 32.08 1.565 ;
      RECT 31.675 5.015 31.845 8.305 ;
      RECT 31.675 7.315 32.08 7.645 ;
      RECT 31.675 6.475 32.08 6.805 ;
      RECT 26.935 6.645 28.24 6.895 ;
      RECT 26.935 6.325 27.115 6.895 ;
      RECT 26.385 6.325 27.115 6.495 ;
      RECT 26.385 5.485 26.555 6.495 ;
      RECT 27.22 5.525 28.965 5.705 ;
      RECT 28.635 4.685 28.965 5.705 ;
      RECT 26.385 5.485 27.445 5.655 ;
      RECT 28.635 4.855 29.455 5.025 ;
      RECT 27.795 4.685 28.125 4.895 ;
      RECT 27.795 4.685 28.965 4.855 ;
      RECT 28.695 3.205 29.025 4.16 ;
      RECT 28.695 3.205 29.375 3.375 ;
      RECT 29.205 1.965 29.375 3.375 ;
      RECT 29.115 1.965 29.445 2.605 ;
      RECT 28.24 3.475 28.515 4.175 ;
      RECT 28.345 1.965 28.515 4.175 ;
      RECT 28.685 2.785 29.035 3.035 ;
      RECT 28.345 2.815 29.035 2.985 ;
      RECT 28.255 1.965 28.515 2.445 ;
      RECT 27.585 5.115 28.465 5.355 ;
      RECT 28.235 5.025 28.465 5.355 ;
      RECT 26.935 5.115 28.465 5.315 ;
      RECT 27.85 5.065 28.465 5.355 ;
      RECT 26.935 4.985 27.105 5.315 ;
      RECT 27.82 5.875 28.07 6.475 ;
      RECT 27.82 5.875 28.295 6.075 ;
      RECT 27.315 3.095 28.07 3.595 ;
      RECT 26.385 2.9 26.645 3.52 ;
      RECT 27.3 3.04 27.315 3.345 ;
      RECT 27.285 3.025 27.305 3.31 ;
      RECT 27.945 2.7 28.175 3.3 ;
      RECT 27.26 2.97 27.28 3.285 ;
      RECT 27.24 3.095 28.175 3.27 ;
      RECT 27.215 3.095 28.175 3.26 ;
      RECT 27.145 3.095 28.175 3.25 ;
      RECT 27.125 3.095 28.175 3.22 ;
      RECT 27.105 2.005 27.275 3.19 ;
      RECT 27.075 3.095 28.175 3.16 ;
      RECT 27.04 3.095 28.175 3.135 ;
      RECT 27.01 3.09 27.4 3.1 ;
      RECT 27.01 3.08 27.375 3.1 ;
      RECT 27.01 3.075 27.36 3.1 ;
      RECT 27.01 3.065 27.345 3.1 ;
      RECT 26.385 2.9 27.275 3.07 ;
      RECT 26.385 3.055 27.335 3.07 ;
      RECT 26.385 3.05 27.325 3.07 ;
      RECT 27.28 2.995 27.29 3.3 ;
      RECT 26.385 3.03 27.31 3.07 ;
      RECT 26.385 3.01 27.295 3.07 ;
      RECT 26.385 2.005 27.275 2.175 ;
      RECT 27.445 2.5 27.775 2.925 ;
      RECT 27.445 2.015 27.665 2.925 ;
      RECT 27.36 5.875 27.57 6.475 ;
      RECT 27.22 5.875 27.57 6.075 ;
      RECT 25.94 3.475 26.215 4.175 ;
      RECT 26.16 1.965 26.215 4.175 ;
      RECT 26.045 2.77 26.215 4.175 ;
      RECT 26.045 1.965 26.215 2.765 ;
      RECT 25.955 1.965 26.215 2.44 ;
      RECT 24.085 3.135 24.335 3.67 ;
      RECT 25.055 3.135 25.77 3.6 ;
      RECT 24.085 3.135 25.875 3.305 ;
      RECT 25.645 2.77 25.875 3.305 ;
      RECT 24.64 2.015 24.895 3.305 ;
      RECT 25.645 2.705 25.705 3.6 ;
      RECT 25.705 2.7 25.875 2.765 ;
      RECT 24.105 2.015 24.895 2.28 ;
      RECT 25.065 5.825 25.74 6.075 ;
      RECT 25.475 5.465 25.74 6.075 ;
      RECT 25.225 6.245 25.555 6.795 ;
      RECT 24.165 6.245 25.555 6.435 ;
      RECT 24.165 5.405 24.335 6.435 ;
      RECT 24.045 5.825 24.335 6.155 ;
      RECT 24.165 5.405 25.105 5.575 ;
      RECT 24.805 4.855 25.105 5.575 ;
      RECT 25.065 2.435 25.475 2.955 ;
      RECT 25.065 2.015 25.265 2.955 ;
      RECT 23.675 2.195 23.845 4.175 ;
      RECT 23.675 2.705 24.47 2.955 ;
      RECT 23.675 2.195 23.925 2.955 ;
      RECT 23.595 2.195 23.925 2.615 ;
      RECT 23.625 6.605 24.185 6.895 ;
      RECT 23.625 4.685 23.875 6.895 ;
      RECT 23.625 4.685 24.085 5.235 ;
      RECT 20.97 7.855 21.14 8.305 ;
      RECT 21.025 6.075 21.195 8.025 ;
      RECT 20.97 5.015 21.14 6.245 ;
      RECT 20.45 5.015 20.62 8.305 ;
      RECT 20.45 7.315 20.855 7.645 ;
      RECT 20.45 6.475 20.855 6.805 ;
      RECT 18.455 1.74 18.625 2.935 ;
      RECT 18.455 1.74 18.92 1.91 ;
      RECT 18.455 6.97 18.92 7.14 ;
      RECT 18.455 5.945 18.625 7.14 ;
      RECT 17.465 1.74 17.635 2.935 ;
      RECT 17.465 1.74 17.93 1.91 ;
      RECT 17.465 6.97 17.93 7.14 ;
      RECT 17.465 5.945 17.635 7.14 ;
      RECT 15.61 2.635 15.78 3.865 ;
      RECT 15.665 0.855 15.835 2.805 ;
      RECT 15.61 0.575 15.78 1.025 ;
      RECT 15.61 7.855 15.78 8.305 ;
      RECT 15.665 6.075 15.835 8.025 ;
      RECT 15.61 5.015 15.78 6.245 ;
      RECT 15.09 0.575 15.26 3.865 ;
      RECT 15.09 2.075 15.495 2.405 ;
      RECT 15.09 1.235 15.495 1.565 ;
      RECT 15.09 5.015 15.26 8.305 ;
      RECT 15.09 7.315 15.495 7.645 ;
      RECT 15.09 6.475 15.495 6.805 ;
      RECT 10.35 6.645 11.655 6.895 ;
      RECT 10.35 6.325 10.53 6.895 ;
      RECT 9.8 6.325 10.53 6.495 ;
      RECT 9.8 5.485 9.97 6.495 ;
      RECT 10.635 5.525 12.38 5.705 ;
      RECT 12.05 4.685 12.38 5.705 ;
      RECT 9.8 5.485 10.86 5.655 ;
      RECT 12.05 4.855 12.87 5.025 ;
      RECT 11.21 4.685 11.54 4.895 ;
      RECT 11.21 4.685 12.38 4.855 ;
      RECT 12.11 3.205 12.44 4.16 ;
      RECT 12.11 3.205 12.79 3.375 ;
      RECT 12.62 1.965 12.79 3.375 ;
      RECT 12.53 1.965 12.86 2.605 ;
      RECT 11.655 3.475 11.93 4.175 ;
      RECT 11.76 1.965 11.93 4.175 ;
      RECT 12.1 2.785 12.45 3.035 ;
      RECT 11.76 2.815 12.45 2.985 ;
      RECT 11.67 1.965 11.93 2.445 ;
      RECT 11 5.115 11.88 5.355 ;
      RECT 11.65 5.025 11.88 5.355 ;
      RECT 10.35 5.115 11.88 5.315 ;
      RECT 11.265 5.065 11.88 5.355 ;
      RECT 10.35 4.985 10.52 5.315 ;
      RECT 11.235 5.875 11.485 6.475 ;
      RECT 11.235 5.875 11.71 6.075 ;
      RECT 10.73 3.095 11.485 3.595 ;
      RECT 9.8 2.9 10.06 3.52 ;
      RECT 10.715 3.04 10.73 3.345 ;
      RECT 10.7 3.025 10.72 3.31 ;
      RECT 11.36 2.7 11.59 3.3 ;
      RECT 10.675 2.97 10.695 3.285 ;
      RECT 10.655 3.095 11.59 3.27 ;
      RECT 10.63 3.095 11.59 3.26 ;
      RECT 10.56 3.095 11.59 3.25 ;
      RECT 10.54 3.095 11.59 3.22 ;
      RECT 10.52 2.005 10.69 3.19 ;
      RECT 10.49 3.095 11.59 3.16 ;
      RECT 10.455 3.095 11.59 3.135 ;
      RECT 10.425 3.09 10.815 3.1 ;
      RECT 10.425 3.08 10.79 3.1 ;
      RECT 10.425 3.075 10.775 3.1 ;
      RECT 10.425 3.065 10.76 3.1 ;
      RECT 9.8 2.9 10.69 3.07 ;
      RECT 9.8 3.055 10.75 3.07 ;
      RECT 9.8 3.05 10.74 3.07 ;
      RECT 10.695 2.995 10.705 3.3 ;
      RECT 9.8 3.03 10.725 3.07 ;
      RECT 9.8 3.01 10.71 3.07 ;
      RECT 9.8 2.005 10.69 2.175 ;
      RECT 10.86 2.5 11.19 2.925 ;
      RECT 10.86 2.015 11.08 2.925 ;
      RECT 10.775 5.875 10.985 6.475 ;
      RECT 10.635 5.875 10.985 6.075 ;
      RECT 9.355 3.475 9.63 4.175 ;
      RECT 9.575 1.965 9.63 4.175 ;
      RECT 9.46 2.77 9.63 4.175 ;
      RECT 9.46 1.965 9.63 2.765 ;
      RECT 9.37 1.965 9.63 2.44 ;
      RECT 7.5 3.135 7.75 3.67 ;
      RECT 8.47 3.135 9.185 3.6 ;
      RECT 7.5 3.135 9.29 3.305 ;
      RECT 9.06 2.77 9.29 3.305 ;
      RECT 8.055 2.015 8.31 3.305 ;
      RECT 9.06 2.705 9.12 3.6 ;
      RECT 9.12 2.7 9.29 2.765 ;
      RECT 7.52 2.015 8.31 2.28 ;
      RECT 8.48 5.825 9.155 6.075 ;
      RECT 8.89 5.465 9.155 6.075 ;
      RECT 8.64 6.245 8.97 6.795 ;
      RECT 7.58 6.245 8.97 6.435 ;
      RECT 7.58 5.405 7.75 6.435 ;
      RECT 7.46 5.825 7.75 6.155 ;
      RECT 7.58 5.405 8.52 5.575 ;
      RECT 8.22 4.855 8.52 5.575 ;
      RECT 8.48 2.435 8.89 2.955 ;
      RECT 8.48 2.015 8.68 2.955 ;
      RECT 7.09 2.195 7.26 4.175 ;
      RECT 7.09 2.705 7.885 2.955 ;
      RECT 7.09 2.195 7.34 2.955 ;
      RECT 7.01 2.195 7.34 2.615 ;
      RECT 7.04 6.605 7.6 6.895 ;
      RECT 7.04 4.685 7.29 6.895 ;
      RECT 7.04 4.685 7.5 5.235 ;
      RECT 4.385 7.855 4.555 8.305 ;
      RECT 4.44 6.075 4.61 8.025 ;
      RECT 4.385 5.015 4.555 6.245 ;
      RECT 3.865 5.015 4.035 8.305 ;
      RECT 3.865 7.315 4.27 7.645 ;
      RECT 3.865 6.475 4.27 6.805 ;
      RECT 1.155 7.855 1.325 8.305 ;
      RECT 1.21 6.075 1.38 8.025 ;
      RECT 1.155 5.015 1.325 6.245 ;
      RECT 0.635 5.015 0.805 8.305 ;
      RECT 0.635 7.315 1.04 7.645 ;
      RECT 0.635 6.475 1.04 6.805 ;
      RECT 85.16 0.575 85.33 1.085 ;
      RECT 85.16 2.395 85.33 3.865 ;
      RECT 85.16 5.015 85.33 6.485 ;
      RECT 85.16 7.795 85.33 8.305 ;
      RECT 84.17 0.575 84.34 1.085 ;
      RECT 84.17 2.395 84.34 3.865 ;
      RECT 84.17 5.015 84.34 6.485 ;
      RECT 84.17 7.795 84.34 8.305 ;
      RECT 82.805 0.575 82.975 3.865 ;
      RECT 82.805 5.015 82.975 8.305 ;
      RECT 82.375 0.575 82.545 1.085 ;
      RECT 82.375 1.655 82.545 3.865 ;
      RECT 82.375 5.015 82.545 7.225 ;
      RECT 82.375 7.795 82.545 8.305 ;
      RECT 81.005 1.66 81.175 2.935 ;
      RECT 81.005 5.945 81.175 7.22 ;
      RECT 79.295 2.785 79.645 3.035 ;
      RECT 78.235 5.875 78.685 6.385 ;
      RECT 76.915 3.835 77.395 4.175 ;
      RECT 76.475 5.825 76.8 6.155 ;
      RECT 76.135 2.345 76.685 2.73 ;
      RECT 74.62 3.835 75.095 4.175 ;
      RECT 74.255 5.825 74.595 6.075 ;
      RECT 72.915 2.785 73.255 3.665 ;
      RECT 71.58 5.015 71.75 8.305 ;
      RECT 71.15 5.015 71.32 7.225 ;
      RECT 71.15 7.795 71.32 8.305 ;
      RECT 69.78 5.945 69.95 7.22 ;
      RECT 68.58 0.575 68.75 1.085 ;
      RECT 68.58 2.395 68.75 3.865 ;
      RECT 68.58 5.015 68.75 6.485 ;
      RECT 68.58 7.795 68.75 8.305 ;
      RECT 67.59 0.575 67.76 1.085 ;
      RECT 67.59 2.395 67.76 3.865 ;
      RECT 67.59 5.015 67.76 6.485 ;
      RECT 67.59 7.795 67.76 8.305 ;
      RECT 66.225 0.575 66.395 3.865 ;
      RECT 66.225 5.015 66.395 8.305 ;
      RECT 65.795 0.575 65.965 1.085 ;
      RECT 65.795 1.655 65.965 3.865 ;
      RECT 65.795 5.015 65.965 7.225 ;
      RECT 65.795 7.795 65.965 8.305 ;
      RECT 64.425 1.66 64.595 2.935 ;
      RECT 64.425 5.945 64.595 7.22 ;
      RECT 62.715 2.785 63.065 3.035 ;
      RECT 61.655 5.875 62.105 6.385 ;
      RECT 60.335 3.835 60.815 4.175 ;
      RECT 59.895 5.825 60.22 6.155 ;
      RECT 59.555 2.345 60.105 2.73 ;
      RECT 58.04 3.835 58.515 4.175 ;
      RECT 57.675 5.825 58.015 6.075 ;
      RECT 56.335 2.785 56.675 3.665 ;
      RECT 55 5.015 55.17 8.305 ;
      RECT 54.57 5.015 54.74 7.225 ;
      RECT 54.57 7.795 54.74 8.305 ;
      RECT 53.2 5.945 53.37 7.22 ;
      RECT 51.995 0.575 52.165 1.085 ;
      RECT 51.995 2.395 52.165 3.865 ;
      RECT 51.995 5.015 52.165 6.485 ;
      RECT 51.995 7.795 52.165 8.305 ;
      RECT 51.005 0.575 51.175 1.085 ;
      RECT 51.005 2.395 51.175 3.865 ;
      RECT 51.005 5.015 51.175 6.485 ;
      RECT 51.005 7.795 51.175 8.305 ;
      RECT 49.64 0.575 49.81 3.865 ;
      RECT 49.64 5.015 49.81 8.305 ;
      RECT 49.21 0.575 49.38 1.085 ;
      RECT 49.21 1.655 49.38 3.865 ;
      RECT 49.21 5.015 49.38 7.225 ;
      RECT 49.21 7.795 49.38 8.305 ;
      RECT 47.84 1.66 48.01 2.935 ;
      RECT 47.84 5.945 48.01 7.22 ;
      RECT 46.13 2.785 46.48 3.035 ;
      RECT 45.07 5.875 45.52 6.385 ;
      RECT 43.75 3.835 44.23 4.175 ;
      RECT 43.31 5.825 43.635 6.155 ;
      RECT 42.97 2.345 43.52 2.73 ;
      RECT 41.455 3.835 41.93 4.175 ;
      RECT 41.09 5.825 41.43 6.075 ;
      RECT 39.75 2.785 40.09 3.665 ;
      RECT 38.415 5.015 38.585 8.305 ;
      RECT 37.985 5.015 38.155 7.225 ;
      RECT 37.985 7.795 38.155 8.305 ;
      RECT 36.615 5.945 36.785 7.22 ;
      RECT 35.41 0.575 35.58 1.085 ;
      RECT 35.41 2.395 35.58 3.865 ;
      RECT 35.41 5.015 35.58 6.485 ;
      RECT 35.41 7.795 35.58 8.305 ;
      RECT 34.42 0.575 34.59 1.085 ;
      RECT 34.42 2.395 34.59 3.865 ;
      RECT 34.42 5.015 34.59 6.485 ;
      RECT 34.42 7.795 34.59 8.305 ;
      RECT 33.055 0.575 33.225 3.865 ;
      RECT 33.055 5.015 33.225 8.305 ;
      RECT 32.625 0.575 32.795 1.085 ;
      RECT 32.625 1.655 32.795 3.865 ;
      RECT 32.625 5.015 32.795 7.225 ;
      RECT 32.625 7.795 32.795 8.305 ;
      RECT 31.255 1.66 31.425 2.935 ;
      RECT 31.255 5.945 31.425 7.22 ;
      RECT 29.545 2.785 29.895 3.035 ;
      RECT 28.485 5.875 28.935 6.385 ;
      RECT 27.165 3.835 27.645 4.175 ;
      RECT 26.725 5.825 27.05 6.155 ;
      RECT 26.385 2.345 26.935 2.73 ;
      RECT 24.87 3.835 25.345 4.175 ;
      RECT 24.505 5.825 24.845 6.075 ;
      RECT 23.165 2.785 23.505 3.665 ;
      RECT 21.83 5.015 22 8.305 ;
      RECT 21.4 5.015 21.57 7.225 ;
      RECT 21.4 7.795 21.57 8.305 ;
      RECT 20.03 5.945 20.2 7.22 ;
      RECT 18.825 0.575 18.995 1.085 ;
      RECT 18.825 2.395 18.995 3.865 ;
      RECT 18.825 5.015 18.995 6.485 ;
      RECT 18.825 7.795 18.995 8.305 ;
      RECT 17.835 0.575 18.005 1.085 ;
      RECT 17.835 2.395 18.005 3.865 ;
      RECT 17.835 5.015 18.005 6.485 ;
      RECT 17.835 7.795 18.005 8.305 ;
      RECT 16.47 0.575 16.64 3.865 ;
      RECT 16.47 5.015 16.64 8.305 ;
      RECT 16.04 0.575 16.21 1.085 ;
      RECT 16.04 1.655 16.21 3.865 ;
      RECT 16.04 5.015 16.21 7.225 ;
      RECT 16.04 7.795 16.21 8.305 ;
      RECT 14.67 1.66 14.84 2.935 ;
      RECT 14.67 5.945 14.84 7.22 ;
      RECT 12.96 2.785 13.31 3.035 ;
      RECT 11.9 5.875 12.35 6.385 ;
      RECT 10.58 3.835 11.06 4.175 ;
      RECT 10.14 5.825 10.465 6.155 ;
      RECT 9.8 2.345 10.35 2.73 ;
      RECT 8.285 3.835 8.76 4.175 ;
      RECT 7.92 5.825 8.26 6.075 ;
      RECT 6.58 2.785 6.92 3.665 ;
      RECT 5.245 5.015 5.415 8.305 ;
      RECT 4.815 5.015 4.985 7.225 ;
      RECT 4.815 7.795 4.985 8.305 ;
      RECT 3.445 5.945 3.615 7.22 ;
      RECT 1.585 5.015 1.755 7.225 ;
      RECT 1.585 7.795 1.755 8.305 ;
      RECT 0.215 5.945 0.385 7.22 ;
  END
END sky130_osu_ring_oscillator_mpr2ca_8_b0r1

MACRO sky130_osu_ring_oscillator_mpr2ca_8_b0r2
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 2.955 0 ;
  SIZE 85.88 BY 8.88 ;
  SYMMETRY X Y R90 ;
  SITE CoreSite ;
  OBS
    LAYER met3 ;
      RECT 74.83 2.735 75.16 3.065 ;
      RECT 74.83 2.75 75.63 3.05 ;
      RECT 74.83 2.73 75.15 3.065 ;
      RECT 69.15 7.97 73.43 8.27 ;
      RECT 73.125 5.795 73.425 8.27 ;
      RECT 69.15 7.03 69.45 8.27 ;
      RECT 68.275 6.995 68.645 7.365 ;
      RECT 68.275 7.03 69.45 7.33 ;
      RECT 74.15 5.795 74.48 6.125 ;
      RECT 72.5 5.795 73.435 6.125 ;
      RECT 72.5 5.81 74.95 6.11 ;
      RECT 72.5 5.795 74.48 6.11 ;
      RECT 74.155 5.79 74.455 6.125 ;
      RECT 72.5 3.765 72.83 6.125 ;
      RECT 72.5 3.765 74.795 4.095 ;
      RECT 72.5 3.765 75.16 4.085 ;
      RECT 74.83 3.755 75.16 4.085 ;
      RECT 72.5 3.77 75.63 4.07 ;
      RECT 74.835 3.705 75.135 4.085 ;
      RECT 74.13 3.075 74.46 3.405 ;
      RECT 73.66 3.09 74.46 3.39 ;
      RECT 74.155 3.06 74.455 3.405 ;
      RECT 73.47 4.775 73.8 5.105 ;
      RECT 73.47 4.79 74.27 5.09 ;
      RECT 72.79 2.39 73.12 2.72 ;
      RECT 72.32 2.41 72.68 2.71 ;
      RECT 72.68 2.405 73.12 2.705 ;
      RECT 72.4 6.49 72.7 6.905 ;
      RECT 72.43 6.475 72.76 6.805 ;
      RECT 71.96 6.49 72.76 6.79 ;
      RECT 58.25 2.735 58.58 3.065 ;
      RECT 58.25 2.75 59.05 3.05 ;
      RECT 58.25 2.73 58.57 3.065 ;
      RECT 52.57 7.97 56.85 8.27 ;
      RECT 56.545 5.795 56.845 8.27 ;
      RECT 52.57 7.03 52.87 8.27 ;
      RECT 51.695 6.995 52.065 7.365 ;
      RECT 51.695 7.03 52.87 7.33 ;
      RECT 57.57 5.795 57.9 6.125 ;
      RECT 55.92 5.795 56.855 6.125 ;
      RECT 55.92 5.81 58.37 6.11 ;
      RECT 55.92 5.795 57.9 6.11 ;
      RECT 57.575 5.79 57.875 6.125 ;
      RECT 55.92 3.765 56.25 6.125 ;
      RECT 55.92 3.765 58.215 4.095 ;
      RECT 55.92 3.765 58.58 4.085 ;
      RECT 58.25 3.755 58.58 4.085 ;
      RECT 55.92 3.77 59.05 4.07 ;
      RECT 58.255 3.705 58.555 4.085 ;
      RECT 57.55 3.075 57.88 3.405 ;
      RECT 57.08 3.09 57.88 3.39 ;
      RECT 57.575 3.06 57.875 3.405 ;
      RECT 56.89 4.775 57.22 5.105 ;
      RECT 56.89 4.79 57.69 5.09 ;
      RECT 56.21 2.39 56.54 2.72 ;
      RECT 55.74 2.41 56.1 2.71 ;
      RECT 56.1 2.405 56.54 2.705 ;
      RECT 55.82 6.49 56.12 6.905 ;
      RECT 55.85 6.475 56.18 6.805 ;
      RECT 55.38 6.49 56.18 6.79 ;
      RECT 41.665 2.735 41.995 3.065 ;
      RECT 41.665 2.75 42.465 3.05 ;
      RECT 41.665 2.73 41.985 3.065 ;
      RECT 35.985 7.97 40.265 8.27 ;
      RECT 39.96 5.795 40.26 8.27 ;
      RECT 35.985 7.03 36.285 8.27 ;
      RECT 35.11 6.995 35.48 7.365 ;
      RECT 35.11 7.03 36.285 7.33 ;
      RECT 40.985 5.795 41.315 6.125 ;
      RECT 39.335 5.795 40.27 6.125 ;
      RECT 39.335 5.81 41.785 6.11 ;
      RECT 39.335 5.795 41.315 6.11 ;
      RECT 40.99 5.79 41.29 6.125 ;
      RECT 39.335 3.765 39.665 6.125 ;
      RECT 39.335 3.765 41.63 4.095 ;
      RECT 39.335 3.765 41.995 4.085 ;
      RECT 41.665 3.755 41.995 4.085 ;
      RECT 39.335 3.77 42.465 4.07 ;
      RECT 41.67 3.705 41.97 4.085 ;
      RECT 40.965 3.075 41.295 3.405 ;
      RECT 40.495 3.09 41.295 3.39 ;
      RECT 40.99 3.06 41.29 3.405 ;
      RECT 40.305 4.775 40.635 5.105 ;
      RECT 40.305 4.79 41.105 5.09 ;
      RECT 39.625 2.39 39.955 2.72 ;
      RECT 39.155 2.41 39.515 2.71 ;
      RECT 39.515 2.405 39.955 2.705 ;
      RECT 39.235 6.49 39.535 6.905 ;
      RECT 39.265 6.475 39.595 6.805 ;
      RECT 38.795 6.49 39.595 6.79 ;
      RECT 25.08 2.735 25.41 3.065 ;
      RECT 25.08 2.75 25.88 3.05 ;
      RECT 25.08 2.73 25.4 3.065 ;
      RECT 19.4 7.97 23.68 8.27 ;
      RECT 23.375 5.795 23.675 8.27 ;
      RECT 19.4 7.03 19.7 8.27 ;
      RECT 18.525 6.995 18.895 7.365 ;
      RECT 18.525 7.03 19.7 7.33 ;
      RECT 24.4 5.795 24.73 6.125 ;
      RECT 22.75 5.795 23.685 6.125 ;
      RECT 22.75 5.81 25.2 6.11 ;
      RECT 22.75 5.795 24.73 6.11 ;
      RECT 24.405 5.79 24.705 6.125 ;
      RECT 22.75 3.765 23.08 6.125 ;
      RECT 22.75 3.765 25.045 4.095 ;
      RECT 22.75 3.765 25.41 4.085 ;
      RECT 25.08 3.755 25.41 4.085 ;
      RECT 22.75 3.77 25.88 4.07 ;
      RECT 25.085 3.705 25.385 4.085 ;
      RECT 24.38 3.075 24.71 3.405 ;
      RECT 23.91 3.09 24.71 3.39 ;
      RECT 24.405 3.06 24.705 3.405 ;
      RECT 23.72 4.775 24.05 5.105 ;
      RECT 23.72 4.79 24.52 5.09 ;
      RECT 23.04 2.39 23.37 2.72 ;
      RECT 22.57 2.41 22.93 2.71 ;
      RECT 22.93 2.405 23.37 2.705 ;
      RECT 22.65 6.49 22.95 6.905 ;
      RECT 22.68 6.475 23.01 6.805 ;
      RECT 22.21 6.49 23.01 6.79 ;
      RECT 8.495 2.735 8.825 3.065 ;
      RECT 8.495 2.75 9.295 3.05 ;
      RECT 8.495 2.73 8.815 3.065 ;
      RECT 2.815 7.97 7.095 8.27 ;
      RECT 6.79 5.795 7.09 8.27 ;
      RECT 2.815 7.03 3.115 8.27 ;
      RECT 1.94 6.995 2.31 7.365 ;
      RECT 1.94 7.03 3.115 7.33 ;
      RECT 7.815 5.795 8.145 6.125 ;
      RECT 6.165 5.795 7.1 6.125 ;
      RECT 6.165 5.81 8.615 6.11 ;
      RECT 6.165 5.795 8.145 6.11 ;
      RECT 7.82 5.79 8.12 6.125 ;
      RECT 6.165 3.765 6.495 6.125 ;
      RECT 6.165 3.765 8.46 4.095 ;
      RECT 6.165 3.765 8.825 4.085 ;
      RECT 8.495 3.755 8.825 4.085 ;
      RECT 6.165 3.77 9.295 4.07 ;
      RECT 8.5 3.705 8.8 4.085 ;
      RECT 7.795 3.075 8.125 3.405 ;
      RECT 7.325 3.09 8.125 3.39 ;
      RECT 7.82 3.06 8.12 3.405 ;
      RECT 7.135 4.775 7.465 5.105 ;
      RECT 7.135 4.79 7.935 5.09 ;
      RECT 6.455 2.39 6.785 2.72 ;
      RECT 5.985 2.41 6.345 2.71 ;
      RECT 6.345 2.405 6.785 2.705 ;
      RECT 6.065 6.49 6.365 6.905 ;
      RECT 6.095 6.475 6.425 6.805 ;
      RECT 5.625 6.49 6.425 6.79 ;
    LAYER via2 ;
      RECT 74.895 2.8 75.095 3 ;
      RECT 74.895 3.82 75.095 4.02 ;
      RECT 74.215 5.86 74.415 6.06 ;
      RECT 74.195 3.14 74.395 3.34 ;
      RECT 73.535 4.84 73.735 5.04 ;
      RECT 73.17 5.86 73.37 6.06 ;
      RECT 72.855 2.455 73.055 2.655 ;
      RECT 72.495 6.54 72.695 6.74 ;
      RECT 68.36 7.08 68.56 7.28 ;
      RECT 58.315 2.8 58.515 3 ;
      RECT 58.315 3.82 58.515 4.02 ;
      RECT 57.635 5.86 57.835 6.06 ;
      RECT 57.615 3.14 57.815 3.34 ;
      RECT 56.955 4.84 57.155 5.04 ;
      RECT 56.59 5.86 56.79 6.06 ;
      RECT 56.275 2.455 56.475 2.655 ;
      RECT 55.915 6.54 56.115 6.74 ;
      RECT 51.78 7.08 51.98 7.28 ;
      RECT 41.73 2.8 41.93 3 ;
      RECT 41.73 3.82 41.93 4.02 ;
      RECT 41.05 5.86 41.25 6.06 ;
      RECT 41.03 3.14 41.23 3.34 ;
      RECT 40.37 4.84 40.57 5.04 ;
      RECT 40.005 5.86 40.205 6.06 ;
      RECT 39.69 2.455 39.89 2.655 ;
      RECT 39.33 6.54 39.53 6.74 ;
      RECT 35.195 7.08 35.395 7.28 ;
      RECT 25.145 2.8 25.345 3 ;
      RECT 25.145 3.82 25.345 4.02 ;
      RECT 24.465 5.86 24.665 6.06 ;
      RECT 24.445 3.14 24.645 3.34 ;
      RECT 23.785 4.84 23.985 5.04 ;
      RECT 23.42 5.86 23.62 6.06 ;
      RECT 23.105 2.455 23.305 2.655 ;
      RECT 22.745 6.54 22.945 6.74 ;
      RECT 18.61 7.08 18.81 7.28 ;
      RECT 8.56 2.8 8.76 3 ;
      RECT 8.56 3.82 8.76 4.02 ;
      RECT 7.88 5.86 8.08 6.06 ;
      RECT 7.86 3.14 8.06 3.34 ;
      RECT 7.2 4.84 7.4 5.04 ;
      RECT 6.835 5.86 7.035 6.06 ;
      RECT 6.52 2.455 6.72 2.655 ;
      RECT 6.16 6.54 6.36 6.74 ;
      RECT 2.025 7.08 2.225 7.28 ;
    LAYER met2 ;
      RECT -1.585 8.6 82.555 8.77 ;
      RECT 82.385 7.3 82.555 8.77 ;
      RECT -1.585 6.255 -1.415 8.77 ;
      RECT 82.35 7.3 82.675 7.625 ;
      RECT -1.625 6.255 -1.345 6.595 ;
      RECT 79.195 6.28 79.515 6.605 ;
      RECT 79.225 5.695 79.395 6.605 ;
      RECT 79.225 5.695 79.4 6.045 ;
      RECT 79.225 5.695 80.2 5.87 ;
      RECT 80.025 1.965 80.2 5.87 ;
      RECT 79.97 1.965 80.32 2.315 ;
      RECT 68.86 8.29 79.04 8.46 ;
      RECT 78.88 2.395 79.04 8.46 ;
      RECT 68.86 6.6 69.03 8.46 ;
      RECT 79.995 6.655 80.32 6.98 ;
      RECT 65.805 6.655 66.13 6.98 ;
      RECT 68.805 6.6 69.085 6.94 ;
      RECT 78.88 6.745 80.32 6.915 ;
      RECT 65.805 6.685 69.085 6.855 ;
      RECT 79.195 2.365 79.515 2.685 ;
      RECT 78.88 2.395 79.515 2.565 ;
      RECT 69.31 7.885 78.395 8.055 ;
      RECT 78.22 3.635 78.395 8.055 ;
      RECT 69.31 5.86 69.48 8.055 ;
      RECT 69.255 5.86 69.535 6.2 ;
      RECT 78.155 5.865 78.48 6.19 ;
      RECT 78.15 3.635 78.475 3.96 ;
      RECT 72.815 2.37 73.095 2.74 ;
      RECT 72.86 1.605 73.03 2.74 ;
      RECT 77.525 1.995 77.85 2.32 ;
      RECT 77.6 1.605 77.77 2.32 ;
      RECT 72.86 1.605 77.77 1.775 ;
      RECT 76.555 4.78 76.815 5.1 ;
      RECT 76.615 2.74 76.755 5.1 ;
      RECT 76.555 2.74 76.815 3.06 ;
      RECT 75.535 5.8 75.795 6.12 ;
      RECT 74.915 5.89 75.795 6.03 ;
      RECT 74.915 3.735 75.055 6.03 ;
      RECT 74.855 3.735 75.135 4.105 ;
      RECT 74.175 5.775 74.455 6.145 ;
      RECT 74.235 3.85 74.375 6.145 ;
      RECT 74.235 3.85 74.715 3.99 ;
      RECT 74.575 2.06 74.715 3.99 ;
      RECT 74.515 2.06 74.775 2.38 ;
      RECT 73.495 4.755 73.775 5.125 ;
      RECT 73.555 2.4 73.695 5.125 ;
      RECT 73.495 2.4 73.755 2.72 ;
      RECT 73.13 5.775 73.41 6.145 ;
      RECT 73.13 5.8 73.415 6.12 ;
      RECT 68.275 6.995 68.645 7.365 ;
      RECT 68.275 6.995 68.65 7.005 ;
      RECT 62.615 6.28 62.935 6.605 ;
      RECT 62.645 5.695 62.815 6.605 ;
      RECT 62.645 5.695 62.82 6.045 ;
      RECT 62.645 5.695 63.62 5.87 ;
      RECT 63.445 1.965 63.62 5.87 ;
      RECT 63.39 1.965 63.74 2.315 ;
      RECT 52.28 8.29 62.46 8.46 ;
      RECT 62.3 2.395 62.46 8.46 ;
      RECT 52.28 6.6 52.45 8.46 ;
      RECT 63.415 6.655 63.74 6.98 ;
      RECT 49.22 6.655 49.545 6.98 ;
      RECT 52.225 6.6 52.505 6.94 ;
      RECT 62.3 6.745 63.74 6.915 ;
      RECT 49.22 6.685 52.505 6.855 ;
      RECT 62.615 2.365 62.935 2.685 ;
      RECT 62.3 2.395 62.935 2.565 ;
      RECT 52.73 7.885 61.815 8.055 ;
      RECT 61.64 3.635 61.815 8.055 ;
      RECT 52.73 5.86 52.9 8.055 ;
      RECT 52.675 5.86 52.955 6.2 ;
      RECT 61.575 5.865 61.9 6.19 ;
      RECT 61.57 3.635 61.895 3.96 ;
      RECT 56.235 2.37 56.515 2.74 ;
      RECT 56.28 1.605 56.45 2.74 ;
      RECT 60.945 1.995 61.27 2.32 ;
      RECT 61.02 1.605 61.19 2.32 ;
      RECT 56.28 1.605 61.19 1.775 ;
      RECT 59.975 4.78 60.235 5.1 ;
      RECT 60.035 2.74 60.175 5.1 ;
      RECT 59.975 2.74 60.235 3.06 ;
      RECT 58.955 5.8 59.215 6.12 ;
      RECT 58.335 5.89 59.215 6.03 ;
      RECT 58.335 3.735 58.475 6.03 ;
      RECT 58.275 3.735 58.555 4.105 ;
      RECT 57.595 5.775 57.875 6.145 ;
      RECT 57.655 3.85 57.795 6.145 ;
      RECT 57.655 3.85 58.135 3.99 ;
      RECT 57.995 2.06 58.135 3.99 ;
      RECT 57.935 2.06 58.195 2.38 ;
      RECT 56.915 4.755 57.195 5.125 ;
      RECT 56.975 2.4 57.115 5.125 ;
      RECT 56.915 2.4 57.175 2.72 ;
      RECT 56.55 5.775 56.83 6.145 ;
      RECT 56.55 5.8 56.835 6.12 ;
      RECT 46.03 6.28 46.35 6.605 ;
      RECT 46.06 5.695 46.23 6.605 ;
      RECT 46.06 5.695 46.235 6.045 ;
      RECT 46.06 5.695 47.035 5.87 ;
      RECT 46.86 1.965 47.035 5.87 ;
      RECT 46.805 1.965 47.155 2.315 ;
      RECT 35.695 8.29 45.875 8.46 ;
      RECT 45.715 2.395 45.875 8.46 ;
      RECT 35.695 6.6 35.865 8.46 ;
      RECT 46.83 6.655 47.155 6.98 ;
      RECT 32.635 6.655 32.96 6.98 ;
      RECT 35.64 6.6 35.92 6.94 ;
      RECT 45.715 6.745 47.155 6.915 ;
      RECT 32.635 6.685 35.92 6.855 ;
      RECT 46.03 2.365 46.35 2.685 ;
      RECT 45.715 2.395 46.35 2.565 ;
      RECT 36.145 7.885 45.23 8.055 ;
      RECT 45.055 3.635 45.23 8.055 ;
      RECT 36.145 5.86 36.315 8.055 ;
      RECT 36.09 5.86 36.37 6.2 ;
      RECT 44.99 5.865 45.315 6.19 ;
      RECT 44.985 3.635 45.31 3.96 ;
      RECT 39.65 2.37 39.93 2.74 ;
      RECT 39.695 1.605 39.865 2.74 ;
      RECT 44.36 1.995 44.685 2.32 ;
      RECT 44.435 1.605 44.605 2.32 ;
      RECT 39.695 1.605 44.605 1.775 ;
      RECT 43.39 4.78 43.65 5.1 ;
      RECT 43.45 2.74 43.59 5.1 ;
      RECT 43.39 2.74 43.65 3.06 ;
      RECT 42.37 5.8 42.63 6.12 ;
      RECT 41.75 5.89 42.63 6.03 ;
      RECT 41.75 3.735 41.89 6.03 ;
      RECT 41.69 3.735 41.97 4.105 ;
      RECT 41.01 5.775 41.29 6.145 ;
      RECT 41.07 3.85 41.21 6.145 ;
      RECT 41.07 3.85 41.55 3.99 ;
      RECT 41.41 2.06 41.55 3.99 ;
      RECT 41.35 2.06 41.61 2.38 ;
      RECT 40.33 4.755 40.61 5.125 ;
      RECT 40.39 2.4 40.53 5.125 ;
      RECT 40.33 2.4 40.59 2.72 ;
      RECT 39.965 5.775 40.245 6.145 ;
      RECT 39.965 5.8 40.25 6.12 ;
      RECT 29.445 6.28 29.765 6.605 ;
      RECT 29.475 5.695 29.645 6.605 ;
      RECT 29.475 5.695 29.65 6.045 ;
      RECT 29.475 5.695 30.45 5.87 ;
      RECT 30.275 1.965 30.45 5.87 ;
      RECT 30.22 1.965 30.57 2.315 ;
      RECT 19.11 8.29 29.29 8.46 ;
      RECT 29.13 2.395 29.29 8.46 ;
      RECT 19.11 6.6 19.28 8.46 ;
      RECT 30.245 6.655 30.57 6.98 ;
      RECT 16.05 6.655 16.375 6.98 ;
      RECT 19.055 6.6 19.335 6.94 ;
      RECT 29.13 6.745 30.57 6.915 ;
      RECT 16.05 6.685 19.335 6.855 ;
      RECT 29.445 2.365 29.765 2.685 ;
      RECT 29.13 2.395 29.765 2.565 ;
      RECT 19.56 7.885 28.645 8.055 ;
      RECT 28.47 3.635 28.645 8.055 ;
      RECT 19.56 5.86 19.73 8.055 ;
      RECT 19.505 5.86 19.785 6.2 ;
      RECT 28.405 5.865 28.73 6.19 ;
      RECT 28.4 3.635 28.725 3.96 ;
      RECT 23.065 2.37 23.345 2.74 ;
      RECT 23.11 1.605 23.28 2.74 ;
      RECT 27.775 1.995 28.1 2.32 ;
      RECT 27.85 1.605 28.02 2.32 ;
      RECT 23.11 1.605 28.02 1.775 ;
      RECT 26.805 4.78 27.065 5.1 ;
      RECT 26.865 2.74 27.005 5.1 ;
      RECT 26.805 2.74 27.065 3.06 ;
      RECT 25.785 5.8 26.045 6.12 ;
      RECT 25.165 5.89 26.045 6.03 ;
      RECT 25.165 3.735 25.305 6.03 ;
      RECT 25.105 3.735 25.385 4.105 ;
      RECT 24.425 5.775 24.705 6.145 ;
      RECT 24.485 3.85 24.625 6.145 ;
      RECT 24.485 3.85 24.965 3.99 ;
      RECT 24.825 2.06 24.965 3.99 ;
      RECT 24.765 2.06 25.025 2.38 ;
      RECT 23.745 4.755 24.025 5.125 ;
      RECT 23.805 2.4 23.945 5.125 ;
      RECT 23.745 2.4 24.005 2.72 ;
      RECT 23.38 5.775 23.66 6.145 ;
      RECT 23.38 5.8 23.665 6.12 ;
      RECT 12.86 6.28 13.18 6.605 ;
      RECT 12.89 5.695 13.06 6.605 ;
      RECT 12.89 5.695 13.065 6.045 ;
      RECT 12.89 5.695 13.865 5.87 ;
      RECT 13.69 1.965 13.865 5.87 ;
      RECT 13.635 1.965 13.985 2.315 ;
      RECT 2.525 8.29 12.705 8.46 ;
      RECT 12.545 2.395 12.705 8.46 ;
      RECT 2.525 6.6 2.695 8.46 ;
      RECT -1.24 6.995 -0.96 7.335 ;
      RECT -1.24 7.06 -0.05 7.23 ;
      RECT -0.22 6.685 -0.05 7.23 ;
      RECT 13.66 6.655 13.985 6.98 ;
      RECT 2.47 6.6 2.75 6.94 ;
      RECT 12.545 6.745 13.985 6.915 ;
      RECT -0.22 6.685 2.75 6.855 ;
      RECT 12.86 2.365 13.18 2.685 ;
      RECT 12.545 2.395 13.18 2.565 ;
      RECT 2.975 7.885 12.06 8.055 ;
      RECT 11.885 3.635 12.06 8.055 ;
      RECT 2.975 5.86 3.145 8.055 ;
      RECT 2.92 5.86 3.2 6.2 ;
      RECT 11.82 5.865 12.145 6.19 ;
      RECT 11.815 3.635 12.14 3.96 ;
      RECT 6.48 2.37 6.76 2.74 ;
      RECT 6.525 1.605 6.695 2.74 ;
      RECT 11.19 1.995 11.515 2.32 ;
      RECT 11.265 1.605 11.435 2.32 ;
      RECT 6.525 1.605 11.435 1.775 ;
      RECT 10.22 4.78 10.48 5.1 ;
      RECT 10.28 2.74 10.42 5.1 ;
      RECT 10.22 2.74 10.48 3.06 ;
      RECT 9.2 5.8 9.46 6.12 ;
      RECT 8.58 5.89 9.46 6.03 ;
      RECT 8.58 3.735 8.72 6.03 ;
      RECT 8.52 3.735 8.8 4.105 ;
      RECT 7.84 5.775 8.12 6.145 ;
      RECT 7.9 3.85 8.04 6.145 ;
      RECT 7.9 3.85 8.38 3.99 ;
      RECT 8.24 2.06 8.38 3.99 ;
      RECT 8.18 2.06 8.44 2.38 ;
      RECT 7.16 4.755 7.44 5.125 ;
      RECT 7.22 2.4 7.36 5.125 ;
      RECT 7.16 2.4 7.42 2.72 ;
      RECT 6.795 5.775 7.075 6.145 ;
      RECT 6.795 5.8 7.08 6.12 ;
      RECT 74.855 2.715 75.135 3.085 ;
      RECT 74.155 3.055 74.435 3.425 ;
      RECT 72.455 6.455 72.735 6.825 ;
      RECT 58.275 2.715 58.555 3.085 ;
      RECT 57.575 3.055 57.855 3.425 ;
      RECT 55.875 6.455 56.155 6.825 ;
      RECT 51.695 6.995 52.065 7.365 ;
      RECT 41.69 2.715 41.97 3.085 ;
      RECT 40.99 3.055 41.27 3.425 ;
      RECT 39.29 6.455 39.57 6.825 ;
      RECT 35.11 6.995 35.48 7.365 ;
      RECT 25.105 2.715 25.385 3.085 ;
      RECT 24.405 3.055 24.685 3.425 ;
      RECT 22.705 6.455 22.985 6.825 ;
      RECT 18.525 6.995 18.895 7.365 ;
      RECT 8.52 2.715 8.8 3.085 ;
      RECT 7.82 3.055 8.1 3.425 ;
      RECT 6.12 6.455 6.4 6.825 ;
      RECT 1.94 6.995 2.31 7.365 ;
    LAYER via1 ;
      RECT 82.44 7.385 82.59 7.535 ;
      RECT 80.085 6.74 80.235 6.89 ;
      RECT 80.07 2.065 80.22 2.215 ;
      RECT 79.28 2.45 79.43 2.6 ;
      RECT 79.28 6.37 79.43 6.52 ;
      RECT 78.245 5.95 78.395 6.1 ;
      RECT 78.24 3.72 78.39 3.87 ;
      RECT 77.615 2.08 77.765 2.23 ;
      RECT 76.61 2.825 76.76 2.975 ;
      RECT 76.61 4.865 76.76 5.015 ;
      RECT 75.59 5.885 75.74 6.035 ;
      RECT 74.91 2.825 75.06 2.975 ;
      RECT 74.91 3.845 75.06 3.995 ;
      RECT 74.57 2.145 74.72 2.295 ;
      RECT 74.23 3.165 74.38 3.315 ;
      RECT 74.23 5.885 74.38 6.035 ;
      RECT 73.55 2.485 73.7 2.635 ;
      RECT 73.55 4.865 73.7 5.015 ;
      RECT 73.21 5.885 73.36 6.035 ;
      RECT 72.87 2.48 73.02 2.63 ;
      RECT 72.53 6.565 72.68 6.715 ;
      RECT 69.32 5.955 69.47 6.105 ;
      RECT 68.87 6.695 69.02 6.845 ;
      RECT 68.385 7.105 68.535 7.255 ;
      RECT 65.895 6.74 66.045 6.89 ;
      RECT 63.505 6.74 63.655 6.89 ;
      RECT 63.49 2.065 63.64 2.215 ;
      RECT 62.7 2.45 62.85 2.6 ;
      RECT 62.7 6.37 62.85 6.52 ;
      RECT 61.665 5.95 61.815 6.1 ;
      RECT 61.66 3.72 61.81 3.87 ;
      RECT 61.035 2.08 61.185 2.23 ;
      RECT 60.03 2.825 60.18 2.975 ;
      RECT 60.03 4.865 60.18 5.015 ;
      RECT 59.01 5.885 59.16 6.035 ;
      RECT 58.33 2.825 58.48 2.975 ;
      RECT 58.33 3.845 58.48 3.995 ;
      RECT 57.99 2.145 58.14 2.295 ;
      RECT 57.65 3.165 57.8 3.315 ;
      RECT 57.65 5.885 57.8 6.035 ;
      RECT 56.97 2.485 57.12 2.635 ;
      RECT 56.97 4.865 57.12 5.015 ;
      RECT 56.63 5.885 56.78 6.035 ;
      RECT 56.29 2.48 56.44 2.63 ;
      RECT 55.95 6.565 56.1 6.715 ;
      RECT 52.74 5.955 52.89 6.105 ;
      RECT 52.29 6.695 52.44 6.845 ;
      RECT 51.805 7.105 51.955 7.255 ;
      RECT 49.31 6.74 49.46 6.89 ;
      RECT 46.92 6.74 47.07 6.89 ;
      RECT 46.905 2.065 47.055 2.215 ;
      RECT 46.115 2.45 46.265 2.6 ;
      RECT 46.115 6.37 46.265 6.52 ;
      RECT 45.08 5.95 45.23 6.1 ;
      RECT 45.075 3.72 45.225 3.87 ;
      RECT 44.45 2.08 44.6 2.23 ;
      RECT 43.445 2.825 43.595 2.975 ;
      RECT 43.445 4.865 43.595 5.015 ;
      RECT 42.425 5.885 42.575 6.035 ;
      RECT 41.745 2.825 41.895 2.975 ;
      RECT 41.745 3.845 41.895 3.995 ;
      RECT 41.405 2.145 41.555 2.295 ;
      RECT 41.065 3.165 41.215 3.315 ;
      RECT 41.065 5.885 41.215 6.035 ;
      RECT 40.385 2.485 40.535 2.635 ;
      RECT 40.385 4.865 40.535 5.015 ;
      RECT 40.045 5.885 40.195 6.035 ;
      RECT 39.705 2.48 39.855 2.63 ;
      RECT 39.365 6.565 39.515 6.715 ;
      RECT 36.155 5.955 36.305 6.105 ;
      RECT 35.705 6.695 35.855 6.845 ;
      RECT 35.22 7.105 35.37 7.255 ;
      RECT 32.725 6.74 32.875 6.89 ;
      RECT 30.335 6.74 30.485 6.89 ;
      RECT 30.32 2.065 30.47 2.215 ;
      RECT 29.53 2.45 29.68 2.6 ;
      RECT 29.53 6.37 29.68 6.52 ;
      RECT 28.495 5.95 28.645 6.1 ;
      RECT 28.49 3.72 28.64 3.87 ;
      RECT 27.865 2.08 28.015 2.23 ;
      RECT 26.86 2.825 27.01 2.975 ;
      RECT 26.86 4.865 27.01 5.015 ;
      RECT 25.84 5.885 25.99 6.035 ;
      RECT 25.16 2.825 25.31 2.975 ;
      RECT 25.16 3.845 25.31 3.995 ;
      RECT 24.82 2.145 24.97 2.295 ;
      RECT 24.48 3.165 24.63 3.315 ;
      RECT 24.48 5.885 24.63 6.035 ;
      RECT 23.8 2.485 23.95 2.635 ;
      RECT 23.8 4.865 23.95 5.015 ;
      RECT 23.46 5.885 23.61 6.035 ;
      RECT 23.12 2.48 23.27 2.63 ;
      RECT 22.78 6.565 22.93 6.715 ;
      RECT 19.57 5.955 19.72 6.105 ;
      RECT 19.12 6.695 19.27 6.845 ;
      RECT 18.635 7.105 18.785 7.255 ;
      RECT 16.14 6.74 16.29 6.89 ;
      RECT 13.75 6.74 13.9 6.89 ;
      RECT 13.735 2.065 13.885 2.215 ;
      RECT 12.945 2.45 13.095 2.6 ;
      RECT 12.945 6.37 13.095 6.52 ;
      RECT 11.91 5.95 12.06 6.1 ;
      RECT 11.905 3.72 12.055 3.87 ;
      RECT 11.28 2.08 11.43 2.23 ;
      RECT 10.275 2.825 10.425 2.975 ;
      RECT 10.275 4.865 10.425 5.015 ;
      RECT 9.255 5.885 9.405 6.035 ;
      RECT 8.575 2.825 8.725 2.975 ;
      RECT 8.575 3.845 8.725 3.995 ;
      RECT 8.235 2.145 8.385 2.295 ;
      RECT 7.895 3.165 8.045 3.315 ;
      RECT 7.895 5.885 8.045 6.035 ;
      RECT 7.215 2.485 7.365 2.635 ;
      RECT 7.215 4.865 7.365 5.015 ;
      RECT 6.875 5.885 7.025 6.035 ;
      RECT 6.535 2.48 6.685 2.63 ;
      RECT 6.195 6.565 6.345 6.715 ;
      RECT 2.985 5.955 3.135 6.105 ;
      RECT 2.535 6.695 2.685 6.845 ;
      RECT 2.05 7.105 2.2 7.255 ;
      RECT -1.175 7.09 -1.025 7.24 ;
      RECT -1.56 6.35 -1.41 6.5 ;
    LAYER met1 ;
      RECT 70.055 0 76.955 1.95 ;
      RECT 53.475 0 60.375 1.95 ;
      RECT 36.89 0 43.79 1.95 ;
      RECT 20.305 0 27.205 1.95 ;
      RECT 3.72 0 10.62 1.95 ;
      RECT 70.055 0 77.145 1.795 ;
      RECT 53.475 0 60.565 1.795 ;
      RECT 36.89 0 43.98 1.795 ;
      RECT 20.305 0 27.395 1.795 ;
      RECT 3.72 0 10.81 1.795 ;
      RECT 69.8 0 77.145 1.655 ;
      RECT 53.22 0 60.565 1.655 ;
      RECT 36.635 0 43.98 1.655 ;
      RECT 20.05 0 27.395 1.655 ;
      RECT 3.465 0 10.81 1.655 ;
      RECT -2.955 0 82.925 0.305 ;
      RECT 76.985 4.15 82.925 4.745 ;
      RECT 77.445 4.135 82.925 4.745 ;
      RECT 66.82 4.13 69.57 4.745 ;
      RECT 60.405 4.15 66.345 4.745 ;
      RECT 50.24 4.13 52.99 4.745 ;
      RECT 43.82 4.15 49.76 4.745 ;
      RECT 33.655 4.13 36.405 4.745 ;
      RECT 27.235 4.15 33.175 4.745 ;
      RECT 17.07 4.13 19.82 4.745 ;
      RECT 10.65 4.15 16.59 4.745 ;
      RECT 0.485 4.13 3.235 4.745 ;
      RECT -2.955 4.13 0.005 4.745 ;
      RECT 66.34 4.13 69.915 4.74 ;
      RECT 49.76 4.13 53.335 4.74 ;
      RECT 33.175 4.13 36.75 4.74 ;
      RECT 16.59 4.13 20.165 4.74 ;
      RECT -2.955 4.13 3.58 4.74 ;
      RECT -2.955 4.19 82.925 4.67 ;
      RECT 76.855 4.15 82.925 4.67 ;
      RECT 60.275 4.15 69.915 4.67 ;
      RECT 43.69 4.15 53.335 4.67 ;
      RECT 27.105 4.15 36.75 4.67 ;
      RECT 10.52 4.15 20.165 4.67 ;
      RECT 60.865 4.135 69.915 4.74 ;
      RECT 44.28 4.135 53.335 4.74 ;
      RECT 27.695 4.135 36.75 4.74 ;
      RECT 11.11 4.135 20.165 4.74 ;
      RECT -2.955 8.575 82.925 8.88 ;
      RECT 69.76 7.18 76.96 8.88 ;
      RECT 67.78 6.315 67.95 8.88 ;
      RECT 53.18 7.18 60.38 8.88 ;
      RECT 51.2 6.315 51.37 8.88 ;
      RECT 36.595 7.18 43.795 8.88 ;
      RECT 34.615 6.315 34.785 8.88 ;
      RECT 20.01 7.18 27.21 8.88 ;
      RECT 18.03 6.315 18.2 8.88 ;
      RECT 3.425 7.18 10.625 8.88 ;
      RECT 1.445 6.315 1.615 8.88 ;
      RECT 70.055 6.91 76.955 8.88 ;
      RECT 53.475 6.91 60.375 8.88 ;
      RECT 36.89 6.91 43.79 8.88 ;
      RECT 20.305 6.91 27.205 8.88 ;
      RECT 3.72 6.91 10.62 8.88 ;
      RECT 72.48 6.51 72.735 8.88 ;
      RECT 55.9 6.51 56.155 8.88 ;
      RECT 39.315 6.51 39.57 8.88 ;
      RECT 22.73 6.51 22.985 8.88 ;
      RECT 6.145 6.51 6.4 8.88 ;
      RECT 72.445 6.51 72.765 6.77 ;
      RECT 55.865 6.51 56.185 6.77 ;
      RECT 39.28 6.51 39.6 6.77 ;
      RECT 22.695 6.51 23.015 6.77 ;
      RECT 6.11 6.51 6.43 6.77 ;
      RECT 71.515 6.57 73.865 6.71 ;
      RECT 73.725 5.845 73.865 6.71 ;
      RECT 54.935 6.57 57.285 6.71 ;
      RECT 57.145 5.845 57.285 6.71 ;
      RECT 38.35 6.57 40.7 6.71 ;
      RECT 40.56 5.845 40.7 6.71 ;
      RECT 21.765 6.57 24.115 6.71 ;
      RECT 23.975 5.845 24.115 6.71 ;
      RECT 5.18 6.57 7.53 6.71 ;
      RECT 7.39 5.845 7.53 6.71 ;
      RECT 71.515 5.845 71.655 6.71 ;
      RECT 54.935 5.845 55.075 6.71 ;
      RECT 38.35 5.845 38.49 6.71 ;
      RECT 21.765 5.845 21.905 6.71 ;
      RECT 5.18 5.845 5.32 6.71 ;
      RECT 67.94 6.285 68.23 6.515 ;
      RECT 51.36 6.285 51.65 6.515 ;
      RECT 34.775 6.285 35.065 6.515 ;
      RECT 18.19 6.285 18.48 6.515 ;
      RECT 1.605 6.285 1.895 6.515 ;
      RECT 67.77 6.315 68.23 6.485 ;
      RECT 51.19 6.315 51.65 6.485 ;
      RECT 34.605 6.315 35.065 6.485 ;
      RECT 18.02 6.315 18.48 6.485 ;
      RECT 1.435 6.315 1.895 6.485 ;
      RECT 73.65 5.845 73.94 6.075 ;
      RECT 71.44 5.845 71.73 6.075 ;
      RECT 57.07 5.845 57.36 6.075 ;
      RECT 54.86 5.845 55.15 6.075 ;
      RECT 40.485 5.845 40.775 6.075 ;
      RECT 38.275 5.845 38.565 6.075 ;
      RECT 23.9 5.845 24.19 6.075 ;
      RECT 21.69 5.845 21.98 6.075 ;
      RECT 7.315 5.845 7.605 6.075 ;
      RECT 5.105 5.845 5.395 6.075 ;
      RECT 82.325 7.765 82.615 7.995 ;
      RECT 82.385 6.285 82.555 7.995 ;
      RECT 82.35 7.3 82.675 7.625 ;
      RECT 82.325 6.285 82.615 6.515 ;
      RECT 82.325 2.365 82.615 2.595 ;
      RECT 82.385 0.885 82.555 2.595 ;
      RECT 82.325 0.885 82.615 1.115 ;
      RECT 81.915 2.735 82.245 2.965 ;
      RECT 81.915 2.765 82.415 2.935 ;
      RECT 81.915 2.395 82.105 2.965 ;
      RECT 81.335 2.365 81.625 2.595 ;
      RECT 81.335 2.395 82.105 2.565 ;
      RECT 81.395 0.885 81.565 2.595 ;
      RECT 81.335 0.885 81.625 1.115 ;
      RECT 81.335 7.765 81.625 7.995 ;
      RECT 81.395 6.285 81.565 7.995 ;
      RECT 81.335 6.285 81.625 6.515 ;
      RECT 81.335 6.325 82.185 6.485 ;
      RECT 82.015 5.915 82.185 6.485 ;
      RECT 81.335 6.32 81.725 6.485 ;
      RECT 81.955 5.915 82.245 6.145 ;
      RECT 81.955 5.945 82.415 6.115 ;
      RECT 80.965 2.735 81.255 2.965 ;
      RECT 80.965 2.765 81.425 2.935 ;
      RECT 81.025 1.655 81.19 2.965 ;
      RECT 79.54 1.625 79.83 1.855 ;
      RECT 79.54 1.655 81.19 1.825 ;
      RECT 79.6 0.885 79.77 1.855 ;
      RECT 79.54 0.885 79.83 1.115 ;
      RECT 79.54 7.765 79.83 7.995 ;
      RECT 79.6 7.025 79.77 7.995 ;
      RECT 79.6 7.12 81.19 7.29 ;
      RECT 81.02 5.915 81.19 7.29 ;
      RECT 79.54 7.025 79.83 7.255 ;
      RECT 80.965 5.915 81.255 6.145 ;
      RECT 80.965 5.945 81.425 6.115 ;
      RECT 77.525 1.995 77.85 2.32 ;
      RECT 79.97 1.965 80.32 2.315 ;
      RECT 77.525 2.025 80.32 2.195 ;
      RECT 79.995 6.655 80.32 6.98 ;
      RECT 79.97 6.655 80.32 6.885 ;
      RECT 79.8 6.685 80.32 6.855 ;
      RECT 79.195 2.365 79.515 2.685 ;
      RECT 79.165 2.365 79.515 2.595 ;
      RECT 78.88 2.395 79.515 2.565 ;
      RECT 79.195 6.28 79.515 6.605 ;
      RECT 79.165 6.285 79.515 6.515 ;
      RECT 78.995 6.315 79.515 6.485 ;
      RECT 78.15 3.635 78.475 3.96 ;
      RECT 78.225 2.735 78.405 3.96 ;
      RECT 78.17 2.735 78.46 2.965 ;
      RECT 78.17 2.765 78.63 2.935 ;
      RECT 78.155 5.865 78.48 6.19 ;
      RECT 78.155 5.945 78.63 6.115 ;
      RECT 76.525 2.77 76.845 3.03 ;
      RECT 76.25 2.83 76.845 2.97 ;
      RECT 74.145 3.11 74.465 3.37 ;
      RECT 76.12 3.125 76.41 3.355 ;
      RECT 74.145 3.17 76.41 3.31 ;
      RECT 75.505 5.83 75.825 6.09 ;
      RECT 75.505 5.89 76.1 6.03 ;
      RECT 74.825 2.77 75.145 3.03 ;
      RECT 70.085 2.785 70.375 3.015 ;
      RECT 70.085 2.83 75.145 2.97 ;
      RECT 74.915 2.49 75.055 3.03 ;
      RECT 74.915 2.49 75.395 2.63 ;
      RECT 75.255 2.105 75.395 2.63 ;
      RECT 75.18 2.105 75.47 2.335 ;
      RECT 74.825 3.79 75.145 4.05 ;
      RECT 74.16 3.805 74.45 4.035 ;
      RECT 71.95 3.805 72.24 4.035 ;
      RECT 71.95 3.85 75.145 3.99 ;
      RECT 73.125 5.83 73.445 6.09 ;
      RECT 74.84 5.845 75.13 6.075 ;
      RECT 72.46 5.845 72.75 6.075 ;
      RECT 72.46 5.89 73.445 6.03 ;
      RECT 74.915 5.55 75.055 6.075 ;
      RECT 73.215 5.55 73.355 6.09 ;
      RECT 73.215 5.55 75.055 5.69 ;
      RECT 72.12 2.445 72.41 2.675 ;
      RECT 72.195 2.15 72.335 2.675 ;
      RECT 74.485 2.09 74.805 2.35 ;
      RECT 74.385 2.105 74.805 2.335 ;
      RECT 72.195 2.15 74.805 2.29 ;
      RECT 73.465 2.43 73.785 2.69 ;
      RECT 73.465 2.49 74.06 2.63 ;
      RECT 73.465 4.81 73.785 5.07 ;
      RECT 70.76 4.825 71.05 5.055 ;
      RECT 70.76 4.87 73.785 5.01 ;
      RECT 72.79 2.39 73.12 2.72 ;
      RECT 72.785 2.425 73.12 2.685 ;
      RECT 73.135 2.445 73.25 2.675 ;
      RECT 72.785 2.44 73.135 2.67 ;
      RECT 72.785 2.49 73.265 2.63 ;
      RECT 72.67 2.49 72.68 2.63 ;
      RECT 72.68 2.485 73.25 2.625 ;
      RECT 69.225 5.89 69.565 6.17 ;
      RECT 66.945 5.915 67.235 6.145 ;
      RECT 66.945 5.945 69.565 6.115 ;
      RECT 68.775 6.63 69.115 6.91 ;
      RECT 68.745 6.655 69.115 6.885 ;
      RECT 68.575 6.685 69.115 6.855 ;
      RECT 68.315 7.765 68.605 7.995 ;
      RECT 68.375 6.995 68.545 7.995 ;
      RECT 68.275 6.995 68.645 7.365 ;
      RECT 65.745 7.765 66.035 7.995 ;
      RECT 65.805 6.285 65.975 7.995 ;
      RECT 65.805 6.655 66.13 6.98 ;
      RECT 65.745 6.285 66.035 6.515 ;
      RECT 65.745 2.365 66.035 2.595 ;
      RECT 65.805 0.885 65.975 2.595 ;
      RECT 65.745 0.885 66.035 1.115 ;
      RECT 65.335 2.735 65.665 2.965 ;
      RECT 65.335 2.765 65.835 2.935 ;
      RECT 65.335 2.395 65.525 2.965 ;
      RECT 64.755 2.365 65.045 2.595 ;
      RECT 64.755 2.395 65.525 2.565 ;
      RECT 64.815 0.885 64.985 2.595 ;
      RECT 64.755 0.885 65.045 1.115 ;
      RECT 64.755 7.765 65.045 7.995 ;
      RECT 64.815 6.285 64.985 7.995 ;
      RECT 64.755 6.285 65.045 6.515 ;
      RECT 64.755 6.325 65.605 6.485 ;
      RECT 65.435 5.915 65.605 6.485 ;
      RECT 64.755 6.32 65.145 6.485 ;
      RECT 65.375 5.915 65.665 6.145 ;
      RECT 65.375 5.945 65.835 6.115 ;
      RECT 64.385 2.735 64.675 2.965 ;
      RECT 64.385 2.765 64.845 2.935 ;
      RECT 64.445 1.655 64.61 2.965 ;
      RECT 62.96 1.625 63.25 1.855 ;
      RECT 62.96 1.655 64.61 1.825 ;
      RECT 63.02 0.885 63.19 1.855 ;
      RECT 62.96 0.885 63.25 1.115 ;
      RECT 62.96 7.765 63.25 7.995 ;
      RECT 63.02 7.025 63.19 7.995 ;
      RECT 63.02 7.12 64.61 7.29 ;
      RECT 64.44 5.915 64.61 7.29 ;
      RECT 62.96 7.025 63.25 7.255 ;
      RECT 64.385 5.915 64.675 6.145 ;
      RECT 64.385 5.945 64.845 6.115 ;
      RECT 60.945 1.995 61.27 2.32 ;
      RECT 63.39 1.965 63.74 2.315 ;
      RECT 60.945 2.025 63.74 2.195 ;
      RECT 63.415 6.655 63.74 6.98 ;
      RECT 63.39 6.655 63.74 6.885 ;
      RECT 63.22 6.685 63.74 6.855 ;
      RECT 62.615 2.365 62.935 2.685 ;
      RECT 62.585 2.365 62.935 2.595 ;
      RECT 62.3 2.395 62.935 2.565 ;
      RECT 62.615 6.28 62.935 6.605 ;
      RECT 62.585 6.285 62.935 6.515 ;
      RECT 62.415 6.315 62.935 6.485 ;
      RECT 61.57 3.635 61.895 3.96 ;
      RECT 61.645 2.735 61.825 3.96 ;
      RECT 61.59 2.735 61.88 2.965 ;
      RECT 61.59 2.765 62.05 2.935 ;
      RECT 61.575 5.865 61.9 6.19 ;
      RECT 61.575 5.945 62.05 6.115 ;
      RECT 59.945 2.77 60.265 3.03 ;
      RECT 59.67 2.83 60.265 2.97 ;
      RECT 57.565 3.11 57.885 3.37 ;
      RECT 59.54 3.125 59.83 3.355 ;
      RECT 57.565 3.17 59.83 3.31 ;
      RECT 58.925 5.83 59.245 6.09 ;
      RECT 58.925 5.89 59.52 6.03 ;
      RECT 58.245 2.77 58.565 3.03 ;
      RECT 53.505 2.785 53.795 3.015 ;
      RECT 53.505 2.83 58.565 2.97 ;
      RECT 58.335 2.49 58.475 3.03 ;
      RECT 58.335 2.49 58.815 2.63 ;
      RECT 58.675 2.105 58.815 2.63 ;
      RECT 58.6 2.105 58.89 2.335 ;
      RECT 58.245 3.79 58.565 4.05 ;
      RECT 57.58 3.805 57.87 4.035 ;
      RECT 55.37 3.805 55.66 4.035 ;
      RECT 55.37 3.85 58.565 3.99 ;
      RECT 56.545 5.83 56.865 6.09 ;
      RECT 58.26 5.845 58.55 6.075 ;
      RECT 55.88 5.845 56.17 6.075 ;
      RECT 55.88 5.89 56.865 6.03 ;
      RECT 58.335 5.55 58.475 6.075 ;
      RECT 56.635 5.55 56.775 6.09 ;
      RECT 56.635 5.55 58.475 5.69 ;
      RECT 55.54 2.445 55.83 2.675 ;
      RECT 55.615 2.15 55.755 2.675 ;
      RECT 57.905 2.09 58.225 2.35 ;
      RECT 57.805 2.105 58.225 2.335 ;
      RECT 55.615 2.15 58.225 2.29 ;
      RECT 56.885 2.43 57.205 2.69 ;
      RECT 56.885 2.49 57.48 2.63 ;
      RECT 56.885 4.81 57.205 5.07 ;
      RECT 54.18 4.825 54.47 5.055 ;
      RECT 54.18 4.87 57.205 5.01 ;
      RECT 56.21 2.39 56.54 2.72 ;
      RECT 56.205 2.425 56.54 2.685 ;
      RECT 56.555 2.445 56.67 2.675 ;
      RECT 56.205 2.44 56.555 2.67 ;
      RECT 56.205 2.49 56.685 2.63 ;
      RECT 56.09 2.49 56.1 2.63 ;
      RECT 56.1 2.485 56.67 2.625 ;
      RECT 52.645 5.89 52.985 6.17 ;
      RECT 50.365 5.915 50.655 6.145 ;
      RECT 50.365 5.945 52.985 6.115 ;
      RECT 52.195 6.63 52.535 6.91 ;
      RECT 52.165 6.655 52.535 6.885 ;
      RECT 51.995 6.685 52.535 6.855 ;
      RECT 51.735 7.765 52.025 7.995 ;
      RECT 51.795 6.995 51.965 7.995 ;
      RECT 51.695 6.995 52.065 7.365 ;
      RECT 49.16 7.765 49.45 7.995 ;
      RECT 49.22 6.285 49.39 7.995 ;
      RECT 49.22 6.655 49.545 6.98 ;
      RECT 49.16 6.285 49.45 6.515 ;
      RECT 49.16 2.365 49.45 2.595 ;
      RECT 49.22 0.885 49.39 2.595 ;
      RECT 49.16 0.885 49.45 1.115 ;
      RECT 48.75 2.735 49.08 2.965 ;
      RECT 48.75 2.765 49.25 2.935 ;
      RECT 48.75 2.395 48.94 2.965 ;
      RECT 48.17 2.365 48.46 2.595 ;
      RECT 48.17 2.395 48.94 2.565 ;
      RECT 48.23 0.885 48.4 2.595 ;
      RECT 48.17 0.885 48.46 1.115 ;
      RECT 48.17 7.765 48.46 7.995 ;
      RECT 48.23 6.285 48.4 7.995 ;
      RECT 48.17 6.285 48.46 6.515 ;
      RECT 48.17 6.325 49.02 6.485 ;
      RECT 48.85 5.915 49.02 6.485 ;
      RECT 48.17 6.32 48.56 6.485 ;
      RECT 48.79 5.915 49.08 6.145 ;
      RECT 48.79 5.945 49.25 6.115 ;
      RECT 47.8 2.735 48.09 2.965 ;
      RECT 47.8 2.765 48.26 2.935 ;
      RECT 47.86 1.655 48.025 2.965 ;
      RECT 46.375 1.625 46.665 1.855 ;
      RECT 46.375 1.655 48.025 1.825 ;
      RECT 46.435 0.885 46.605 1.855 ;
      RECT 46.375 0.885 46.665 1.115 ;
      RECT 46.375 7.765 46.665 7.995 ;
      RECT 46.435 7.025 46.605 7.995 ;
      RECT 46.435 7.12 48.025 7.29 ;
      RECT 47.855 5.915 48.025 7.29 ;
      RECT 46.375 7.025 46.665 7.255 ;
      RECT 47.8 5.915 48.09 6.145 ;
      RECT 47.8 5.945 48.26 6.115 ;
      RECT 44.36 1.995 44.685 2.32 ;
      RECT 46.805 1.965 47.155 2.315 ;
      RECT 44.36 2.025 47.155 2.195 ;
      RECT 46.83 6.655 47.155 6.98 ;
      RECT 46.805 6.655 47.155 6.885 ;
      RECT 46.635 6.685 47.155 6.855 ;
      RECT 46.03 2.365 46.35 2.685 ;
      RECT 46 2.365 46.35 2.595 ;
      RECT 45.715 2.395 46.35 2.565 ;
      RECT 46.03 6.28 46.35 6.605 ;
      RECT 46 6.285 46.35 6.515 ;
      RECT 45.83 6.315 46.35 6.485 ;
      RECT 44.985 3.635 45.31 3.96 ;
      RECT 45.06 2.735 45.24 3.96 ;
      RECT 45.005 2.735 45.295 2.965 ;
      RECT 45.005 2.765 45.465 2.935 ;
      RECT 44.99 5.865 45.315 6.19 ;
      RECT 44.99 5.945 45.465 6.115 ;
      RECT 43.36 2.77 43.68 3.03 ;
      RECT 43.085 2.83 43.68 2.97 ;
      RECT 40.98 3.11 41.3 3.37 ;
      RECT 42.955 3.125 43.245 3.355 ;
      RECT 40.98 3.17 43.245 3.31 ;
      RECT 42.34 5.83 42.66 6.09 ;
      RECT 42.34 5.89 42.935 6.03 ;
      RECT 41.66 2.77 41.98 3.03 ;
      RECT 36.92 2.785 37.21 3.015 ;
      RECT 36.92 2.83 41.98 2.97 ;
      RECT 41.75 2.49 41.89 3.03 ;
      RECT 41.75 2.49 42.23 2.63 ;
      RECT 42.09 2.105 42.23 2.63 ;
      RECT 42.015 2.105 42.305 2.335 ;
      RECT 41.66 3.79 41.98 4.05 ;
      RECT 40.995 3.805 41.285 4.035 ;
      RECT 38.785 3.805 39.075 4.035 ;
      RECT 38.785 3.85 41.98 3.99 ;
      RECT 39.96 5.83 40.28 6.09 ;
      RECT 41.675 5.845 41.965 6.075 ;
      RECT 39.295 5.845 39.585 6.075 ;
      RECT 39.295 5.89 40.28 6.03 ;
      RECT 41.75 5.55 41.89 6.075 ;
      RECT 40.05 5.55 40.19 6.09 ;
      RECT 40.05 5.55 41.89 5.69 ;
      RECT 38.955 2.445 39.245 2.675 ;
      RECT 39.03 2.15 39.17 2.675 ;
      RECT 41.32 2.09 41.64 2.35 ;
      RECT 41.22 2.105 41.64 2.335 ;
      RECT 39.03 2.15 41.64 2.29 ;
      RECT 40.3 2.43 40.62 2.69 ;
      RECT 40.3 2.49 40.895 2.63 ;
      RECT 40.3 4.81 40.62 5.07 ;
      RECT 37.595 4.825 37.885 5.055 ;
      RECT 37.595 4.87 40.62 5.01 ;
      RECT 39.625 2.39 39.955 2.72 ;
      RECT 39.62 2.425 39.955 2.685 ;
      RECT 39.97 2.445 40.085 2.675 ;
      RECT 39.62 2.44 39.97 2.67 ;
      RECT 39.62 2.49 40.1 2.63 ;
      RECT 39.505 2.49 39.515 2.63 ;
      RECT 39.515 2.485 40.085 2.625 ;
      RECT 36.06 5.89 36.4 6.17 ;
      RECT 33.78 5.915 34.07 6.145 ;
      RECT 33.78 5.945 36.4 6.115 ;
      RECT 35.61 6.63 35.95 6.91 ;
      RECT 35.58 6.655 35.95 6.885 ;
      RECT 35.41 6.685 35.95 6.855 ;
      RECT 35.15 7.765 35.44 7.995 ;
      RECT 35.21 6.995 35.38 7.995 ;
      RECT 35.11 6.995 35.48 7.365 ;
      RECT 32.575 7.765 32.865 7.995 ;
      RECT 32.635 6.285 32.805 7.995 ;
      RECT 32.635 6.655 32.96 6.98 ;
      RECT 32.575 6.285 32.865 6.515 ;
      RECT 32.575 2.365 32.865 2.595 ;
      RECT 32.635 0.885 32.805 2.595 ;
      RECT 32.575 0.885 32.865 1.115 ;
      RECT 32.165 2.735 32.495 2.965 ;
      RECT 32.165 2.765 32.665 2.935 ;
      RECT 32.165 2.395 32.355 2.965 ;
      RECT 31.585 2.365 31.875 2.595 ;
      RECT 31.585 2.395 32.355 2.565 ;
      RECT 31.645 0.885 31.815 2.595 ;
      RECT 31.585 0.885 31.875 1.115 ;
      RECT 31.585 7.765 31.875 7.995 ;
      RECT 31.645 6.285 31.815 7.995 ;
      RECT 31.585 6.285 31.875 6.515 ;
      RECT 31.585 6.325 32.435 6.485 ;
      RECT 32.265 5.915 32.435 6.485 ;
      RECT 31.585 6.32 31.975 6.485 ;
      RECT 32.205 5.915 32.495 6.145 ;
      RECT 32.205 5.945 32.665 6.115 ;
      RECT 31.215 2.735 31.505 2.965 ;
      RECT 31.215 2.765 31.675 2.935 ;
      RECT 31.275 1.655 31.44 2.965 ;
      RECT 29.79 1.625 30.08 1.855 ;
      RECT 29.79 1.655 31.44 1.825 ;
      RECT 29.85 0.885 30.02 1.855 ;
      RECT 29.79 0.885 30.08 1.115 ;
      RECT 29.79 7.765 30.08 7.995 ;
      RECT 29.85 7.025 30.02 7.995 ;
      RECT 29.85 7.12 31.44 7.29 ;
      RECT 31.27 5.915 31.44 7.29 ;
      RECT 29.79 7.025 30.08 7.255 ;
      RECT 31.215 5.915 31.505 6.145 ;
      RECT 31.215 5.945 31.675 6.115 ;
      RECT 27.775 1.995 28.1 2.32 ;
      RECT 30.22 1.965 30.57 2.315 ;
      RECT 27.775 2.025 30.57 2.195 ;
      RECT 30.245 6.655 30.57 6.98 ;
      RECT 30.22 6.655 30.57 6.885 ;
      RECT 30.05 6.685 30.57 6.855 ;
      RECT 29.445 2.365 29.765 2.685 ;
      RECT 29.415 2.365 29.765 2.595 ;
      RECT 29.13 2.395 29.765 2.565 ;
      RECT 29.445 6.28 29.765 6.605 ;
      RECT 29.415 6.285 29.765 6.515 ;
      RECT 29.245 6.315 29.765 6.485 ;
      RECT 28.4 3.635 28.725 3.96 ;
      RECT 28.475 2.735 28.655 3.96 ;
      RECT 28.42 2.735 28.71 2.965 ;
      RECT 28.42 2.765 28.88 2.935 ;
      RECT 28.405 5.865 28.73 6.19 ;
      RECT 28.405 5.945 28.88 6.115 ;
      RECT 26.775 2.77 27.095 3.03 ;
      RECT 26.5 2.83 27.095 2.97 ;
      RECT 24.395 3.11 24.715 3.37 ;
      RECT 26.37 3.125 26.66 3.355 ;
      RECT 24.395 3.17 26.66 3.31 ;
      RECT 25.755 5.83 26.075 6.09 ;
      RECT 25.755 5.89 26.35 6.03 ;
      RECT 25.075 2.77 25.395 3.03 ;
      RECT 20.335 2.785 20.625 3.015 ;
      RECT 20.335 2.83 25.395 2.97 ;
      RECT 25.165 2.49 25.305 3.03 ;
      RECT 25.165 2.49 25.645 2.63 ;
      RECT 25.505 2.105 25.645 2.63 ;
      RECT 25.43 2.105 25.72 2.335 ;
      RECT 25.075 3.79 25.395 4.05 ;
      RECT 24.41 3.805 24.7 4.035 ;
      RECT 22.2 3.805 22.49 4.035 ;
      RECT 22.2 3.85 25.395 3.99 ;
      RECT 23.375 5.83 23.695 6.09 ;
      RECT 25.09 5.845 25.38 6.075 ;
      RECT 22.71 5.845 23 6.075 ;
      RECT 22.71 5.89 23.695 6.03 ;
      RECT 25.165 5.55 25.305 6.075 ;
      RECT 23.465 5.55 23.605 6.09 ;
      RECT 23.465 5.55 25.305 5.69 ;
      RECT 22.37 2.445 22.66 2.675 ;
      RECT 22.445 2.15 22.585 2.675 ;
      RECT 24.735 2.09 25.055 2.35 ;
      RECT 24.635 2.105 25.055 2.335 ;
      RECT 22.445 2.15 25.055 2.29 ;
      RECT 23.715 2.43 24.035 2.69 ;
      RECT 23.715 2.49 24.31 2.63 ;
      RECT 23.715 4.81 24.035 5.07 ;
      RECT 21.01 4.825 21.3 5.055 ;
      RECT 21.01 4.87 24.035 5.01 ;
      RECT 23.04 2.39 23.37 2.72 ;
      RECT 23.035 2.425 23.37 2.685 ;
      RECT 23.385 2.445 23.5 2.675 ;
      RECT 23.035 2.44 23.385 2.67 ;
      RECT 23.035 2.49 23.515 2.63 ;
      RECT 22.92 2.49 22.93 2.63 ;
      RECT 22.93 2.485 23.5 2.625 ;
      RECT 19.475 5.89 19.815 6.17 ;
      RECT 17.195 5.915 17.485 6.145 ;
      RECT 17.195 5.945 19.815 6.115 ;
      RECT 19.025 6.63 19.365 6.91 ;
      RECT 18.995 6.655 19.365 6.885 ;
      RECT 18.825 6.685 19.365 6.855 ;
      RECT 18.565 7.765 18.855 7.995 ;
      RECT 18.625 6.995 18.795 7.995 ;
      RECT 18.525 6.995 18.895 7.365 ;
      RECT 15.99 7.765 16.28 7.995 ;
      RECT 16.05 6.285 16.22 7.995 ;
      RECT 16.05 6.655 16.375 6.98 ;
      RECT 15.99 6.285 16.28 6.515 ;
      RECT 15.99 2.365 16.28 2.595 ;
      RECT 16.05 0.885 16.22 2.595 ;
      RECT 15.99 0.885 16.28 1.115 ;
      RECT 15.58 2.735 15.91 2.965 ;
      RECT 15.58 2.765 16.08 2.935 ;
      RECT 15.58 2.395 15.77 2.965 ;
      RECT 15 2.365 15.29 2.595 ;
      RECT 15 2.395 15.77 2.565 ;
      RECT 15.06 0.885 15.23 2.595 ;
      RECT 15 0.885 15.29 1.115 ;
      RECT 15 7.765 15.29 7.995 ;
      RECT 15.06 6.285 15.23 7.995 ;
      RECT 15 6.285 15.29 6.515 ;
      RECT 15 6.325 15.85 6.485 ;
      RECT 15.68 5.915 15.85 6.485 ;
      RECT 15 6.32 15.39 6.485 ;
      RECT 15.62 5.915 15.91 6.145 ;
      RECT 15.62 5.945 16.08 6.115 ;
      RECT 14.63 2.735 14.92 2.965 ;
      RECT 14.63 2.765 15.09 2.935 ;
      RECT 14.69 1.655 14.855 2.965 ;
      RECT 13.205 1.625 13.495 1.855 ;
      RECT 13.205 1.655 14.855 1.825 ;
      RECT 13.265 0.885 13.435 1.855 ;
      RECT 13.205 0.885 13.495 1.115 ;
      RECT 13.205 7.765 13.495 7.995 ;
      RECT 13.265 7.025 13.435 7.995 ;
      RECT 13.265 7.12 14.855 7.29 ;
      RECT 14.685 5.915 14.855 7.29 ;
      RECT 13.205 7.025 13.495 7.255 ;
      RECT 14.63 5.915 14.92 6.145 ;
      RECT 14.63 5.945 15.09 6.115 ;
      RECT 11.19 1.995 11.515 2.32 ;
      RECT 13.635 1.965 13.985 2.315 ;
      RECT 11.19 2.025 13.985 2.195 ;
      RECT 13.66 6.655 13.985 6.98 ;
      RECT 13.635 6.655 13.985 6.885 ;
      RECT 13.465 6.685 13.985 6.855 ;
      RECT 12.86 2.365 13.18 2.685 ;
      RECT 12.83 2.365 13.18 2.595 ;
      RECT 12.545 2.395 13.18 2.565 ;
      RECT 12.86 6.28 13.18 6.605 ;
      RECT 12.83 6.285 13.18 6.515 ;
      RECT 12.66 6.315 13.18 6.485 ;
      RECT 11.815 3.635 12.14 3.96 ;
      RECT 11.89 2.735 12.07 3.96 ;
      RECT 11.835 2.735 12.125 2.965 ;
      RECT 11.835 2.765 12.295 2.935 ;
      RECT 11.82 5.865 12.145 6.19 ;
      RECT 11.82 5.945 12.295 6.115 ;
      RECT 10.19 2.77 10.51 3.03 ;
      RECT 9.915 2.83 10.51 2.97 ;
      RECT 7.81 3.11 8.13 3.37 ;
      RECT 9.785 3.125 10.075 3.355 ;
      RECT 7.81 3.17 10.075 3.31 ;
      RECT 9.17 5.83 9.49 6.09 ;
      RECT 9.17 5.89 9.765 6.03 ;
      RECT 8.49 2.77 8.81 3.03 ;
      RECT 3.75 2.785 4.04 3.015 ;
      RECT 3.75 2.83 8.81 2.97 ;
      RECT 8.58 2.49 8.72 3.03 ;
      RECT 8.58 2.49 9.06 2.63 ;
      RECT 8.92 2.105 9.06 2.63 ;
      RECT 8.845 2.105 9.135 2.335 ;
      RECT 8.49 3.79 8.81 4.05 ;
      RECT 7.825 3.805 8.115 4.035 ;
      RECT 5.615 3.805 5.905 4.035 ;
      RECT 5.615 3.85 8.81 3.99 ;
      RECT 6.79 5.83 7.11 6.09 ;
      RECT 8.505 5.845 8.795 6.075 ;
      RECT 6.125 5.845 6.415 6.075 ;
      RECT 6.125 5.89 7.11 6.03 ;
      RECT 8.58 5.55 8.72 6.075 ;
      RECT 6.88 5.55 7.02 6.09 ;
      RECT 6.88 5.55 8.72 5.69 ;
      RECT 5.785 2.445 6.075 2.675 ;
      RECT 5.86 2.15 6 2.675 ;
      RECT 8.15 2.09 8.47 2.35 ;
      RECT 8.05 2.105 8.47 2.335 ;
      RECT 5.86 2.15 8.47 2.29 ;
      RECT 7.13 2.43 7.45 2.69 ;
      RECT 7.13 2.49 7.725 2.63 ;
      RECT 7.13 4.81 7.45 5.07 ;
      RECT 4.425 4.825 4.715 5.055 ;
      RECT 4.425 4.87 7.45 5.01 ;
      RECT 6.455 2.39 6.785 2.72 ;
      RECT 6.45 2.425 6.785 2.685 ;
      RECT 6.8 2.445 6.915 2.675 ;
      RECT 6.45 2.44 6.8 2.67 ;
      RECT 6.45 2.49 6.93 2.63 ;
      RECT 6.335 2.49 6.345 2.63 ;
      RECT 6.345 2.485 6.915 2.625 ;
      RECT 2.89 5.89 3.23 6.17 ;
      RECT 0.61 5.915 0.9 6.145 ;
      RECT 0.61 5.945 3.23 6.115 ;
      RECT 2.44 6.63 2.78 6.91 ;
      RECT 2.41 6.655 2.78 6.885 ;
      RECT 2.24 6.685 2.78 6.855 ;
      RECT 1.98 7.765 2.27 7.995 ;
      RECT 2.04 6.995 2.21 7.995 ;
      RECT 1.94 6.995 2.31 7.365 ;
      RECT -0.82 6.655 -0.53 6.885 ;
      RECT -0.99 6.685 -0.53 6.855 ;
      RECT -1.25 7.765 -0.96 7.995 ;
      RECT -1.19 7.025 -1.02 7.995 ;
      RECT -1.27 7.025 -0.93 7.305 ;
      RECT -1.655 6.285 -1.315 6.565 ;
      RECT -1.795 6.315 -1.315 6.485 ;
      RECT -2.62 5.915 -2.33 6.145 ;
      RECT -2.62 5.945 -2.16 6.115 ;
      RECT 76.2 4.81 76.845 5.07 ;
      RECT 74.145 5.83 74.465 6.09 ;
      RECT 59.62 4.81 60.265 5.07 ;
      RECT 57.565 5.83 57.885 6.09 ;
      RECT 43.035 4.81 43.68 5.07 ;
      RECT 40.98 5.83 41.3 6.09 ;
      RECT 26.45 4.81 27.095 5.07 ;
      RECT 24.395 5.83 24.715 6.09 ;
      RECT 9.865 4.81 10.51 5.07 ;
      RECT 7.81 5.83 8.13 6.09 ;
    LAYER mcon ;
      RECT 82.385 0.915 82.555 1.085 ;
      RECT 82.385 2.395 82.555 2.565 ;
      RECT 82.385 6.315 82.555 6.485 ;
      RECT 82.385 7.795 82.555 7.965 ;
      RECT 82.035 0.105 82.205 0.275 ;
      RECT 82.035 4.165 82.205 4.335 ;
      RECT 82.035 4.545 82.205 4.715 ;
      RECT 82.035 8.605 82.205 8.775 ;
      RECT 82.015 2.765 82.185 2.935 ;
      RECT 82.015 5.945 82.185 6.115 ;
      RECT 81.395 0.915 81.565 1.085 ;
      RECT 81.395 2.395 81.565 2.565 ;
      RECT 81.395 6.315 81.565 6.485 ;
      RECT 81.395 7.795 81.565 7.965 ;
      RECT 81.045 0.105 81.215 0.275 ;
      RECT 81.045 4.165 81.215 4.335 ;
      RECT 81.045 4.545 81.215 4.715 ;
      RECT 81.045 8.605 81.215 8.775 ;
      RECT 81.025 2.765 81.195 2.935 ;
      RECT 81.025 5.945 81.195 6.115 ;
      RECT 80.34 0.105 80.51 0.275 ;
      RECT 80.34 4.165 80.51 4.335 ;
      RECT 80.34 4.545 80.51 4.715 ;
      RECT 80.34 8.605 80.51 8.775 ;
      RECT 80.03 2.025 80.2 2.195 ;
      RECT 80.03 6.685 80.2 6.855 ;
      RECT 79.66 0.105 79.83 0.275 ;
      RECT 79.66 8.605 79.83 8.775 ;
      RECT 79.6 0.915 79.77 1.085 ;
      RECT 79.6 1.655 79.77 1.825 ;
      RECT 79.6 7.055 79.77 7.225 ;
      RECT 79.6 7.795 79.77 7.965 ;
      RECT 79.225 2.395 79.395 2.565 ;
      RECT 79.225 6.315 79.395 6.485 ;
      RECT 78.98 0.105 79.15 0.275 ;
      RECT 78.98 8.605 79.15 8.775 ;
      RECT 78.3 0.105 78.47 0.275 ;
      RECT 78.3 8.605 78.47 8.775 ;
      RECT 78.23 2.765 78.4 2.935 ;
      RECT 78.23 5.945 78.4 6.115 ;
      RECT 76.64 1.625 76.81 1.795 ;
      RECT 76.64 4.345 76.81 4.515 ;
      RECT 76.64 7.065 76.81 7.235 ;
      RECT 76.6 2.815 76.77 2.985 ;
      RECT 76.26 4.855 76.43 5.025 ;
      RECT 76.18 1.625 76.35 1.795 ;
      RECT 76.18 3.155 76.35 3.325 ;
      RECT 76.18 4.345 76.35 4.515 ;
      RECT 76.18 7.065 76.35 7.235 ;
      RECT 75.72 1.625 75.89 1.795 ;
      RECT 75.72 4.345 75.89 4.515 ;
      RECT 75.72 7.065 75.89 7.235 ;
      RECT 75.58 5.875 75.75 6.045 ;
      RECT 75.26 1.625 75.43 1.795 ;
      RECT 75.26 4.345 75.43 4.515 ;
      RECT 75.26 7.065 75.43 7.235 ;
      RECT 75.24 2.135 75.41 2.305 ;
      RECT 74.9 5.875 75.07 6.045 ;
      RECT 74.8 1.625 74.97 1.795 ;
      RECT 74.8 4.345 74.97 4.515 ;
      RECT 74.8 7.065 74.97 7.235 ;
      RECT 74.445 2.135 74.615 2.305 ;
      RECT 74.34 1.625 74.51 1.795 ;
      RECT 74.34 4.345 74.51 4.515 ;
      RECT 74.34 7.065 74.51 7.235 ;
      RECT 74.22 3.835 74.39 4.005 ;
      RECT 74.22 5.875 74.39 6.045 ;
      RECT 73.88 1.625 74.05 1.795 ;
      RECT 73.88 4.345 74.05 4.515 ;
      RECT 73.88 7.065 74.05 7.235 ;
      RECT 73.71 5.875 73.88 6.045 ;
      RECT 73.54 2.475 73.71 2.645 ;
      RECT 73.42 1.625 73.59 1.795 ;
      RECT 73.42 4.345 73.59 4.515 ;
      RECT 73.42 7.065 73.59 7.235 ;
      RECT 72.96 1.625 73.13 1.795 ;
      RECT 72.96 4.345 73.13 4.515 ;
      RECT 72.96 7.065 73.13 7.235 ;
      RECT 72.52 5.875 72.69 6.045 ;
      RECT 72.5 1.625 72.67 1.795 ;
      RECT 72.5 4.345 72.67 4.515 ;
      RECT 72.5 7.065 72.67 7.235 ;
      RECT 72.18 2.475 72.35 2.645 ;
      RECT 72.04 1.625 72.21 1.795 ;
      RECT 72.04 4.345 72.21 4.515 ;
      RECT 72.04 7.065 72.21 7.235 ;
      RECT 72.01 3.835 72.18 4.005 ;
      RECT 71.58 1.625 71.75 1.795 ;
      RECT 71.58 4.345 71.75 4.515 ;
      RECT 71.58 7.065 71.75 7.235 ;
      RECT 71.5 5.875 71.67 6.045 ;
      RECT 71.12 1.625 71.29 1.795 ;
      RECT 71.12 4.345 71.29 4.515 ;
      RECT 71.12 7.065 71.29 7.235 ;
      RECT 70.82 4.855 70.99 5.025 ;
      RECT 70.66 1.625 70.83 1.795 ;
      RECT 70.66 4.345 70.83 4.515 ;
      RECT 70.66 7.065 70.83 7.235 ;
      RECT 70.2 1.625 70.37 1.795 ;
      RECT 70.2 4.345 70.37 4.515 ;
      RECT 70.2 7.065 70.37 7.235 ;
      RECT 70.145 2.815 70.315 2.985 ;
      RECT 69.115 4.545 69.285 4.715 ;
      RECT 69.115 8.605 69.285 8.775 ;
      RECT 68.805 6.685 68.975 6.855 ;
      RECT 68.435 8.605 68.605 8.775 ;
      RECT 68.375 7.055 68.545 7.225 ;
      RECT 68.375 7.795 68.545 7.965 ;
      RECT 68 6.315 68.17 6.485 ;
      RECT 67.755 8.605 67.925 8.775 ;
      RECT 67.075 8.605 67.245 8.775 ;
      RECT 67.005 5.945 67.175 6.115 ;
      RECT 65.805 0.915 65.975 1.085 ;
      RECT 65.805 2.395 65.975 2.565 ;
      RECT 65.805 6.315 65.975 6.485 ;
      RECT 65.805 7.795 65.975 7.965 ;
      RECT 65.455 0.105 65.625 0.275 ;
      RECT 65.455 4.165 65.625 4.335 ;
      RECT 65.455 4.545 65.625 4.715 ;
      RECT 65.455 8.605 65.625 8.775 ;
      RECT 65.435 2.765 65.605 2.935 ;
      RECT 65.435 5.945 65.605 6.115 ;
      RECT 64.815 0.915 64.985 1.085 ;
      RECT 64.815 2.395 64.985 2.565 ;
      RECT 64.815 6.315 64.985 6.485 ;
      RECT 64.815 7.795 64.985 7.965 ;
      RECT 64.465 0.105 64.635 0.275 ;
      RECT 64.465 4.165 64.635 4.335 ;
      RECT 64.465 4.545 64.635 4.715 ;
      RECT 64.465 8.605 64.635 8.775 ;
      RECT 64.445 2.765 64.615 2.935 ;
      RECT 64.445 5.945 64.615 6.115 ;
      RECT 63.76 0.105 63.93 0.275 ;
      RECT 63.76 4.165 63.93 4.335 ;
      RECT 63.76 4.545 63.93 4.715 ;
      RECT 63.76 8.605 63.93 8.775 ;
      RECT 63.45 2.025 63.62 2.195 ;
      RECT 63.45 6.685 63.62 6.855 ;
      RECT 63.08 0.105 63.25 0.275 ;
      RECT 63.08 8.605 63.25 8.775 ;
      RECT 63.02 0.915 63.19 1.085 ;
      RECT 63.02 1.655 63.19 1.825 ;
      RECT 63.02 7.055 63.19 7.225 ;
      RECT 63.02 7.795 63.19 7.965 ;
      RECT 62.645 2.395 62.815 2.565 ;
      RECT 62.645 6.315 62.815 6.485 ;
      RECT 62.4 0.105 62.57 0.275 ;
      RECT 62.4 8.605 62.57 8.775 ;
      RECT 61.72 0.105 61.89 0.275 ;
      RECT 61.72 8.605 61.89 8.775 ;
      RECT 61.65 2.765 61.82 2.935 ;
      RECT 61.65 5.945 61.82 6.115 ;
      RECT 60.06 1.625 60.23 1.795 ;
      RECT 60.06 4.345 60.23 4.515 ;
      RECT 60.06 7.065 60.23 7.235 ;
      RECT 60.02 2.815 60.19 2.985 ;
      RECT 59.68 4.855 59.85 5.025 ;
      RECT 59.6 1.625 59.77 1.795 ;
      RECT 59.6 3.155 59.77 3.325 ;
      RECT 59.6 4.345 59.77 4.515 ;
      RECT 59.6 7.065 59.77 7.235 ;
      RECT 59.14 1.625 59.31 1.795 ;
      RECT 59.14 4.345 59.31 4.515 ;
      RECT 59.14 7.065 59.31 7.235 ;
      RECT 59 5.875 59.17 6.045 ;
      RECT 58.68 1.625 58.85 1.795 ;
      RECT 58.68 4.345 58.85 4.515 ;
      RECT 58.68 7.065 58.85 7.235 ;
      RECT 58.66 2.135 58.83 2.305 ;
      RECT 58.32 5.875 58.49 6.045 ;
      RECT 58.22 1.625 58.39 1.795 ;
      RECT 58.22 4.345 58.39 4.515 ;
      RECT 58.22 7.065 58.39 7.235 ;
      RECT 57.865 2.135 58.035 2.305 ;
      RECT 57.76 1.625 57.93 1.795 ;
      RECT 57.76 4.345 57.93 4.515 ;
      RECT 57.76 7.065 57.93 7.235 ;
      RECT 57.64 3.835 57.81 4.005 ;
      RECT 57.64 5.875 57.81 6.045 ;
      RECT 57.3 1.625 57.47 1.795 ;
      RECT 57.3 4.345 57.47 4.515 ;
      RECT 57.3 7.065 57.47 7.235 ;
      RECT 57.13 5.875 57.3 6.045 ;
      RECT 56.96 2.475 57.13 2.645 ;
      RECT 56.84 1.625 57.01 1.795 ;
      RECT 56.84 4.345 57.01 4.515 ;
      RECT 56.84 7.065 57.01 7.235 ;
      RECT 56.38 1.625 56.55 1.795 ;
      RECT 56.38 4.345 56.55 4.515 ;
      RECT 56.38 7.065 56.55 7.235 ;
      RECT 55.94 5.875 56.11 6.045 ;
      RECT 55.92 1.625 56.09 1.795 ;
      RECT 55.92 4.345 56.09 4.515 ;
      RECT 55.92 7.065 56.09 7.235 ;
      RECT 55.6 2.475 55.77 2.645 ;
      RECT 55.46 1.625 55.63 1.795 ;
      RECT 55.46 4.345 55.63 4.515 ;
      RECT 55.46 7.065 55.63 7.235 ;
      RECT 55.43 3.835 55.6 4.005 ;
      RECT 55 1.625 55.17 1.795 ;
      RECT 55 4.345 55.17 4.515 ;
      RECT 55 7.065 55.17 7.235 ;
      RECT 54.92 5.875 55.09 6.045 ;
      RECT 54.54 1.625 54.71 1.795 ;
      RECT 54.54 4.345 54.71 4.515 ;
      RECT 54.54 7.065 54.71 7.235 ;
      RECT 54.24 4.855 54.41 5.025 ;
      RECT 54.08 1.625 54.25 1.795 ;
      RECT 54.08 4.345 54.25 4.515 ;
      RECT 54.08 7.065 54.25 7.235 ;
      RECT 53.62 1.625 53.79 1.795 ;
      RECT 53.62 4.345 53.79 4.515 ;
      RECT 53.62 7.065 53.79 7.235 ;
      RECT 53.565 2.815 53.735 2.985 ;
      RECT 52.535 4.545 52.705 4.715 ;
      RECT 52.535 8.605 52.705 8.775 ;
      RECT 52.225 6.685 52.395 6.855 ;
      RECT 51.855 8.605 52.025 8.775 ;
      RECT 51.795 7.055 51.965 7.225 ;
      RECT 51.795 7.795 51.965 7.965 ;
      RECT 51.42 6.315 51.59 6.485 ;
      RECT 51.175 8.605 51.345 8.775 ;
      RECT 50.495 8.605 50.665 8.775 ;
      RECT 50.425 5.945 50.595 6.115 ;
      RECT 49.22 0.915 49.39 1.085 ;
      RECT 49.22 2.395 49.39 2.565 ;
      RECT 49.22 6.315 49.39 6.485 ;
      RECT 49.22 7.795 49.39 7.965 ;
      RECT 48.87 0.105 49.04 0.275 ;
      RECT 48.87 4.165 49.04 4.335 ;
      RECT 48.87 4.545 49.04 4.715 ;
      RECT 48.87 8.605 49.04 8.775 ;
      RECT 48.85 2.765 49.02 2.935 ;
      RECT 48.85 5.945 49.02 6.115 ;
      RECT 48.23 0.915 48.4 1.085 ;
      RECT 48.23 2.395 48.4 2.565 ;
      RECT 48.23 6.315 48.4 6.485 ;
      RECT 48.23 7.795 48.4 7.965 ;
      RECT 47.88 0.105 48.05 0.275 ;
      RECT 47.88 4.165 48.05 4.335 ;
      RECT 47.88 4.545 48.05 4.715 ;
      RECT 47.88 8.605 48.05 8.775 ;
      RECT 47.86 2.765 48.03 2.935 ;
      RECT 47.86 5.945 48.03 6.115 ;
      RECT 47.175 0.105 47.345 0.275 ;
      RECT 47.175 4.165 47.345 4.335 ;
      RECT 47.175 4.545 47.345 4.715 ;
      RECT 47.175 8.605 47.345 8.775 ;
      RECT 46.865 2.025 47.035 2.195 ;
      RECT 46.865 6.685 47.035 6.855 ;
      RECT 46.495 0.105 46.665 0.275 ;
      RECT 46.495 8.605 46.665 8.775 ;
      RECT 46.435 0.915 46.605 1.085 ;
      RECT 46.435 1.655 46.605 1.825 ;
      RECT 46.435 7.055 46.605 7.225 ;
      RECT 46.435 7.795 46.605 7.965 ;
      RECT 46.06 2.395 46.23 2.565 ;
      RECT 46.06 6.315 46.23 6.485 ;
      RECT 45.815 0.105 45.985 0.275 ;
      RECT 45.815 8.605 45.985 8.775 ;
      RECT 45.135 0.105 45.305 0.275 ;
      RECT 45.135 8.605 45.305 8.775 ;
      RECT 45.065 2.765 45.235 2.935 ;
      RECT 45.065 5.945 45.235 6.115 ;
      RECT 43.475 1.625 43.645 1.795 ;
      RECT 43.475 4.345 43.645 4.515 ;
      RECT 43.475 7.065 43.645 7.235 ;
      RECT 43.435 2.815 43.605 2.985 ;
      RECT 43.095 4.855 43.265 5.025 ;
      RECT 43.015 1.625 43.185 1.795 ;
      RECT 43.015 3.155 43.185 3.325 ;
      RECT 43.015 4.345 43.185 4.515 ;
      RECT 43.015 7.065 43.185 7.235 ;
      RECT 42.555 1.625 42.725 1.795 ;
      RECT 42.555 4.345 42.725 4.515 ;
      RECT 42.555 7.065 42.725 7.235 ;
      RECT 42.415 5.875 42.585 6.045 ;
      RECT 42.095 1.625 42.265 1.795 ;
      RECT 42.095 4.345 42.265 4.515 ;
      RECT 42.095 7.065 42.265 7.235 ;
      RECT 42.075 2.135 42.245 2.305 ;
      RECT 41.735 5.875 41.905 6.045 ;
      RECT 41.635 1.625 41.805 1.795 ;
      RECT 41.635 4.345 41.805 4.515 ;
      RECT 41.635 7.065 41.805 7.235 ;
      RECT 41.28 2.135 41.45 2.305 ;
      RECT 41.175 1.625 41.345 1.795 ;
      RECT 41.175 4.345 41.345 4.515 ;
      RECT 41.175 7.065 41.345 7.235 ;
      RECT 41.055 3.835 41.225 4.005 ;
      RECT 41.055 5.875 41.225 6.045 ;
      RECT 40.715 1.625 40.885 1.795 ;
      RECT 40.715 4.345 40.885 4.515 ;
      RECT 40.715 7.065 40.885 7.235 ;
      RECT 40.545 5.875 40.715 6.045 ;
      RECT 40.375 2.475 40.545 2.645 ;
      RECT 40.255 1.625 40.425 1.795 ;
      RECT 40.255 4.345 40.425 4.515 ;
      RECT 40.255 7.065 40.425 7.235 ;
      RECT 39.795 1.625 39.965 1.795 ;
      RECT 39.795 4.345 39.965 4.515 ;
      RECT 39.795 7.065 39.965 7.235 ;
      RECT 39.355 5.875 39.525 6.045 ;
      RECT 39.335 1.625 39.505 1.795 ;
      RECT 39.335 4.345 39.505 4.515 ;
      RECT 39.335 7.065 39.505 7.235 ;
      RECT 39.015 2.475 39.185 2.645 ;
      RECT 38.875 1.625 39.045 1.795 ;
      RECT 38.875 4.345 39.045 4.515 ;
      RECT 38.875 7.065 39.045 7.235 ;
      RECT 38.845 3.835 39.015 4.005 ;
      RECT 38.415 1.625 38.585 1.795 ;
      RECT 38.415 4.345 38.585 4.515 ;
      RECT 38.415 7.065 38.585 7.235 ;
      RECT 38.335 5.875 38.505 6.045 ;
      RECT 37.955 1.625 38.125 1.795 ;
      RECT 37.955 4.345 38.125 4.515 ;
      RECT 37.955 7.065 38.125 7.235 ;
      RECT 37.655 4.855 37.825 5.025 ;
      RECT 37.495 1.625 37.665 1.795 ;
      RECT 37.495 4.345 37.665 4.515 ;
      RECT 37.495 7.065 37.665 7.235 ;
      RECT 37.035 1.625 37.205 1.795 ;
      RECT 37.035 4.345 37.205 4.515 ;
      RECT 37.035 7.065 37.205 7.235 ;
      RECT 36.98 2.815 37.15 2.985 ;
      RECT 35.95 4.545 36.12 4.715 ;
      RECT 35.95 8.605 36.12 8.775 ;
      RECT 35.64 6.685 35.81 6.855 ;
      RECT 35.27 8.605 35.44 8.775 ;
      RECT 35.21 7.055 35.38 7.225 ;
      RECT 35.21 7.795 35.38 7.965 ;
      RECT 34.835 6.315 35.005 6.485 ;
      RECT 34.59 8.605 34.76 8.775 ;
      RECT 33.91 8.605 34.08 8.775 ;
      RECT 33.84 5.945 34.01 6.115 ;
      RECT 32.635 0.915 32.805 1.085 ;
      RECT 32.635 2.395 32.805 2.565 ;
      RECT 32.635 6.315 32.805 6.485 ;
      RECT 32.635 7.795 32.805 7.965 ;
      RECT 32.285 0.105 32.455 0.275 ;
      RECT 32.285 4.165 32.455 4.335 ;
      RECT 32.285 4.545 32.455 4.715 ;
      RECT 32.285 8.605 32.455 8.775 ;
      RECT 32.265 2.765 32.435 2.935 ;
      RECT 32.265 5.945 32.435 6.115 ;
      RECT 31.645 0.915 31.815 1.085 ;
      RECT 31.645 2.395 31.815 2.565 ;
      RECT 31.645 6.315 31.815 6.485 ;
      RECT 31.645 7.795 31.815 7.965 ;
      RECT 31.295 0.105 31.465 0.275 ;
      RECT 31.295 4.165 31.465 4.335 ;
      RECT 31.295 4.545 31.465 4.715 ;
      RECT 31.295 8.605 31.465 8.775 ;
      RECT 31.275 2.765 31.445 2.935 ;
      RECT 31.275 5.945 31.445 6.115 ;
      RECT 30.59 0.105 30.76 0.275 ;
      RECT 30.59 4.165 30.76 4.335 ;
      RECT 30.59 4.545 30.76 4.715 ;
      RECT 30.59 8.605 30.76 8.775 ;
      RECT 30.28 2.025 30.45 2.195 ;
      RECT 30.28 6.685 30.45 6.855 ;
      RECT 29.91 0.105 30.08 0.275 ;
      RECT 29.91 8.605 30.08 8.775 ;
      RECT 29.85 0.915 30.02 1.085 ;
      RECT 29.85 1.655 30.02 1.825 ;
      RECT 29.85 7.055 30.02 7.225 ;
      RECT 29.85 7.795 30.02 7.965 ;
      RECT 29.475 2.395 29.645 2.565 ;
      RECT 29.475 6.315 29.645 6.485 ;
      RECT 29.23 0.105 29.4 0.275 ;
      RECT 29.23 8.605 29.4 8.775 ;
      RECT 28.55 0.105 28.72 0.275 ;
      RECT 28.55 8.605 28.72 8.775 ;
      RECT 28.48 2.765 28.65 2.935 ;
      RECT 28.48 5.945 28.65 6.115 ;
      RECT 26.89 1.625 27.06 1.795 ;
      RECT 26.89 4.345 27.06 4.515 ;
      RECT 26.89 7.065 27.06 7.235 ;
      RECT 26.85 2.815 27.02 2.985 ;
      RECT 26.51 4.855 26.68 5.025 ;
      RECT 26.43 1.625 26.6 1.795 ;
      RECT 26.43 3.155 26.6 3.325 ;
      RECT 26.43 4.345 26.6 4.515 ;
      RECT 26.43 7.065 26.6 7.235 ;
      RECT 25.97 1.625 26.14 1.795 ;
      RECT 25.97 4.345 26.14 4.515 ;
      RECT 25.97 7.065 26.14 7.235 ;
      RECT 25.83 5.875 26 6.045 ;
      RECT 25.51 1.625 25.68 1.795 ;
      RECT 25.51 4.345 25.68 4.515 ;
      RECT 25.51 7.065 25.68 7.235 ;
      RECT 25.49 2.135 25.66 2.305 ;
      RECT 25.15 5.875 25.32 6.045 ;
      RECT 25.05 1.625 25.22 1.795 ;
      RECT 25.05 4.345 25.22 4.515 ;
      RECT 25.05 7.065 25.22 7.235 ;
      RECT 24.695 2.135 24.865 2.305 ;
      RECT 24.59 1.625 24.76 1.795 ;
      RECT 24.59 4.345 24.76 4.515 ;
      RECT 24.59 7.065 24.76 7.235 ;
      RECT 24.47 3.835 24.64 4.005 ;
      RECT 24.47 5.875 24.64 6.045 ;
      RECT 24.13 1.625 24.3 1.795 ;
      RECT 24.13 4.345 24.3 4.515 ;
      RECT 24.13 7.065 24.3 7.235 ;
      RECT 23.96 5.875 24.13 6.045 ;
      RECT 23.79 2.475 23.96 2.645 ;
      RECT 23.67 1.625 23.84 1.795 ;
      RECT 23.67 4.345 23.84 4.515 ;
      RECT 23.67 7.065 23.84 7.235 ;
      RECT 23.21 1.625 23.38 1.795 ;
      RECT 23.21 4.345 23.38 4.515 ;
      RECT 23.21 7.065 23.38 7.235 ;
      RECT 22.77 5.875 22.94 6.045 ;
      RECT 22.75 1.625 22.92 1.795 ;
      RECT 22.75 4.345 22.92 4.515 ;
      RECT 22.75 7.065 22.92 7.235 ;
      RECT 22.43 2.475 22.6 2.645 ;
      RECT 22.29 1.625 22.46 1.795 ;
      RECT 22.29 4.345 22.46 4.515 ;
      RECT 22.29 7.065 22.46 7.235 ;
      RECT 22.26 3.835 22.43 4.005 ;
      RECT 21.83 1.625 22 1.795 ;
      RECT 21.83 4.345 22 4.515 ;
      RECT 21.83 7.065 22 7.235 ;
      RECT 21.75 5.875 21.92 6.045 ;
      RECT 21.37 1.625 21.54 1.795 ;
      RECT 21.37 4.345 21.54 4.515 ;
      RECT 21.37 7.065 21.54 7.235 ;
      RECT 21.07 4.855 21.24 5.025 ;
      RECT 20.91 1.625 21.08 1.795 ;
      RECT 20.91 4.345 21.08 4.515 ;
      RECT 20.91 7.065 21.08 7.235 ;
      RECT 20.45 1.625 20.62 1.795 ;
      RECT 20.45 4.345 20.62 4.515 ;
      RECT 20.45 7.065 20.62 7.235 ;
      RECT 20.395 2.815 20.565 2.985 ;
      RECT 19.365 4.545 19.535 4.715 ;
      RECT 19.365 8.605 19.535 8.775 ;
      RECT 19.055 6.685 19.225 6.855 ;
      RECT 18.685 8.605 18.855 8.775 ;
      RECT 18.625 7.055 18.795 7.225 ;
      RECT 18.625 7.795 18.795 7.965 ;
      RECT 18.25 6.315 18.42 6.485 ;
      RECT 18.005 8.605 18.175 8.775 ;
      RECT 17.325 8.605 17.495 8.775 ;
      RECT 17.255 5.945 17.425 6.115 ;
      RECT 16.05 0.915 16.22 1.085 ;
      RECT 16.05 2.395 16.22 2.565 ;
      RECT 16.05 6.315 16.22 6.485 ;
      RECT 16.05 7.795 16.22 7.965 ;
      RECT 15.7 0.105 15.87 0.275 ;
      RECT 15.7 4.165 15.87 4.335 ;
      RECT 15.7 4.545 15.87 4.715 ;
      RECT 15.7 8.605 15.87 8.775 ;
      RECT 15.68 2.765 15.85 2.935 ;
      RECT 15.68 5.945 15.85 6.115 ;
      RECT 15.06 0.915 15.23 1.085 ;
      RECT 15.06 2.395 15.23 2.565 ;
      RECT 15.06 6.315 15.23 6.485 ;
      RECT 15.06 7.795 15.23 7.965 ;
      RECT 14.71 0.105 14.88 0.275 ;
      RECT 14.71 4.165 14.88 4.335 ;
      RECT 14.71 4.545 14.88 4.715 ;
      RECT 14.71 8.605 14.88 8.775 ;
      RECT 14.69 2.765 14.86 2.935 ;
      RECT 14.69 5.945 14.86 6.115 ;
      RECT 14.005 0.105 14.175 0.275 ;
      RECT 14.005 4.165 14.175 4.335 ;
      RECT 14.005 4.545 14.175 4.715 ;
      RECT 14.005 8.605 14.175 8.775 ;
      RECT 13.695 2.025 13.865 2.195 ;
      RECT 13.695 6.685 13.865 6.855 ;
      RECT 13.325 0.105 13.495 0.275 ;
      RECT 13.325 8.605 13.495 8.775 ;
      RECT 13.265 0.915 13.435 1.085 ;
      RECT 13.265 1.655 13.435 1.825 ;
      RECT 13.265 7.055 13.435 7.225 ;
      RECT 13.265 7.795 13.435 7.965 ;
      RECT 12.89 2.395 13.06 2.565 ;
      RECT 12.89 6.315 13.06 6.485 ;
      RECT 12.645 0.105 12.815 0.275 ;
      RECT 12.645 8.605 12.815 8.775 ;
      RECT 11.965 0.105 12.135 0.275 ;
      RECT 11.965 8.605 12.135 8.775 ;
      RECT 11.895 2.765 12.065 2.935 ;
      RECT 11.895 5.945 12.065 6.115 ;
      RECT 10.305 1.625 10.475 1.795 ;
      RECT 10.305 4.345 10.475 4.515 ;
      RECT 10.305 7.065 10.475 7.235 ;
      RECT 10.265 2.815 10.435 2.985 ;
      RECT 9.925 4.855 10.095 5.025 ;
      RECT 9.845 1.625 10.015 1.795 ;
      RECT 9.845 3.155 10.015 3.325 ;
      RECT 9.845 4.345 10.015 4.515 ;
      RECT 9.845 7.065 10.015 7.235 ;
      RECT 9.385 1.625 9.555 1.795 ;
      RECT 9.385 4.345 9.555 4.515 ;
      RECT 9.385 7.065 9.555 7.235 ;
      RECT 9.245 5.875 9.415 6.045 ;
      RECT 8.925 1.625 9.095 1.795 ;
      RECT 8.925 4.345 9.095 4.515 ;
      RECT 8.925 7.065 9.095 7.235 ;
      RECT 8.905 2.135 9.075 2.305 ;
      RECT 8.565 5.875 8.735 6.045 ;
      RECT 8.465 1.625 8.635 1.795 ;
      RECT 8.465 4.345 8.635 4.515 ;
      RECT 8.465 7.065 8.635 7.235 ;
      RECT 8.11 2.135 8.28 2.305 ;
      RECT 8.005 1.625 8.175 1.795 ;
      RECT 8.005 4.345 8.175 4.515 ;
      RECT 8.005 7.065 8.175 7.235 ;
      RECT 7.885 3.835 8.055 4.005 ;
      RECT 7.885 5.875 8.055 6.045 ;
      RECT 7.545 1.625 7.715 1.795 ;
      RECT 7.545 4.345 7.715 4.515 ;
      RECT 7.545 7.065 7.715 7.235 ;
      RECT 7.375 5.875 7.545 6.045 ;
      RECT 7.205 2.475 7.375 2.645 ;
      RECT 7.085 1.625 7.255 1.795 ;
      RECT 7.085 4.345 7.255 4.515 ;
      RECT 7.085 7.065 7.255 7.235 ;
      RECT 6.625 1.625 6.795 1.795 ;
      RECT 6.625 4.345 6.795 4.515 ;
      RECT 6.625 7.065 6.795 7.235 ;
      RECT 6.185 5.875 6.355 6.045 ;
      RECT 6.165 1.625 6.335 1.795 ;
      RECT 6.165 4.345 6.335 4.515 ;
      RECT 6.165 7.065 6.335 7.235 ;
      RECT 5.845 2.475 6.015 2.645 ;
      RECT 5.705 1.625 5.875 1.795 ;
      RECT 5.705 4.345 5.875 4.515 ;
      RECT 5.705 7.065 5.875 7.235 ;
      RECT 5.675 3.835 5.845 4.005 ;
      RECT 5.245 1.625 5.415 1.795 ;
      RECT 5.245 4.345 5.415 4.515 ;
      RECT 5.245 7.065 5.415 7.235 ;
      RECT 5.165 5.875 5.335 6.045 ;
      RECT 4.785 1.625 4.955 1.795 ;
      RECT 4.785 4.345 4.955 4.515 ;
      RECT 4.785 7.065 4.955 7.235 ;
      RECT 4.485 4.855 4.655 5.025 ;
      RECT 4.325 1.625 4.495 1.795 ;
      RECT 4.325 4.345 4.495 4.515 ;
      RECT 4.325 7.065 4.495 7.235 ;
      RECT 3.865 1.625 4.035 1.795 ;
      RECT 3.865 4.345 4.035 4.515 ;
      RECT 3.865 7.065 4.035 7.235 ;
      RECT 3.81 2.815 3.98 2.985 ;
      RECT 2.78 4.545 2.95 4.715 ;
      RECT 2.78 8.605 2.95 8.775 ;
      RECT 2.47 6.685 2.64 6.855 ;
      RECT 2.1 8.605 2.27 8.775 ;
      RECT 2.04 7.055 2.21 7.225 ;
      RECT 2.04 7.795 2.21 7.965 ;
      RECT 1.665 6.315 1.835 6.485 ;
      RECT 1.42 8.605 1.59 8.775 ;
      RECT 0.74 8.605 0.91 8.775 ;
      RECT 0.67 5.945 0.84 6.115 ;
      RECT -0.45 4.545 -0.28 4.715 ;
      RECT -0.45 8.605 -0.28 8.775 ;
      RECT -0.76 6.685 -0.59 6.855 ;
      RECT -1.13 8.605 -0.96 8.775 ;
      RECT -1.19 7.055 -1.02 7.225 ;
      RECT -1.19 7.795 -1.02 7.965 ;
      RECT -1.565 6.315 -1.395 6.485 ;
      RECT -1.81 8.605 -1.64 8.775 ;
      RECT -2.49 8.605 -2.32 8.775 ;
      RECT -2.56 5.945 -2.39 6.115 ;
    LAYER li ;
      RECT 70.14 0 70.4 2.615 ;
      RECT 53.56 0 53.82 2.615 ;
      RECT 36.975 0 37.235 2.615 ;
      RECT 20.39 0 20.65 2.615 ;
      RECT 3.805 0 4.065 2.615 ;
      RECT 76.59 0 76.86 2.605 ;
      RECT 75.68 0 75.92 2.605 ;
      RECT 60.01 0 60.28 2.605 ;
      RECT 59.1 0 59.34 2.605 ;
      RECT 43.425 0 43.695 2.605 ;
      RECT 42.515 0 42.755 2.605 ;
      RECT 26.84 0 27.11 2.605 ;
      RECT 25.93 0 26.17 2.605 ;
      RECT 10.255 0 10.525 2.605 ;
      RECT 9.345 0 9.585 2.605 ;
      RECT 74.81 0 75.06 2.335 ;
      RECT 58.23 0 58.48 2.335 ;
      RECT 41.645 0 41.895 2.335 ;
      RECT 25.06 0 25.31 2.335 ;
      RECT 8.475 0 8.725 2.335 ;
      RECT 72.43 0 72.76 2.255 ;
      RECT 55.85 0 56.18 2.255 ;
      RECT 39.265 0 39.595 2.255 ;
      RECT 22.68 0 23.01 2.255 ;
      RECT 6.095 0 6.425 2.255 ;
      RECT 70.055 0 77.145 1.795 ;
      RECT 53.475 0 60.565 1.795 ;
      RECT 36.89 0 43.98 1.795 ;
      RECT 20.305 0 27.395 1.795 ;
      RECT 3.72 0 10.81 1.795 ;
      RECT 69.8 0 77.145 1.655 ;
      RECT 53.22 0 60.565 1.655 ;
      RECT 36.635 0 43.98 1.655 ;
      RECT 20.05 0 27.395 1.655 ;
      RECT 3.465 0 10.81 1.655 ;
      RECT 81.955 0 82.125 0.935 ;
      RECT 80.965 0 81.135 0.935 ;
      RECT 78.22 0 78.39 0.935 ;
      RECT 65.375 0 65.545 0.935 ;
      RECT 64.385 0 64.555 0.935 ;
      RECT 61.64 0 61.81 0.935 ;
      RECT 48.79 0 48.96 0.935 ;
      RECT 47.8 0 47.97 0.935 ;
      RECT 45.055 0 45.225 0.935 ;
      RECT 32.205 0 32.375 0.935 ;
      RECT 31.215 0 31.385 0.935 ;
      RECT 28.47 0 28.64 0.935 ;
      RECT 15.62 0 15.79 0.935 ;
      RECT 14.63 0 14.8 0.935 ;
      RECT 11.885 0 12.055 0.935 ;
      RECT -2.955 0 82.925 0.305 ;
      RECT -0.76 4.13 -0.59 8.305 ;
      RECT 81.955 3.405 82.125 5.475 ;
      RECT 80.965 3.405 81.135 5.475 ;
      RECT 78.22 3.405 78.39 5.475 ;
      RECT 66.995 4.13 67.165 5.475 ;
      RECT 65.375 3.405 65.545 5.475 ;
      RECT 64.385 3.405 64.555 5.475 ;
      RECT 61.64 3.405 61.81 5.475 ;
      RECT 50.415 4.13 50.585 5.475 ;
      RECT 48.79 3.405 48.96 5.475 ;
      RECT 47.8 3.405 47.97 5.475 ;
      RECT 45.055 3.405 45.225 5.475 ;
      RECT 33.83 4.13 34 5.475 ;
      RECT 32.205 3.405 32.375 5.475 ;
      RECT 31.215 3.405 31.385 5.475 ;
      RECT 28.47 3.405 28.64 5.475 ;
      RECT 17.245 4.13 17.415 5.475 ;
      RECT 15.62 3.405 15.79 5.475 ;
      RECT 14.63 3.405 14.8 5.475 ;
      RECT 11.885 3.405 12.055 5.475 ;
      RECT 0.66 4.13 0.83 5.475 ;
      RECT -2.57 4.13 -2.4 5.475 ;
      RECT 73.41 3.69 73.675 5.295 ;
      RECT 56.83 3.69 57.095 5.295 ;
      RECT 40.245 3.69 40.51 5.295 ;
      RECT 23.66 3.69 23.925 5.295 ;
      RECT 7.075 3.69 7.34 5.295 ;
      RECT 71.25 3.84 71.58 5.235 ;
      RECT 54.67 3.84 55 5.235 ;
      RECT 38.085 3.84 38.415 5.235 ;
      RECT 21.5 3.84 21.83 5.235 ;
      RECT 4.915 3.84 5.245 5.235 ;
      RECT 72.25 4.345 72.53 5.185 ;
      RECT 55.67 4.345 55.95 5.185 ;
      RECT 39.085 4.345 39.365 5.185 ;
      RECT 22.5 4.345 22.78 5.185 ;
      RECT 5.915 4.345 6.195 5.185 ;
      RECT 74.225 4.345 74.6 4.895 ;
      RECT 57.645 4.345 58.02 4.895 ;
      RECT 41.06 4.345 41.435 4.895 ;
      RECT 24.475 4.345 24.85 4.895 ;
      RECT 7.89 4.345 8.265 4.895 ;
      RECT 76.985 4.135 82.925 4.745 ;
      RECT 66.82 4.13 69.57 4.745 ;
      RECT 60.405 4.135 66.345 4.745 ;
      RECT 50.24 4.13 52.99 4.745 ;
      RECT 43.82 4.135 49.76 4.745 ;
      RECT 33.655 4.13 36.405 4.745 ;
      RECT 27.235 4.135 33.175 4.745 ;
      RECT 17.07 4.13 19.82 4.745 ;
      RECT 10.65 4.135 16.59 4.745 ;
      RECT 0.485 4.13 3.235 4.745 ;
      RECT -2.955 4.13 0.005 4.745 ;
      RECT 66.34 4.13 69.915 4.74 ;
      RECT 49.76 4.13 53.335 4.74 ;
      RECT 33.175 4.13 36.75 4.74 ;
      RECT 16.59 4.13 20.165 4.74 ;
      RECT -2.955 4.13 3.58 4.74 ;
      RECT 76.855 4.135 82.925 4.67 ;
      RECT 60.275 4.135 69.915 4.67 ;
      RECT 43.69 4.135 53.335 4.67 ;
      RECT 27.105 4.135 36.75 4.67 ;
      RECT 10.52 4.135 20.165 4.67 ;
      RECT -2.955 4.345 82.925 4.515 ;
      RECT 76.53 3.205 76.86 4.515 ;
      RECT 74.79 3.8 75.045 4.515 ;
      RECT 73.36 3.69 73.965 4.515 ;
      RECT 72.49 3.8 72.705 4.515 ;
      RECT 71.06 3.84 71.675 4.515 ;
      RECT 71.48 3.475 71.675 4.515 ;
      RECT 70.14 3.835 70.4 4.515 ;
      RECT 59.95 3.205 60.28 4.515 ;
      RECT 58.21 3.8 58.465 4.515 ;
      RECT 56.78 3.69 57.385 4.515 ;
      RECT 55.91 3.8 56.125 4.515 ;
      RECT 54.48 3.84 55.095 4.515 ;
      RECT 54.9 3.475 55.095 4.515 ;
      RECT 53.56 3.835 53.82 4.515 ;
      RECT 43.365 3.205 43.695 4.515 ;
      RECT 41.625 3.8 41.88 4.515 ;
      RECT 40.195 3.69 40.8 4.515 ;
      RECT 39.325 3.8 39.54 4.515 ;
      RECT 37.895 3.84 38.51 4.515 ;
      RECT 38.315 3.475 38.51 4.515 ;
      RECT 36.975 3.835 37.235 4.515 ;
      RECT 26.78 3.205 27.11 4.515 ;
      RECT 25.04 3.8 25.295 4.515 ;
      RECT 23.61 3.69 24.215 4.515 ;
      RECT 22.74 3.8 22.955 4.515 ;
      RECT 21.31 3.84 21.925 4.515 ;
      RECT 21.73 3.475 21.925 4.515 ;
      RECT 20.39 3.835 20.65 4.515 ;
      RECT 10.195 3.205 10.525 4.515 ;
      RECT 8.455 3.8 8.71 4.515 ;
      RECT 7.025 3.69 7.63 4.515 ;
      RECT 6.155 3.8 6.37 4.515 ;
      RECT 4.725 3.84 5.34 4.515 ;
      RECT 5.145 3.475 5.34 4.515 ;
      RECT 3.805 3.835 4.065 4.515 ;
      RECT 73.79 3.42 73.975 3.79 ;
      RECT 57.21 3.42 57.395 3.79 ;
      RECT 40.625 3.42 40.81 3.79 ;
      RECT 24.04 3.42 24.225 3.79 ;
      RECT 7.455 3.42 7.64 3.79 ;
      RECT 73.79 3.42 74.12 3.665 ;
      RECT 71.48 3.475 71.81 3.665 ;
      RECT 57.21 3.42 57.54 3.665 ;
      RECT 54.9 3.475 55.23 3.665 ;
      RECT 40.625 3.42 40.955 3.665 ;
      RECT 38.315 3.475 38.645 3.665 ;
      RECT 24.04 3.42 24.37 3.665 ;
      RECT 21.73 3.475 22.06 3.665 ;
      RECT 7.455 3.42 7.785 3.665 ;
      RECT 5.145 3.475 5.475 3.665 ;
      RECT -2.955 8.575 82.925 8.88 ;
      RECT 81.955 7.945 82.125 8.88 ;
      RECT 80.965 7.945 81.135 8.88 ;
      RECT 78.22 7.945 78.39 8.88 ;
      RECT 69.76 7.18 76.96 8.88 ;
      RECT 66.995 7.945 67.165 8.88 ;
      RECT 65.375 7.945 65.545 8.88 ;
      RECT 64.385 7.945 64.555 8.88 ;
      RECT 61.64 7.945 61.81 8.88 ;
      RECT 53.18 7.18 60.38 8.88 ;
      RECT 50.415 7.945 50.585 8.88 ;
      RECT 48.79 7.945 48.96 8.88 ;
      RECT 47.8 7.945 47.97 8.88 ;
      RECT 45.055 7.945 45.225 8.88 ;
      RECT 36.595 7.18 43.795 8.88 ;
      RECT 33.83 7.945 34 8.88 ;
      RECT 32.205 7.945 32.375 8.88 ;
      RECT 31.215 7.945 31.385 8.88 ;
      RECT 28.47 7.945 28.64 8.88 ;
      RECT 20.01 7.18 27.21 8.88 ;
      RECT 17.245 7.945 17.415 8.88 ;
      RECT 15.62 7.945 15.79 8.88 ;
      RECT 14.63 7.945 14.8 8.88 ;
      RECT 11.885 7.945 12.055 8.88 ;
      RECT 3.425 7.18 10.625 8.88 ;
      RECT 0.66 7.945 0.83 8.88 ;
      RECT -2.57 7.945 -2.4 8.88 ;
      RECT 70.055 7.065 76.955 8.88 ;
      RECT 53.475 7.065 60.375 8.88 ;
      RECT 36.89 7.065 43.79 8.88 ;
      RECT 20.305 7.065 27.205 8.88 ;
      RECT 3.72 7.065 10.62 8.88 ;
      RECT 75.49 6.555 75.94 8.88 ;
      RECT 73.4 6.665 73.73 8.88 ;
      RECT 71.33 6.605 71.58 8.88 ;
      RECT 58.91 6.555 59.36 8.88 ;
      RECT 56.82 6.665 57.15 8.88 ;
      RECT 54.75 6.605 55 8.88 ;
      RECT 42.325 6.555 42.775 8.88 ;
      RECT 40.235 6.665 40.565 8.88 ;
      RECT 38.165 6.605 38.415 8.88 ;
      RECT 25.74 6.555 26.19 8.88 ;
      RECT 23.65 6.665 23.98 8.88 ;
      RECT 21.58 6.605 21.83 8.88 ;
      RECT 9.155 6.555 9.605 8.88 ;
      RECT 7.065 6.665 7.395 8.88 ;
      RECT 4.995 6.605 5.245 8.88 ;
      RECT 82.015 1.74 82.185 2.935 ;
      RECT 82.015 1.74 82.48 1.91 ;
      RECT 82.015 6.97 82.48 7.14 ;
      RECT 82.015 5.945 82.185 7.14 ;
      RECT 81.025 1.74 81.195 2.935 ;
      RECT 81.025 1.74 81.49 1.91 ;
      RECT 81.025 6.97 81.49 7.14 ;
      RECT 81.025 5.945 81.195 7.14 ;
      RECT 79.17 2.635 79.34 3.865 ;
      RECT 79.225 0.855 79.395 2.805 ;
      RECT 79.17 0.575 79.34 1.025 ;
      RECT 79.17 7.855 79.34 8.305 ;
      RECT 79.225 6.075 79.395 8.025 ;
      RECT 79.17 5.015 79.34 6.245 ;
      RECT 78.65 0.575 78.82 3.865 ;
      RECT 78.65 2.075 79.055 2.405 ;
      RECT 78.65 1.235 79.055 1.565 ;
      RECT 78.65 5.015 78.82 8.305 ;
      RECT 78.65 7.315 79.055 7.645 ;
      RECT 78.65 6.475 79.055 6.805 ;
      RECT 73.91 6.645 75.215 6.895 ;
      RECT 73.91 6.325 74.09 6.895 ;
      RECT 73.36 6.325 74.09 6.495 ;
      RECT 73.36 5.485 73.53 6.495 ;
      RECT 74.195 5.525 75.94 5.705 ;
      RECT 75.61 4.685 75.94 5.705 ;
      RECT 73.36 5.485 74.42 5.655 ;
      RECT 75.61 4.855 76.43 5.025 ;
      RECT 74.77 4.685 75.1 4.895 ;
      RECT 74.77 4.685 75.94 4.855 ;
      RECT 75.67 3.205 76 4.16 ;
      RECT 75.67 3.205 76.35 3.375 ;
      RECT 76.18 1.965 76.35 3.375 ;
      RECT 76.09 1.965 76.42 2.605 ;
      RECT 75.215 3.475 75.49 4.175 ;
      RECT 75.32 1.965 75.49 4.175 ;
      RECT 75.66 2.785 76.01 3.035 ;
      RECT 75.32 2.815 76.01 2.985 ;
      RECT 75.23 1.965 75.49 2.445 ;
      RECT 74.56 5.115 75.44 5.355 ;
      RECT 75.21 5.025 75.44 5.355 ;
      RECT 73.91 5.115 75.44 5.315 ;
      RECT 74.825 5.065 75.44 5.355 ;
      RECT 73.91 4.985 74.08 5.315 ;
      RECT 74.795 5.875 75.045 6.475 ;
      RECT 74.795 5.875 75.27 6.075 ;
      RECT 74.29 3.095 75.045 3.595 ;
      RECT 73.36 2.9 73.62 3.52 ;
      RECT 74.275 3.04 74.29 3.345 ;
      RECT 74.26 3.025 74.28 3.31 ;
      RECT 74.92 2.7 75.15 3.3 ;
      RECT 74.235 2.97 74.255 3.285 ;
      RECT 74.215 3.095 75.15 3.27 ;
      RECT 74.19 3.095 75.15 3.26 ;
      RECT 74.12 3.095 75.15 3.25 ;
      RECT 74.1 3.095 75.15 3.22 ;
      RECT 74.08 2.005 74.25 3.19 ;
      RECT 74.05 3.095 75.15 3.16 ;
      RECT 74.015 3.095 75.15 3.135 ;
      RECT 73.985 3.09 74.375 3.1 ;
      RECT 73.985 3.08 74.35 3.1 ;
      RECT 73.985 3.075 74.335 3.1 ;
      RECT 73.985 3.065 74.32 3.1 ;
      RECT 73.36 2.9 74.25 3.07 ;
      RECT 73.36 3.055 74.31 3.07 ;
      RECT 73.36 3.05 74.3 3.07 ;
      RECT 74.255 2.995 74.265 3.3 ;
      RECT 73.36 3.03 74.285 3.07 ;
      RECT 73.36 3.01 74.27 3.07 ;
      RECT 73.36 2.005 74.25 2.175 ;
      RECT 74.42 2.5 74.75 2.925 ;
      RECT 74.42 2.015 74.64 2.925 ;
      RECT 74.335 5.875 74.545 6.475 ;
      RECT 74.195 5.875 74.545 6.075 ;
      RECT 72.915 3.475 73.19 4.175 ;
      RECT 73.135 1.965 73.19 4.175 ;
      RECT 73.02 2.77 73.19 4.175 ;
      RECT 73.02 1.965 73.19 2.765 ;
      RECT 72.93 1.965 73.19 2.44 ;
      RECT 71.06 3.135 71.31 3.67 ;
      RECT 72.03 3.135 72.745 3.6 ;
      RECT 71.06 3.135 72.85 3.305 ;
      RECT 72.62 2.77 72.85 3.305 ;
      RECT 71.615 2.015 71.87 3.305 ;
      RECT 72.62 2.705 72.68 3.6 ;
      RECT 72.68 2.7 72.85 2.765 ;
      RECT 71.08 2.015 71.87 2.28 ;
      RECT 72.04 5.825 72.715 6.075 ;
      RECT 72.45 5.465 72.715 6.075 ;
      RECT 72.2 6.245 72.53 6.795 ;
      RECT 71.14 6.245 72.53 6.435 ;
      RECT 71.14 5.405 71.31 6.435 ;
      RECT 71.02 5.825 71.31 6.155 ;
      RECT 71.14 5.405 72.08 5.575 ;
      RECT 71.78 4.855 72.08 5.575 ;
      RECT 72.04 2.435 72.45 2.955 ;
      RECT 72.04 2.015 72.24 2.955 ;
      RECT 70.65 2.195 70.82 4.175 ;
      RECT 70.65 2.705 71.445 2.955 ;
      RECT 70.65 2.195 70.9 2.955 ;
      RECT 70.57 2.195 70.9 2.615 ;
      RECT 70.6 6.605 71.16 6.895 ;
      RECT 70.6 4.685 70.85 6.895 ;
      RECT 70.6 4.685 71.06 5.235 ;
      RECT 67.945 7.855 68.115 8.305 ;
      RECT 68 6.075 68.17 8.025 ;
      RECT 67.945 5.015 68.115 6.245 ;
      RECT 67.425 5.015 67.595 8.305 ;
      RECT 67.425 7.315 67.83 7.645 ;
      RECT 67.425 6.475 67.83 6.805 ;
      RECT 65.435 1.74 65.605 2.935 ;
      RECT 65.435 1.74 65.9 1.91 ;
      RECT 65.435 6.97 65.9 7.14 ;
      RECT 65.435 5.945 65.605 7.14 ;
      RECT 64.445 1.74 64.615 2.935 ;
      RECT 64.445 1.74 64.91 1.91 ;
      RECT 64.445 6.97 64.91 7.14 ;
      RECT 64.445 5.945 64.615 7.14 ;
      RECT 62.59 2.635 62.76 3.865 ;
      RECT 62.645 0.855 62.815 2.805 ;
      RECT 62.59 0.575 62.76 1.025 ;
      RECT 62.59 7.855 62.76 8.305 ;
      RECT 62.645 6.075 62.815 8.025 ;
      RECT 62.59 5.015 62.76 6.245 ;
      RECT 62.07 0.575 62.24 3.865 ;
      RECT 62.07 2.075 62.475 2.405 ;
      RECT 62.07 1.235 62.475 1.565 ;
      RECT 62.07 5.015 62.24 8.305 ;
      RECT 62.07 7.315 62.475 7.645 ;
      RECT 62.07 6.475 62.475 6.805 ;
      RECT 57.33 6.645 58.635 6.895 ;
      RECT 57.33 6.325 57.51 6.895 ;
      RECT 56.78 6.325 57.51 6.495 ;
      RECT 56.78 5.485 56.95 6.495 ;
      RECT 57.615 5.525 59.36 5.705 ;
      RECT 59.03 4.685 59.36 5.705 ;
      RECT 56.78 5.485 57.84 5.655 ;
      RECT 59.03 4.855 59.85 5.025 ;
      RECT 58.19 4.685 58.52 4.895 ;
      RECT 58.19 4.685 59.36 4.855 ;
      RECT 59.09 3.205 59.42 4.16 ;
      RECT 59.09 3.205 59.77 3.375 ;
      RECT 59.6 1.965 59.77 3.375 ;
      RECT 59.51 1.965 59.84 2.605 ;
      RECT 58.635 3.475 58.91 4.175 ;
      RECT 58.74 1.965 58.91 4.175 ;
      RECT 59.08 2.785 59.43 3.035 ;
      RECT 58.74 2.815 59.43 2.985 ;
      RECT 58.65 1.965 58.91 2.445 ;
      RECT 57.98 5.115 58.86 5.355 ;
      RECT 58.63 5.025 58.86 5.355 ;
      RECT 57.33 5.115 58.86 5.315 ;
      RECT 58.245 5.065 58.86 5.355 ;
      RECT 57.33 4.985 57.5 5.315 ;
      RECT 58.215 5.875 58.465 6.475 ;
      RECT 58.215 5.875 58.69 6.075 ;
      RECT 57.71 3.095 58.465 3.595 ;
      RECT 56.78 2.9 57.04 3.52 ;
      RECT 57.695 3.04 57.71 3.345 ;
      RECT 57.68 3.025 57.7 3.31 ;
      RECT 58.34 2.7 58.57 3.3 ;
      RECT 57.655 2.97 57.675 3.285 ;
      RECT 57.635 3.095 58.57 3.27 ;
      RECT 57.61 3.095 58.57 3.26 ;
      RECT 57.54 3.095 58.57 3.25 ;
      RECT 57.52 3.095 58.57 3.22 ;
      RECT 57.5 2.005 57.67 3.19 ;
      RECT 57.47 3.095 58.57 3.16 ;
      RECT 57.435 3.095 58.57 3.135 ;
      RECT 57.405 3.09 57.795 3.1 ;
      RECT 57.405 3.08 57.77 3.1 ;
      RECT 57.405 3.075 57.755 3.1 ;
      RECT 57.405 3.065 57.74 3.1 ;
      RECT 56.78 2.9 57.67 3.07 ;
      RECT 56.78 3.055 57.73 3.07 ;
      RECT 56.78 3.05 57.72 3.07 ;
      RECT 57.675 2.995 57.685 3.3 ;
      RECT 56.78 3.03 57.705 3.07 ;
      RECT 56.78 3.01 57.69 3.07 ;
      RECT 56.78 2.005 57.67 2.175 ;
      RECT 57.84 2.5 58.17 2.925 ;
      RECT 57.84 2.015 58.06 2.925 ;
      RECT 57.755 5.875 57.965 6.475 ;
      RECT 57.615 5.875 57.965 6.075 ;
      RECT 56.335 3.475 56.61 4.175 ;
      RECT 56.555 1.965 56.61 4.175 ;
      RECT 56.44 2.77 56.61 4.175 ;
      RECT 56.44 1.965 56.61 2.765 ;
      RECT 56.35 1.965 56.61 2.44 ;
      RECT 54.48 3.135 54.73 3.67 ;
      RECT 55.45 3.135 56.165 3.6 ;
      RECT 54.48 3.135 56.27 3.305 ;
      RECT 56.04 2.77 56.27 3.305 ;
      RECT 55.035 2.015 55.29 3.305 ;
      RECT 56.04 2.705 56.1 3.6 ;
      RECT 56.1 2.7 56.27 2.765 ;
      RECT 54.5 2.015 55.29 2.28 ;
      RECT 55.46 5.825 56.135 6.075 ;
      RECT 55.87 5.465 56.135 6.075 ;
      RECT 55.62 6.245 55.95 6.795 ;
      RECT 54.56 6.245 55.95 6.435 ;
      RECT 54.56 5.405 54.73 6.435 ;
      RECT 54.44 5.825 54.73 6.155 ;
      RECT 54.56 5.405 55.5 5.575 ;
      RECT 55.2 4.855 55.5 5.575 ;
      RECT 55.46 2.435 55.87 2.955 ;
      RECT 55.46 2.015 55.66 2.955 ;
      RECT 54.07 2.195 54.24 4.175 ;
      RECT 54.07 2.705 54.865 2.955 ;
      RECT 54.07 2.195 54.32 2.955 ;
      RECT 53.99 2.195 54.32 2.615 ;
      RECT 54.02 6.605 54.58 6.895 ;
      RECT 54.02 4.685 54.27 6.895 ;
      RECT 54.02 4.685 54.48 5.235 ;
      RECT 51.365 7.855 51.535 8.305 ;
      RECT 51.42 6.075 51.59 8.025 ;
      RECT 51.365 5.015 51.535 6.245 ;
      RECT 50.845 5.015 51.015 8.305 ;
      RECT 50.845 7.315 51.25 7.645 ;
      RECT 50.845 6.475 51.25 6.805 ;
      RECT 48.85 1.74 49.02 2.935 ;
      RECT 48.85 1.74 49.315 1.91 ;
      RECT 48.85 6.97 49.315 7.14 ;
      RECT 48.85 5.945 49.02 7.14 ;
      RECT 47.86 1.74 48.03 2.935 ;
      RECT 47.86 1.74 48.325 1.91 ;
      RECT 47.86 6.97 48.325 7.14 ;
      RECT 47.86 5.945 48.03 7.14 ;
      RECT 46.005 2.635 46.175 3.865 ;
      RECT 46.06 0.855 46.23 2.805 ;
      RECT 46.005 0.575 46.175 1.025 ;
      RECT 46.005 7.855 46.175 8.305 ;
      RECT 46.06 6.075 46.23 8.025 ;
      RECT 46.005 5.015 46.175 6.245 ;
      RECT 45.485 0.575 45.655 3.865 ;
      RECT 45.485 2.075 45.89 2.405 ;
      RECT 45.485 1.235 45.89 1.565 ;
      RECT 45.485 5.015 45.655 8.305 ;
      RECT 45.485 7.315 45.89 7.645 ;
      RECT 45.485 6.475 45.89 6.805 ;
      RECT 40.745 6.645 42.05 6.895 ;
      RECT 40.745 6.325 40.925 6.895 ;
      RECT 40.195 6.325 40.925 6.495 ;
      RECT 40.195 5.485 40.365 6.495 ;
      RECT 41.03 5.525 42.775 5.705 ;
      RECT 42.445 4.685 42.775 5.705 ;
      RECT 40.195 5.485 41.255 5.655 ;
      RECT 42.445 4.855 43.265 5.025 ;
      RECT 41.605 4.685 41.935 4.895 ;
      RECT 41.605 4.685 42.775 4.855 ;
      RECT 42.505 3.205 42.835 4.16 ;
      RECT 42.505 3.205 43.185 3.375 ;
      RECT 43.015 1.965 43.185 3.375 ;
      RECT 42.925 1.965 43.255 2.605 ;
      RECT 42.05 3.475 42.325 4.175 ;
      RECT 42.155 1.965 42.325 4.175 ;
      RECT 42.495 2.785 42.845 3.035 ;
      RECT 42.155 2.815 42.845 2.985 ;
      RECT 42.065 1.965 42.325 2.445 ;
      RECT 41.395 5.115 42.275 5.355 ;
      RECT 42.045 5.025 42.275 5.355 ;
      RECT 40.745 5.115 42.275 5.315 ;
      RECT 41.66 5.065 42.275 5.355 ;
      RECT 40.745 4.985 40.915 5.315 ;
      RECT 41.63 5.875 41.88 6.475 ;
      RECT 41.63 5.875 42.105 6.075 ;
      RECT 41.125 3.095 41.88 3.595 ;
      RECT 40.195 2.9 40.455 3.52 ;
      RECT 41.11 3.04 41.125 3.345 ;
      RECT 41.095 3.025 41.115 3.31 ;
      RECT 41.755 2.7 41.985 3.3 ;
      RECT 41.07 2.97 41.09 3.285 ;
      RECT 41.05 3.095 41.985 3.27 ;
      RECT 41.025 3.095 41.985 3.26 ;
      RECT 40.955 3.095 41.985 3.25 ;
      RECT 40.935 3.095 41.985 3.22 ;
      RECT 40.915 2.005 41.085 3.19 ;
      RECT 40.885 3.095 41.985 3.16 ;
      RECT 40.85 3.095 41.985 3.135 ;
      RECT 40.82 3.09 41.21 3.1 ;
      RECT 40.82 3.08 41.185 3.1 ;
      RECT 40.82 3.075 41.17 3.1 ;
      RECT 40.82 3.065 41.155 3.1 ;
      RECT 40.195 2.9 41.085 3.07 ;
      RECT 40.195 3.055 41.145 3.07 ;
      RECT 40.195 3.05 41.135 3.07 ;
      RECT 41.09 2.995 41.1 3.3 ;
      RECT 40.195 3.03 41.12 3.07 ;
      RECT 40.195 3.01 41.105 3.07 ;
      RECT 40.195 2.005 41.085 2.175 ;
      RECT 41.255 2.5 41.585 2.925 ;
      RECT 41.255 2.015 41.475 2.925 ;
      RECT 41.17 5.875 41.38 6.475 ;
      RECT 41.03 5.875 41.38 6.075 ;
      RECT 39.75 3.475 40.025 4.175 ;
      RECT 39.97 1.965 40.025 4.175 ;
      RECT 39.855 2.77 40.025 4.175 ;
      RECT 39.855 1.965 40.025 2.765 ;
      RECT 39.765 1.965 40.025 2.44 ;
      RECT 37.895 3.135 38.145 3.67 ;
      RECT 38.865 3.135 39.58 3.6 ;
      RECT 37.895 3.135 39.685 3.305 ;
      RECT 39.455 2.77 39.685 3.305 ;
      RECT 38.45 2.015 38.705 3.305 ;
      RECT 39.455 2.705 39.515 3.6 ;
      RECT 39.515 2.7 39.685 2.765 ;
      RECT 37.915 2.015 38.705 2.28 ;
      RECT 38.875 5.825 39.55 6.075 ;
      RECT 39.285 5.465 39.55 6.075 ;
      RECT 39.035 6.245 39.365 6.795 ;
      RECT 37.975 6.245 39.365 6.435 ;
      RECT 37.975 5.405 38.145 6.435 ;
      RECT 37.855 5.825 38.145 6.155 ;
      RECT 37.975 5.405 38.915 5.575 ;
      RECT 38.615 4.855 38.915 5.575 ;
      RECT 38.875 2.435 39.285 2.955 ;
      RECT 38.875 2.015 39.075 2.955 ;
      RECT 37.485 2.195 37.655 4.175 ;
      RECT 37.485 2.705 38.28 2.955 ;
      RECT 37.485 2.195 37.735 2.955 ;
      RECT 37.405 2.195 37.735 2.615 ;
      RECT 37.435 6.605 37.995 6.895 ;
      RECT 37.435 4.685 37.685 6.895 ;
      RECT 37.435 4.685 37.895 5.235 ;
      RECT 34.78 7.855 34.95 8.305 ;
      RECT 34.835 6.075 35.005 8.025 ;
      RECT 34.78 5.015 34.95 6.245 ;
      RECT 34.26 5.015 34.43 8.305 ;
      RECT 34.26 7.315 34.665 7.645 ;
      RECT 34.26 6.475 34.665 6.805 ;
      RECT 32.265 1.74 32.435 2.935 ;
      RECT 32.265 1.74 32.73 1.91 ;
      RECT 32.265 6.97 32.73 7.14 ;
      RECT 32.265 5.945 32.435 7.14 ;
      RECT 31.275 1.74 31.445 2.935 ;
      RECT 31.275 1.74 31.74 1.91 ;
      RECT 31.275 6.97 31.74 7.14 ;
      RECT 31.275 5.945 31.445 7.14 ;
      RECT 29.42 2.635 29.59 3.865 ;
      RECT 29.475 0.855 29.645 2.805 ;
      RECT 29.42 0.575 29.59 1.025 ;
      RECT 29.42 7.855 29.59 8.305 ;
      RECT 29.475 6.075 29.645 8.025 ;
      RECT 29.42 5.015 29.59 6.245 ;
      RECT 28.9 0.575 29.07 3.865 ;
      RECT 28.9 2.075 29.305 2.405 ;
      RECT 28.9 1.235 29.305 1.565 ;
      RECT 28.9 5.015 29.07 8.305 ;
      RECT 28.9 7.315 29.305 7.645 ;
      RECT 28.9 6.475 29.305 6.805 ;
      RECT 24.16 6.645 25.465 6.895 ;
      RECT 24.16 6.325 24.34 6.895 ;
      RECT 23.61 6.325 24.34 6.495 ;
      RECT 23.61 5.485 23.78 6.495 ;
      RECT 24.445 5.525 26.19 5.705 ;
      RECT 25.86 4.685 26.19 5.705 ;
      RECT 23.61 5.485 24.67 5.655 ;
      RECT 25.86 4.855 26.68 5.025 ;
      RECT 25.02 4.685 25.35 4.895 ;
      RECT 25.02 4.685 26.19 4.855 ;
      RECT 25.92 3.205 26.25 4.16 ;
      RECT 25.92 3.205 26.6 3.375 ;
      RECT 26.43 1.965 26.6 3.375 ;
      RECT 26.34 1.965 26.67 2.605 ;
      RECT 25.465 3.475 25.74 4.175 ;
      RECT 25.57 1.965 25.74 4.175 ;
      RECT 25.91 2.785 26.26 3.035 ;
      RECT 25.57 2.815 26.26 2.985 ;
      RECT 25.48 1.965 25.74 2.445 ;
      RECT 24.81 5.115 25.69 5.355 ;
      RECT 25.46 5.025 25.69 5.355 ;
      RECT 24.16 5.115 25.69 5.315 ;
      RECT 25.075 5.065 25.69 5.355 ;
      RECT 24.16 4.985 24.33 5.315 ;
      RECT 25.045 5.875 25.295 6.475 ;
      RECT 25.045 5.875 25.52 6.075 ;
      RECT 24.54 3.095 25.295 3.595 ;
      RECT 23.61 2.9 23.87 3.52 ;
      RECT 24.525 3.04 24.54 3.345 ;
      RECT 24.51 3.025 24.53 3.31 ;
      RECT 25.17 2.7 25.4 3.3 ;
      RECT 24.485 2.97 24.505 3.285 ;
      RECT 24.465 3.095 25.4 3.27 ;
      RECT 24.44 3.095 25.4 3.26 ;
      RECT 24.37 3.095 25.4 3.25 ;
      RECT 24.35 3.095 25.4 3.22 ;
      RECT 24.33 2.005 24.5 3.19 ;
      RECT 24.3 3.095 25.4 3.16 ;
      RECT 24.265 3.095 25.4 3.135 ;
      RECT 24.235 3.09 24.625 3.1 ;
      RECT 24.235 3.08 24.6 3.1 ;
      RECT 24.235 3.075 24.585 3.1 ;
      RECT 24.235 3.065 24.57 3.1 ;
      RECT 23.61 2.9 24.5 3.07 ;
      RECT 23.61 3.055 24.56 3.07 ;
      RECT 23.61 3.05 24.55 3.07 ;
      RECT 24.505 2.995 24.515 3.3 ;
      RECT 23.61 3.03 24.535 3.07 ;
      RECT 23.61 3.01 24.52 3.07 ;
      RECT 23.61 2.005 24.5 2.175 ;
      RECT 24.67 2.5 25 2.925 ;
      RECT 24.67 2.015 24.89 2.925 ;
      RECT 24.585 5.875 24.795 6.475 ;
      RECT 24.445 5.875 24.795 6.075 ;
      RECT 23.165 3.475 23.44 4.175 ;
      RECT 23.385 1.965 23.44 4.175 ;
      RECT 23.27 2.77 23.44 4.175 ;
      RECT 23.27 1.965 23.44 2.765 ;
      RECT 23.18 1.965 23.44 2.44 ;
      RECT 21.31 3.135 21.56 3.67 ;
      RECT 22.28 3.135 22.995 3.6 ;
      RECT 21.31 3.135 23.1 3.305 ;
      RECT 22.87 2.77 23.1 3.305 ;
      RECT 21.865 2.015 22.12 3.305 ;
      RECT 22.87 2.705 22.93 3.6 ;
      RECT 22.93 2.7 23.1 2.765 ;
      RECT 21.33 2.015 22.12 2.28 ;
      RECT 22.29 5.825 22.965 6.075 ;
      RECT 22.7 5.465 22.965 6.075 ;
      RECT 22.45 6.245 22.78 6.795 ;
      RECT 21.39 6.245 22.78 6.435 ;
      RECT 21.39 5.405 21.56 6.435 ;
      RECT 21.27 5.825 21.56 6.155 ;
      RECT 21.39 5.405 22.33 5.575 ;
      RECT 22.03 4.855 22.33 5.575 ;
      RECT 22.29 2.435 22.7 2.955 ;
      RECT 22.29 2.015 22.49 2.955 ;
      RECT 20.9 2.195 21.07 4.175 ;
      RECT 20.9 2.705 21.695 2.955 ;
      RECT 20.9 2.195 21.15 2.955 ;
      RECT 20.82 2.195 21.15 2.615 ;
      RECT 20.85 6.605 21.41 6.895 ;
      RECT 20.85 4.685 21.1 6.895 ;
      RECT 20.85 4.685 21.31 5.235 ;
      RECT 18.195 7.855 18.365 8.305 ;
      RECT 18.25 6.075 18.42 8.025 ;
      RECT 18.195 5.015 18.365 6.245 ;
      RECT 17.675 5.015 17.845 8.305 ;
      RECT 17.675 7.315 18.08 7.645 ;
      RECT 17.675 6.475 18.08 6.805 ;
      RECT 15.68 1.74 15.85 2.935 ;
      RECT 15.68 1.74 16.145 1.91 ;
      RECT 15.68 6.97 16.145 7.14 ;
      RECT 15.68 5.945 15.85 7.14 ;
      RECT 14.69 1.74 14.86 2.935 ;
      RECT 14.69 1.74 15.155 1.91 ;
      RECT 14.69 6.97 15.155 7.14 ;
      RECT 14.69 5.945 14.86 7.14 ;
      RECT 12.835 2.635 13.005 3.865 ;
      RECT 12.89 0.855 13.06 2.805 ;
      RECT 12.835 0.575 13.005 1.025 ;
      RECT 12.835 7.855 13.005 8.305 ;
      RECT 12.89 6.075 13.06 8.025 ;
      RECT 12.835 5.015 13.005 6.245 ;
      RECT 12.315 0.575 12.485 3.865 ;
      RECT 12.315 2.075 12.72 2.405 ;
      RECT 12.315 1.235 12.72 1.565 ;
      RECT 12.315 5.015 12.485 8.305 ;
      RECT 12.315 7.315 12.72 7.645 ;
      RECT 12.315 6.475 12.72 6.805 ;
      RECT 7.575 6.645 8.88 6.895 ;
      RECT 7.575 6.325 7.755 6.895 ;
      RECT 7.025 6.325 7.755 6.495 ;
      RECT 7.025 5.485 7.195 6.495 ;
      RECT 7.86 5.525 9.605 5.705 ;
      RECT 9.275 4.685 9.605 5.705 ;
      RECT 7.025 5.485 8.085 5.655 ;
      RECT 9.275 4.855 10.095 5.025 ;
      RECT 8.435 4.685 8.765 4.895 ;
      RECT 8.435 4.685 9.605 4.855 ;
      RECT 9.335 3.205 9.665 4.16 ;
      RECT 9.335 3.205 10.015 3.375 ;
      RECT 9.845 1.965 10.015 3.375 ;
      RECT 9.755 1.965 10.085 2.605 ;
      RECT 8.88 3.475 9.155 4.175 ;
      RECT 8.985 1.965 9.155 4.175 ;
      RECT 9.325 2.785 9.675 3.035 ;
      RECT 8.985 2.815 9.675 2.985 ;
      RECT 8.895 1.965 9.155 2.445 ;
      RECT 8.225 5.115 9.105 5.355 ;
      RECT 8.875 5.025 9.105 5.355 ;
      RECT 7.575 5.115 9.105 5.315 ;
      RECT 8.49 5.065 9.105 5.355 ;
      RECT 7.575 4.985 7.745 5.315 ;
      RECT 8.46 5.875 8.71 6.475 ;
      RECT 8.46 5.875 8.935 6.075 ;
      RECT 7.955 3.095 8.71 3.595 ;
      RECT 7.025 2.9 7.285 3.52 ;
      RECT 7.94 3.04 7.955 3.345 ;
      RECT 7.925 3.025 7.945 3.31 ;
      RECT 8.585 2.7 8.815 3.3 ;
      RECT 7.9 2.97 7.92 3.285 ;
      RECT 7.88 3.095 8.815 3.27 ;
      RECT 7.855 3.095 8.815 3.26 ;
      RECT 7.785 3.095 8.815 3.25 ;
      RECT 7.765 3.095 8.815 3.22 ;
      RECT 7.745 2.005 7.915 3.19 ;
      RECT 7.715 3.095 8.815 3.16 ;
      RECT 7.68 3.095 8.815 3.135 ;
      RECT 7.65 3.09 8.04 3.1 ;
      RECT 7.65 3.08 8.015 3.1 ;
      RECT 7.65 3.075 8 3.1 ;
      RECT 7.65 3.065 7.985 3.1 ;
      RECT 7.025 2.9 7.915 3.07 ;
      RECT 7.025 3.055 7.975 3.07 ;
      RECT 7.025 3.05 7.965 3.07 ;
      RECT 7.92 2.995 7.93 3.3 ;
      RECT 7.025 3.03 7.95 3.07 ;
      RECT 7.025 3.01 7.935 3.07 ;
      RECT 7.025 2.005 7.915 2.175 ;
      RECT 8.085 2.5 8.415 2.925 ;
      RECT 8.085 2.015 8.305 2.925 ;
      RECT 8 5.875 8.21 6.475 ;
      RECT 7.86 5.875 8.21 6.075 ;
      RECT 6.58 3.475 6.855 4.175 ;
      RECT 6.8 1.965 6.855 4.175 ;
      RECT 6.685 2.77 6.855 4.175 ;
      RECT 6.685 1.965 6.855 2.765 ;
      RECT 6.595 1.965 6.855 2.44 ;
      RECT 4.725 3.135 4.975 3.67 ;
      RECT 5.695 3.135 6.41 3.6 ;
      RECT 4.725 3.135 6.515 3.305 ;
      RECT 6.285 2.77 6.515 3.305 ;
      RECT 5.28 2.015 5.535 3.305 ;
      RECT 6.285 2.705 6.345 3.6 ;
      RECT 6.345 2.7 6.515 2.765 ;
      RECT 4.745 2.015 5.535 2.28 ;
      RECT 5.705 5.825 6.38 6.075 ;
      RECT 6.115 5.465 6.38 6.075 ;
      RECT 5.865 6.245 6.195 6.795 ;
      RECT 4.805 6.245 6.195 6.435 ;
      RECT 4.805 5.405 4.975 6.435 ;
      RECT 4.685 5.825 4.975 6.155 ;
      RECT 4.805 5.405 5.745 5.575 ;
      RECT 5.445 4.855 5.745 5.575 ;
      RECT 5.705 2.435 6.115 2.955 ;
      RECT 5.705 2.015 5.905 2.955 ;
      RECT 4.315 2.195 4.485 4.175 ;
      RECT 4.315 2.705 5.11 2.955 ;
      RECT 4.315 2.195 4.565 2.955 ;
      RECT 4.235 2.195 4.565 2.615 ;
      RECT 4.265 6.605 4.825 6.895 ;
      RECT 4.265 4.685 4.515 6.895 ;
      RECT 4.265 4.685 4.725 5.235 ;
      RECT 1.61 7.855 1.78 8.305 ;
      RECT 1.665 6.075 1.835 8.025 ;
      RECT 1.61 5.015 1.78 6.245 ;
      RECT 1.09 5.015 1.26 8.305 ;
      RECT 1.09 7.315 1.495 7.645 ;
      RECT 1.09 6.475 1.495 6.805 ;
      RECT -1.62 7.855 -1.45 8.305 ;
      RECT -1.565 6.075 -1.395 8.025 ;
      RECT -1.62 5.015 -1.45 6.245 ;
      RECT -2.14 5.015 -1.97 8.305 ;
      RECT -2.14 7.315 -1.735 7.645 ;
      RECT -2.14 6.475 -1.735 6.805 ;
      RECT 82.385 0.575 82.555 1.085 ;
      RECT 82.385 2.395 82.555 3.865 ;
      RECT 82.385 5.015 82.555 6.485 ;
      RECT 82.385 7.795 82.555 8.305 ;
      RECT 81.395 0.575 81.565 1.085 ;
      RECT 81.395 2.395 81.565 3.865 ;
      RECT 81.395 5.015 81.565 6.485 ;
      RECT 81.395 7.795 81.565 8.305 ;
      RECT 80.03 0.575 80.2 3.865 ;
      RECT 80.03 5.015 80.2 8.305 ;
      RECT 79.6 0.575 79.77 1.085 ;
      RECT 79.6 1.655 79.77 3.865 ;
      RECT 79.6 5.015 79.77 7.225 ;
      RECT 79.6 7.795 79.77 8.305 ;
      RECT 78.23 1.66 78.4 2.935 ;
      RECT 78.23 5.945 78.4 7.22 ;
      RECT 76.52 2.785 76.87 3.035 ;
      RECT 75.46 5.875 75.91 6.385 ;
      RECT 74.14 3.835 74.62 4.175 ;
      RECT 73.7 5.825 74.025 6.155 ;
      RECT 73.36 2.345 73.91 2.73 ;
      RECT 71.845 3.835 72.32 4.175 ;
      RECT 71.48 5.825 71.82 6.075 ;
      RECT 70.14 2.785 70.48 3.665 ;
      RECT 68.805 5.015 68.975 8.305 ;
      RECT 68.375 5.015 68.545 7.225 ;
      RECT 68.375 7.795 68.545 8.305 ;
      RECT 67.005 5.945 67.175 7.22 ;
      RECT 65.805 0.575 65.975 1.085 ;
      RECT 65.805 2.395 65.975 3.865 ;
      RECT 65.805 5.015 65.975 6.485 ;
      RECT 65.805 7.795 65.975 8.305 ;
      RECT 64.815 0.575 64.985 1.085 ;
      RECT 64.815 2.395 64.985 3.865 ;
      RECT 64.815 5.015 64.985 6.485 ;
      RECT 64.815 7.795 64.985 8.305 ;
      RECT 63.45 0.575 63.62 3.865 ;
      RECT 63.45 5.015 63.62 8.305 ;
      RECT 63.02 0.575 63.19 1.085 ;
      RECT 63.02 1.655 63.19 3.865 ;
      RECT 63.02 5.015 63.19 7.225 ;
      RECT 63.02 7.795 63.19 8.305 ;
      RECT 61.65 1.66 61.82 2.935 ;
      RECT 61.65 5.945 61.82 7.22 ;
      RECT 59.94 2.785 60.29 3.035 ;
      RECT 58.88 5.875 59.33 6.385 ;
      RECT 57.56 3.835 58.04 4.175 ;
      RECT 57.12 5.825 57.445 6.155 ;
      RECT 56.78 2.345 57.33 2.73 ;
      RECT 55.265 3.835 55.74 4.175 ;
      RECT 54.9 5.825 55.24 6.075 ;
      RECT 53.56 2.785 53.9 3.665 ;
      RECT 52.225 5.015 52.395 8.305 ;
      RECT 51.795 5.015 51.965 7.225 ;
      RECT 51.795 7.795 51.965 8.305 ;
      RECT 50.425 5.945 50.595 7.22 ;
      RECT 49.22 0.575 49.39 1.085 ;
      RECT 49.22 2.395 49.39 3.865 ;
      RECT 49.22 5.015 49.39 6.485 ;
      RECT 49.22 7.795 49.39 8.305 ;
      RECT 48.23 0.575 48.4 1.085 ;
      RECT 48.23 2.395 48.4 3.865 ;
      RECT 48.23 5.015 48.4 6.485 ;
      RECT 48.23 7.795 48.4 8.305 ;
      RECT 46.865 0.575 47.035 3.865 ;
      RECT 46.865 5.015 47.035 8.305 ;
      RECT 46.435 0.575 46.605 1.085 ;
      RECT 46.435 1.655 46.605 3.865 ;
      RECT 46.435 5.015 46.605 7.225 ;
      RECT 46.435 7.795 46.605 8.305 ;
      RECT 45.065 1.66 45.235 2.935 ;
      RECT 45.065 5.945 45.235 7.22 ;
      RECT 43.355 2.785 43.705 3.035 ;
      RECT 42.295 5.875 42.745 6.385 ;
      RECT 40.975 3.835 41.455 4.175 ;
      RECT 40.535 5.825 40.86 6.155 ;
      RECT 40.195 2.345 40.745 2.73 ;
      RECT 38.68 3.835 39.155 4.175 ;
      RECT 38.315 5.825 38.655 6.075 ;
      RECT 36.975 2.785 37.315 3.665 ;
      RECT 35.64 5.015 35.81 8.305 ;
      RECT 35.21 5.015 35.38 7.225 ;
      RECT 35.21 7.795 35.38 8.305 ;
      RECT 33.84 5.945 34.01 7.22 ;
      RECT 32.635 0.575 32.805 1.085 ;
      RECT 32.635 2.395 32.805 3.865 ;
      RECT 32.635 5.015 32.805 6.485 ;
      RECT 32.635 7.795 32.805 8.305 ;
      RECT 31.645 0.575 31.815 1.085 ;
      RECT 31.645 2.395 31.815 3.865 ;
      RECT 31.645 5.015 31.815 6.485 ;
      RECT 31.645 7.795 31.815 8.305 ;
      RECT 30.28 0.575 30.45 3.865 ;
      RECT 30.28 5.015 30.45 8.305 ;
      RECT 29.85 0.575 30.02 1.085 ;
      RECT 29.85 1.655 30.02 3.865 ;
      RECT 29.85 5.015 30.02 7.225 ;
      RECT 29.85 7.795 30.02 8.305 ;
      RECT 28.48 1.66 28.65 2.935 ;
      RECT 28.48 5.945 28.65 7.22 ;
      RECT 26.77 2.785 27.12 3.035 ;
      RECT 25.71 5.875 26.16 6.385 ;
      RECT 24.39 3.835 24.87 4.175 ;
      RECT 23.95 5.825 24.275 6.155 ;
      RECT 23.61 2.345 24.16 2.73 ;
      RECT 22.095 3.835 22.57 4.175 ;
      RECT 21.73 5.825 22.07 6.075 ;
      RECT 20.39 2.785 20.73 3.665 ;
      RECT 19.055 5.015 19.225 8.305 ;
      RECT 18.625 5.015 18.795 7.225 ;
      RECT 18.625 7.795 18.795 8.305 ;
      RECT 17.255 5.945 17.425 7.22 ;
      RECT 16.05 0.575 16.22 1.085 ;
      RECT 16.05 2.395 16.22 3.865 ;
      RECT 16.05 5.015 16.22 6.485 ;
      RECT 16.05 7.795 16.22 8.305 ;
      RECT 15.06 0.575 15.23 1.085 ;
      RECT 15.06 2.395 15.23 3.865 ;
      RECT 15.06 5.015 15.23 6.485 ;
      RECT 15.06 7.795 15.23 8.305 ;
      RECT 13.695 0.575 13.865 3.865 ;
      RECT 13.695 5.015 13.865 8.305 ;
      RECT 13.265 0.575 13.435 1.085 ;
      RECT 13.265 1.655 13.435 3.865 ;
      RECT 13.265 5.015 13.435 7.225 ;
      RECT 13.265 7.795 13.435 8.305 ;
      RECT 11.895 1.66 12.065 2.935 ;
      RECT 11.895 5.945 12.065 7.22 ;
      RECT 10.185 2.785 10.535 3.035 ;
      RECT 9.125 5.875 9.575 6.385 ;
      RECT 7.805 3.835 8.285 4.175 ;
      RECT 7.365 5.825 7.69 6.155 ;
      RECT 7.025 2.345 7.575 2.73 ;
      RECT 5.51 3.835 5.985 4.175 ;
      RECT 5.145 5.825 5.485 6.075 ;
      RECT 3.805 2.785 4.145 3.665 ;
      RECT 2.47 5.015 2.64 8.305 ;
      RECT 2.04 5.015 2.21 7.225 ;
      RECT 2.04 7.795 2.21 8.305 ;
      RECT 0.67 5.945 0.84 7.22 ;
      RECT -1.19 5.015 -1.02 7.225 ;
      RECT -1.19 7.795 -1.02 8.305 ;
      RECT -2.56 5.945 -2.39 7.22 ;
  END
END sky130_osu_ring_oscillator_mpr2ca_8_b0r2

MACRO sky130_osu_ring_oscillator_mpr2ct_8_b0r1
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 3.44 0 ;
  SIZE 88.91 BY 8.88 ;
  SYMMETRY X Y R90 ;
  SITE CoreSite ;
  OBS
    LAYER met3 ;
      RECT 71.5 7.435 77.515 7.735 ;
      RECT 77.215 5.805 77.515 7.735 ;
      RECT 76.16 5.785 76.46 7.735 ;
      RECT 75.13 6.48 75.43 7.735 ;
      RECT 71.5 7.035 71.8 7.735 ;
      RECT 70.365 7 70.735 7.37 ;
      RECT 70.365 7.035 71.8 7.335 ;
      RECT 75.1 6.48 75.43 6.81 ;
      RECT 74.63 6.495 75.43 6.795 ;
      RECT 75.01 6.455 75.31 6.795 ;
      RECT 77.14 5.805 77.515 6.17 ;
      RECT 77.205 5.765 77.505 6.17 ;
      RECT 76.12 5.785 76.46 6.135 ;
      RECT 76.135 5.745 76.435 6.135 ;
      RECT 76.11 5.79 76.46 6.12 ;
      RECT 77.14 5.805 77.95 6.105 ;
      RECT 75.64 5.805 76.46 6.105 ;
      RECT 77.15 5.79 77.505 6.17 ;
      RECT 76.8 3.755 77.13 4.085 ;
      RECT 76.8 3.77 77.6 4.07 ;
      RECT 76.815 3.725 77.115 4.085 ;
      RECT 76.46 3.075 76.79 3.405 ;
      RECT 76.46 3.09 77.26 3.39 ;
      RECT 76.545 3.065 76.845 3.39 ;
      RECT 75.78 4.155 76.11 4.485 ;
      RECT 73.74 4.155 74.07 4.485 ;
      RECT 73.74 4.17 76.11 4.47 ;
      RECT 75.43 3.415 75.76 3.745 ;
      RECT 74.97 3.43 75.77 3.73 ;
      RECT 75.1 2.225 75.43 2.555 ;
      RECT 74.63 2.24 75.43 2.54 ;
      RECT 75.09 2.235 75.43 2.54 ;
      RECT 74.42 5.79 74.75 6.12 ;
      RECT 73.95 5.805 74.75 6.105 ;
      RECT 54.28 7.435 60.295 7.735 ;
      RECT 59.995 5.805 60.295 7.735 ;
      RECT 58.94 5.785 59.24 7.735 ;
      RECT 57.91 6.48 58.21 7.735 ;
      RECT 54.28 7.035 54.58 7.735 ;
      RECT 53.145 7 53.515 7.37 ;
      RECT 53.145 7.035 54.58 7.335 ;
      RECT 57.88 6.48 58.21 6.81 ;
      RECT 57.41 6.495 58.21 6.795 ;
      RECT 57.79 6.455 58.09 6.795 ;
      RECT 59.92 5.805 60.295 6.17 ;
      RECT 59.985 5.765 60.285 6.17 ;
      RECT 58.9 5.785 59.24 6.135 ;
      RECT 58.915 5.745 59.215 6.135 ;
      RECT 58.89 5.79 59.24 6.12 ;
      RECT 59.92 5.805 60.73 6.105 ;
      RECT 58.42 5.805 59.24 6.105 ;
      RECT 59.93 5.79 60.285 6.17 ;
      RECT 59.58 3.755 59.91 4.085 ;
      RECT 59.58 3.77 60.38 4.07 ;
      RECT 59.595 3.725 59.895 4.085 ;
      RECT 59.24 3.075 59.57 3.405 ;
      RECT 59.24 3.09 60.04 3.39 ;
      RECT 59.325 3.065 59.625 3.39 ;
      RECT 58.56 4.155 58.89 4.485 ;
      RECT 56.52 4.155 56.85 4.485 ;
      RECT 56.52 4.17 58.89 4.47 ;
      RECT 58.21 3.415 58.54 3.745 ;
      RECT 57.75 3.43 58.55 3.73 ;
      RECT 57.88 2.225 58.21 2.555 ;
      RECT 57.41 2.24 58.21 2.54 ;
      RECT 57.87 2.235 58.21 2.54 ;
      RECT 57.2 5.79 57.53 6.12 ;
      RECT 56.73 5.805 57.53 6.105 ;
      RECT 37.06 7.435 43.075 7.735 ;
      RECT 42.775 5.805 43.075 7.735 ;
      RECT 41.72 5.785 42.02 7.735 ;
      RECT 40.69 6.48 40.99 7.735 ;
      RECT 37.06 7.035 37.36 7.735 ;
      RECT 35.925 7 36.295 7.37 ;
      RECT 35.925 7.035 37.36 7.335 ;
      RECT 40.66 6.48 40.99 6.81 ;
      RECT 40.19 6.495 40.99 6.795 ;
      RECT 40.57 6.455 40.87 6.795 ;
      RECT 42.7 5.805 43.075 6.17 ;
      RECT 42.765 5.765 43.065 6.17 ;
      RECT 41.68 5.785 42.02 6.135 ;
      RECT 41.695 5.745 41.995 6.135 ;
      RECT 41.67 5.79 42.02 6.12 ;
      RECT 42.7 5.805 43.51 6.105 ;
      RECT 41.2 5.805 42.02 6.105 ;
      RECT 42.71 5.79 43.065 6.17 ;
      RECT 42.36 3.755 42.69 4.085 ;
      RECT 42.36 3.77 43.16 4.07 ;
      RECT 42.375 3.725 42.675 4.085 ;
      RECT 42.02 3.075 42.35 3.405 ;
      RECT 42.02 3.09 42.82 3.39 ;
      RECT 42.105 3.065 42.405 3.39 ;
      RECT 41.34 4.155 41.67 4.485 ;
      RECT 39.3 4.155 39.63 4.485 ;
      RECT 39.3 4.17 41.67 4.47 ;
      RECT 40.99 3.415 41.32 3.745 ;
      RECT 40.53 3.43 41.33 3.73 ;
      RECT 40.66 2.225 40.99 2.555 ;
      RECT 40.19 2.24 40.99 2.54 ;
      RECT 40.65 2.235 40.99 2.54 ;
      RECT 39.98 5.79 40.31 6.12 ;
      RECT 39.51 5.805 40.31 6.105 ;
      RECT 19.84 7.435 25.855 7.735 ;
      RECT 25.555 5.805 25.855 7.735 ;
      RECT 24.5 5.785 24.8 7.735 ;
      RECT 23.47 6.48 23.77 7.735 ;
      RECT 19.84 7.035 20.14 7.735 ;
      RECT 18.705 7 19.075 7.37 ;
      RECT 18.705 7.035 20.14 7.335 ;
      RECT 23.44 6.48 23.77 6.81 ;
      RECT 22.97 6.495 23.77 6.795 ;
      RECT 23.35 6.455 23.65 6.795 ;
      RECT 25.48 5.805 25.855 6.17 ;
      RECT 25.545 5.765 25.845 6.17 ;
      RECT 24.46 5.785 24.8 6.135 ;
      RECT 24.475 5.745 24.775 6.135 ;
      RECT 24.45 5.79 24.8 6.12 ;
      RECT 25.48 5.805 26.29 6.105 ;
      RECT 23.98 5.805 24.8 6.105 ;
      RECT 25.49 5.79 25.845 6.17 ;
      RECT 25.14 3.755 25.47 4.085 ;
      RECT 25.14 3.77 25.94 4.07 ;
      RECT 25.155 3.725 25.455 4.085 ;
      RECT 24.8 3.075 25.13 3.405 ;
      RECT 24.8 3.09 25.6 3.39 ;
      RECT 24.885 3.065 25.185 3.39 ;
      RECT 24.12 4.155 24.45 4.485 ;
      RECT 22.08 4.155 22.41 4.485 ;
      RECT 22.08 4.17 24.45 4.47 ;
      RECT 23.77 3.415 24.1 3.745 ;
      RECT 23.31 3.43 24.11 3.73 ;
      RECT 23.44 2.225 23.77 2.555 ;
      RECT 22.97 2.24 23.77 2.54 ;
      RECT 23.43 2.235 23.77 2.54 ;
      RECT 22.76 5.79 23.09 6.12 ;
      RECT 22.29 5.805 23.09 6.105 ;
      RECT 2.62 7.435 8.635 7.735 ;
      RECT 8.335 5.805 8.635 7.735 ;
      RECT 7.28 5.785 7.58 7.735 ;
      RECT 6.25 6.48 6.55 7.735 ;
      RECT 2.62 7.035 2.92 7.735 ;
      RECT 1.485 7 1.855 7.37 ;
      RECT 1.485 7.035 2.92 7.335 ;
      RECT 6.22 6.48 6.55 6.81 ;
      RECT 5.75 6.495 6.55 6.795 ;
      RECT 6.13 6.455 6.43 6.795 ;
      RECT 8.26 5.805 8.635 6.17 ;
      RECT 8.325 5.765 8.625 6.17 ;
      RECT 7.24 5.785 7.58 6.135 ;
      RECT 7.255 5.745 7.555 6.135 ;
      RECT 7.23 5.79 7.58 6.12 ;
      RECT 8.26 5.805 9.07 6.105 ;
      RECT 6.76 5.805 7.58 6.105 ;
      RECT 8.27 5.79 8.625 6.17 ;
      RECT 7.92 3.755 8.25 4.085 ;
      RECT 7.92 3.77 8.72 4.07 ;
      RECT 7.935 3.725 8.235 4.085 ;
      RECT 7.58 3.075 7.91 3.405 ;
      RECT 7.58 3.09 8.38 3.39 ;
      RECT 7.665 3.065 7.965 3.39 ;
      RECT 6.9 4.155 7.23 4.485 ;
      RECT 4.86 4.155 5.19 4.485 ;
      RECT 4.86 4.17 7.23 4.47 ;
      RECT 6.55 3.415 6.88 3.745 ;
      RECT 6.09 3.43 6.89 3.73 ;
      RECT 6.22 2.225 6.55 2.555 ;
      RECT 5.75 2.24 6.55 2.54 ;
      RECT 6.21 2.235 6.55 2.54 ;
      RECT 5.54 5.79 5.87 6.12 ;
      RECT 5.07 5.805 5.87 6.105 ;
    LAYER via2 ;
      RECT 77.215 5.855 77.415 6.055 ;
      RECT 76.865 3.82 77.065 4.02 ;
      RECT 76.525 3.14 76.725 3.34 ;
      RECT 76.175 5.855 76.375 6.055 ;
      RECT 75.845 4.22 76.045 4.42 ;
      RECT 75.495 3.48 75.695 3.68 ;
      RECT 75.165 2.29 75.365 2.49 ;
      RECT 75.165 6.545 75.365 6.745 ;
      RECT 74.485 5.855 74.685 6.055 ;
      RECT 73.805 4.22 74.005 4.42 ;
      RECT 70.45 7.085 70.65 7.285 ;
      RECT 59.995 5.855 60.195 6.055 ;
      RECT 59.645 3.82 59.845 4.02 ;
      RECT 59.305 3.14 59.505 3.34 ;
      RECT 58.955 5.855 59.155 6.055 ;
      RECT 58.625 4.22 58.825 4.42 ;
      RECT 58.275 3.48 58.475 3.68 ;
      RECT 57.945 2.29 58.145 2.49 ;
      RECT 57.945 6.545 58.145 6.745 ;
      RECT 57.265 5.855 57.465 6.055 ;
      RECT 56.585 4.22 56.785 4.42 ;
      RECT 53.23 7.085 53.43 7.285 ;
      RECT 42.775 5.855 42.975 6.055 ;
      RECT 42.425 3.82 42.625 4.02 ;
      RECT 42.085 3.14 42.285 3.34 ;
      RECT 41.735 5.855 41.935 6.055 ;
      RECT 41.405 4.22 41.605 4.42 ;
      RECT 41.055 3.48 41.255 3.68 ;
      RECT 40.725 2.29 40.925 2.49 ;
      RECT 40.725 6.545 40.925 6.745 ;
      RECT 40.045 5.855 40.245 6.055 ;
      RECT 39.365 4.22 39.565 4.42 ;
      RECT 36.01 7.085 36.21 7.285 ;
      RECT 25.555 5.855 25.755 6.055 ;
      RECT 25.205 3.82 25.405 4.02 ;
      RECT 24.865 3.14 25.065 3.34 ;
      RECT 24.515 5.855 24.715 6.055 ;
      RECT 24.185 4.22 24.385 4.42 ;
      RECT 23.835 3.48 24.035 3.68 ;
      RECT 23.505 2.29 23.705 2.49 ;
      RECT 23.505 6.545 23.705 6.745 ;
      RECT 22.825 5.855 23.025 6.055 ;
      RECT 22.145 4.22 22.345 4.42 ;
      RECT 18.79 7.085 18.99 7.285 ;
      RECT 8.335 5.855 8.535 6.055 ;
      RECT 7.985 3.82 8.185 4.02 ;
      RECT 7.645 3.14 7.845 3.34 ;
      RECT 7.295 5.855 7.495 6.055 ;
      RECT 6.965 4.22 7.165 4.42 ;
      RECT 6.615 3.48 6.815 3.68 ;
      RECT 6.285 2.29 6.485 2.49 ;
      RECT 6.285 6.545 6.485 6.745 ;
      RECT 5.605 5.855 5.805 6.055 ;
      RECT 4.925 4.22 5.125 4.42 ;
      RECT 1.57 7.085 1.77 7.285 ;
    LAYER met2 ;
      RECT -2.21 8.6 85.1 8.77 ;
      RECT 84.93 7.3 85.1 8.77 ;
      RECT -2.21 6.255 -2.04 8.77 ;
      RECT 84.895 7.3 85.22 7.625 ;
      RECT -2.265 6.255 -1.985 6.595 ;
      RECT 81.74 6.28 82.06 6.605 ;
      RECT 81.77 5.695 81.94 6.605 ;
      RECT 81.77 5.695 81.945 6.045 ;
      RECT 81.77 5.695 82.745 5.87 ;
      RECT 82.57 1.965 82.745 5.87 ;
      RECT 76.485 3.055 76.765 3.425 ;
      RECT 76.555 2.345 76.73 3.425 ;
      RECT 76.555 2.345 79.775 2.52 ;
      RECT 79.6 2.025 79.775 2.52 ;
      RECT 80.07 1.995 80.395 2.32 ;
      RECT 82.515 1.965 82.865 2.315 ;
      RECT 79.6 2.025 82.865 2.195 ;
      RECT 70.89 8.29 81.585 8.46 ;
      RECT 81.425 2.395 81.585 8.46 ;
      RECT 70.89 6.545 71.06 8.46 ;
      RECT 82.54 6.655 82.865 6.98 ;
      RECT 67.71 6.655 68.035 6.98 ;
      RECT 81.425 6.745 82.865 6.915 ;
      RECT 70.84 6.545 71.12 6.885 ;
      RECT 67.71 6.685 71.12 6.855 ;
      RECT 81.74 2.365 82.06 2.685 ;
      RECT 81.425 2.395 82.06 2.565 ;
      RECT 71.395 7.55 80.945 7.72 ;
      RECT 80.775 5.855 80.945 7.72 ;
      RECT 71.395 5.86 71.565 7.72 ;
      RECT 71.34 5.86 71.62 6.2 ;
      RECT 80.695 5.855 81.02 6.18 ;
      RECT 80.765 3.495 80.935 6.18 ;
      RECT 80.695 3.495 81.02 3.82 ;
      RECT 78.195 6.48 78.455 6.8 ;
      RECT 78.255 2.74 78.395 6.8 ;
      RECT 78.195 2.74 78.455 3.06 ;
      RECT 77.515 4.78 77.775 5.1 ;
      RECT 77.575 3.76 77.715 5.1 ;
      RECT 77.515 3.76 77.775 4.08 ;
      RECT 76.495 6.48 76.755 6.8 ;
      RECT 76.555 5.21 76.695 6.8 ;
      RECT 75.875 5.21 76.695 5.35 ;
      RECT 75.875 2.74 76.015 5.35 ;
      RECT 75.805 4.135 76.085 4.505 ;
      RECT 75.815 2.74 76.075 3.06 ;
      RECT 73.765 4.135 74.045 4.505 ;
      RECT 73.835 2.4 73.975 4.505 ;
      RECT 73.775 2.4 74.035 2.72 ;
      RECT 73.095 4.78 73.355 5.1 ;
      RECT 73.155 2.74 73.295 5.1 ;
      RECT 73.095 2.74 73.355 3.06 ;
      RECT 64.52 6.28 64.84 6.605 ;
      RECT 64.55 5.695 64.72 6.605 ;
      RECT 64.55 5.695 64.725 6.045 ;
      RECT 64.55 5.695 65.525 5.87 ;
      RECT 65.35 1.965 65.525 5.87 ;
      RECT 59.265 3.055 59.545 3.425 ;
      RECT 59.335 2.345 59.51 3.425 ;
      RECT 59.335 2.345 62.555 2.52 ;
      RECT 62.38 2.025 62.555 2.52 ;
      RECT 62.85 1.995 63.175 2.32 ;
      RECT 65.295 1.965 65.645 2.315 ;
      RECT 62.38 2.025 65.645 2.195 ;
      RECT 53.67 8.29 64.365 8.46 ;
      RECT 64.205 2.395 64.365 8.46 ;
      RECT 53.67 6.545 53.84 8.46 ;
      RECT 65.32 6.655 65.645 6.98 ;
      RECT 50.49 6.655 50.815 6.98 ;
      RECT 64.205 6.745 65.645 6.915 ;
      RECT 53.62 6.545 53.9 6.885 ;
      RECT 50.49 6.685 53.9 6.855 ;
      RECT 64.52 2.365 64.84 2.685 ;
      RECT 64.205 2.395 64.84 2.565 ;
      RECT 54.175 7.55 63.725 7.72 ;
      RECT 63.555 5.855 63.725 7.72 ;
      RECT 54.175 5.86 54.345 7.72 ;
      RECT 54.12 5.86 54.4 6.2 ;
      RECT 63.475 5.855 63.8 6.18 ;
      RECT 63.545 3.495 63.715 6.18 ;
      RECT 63.475 3.495 63.8 3.82 ;
      RECT 60.975 6.48 61.235 6.8 ;
      RECT 61.035 2.74 61.175 6.8 ;
      RECT 60.975 2.74 61.235 3.06 ;
      RECT 60.295 4.78 60.555 5.1 ;
      RECT 60.355 3.76 60.495 5.1 ;
      RECT 60.295 3.76 60.555 4.08 ;
      RECT 59.275 6.48 59.535 6.8 ;
      RECT 59.335 5.21 59.475 6.8 ;
      RECT 58.655 5.21 59.475 5.35 ;
      RECT 58.655 2.74 58.795 5.35 ;
      RECT 58.585 4.135 58.865 4.505 ;
      RECT 58.595 2.74 58.855 3.06 ;
      RECT 56.545 4.135 56.825 4.505 ;
      RECT 56.615 2.4 56.755 4.505 ;
      RECT 56.555 2.4 56.815 2.72 ;
      RECT 55.875 4.78 56.135 5.1 ;
      RECT 55.935 2.74 56.075 5.1 ;
      RECT 55.875 2.74 56.135 3.06 ;
      RECT 47.3 6.28 47.62 6.605 ;
      RECT 47.33 5.695 47.5 6.605 ;
      RECT 47.33 5.695 47.505 6.045 ;
      RECT 47.33 5.695 48.305 5.87 ;
      RECT 48.13 1.965 48.305 5.87 ;
      RECT 42.045 3.055 42.325 3.425 ;
      RECT 42.115 2.345 42.29 3.425 ;
      RECT 42.115 2.345 45.335 2.52 ;
      RECT 45.16 2.025 45.335 2.52 ;
      RECT 45.63 1.995 45.955 2.32 ;
      RECT 48.075 1.965 48.425 2.315 ;
      RECT 45.16 2.025 48.425 2.195 ;
      RECT 36.45 8.29 47.145 8.46 ;
      RECT 46.985 2.395 47.145 8.46 ;
      RECT 36.45 6.545 36.62 8.46 ;
      RECT 48.1 6.655 48.425 6.98 ;
      RECT 33.27 6.655 33.595 6.98 ;
      RECT 46.985 6.745 48.425 6.915 ;
      RECT 36.4 6.545 36.68 6.885 ;
      RECT 33.27 6.685 36.69 6.855 ;
      RECT 47.3 2.365 47.62 2.685 ;
      RECT 46.985 2.395 47.62 2.565 ;
      RECT 36.955 7.55 46.505 7.72 ;
      RECT 46.335 5.855 46.505 7.72 ;
      RECT 36.955 5.86 37.125 7.72 ;
      RECT 36.9 5.86 37.18 6.2 ;
      RECT 46.255 5.855 46.58 6.18 ;
      RECT 46.325 3.495 46.495 6.18 ;
      RECT 46.255 3.495 46.58 3.82 ;
      RECT 43.755 6.48 44.015 6.8 ;
      RECT 43.815 2.74 43.955 6.8 ;
      RECT 43.755 2.74 44.015 3.06 ;
      RECT 43.075 4.78 43.335 5.1 ;
      RECT 43.135 3.76 43.275 5.1 ;
      RECT 43.075 3.76 43.335 4.08 ;
      RECT 42.055 6.48 42.315 6.8 ;
      RECT 42.115 5.21 42.255 6.8 ;
      RECT 41.435 5.21 42.255 5.35 ;
      RECT 41.435 2.74 41.575 5.35 ;
      RECT 41.365 4.135 41.645 4.505 ;
      RECT 41.375 2.74 41.635 3.06 ;
      RECT 39.325 4.135 39.605 4.505 ;
      RECT 39.395 2.4 39.535 4.505 ;
      RECT 39.335 2.4 39.595 2.72 ;
      RECT 38.655 4.78 38.915 5.1 ;
      RECT 38.715 2.74 38.855 5.1 ;
      RECT 38.655 2.74 38.915 3.06 ;
      RECT 30.08 6.28 30.4 6.605 ;
      RECT 30.11 5.695 30.28 6.605 ;
      RECT 30.11 5.695 30.285 6.045 ;
      RECT 30.11 5.695 31.085 5.87 ;
      RECT 30.91 1.965 31.085 5.87 ;
      RECT 24.825 3.055 25.105 3.425 ;
      RECT 24.895 2.345 25.07 3.425 ;
      RECT 24.895 2.345 28.115 2.52 ;
      RECT 27.94 2.025 28.115 2.52 ;
      RECT 28.41 1.995 28.735 2.32 ;
      RECT 30.855 1.965 31.205 2.315 ;
      RECT 27.94 2.025 31.205 2.195 ;
      RECT 19.23 8.29 29.925 8.46 ;
      RECT 29.765 2.395 29.925 8.46 ;
      RECT 19.23 6.545 19.4 8.46 ;
      RECT 30.88 6.655 31.205 6.98 ;
      RECT 16.05 6.655 16.375 6.98 ;
      RECT 29.765 6.745 31.205 6.915 ;
      RECT 19.18 6.545 19.46 6.885 ;
      RECT 16.05 6.685 19.46 6.855 ;
      RECT 30.08 2.365 30.4 2.685 ;
      RECT 29.765 2.395 30.4 2.565 ;
      RECT 19.735 7.55 29.285 7.72 ;
      RECT 29.115 5.855 29.285 7.72 ;
      RECT 19.735 5.86 19.905 7.72 ;
      RECT 19.68 5.86 19.96 6.2 ;
      RECT 29.035 5.855 29.36 6.18 ;
      RECT 29.105 3.495 29.275 6.18 ;
      RECT 29.035 3.495 29.36 3.82 ;
      RECT 26.535 6.48 26.795 6.8 ;
      RECT 26.595 2.74 26.735 6.8 ;
      RECT 26.535 2.74 26.795 3.06 ;
      RECT 25.855 4.78 26.115 5.1 ;
      RECT 25.915 3.76 26.055 5.1 ;
      RECT 25.855 3.76 26.115 4.08 ;
      RECT 24.835 6.48 25.095 6.8 ;
      RECT 24.895 5.21 25.035 6.8 ;
      RECT 24.215 5.21 25.035 5.35 ;
      RECT 24.215 2.74 24.355 5.35 ;
      RECT 24.145 4.135 24.425 4.505 ;
      RECT 24.155 2.74 24.415 3.06 ;
      RECT 22.105 4.135 22.385 4.505 ;
      RECT 22.175 2.4 22.315 4.505 ;
      RECT 22.115 2.4 22.375 2.72 ;
      RECT 21.435 4.78 21.695 5.1 ;
      RECT 21.495 2.74 21.635 5.1 ;
      RECT 21.435 2.74 21.695 3.06 ;
      RECT 12.86 6.28 13.18 6.605 ;
      RECT 12.89 5.695 13.06 6.605 ;
      RECT 12.89 5.695 13.065 6.045 ;
      RECT 12.89 5.695 13.865 5.87 ;
      RECT 13.69 1.965 13.865 5.87 ;
      RECT 7.605 3.055 7.885 3.425 ;
      RECT 7.675 2.345 7.85 3.425 ;
      RECT 7.675 2.345 10.895 2.52 ;
      RECT 10.72 2.025 10.895 2.52 ;
      RECT 11.19 1.995 11.515 2.32 ;
      RECT 13.635 1.965 13.985 2.315 ;
      RECT 10.72 2.025 13.985 2.195 ;
      RECT 2.01 8.29 12.705 8.46 ;
      RECT 12.545 2.395 12.705 8.46 ;
      RECT 2.01 6.545 2.18 8.46 ;
      RECT -1.89 6.995 -1.61 7.335 ;
      RECT -1.89 7.06 -0.68 7.23 ;
      RECT -0.85 6.685 -0.68 7.23 ;
      RECT 13.66 6.655 13.985 6.98 ;
      RECT 12.545 6.745 13.985 6.915 ;
      RECT 1.96 6.545 2.24 6.885 ;
      RECT -0.85 6.685 2.24 6.855 ;
      RECT 12.86 2.365 13.18 2.685 ;
      RECT 12.545 2.395 13.18 2.565 ;
      RECT 2.515 7.55 12.065 7.72 ;
      RECT 11.895 5.855 12.065 7.72 ;
      RECT 2.515 5.86 2.685 7.72 ;
      RECT 2.46 5.86 2.74 6.2 ;
      RECT 11.815 5.855 12.14 6.18 ;
      RECT 11.885 3.495 12.055 6.18 ;
      RECT 11.815 3.495 12.14 3.82 ;
      RECT 9.315 6.48 9.575 6.8 ;
      RECT 9.375 2.74 9.515 6.8 ;
      RECT 9.315 2.74 9.575 3.06 ;
      RECT 8.635 4.78 8.895 5.1 ;
      RECT 8.695 3.76 8.835 5.1 ;
      RECT 8.635 3.76 8.895 4.08 ;
      RECT 7.615 6.48 7.875 6.8 ;
      RECT 7.675 5.21 7.815 6.8 ;
      RECT 6.995 5.21 7.815 5.35 ;
      RECT 6.995 2.74 7.135 5.35 ;
      RECT 6.925 4.135 7.205 4.505 ;
      RECT 6.935 2.74 7.195 3.06 ;
      RECT 4.885 4.135 5.165 4.505 ;
      RECT 4.955 2.4 5.095 4.505 ;
      RECT 4.895 2.4 5.155 2.72 ;
      RECT 4.215 4.78 4.475 5.1 ;
      RECT 4.275 2.74 4.415 5.1 ;
      RECT 4.215 2.74 4.475 3.06 ;
      RECT 77.175 5.77 77.455 6.14 ;
      RECT 76.825 3.735 77.105 4.105 ;
      RECT 76.135 5.77 76.415 6.14 ;
      RECT 75.455 3.395 75.735 3.765 ;
      RECT 75.125 2.205 75.405 2.575 ;
      RECT 75.125 6.46 75.405 6.83 ;
      RECT 74.445 5.77 74.725 6.14 ;
      RECT 70.365 7 70.735 7.37 ;
      RECT 59.955 5.77 60.235 6.14 ;
      RECT 59.605 3.735 59.885 4.105 ;
      RECT 58.915 5.77 59.195 6.14 ;
      RECT 58.235 3.395 58.515 3.765 ;
      RECT 57.905 2.205 58.185 2.575 ;
      RECT 57.905 6.46 58.185 6.83 ;
      RECT 57.225 5.77 57.505 6.14 ;
      RECT 53.145 7 53.515 7.37 ;
      RECT 42.735 5.77 43.015 6.14 ;
      RECT 42.385 3.735 42.665 4.105 ;
      RECT 41.695 5.77 41.975 6.14 ;
      RECT 41.015 3.395 41.295 3.765 ;
      RECT 40.685 2.205 40.965 2.575 ;
      RECT 40.685 6.46 40.965 6.83 ;
      RECT 40.005 5.77 40.285 6.14 ;
      RECT 35.925 7 36.295 7.37 ;
      RECT 25.515 5.77 25.795 6.14 ;
      RECT 25.165 3.735 25.445 4.105 ;
      RECT 24.475 5.77 24.755 6.14 ;
      RECT 23.795 3.395 24.075 3.765 ;
      RECT 23.465 2.205 23.745 2.575 ;
      RECT 23.465 6.46 23.745 6.83 ;
      RECT 22.785 5.77 23.065 6.14 ;
      RECT 18.705 7 19.075 7.37 ;
      RECT 8.295 5.77 8.575 6.14 ;
      RECT 7.945 3.735 8.225 4.105 ;
      RECT 7.255 5.77 7.535 6.14 ;
      RECT 6.575 3.395 6.855 3.765 ;
      RECT 6.245 2.205 6.525 2.575 ;
      RECT 6.245 6.46 6.525 6.83 ;
      RECT 5.565 5.77 5.845 6.14 ;
      RECT 1.485 7 1.855 7.37 ;
    LAYER via1 ;
      RECT 84.985 7.385 85.135 7.535 ;
      RECT 82.63 6.74 82.78 6.89 ;
      RECT 82.615 2.065 82.765 2.215 ;
      RECT 81.825 2.45 81.975 2.6 ;
      RECT 81.825 6.37 81.975 6.52 ;
      RECT 80.785 3.58 80.935 3.73 ;
      RECT 80.785 5.94 80.935 6.09 ;
      RECT 80.16 2.08 80.31 2.23 ;
      RECT 78.25 2.825 78.4 2.975 ;
      RECT 78.25 6.565 78.4 6.715 ;
      RECT 77.57 3.845 77.72 3.995 ;
      RECT 77.57 4.865 77.72 5.015 ;
      RECT 77.23 5.885 77.38 6.035 ;
      RECT 76.89 3.845 77.04 3.995 ;
      RECT 76.55 3.165 76.7 3.315 ;
      RECT 76.55 6.565 76.7 6.715 ;
      RECT 76.2 5.885 76.35 6.035 ;
      RECT 75.87 2.825 76.02 2.975 ;
      RECT 75.53 3.505 75.68 3.655 ;
      RECT 75.19 2.315 75.34 2.465 ;
      RECT 75.19 6.565 75.34 6.715 ;
      RECT 74.51 5.885 74.66 6.035 ;
      RECT 73.83 2.485 73.98 2.635 ;
      RECT 73.15 2.825 73.3 2.975 ;
      RECT 73.15 4.865 73.3 5.015 ;
      RECT 71.405 5.955 71.555 6.105 ;
      RECT 70.905 6.64 71.055 6.79 ;
      RECT 70.475 7.11 70.625 7.26 ;
      RECT 67.8 6.74 67.95 6.89 ;
      RECT 65.41 6.74 65.56 6.89 ;
      RECT 65.395 2.065 65.545 2.215 ;
      RECT 64.605 2.45 64.755 2.6 ;
      RECT 64.605 6.37 64.755 6.52 ;
      RECT 63.565 3.58 63.715 3.73 ;
      RECT 63.565 5.94 63.715 6.09 ;
      RECT 62.94 2.08 63.09 2.23 ;
      RECT 61.03 2.825 61.18 2.975 ;
      RECT 61.03 6.565 61.18 6.715 ;
      RECT 60.35 3.845 60.5 3.995 ;
      RECT 60.35 4.865 60.5 5.015 ;
      RECT 60.01 5.885 60.16 6.035 ;
      RECT 59.67 3.845 59.82 3.995 ;
      RECT 59.33 3.165 59.48 3.315 ;
      RECT 59.33 6.565 59.48 6.715 ;
      RECT 58.98 5.885 59.13 6.035 ;
      RECT 58.65 2.825 58.8 2.975 ;
      RECT 58.31 3.505 58.46 3.655 ;
      RECT 57.97 2.315 58.12 2.465 ;
      RECT 57.97 6.565 58.12 6.715 ;
      RECT 57.29 5.885 57.44 6.035 ;
      RECT 56.61 2.485 56.76 2.635 ;
      RECT 55.93 2.825 56.08 2.975 ;
      RECT 55.93 4.865 56.08 5.015 ;
      RECT 54.185 5.955 54.335 6.105 ;
      RECT 53.685 6.64 53.835 6.79 ;
      RECT 53.255 7.11 53.405 7.26 ;
      RECT 50.58 6.74 50.73 6.89 ;
      RECT 48.19 6.74 48.34 6.89 ;
      RECT 48.175 2.065 48.325 2.215 ;
      RECT 47.385 2.45 47.535 2.6 ;
      RECT 47.385 6.37 47.535 6.52 ;
      RECT 46.345 3.58 46.495 3.73 ;
      RECT 46.345 5.94 46.495 6.09 ;
      RECT 45.72 2.08 45.87 2.23 ;
      RECT 43.81 2.825 43.96 2.975 ;
      RECT 43.81 6.565 43.96 6.715 ;
      RECT 43.13 3.845 43.28 3.995 ;
      RECT 43.13 4.865 43.28 5.015 ;
      RECT 42.79 5.885 42.94 6.035 ;
      RECT 42.45 3.845 42.6 3.995 ;
      RECT 42.11 3.165 42.26 3.315 ;
      RECT 42.11 6.565 42.26 6.715 ;
      RECT 41.76 5.885 41.91 6.035 ;
      RECT 41.43 2.825 41.58 2.975 ;
      RECT 41.09 3.505 41.24 3.655 ;
      RECT 40.75 2.315 40.9 2.465 ;
      RECT 40.75 6.565 40.9 6.715 ;
      RECT 40.07 5.885 40.22 6.035 ;
      RECT 39.39 2.485 39.54 2.635 ;
      RECT 38.71 2.825 38.86 2.975 ;
      RECT 38.71 4.865 38.86 5.015 ;
      RECT 36.965 5.955 37.115 6.105 ;
      RECT 36.465 6.64 36.615 6.79 ;
      RECT 36.035 7.11 36.185 7.26 ;
      RECT 33.36 6.74 33.51 6.89 ;
      RECT 30.97 6.74 31.12 6.89 ;
      RECT 30.955 2.065 31.105 2.215 ;
      RECT 30.165 2.45 30.315 2.6 ;
      RECT 30.165 6.37 30.315 6.52 ;
      RECT 29.125 3.58 29.275 3.73 ;
      RECT 29.125 5.94 29.275 6.09 ;
      RECT 28.5 2.08 28.65 2.23 ;
      RECT 26.59 2.825 26.74 2.975 ;
      RECT 26.59 6.565 26.74 6.715 ;
      RECT 25.91 3.845 26.06 3.995 ;
      RECT 25.91 4.865 26.06 5.015 ;
      RECT 25.57 5.885 25.72 6.035 ;
      RECT 25.23 3.845 25.38 3.995 ;
      RECT 24.89 3.165 25.04 3.315 ;
      RECT 24.89 6.565 25.04 6.715 ;
      RECT 24.54 5.885 24.69 6.035 ;
      RECT 24.21 2.825 24.36 2.975 ;
      RECT 23.87 3.505 24.02 3.655 ;
      RECT 23.53 2.315 23.68 2.465 ;
      RECT 23.53 6.565 23.68 6.715 ;
      RECT 22.85 5.885 23 6.035 ;
      RECT 22.17 2.485 22.32 2.635 ;
      RECT 21.49 2.825 21.64 2.975 ;
      RECT 21.49 4.865 21.64 5.015 ;
      RECT 19.745 5.955 19.895 6.105 ;
      RECT 19.245 6.64 19.395 6.79 ;
      RECT 18.815 7.11 18.965 7.26 ;
      RECT 16.14 6.74 16.29 6.89 ;
      RECT 13.75 6.74 13.9 6.89 ;
      RECT 13.735 2.065 13.885 2.215 ;
      RECT 12.945 2.45 13.095 2.6 ;
      RECT 12.945 6.37 13.095 6.52 ;
      RECT 11.905 3.58 12.055 3.73 ;
      RECT 11.905 5.94 12.055 6.09 ;
      RECT 11.28 2.08 11.43 2.23 ;
      RECT 9.37 2.825 9.52 2.975 ;
      RECT 9.37 6.565 9.52 6.715 ;
      RECT 8.69 3.845 8.84 3.995 ;
      RECT 8.69 4.865 8.84 5.015 ;
      RECT 8.35 5.885 8.5 6.035 ;
      RECT 8.01 3.845 8.16 3.995 ;
      RECT 7.67 3.165 7.82 3.315 ;
      RECT 7.67 6.565 7.82 6.715 ;
      RECT 7.32 5.885 7.47 6.035 ;
      RECT 6.99 2.825 7.14 2.975 ;
      RECT 6.65 3.505 6.8 3.655 ;
      RECT 6.31 2.315 6.46 2.465 ;
      RECT 6.31 6.565 6.46 6.715 ;
      RECT 5.63 5.885 5.78 6.035 ;
      RECT 4.95 2.485 5.1 2.635 ;
      RECT 4.27 2.825 4.42 2.975 ;
      RECT 4.27 4.865 4.42 5.015 ;
      RECT 2.525 5.955 2.675 6.105 ;
      RECT 2.025 6.64 2.175 6.79 ;
      RECT 1.595 7.11 1.745 7.26 ;
      RECT -1.825 7.09 -1.675 7.24 ;
      RECT -2.2 6.35 -2.05 6.5 ;
    LAYER met1 ;
      RECT 72.035 0 79.395 1.95 ;
      RECT 54.815 0 62.175 1.95 ;
      RECT 37.595 0 44.955 1.95 ;
      RECT 20.375 0 27.735 1.95 ;
      RECT 3.155 0 10.515 1.95 ;
      RECT 72.035 0 79.69 1.795 ;
      RECT 54.815 0 62.47 1.795 ;
      RECT 37.595 0 45.25 1.795 ;
      RECT 20.375 0 28.03 1.795 ;
      RECT 3.155 0 10.81 1.795 ;
      RECT 72.03 0 79.69 1.635 ;
      RECT 54.81 0 62.47 1.635 ;
      RECT 37.59 0 45.25 1.635 ;
      RECT 20.37 0 28.03 1.635 ;
      RECT 3.15 0 10.81 1.635 ;
      RECT -3.385 0 85.47 0.305 ;
      RECT 79.485 4.135 85.47 4.745 ;
      RECT 68.905 4.13 71.655 4.745 ;
      RECT 62.265 4.135 68.25 4.745 ;
      RECT 51.685 4.13 54.435 4.745 ;
      RECT 45.045 4.135 51.03 4.745 ;
      RECT 34.465 4.13 37.215 4.745 ;
      RECT 27.825 4.135 33.81 4.745 ;
      RECT 17.245 4.13 19.995 4.745 ;
      RECT 10.605 4.135 16.59 4.745 ;
      RECT 0.025 4.13 2.775 4.745 ;
      RECT -3.385 4.13 -0.635 4.745 ;
      RECT 62.265 4.19 72.41 4.74 ;
      RECT 45.045 4.19 55.19 4.74 ;
      RECT 27.825 4.19 37.97 4.74 ;
      RECT 10.605 4.19 20.75 4.74 ;
      RECT -3.385 4.19 3.53 4.74 ;
      RECT -3.385 4.19 85.47 4.67 ;
      RECT 79.48 4.135 85.47 4.67 ;
      RECT 62.26 4.135 72.39 4.67 ;
      RECT 68.245 4.13 72.39 4.74 ;
      RECT 45.04 4.135 55.17 4.67 ;
      RECT 51.025 4.13 55.17 4.74 ;
      RECT 27.82 4.135 37.95 4.67 ;
      RECT 33.805 4.13 37.95 4.74 ;
      RECT 10.6 4.135 20.73 4.67 ;
      RECT 16.585 4.13 20.73 4.74 ;
      RECT -3.385 4.13 3.51 4.74 ;
      RECT -3.385 8.575 85.47 8.88 ;
      RECT 72.305 7.18 79.505 8.88 ;
      RECT 69.625 6.315 69.795 8.88 ;
      RECT 55.085 7.18 62.285 8.88 ;
      RECT 52.405 6.315 52.575 8.88 ;
      RECT 37.865 7.18 45.065 8.88 ;
      RECT 35.185 6.315 35.355 8.88 ;
      RECT 20.645 7.18 27.845 8.88 ;
      RECT 17.965 6.315 18.135 8.88 ;
      RECT 3.425 7.18 10.625 8.88 ;
      RECT 0.745 6.315 0.915 8.88 ;
      RECT 72.035 6.91 79.395 7.39 ;
      RECT 54.815 6.91 62.175 7.39 ;
      RECT 37.595 6.91 44.955 7.39 ;
      RECT 20.375 6.91 27.735 7.39 ;
      RECT 3.155 6.91 10.515 7.39 ;
      RECT 70.025 6.285 70.315 6.515 ;
      RECT 52.805 6.285 53.095 6.515 ;
      RECT 35.585 6.285 35.875 6.515 ;
      RECT 18.365 6.285 18.655 6.515 ;
      RECT 1.145 6.285 1.435 6.515 ;
      RECT 69.625 6.315 70.315 6.485 ;
      RECT 52.405 6.315 53.095 6.485 ;
      RECT 35.185 6.315 35.875 6.485 ;
      RECT 17.965 6.315 18.655 6.485 ;
      RECT 0.745 6.315 1.435 6.485 ;
      RECT 84.87 7.765 85.16 7.995 ;
      RECT 84.93 6.285 85.1 7.995 ;
      RECT 84.895 7.3 85.22 7.625 ;
      RECT 84.87 6.285 85.16 6.515 ;
      RECT 84.87 2.365 85.16 2.595 ;
      RECT 84.93 0.885 85.1 2.595 ;
      RECT 84.87 0.885 85.16 1.115 ;
      RECT 84.46 2.735 84.79 2.965 ;
      RECT 84.46 2.765 84.96 2.935 ;
      RECT 84.46 2.395 84.65 2.965 ;
      RECT 83.88 2.365 84.17 2.595 ;
      RECT 83.88 2.395 84.65 2.565 ;
      RECT 83.94 0.885 84.11 2.595 ;
      RECT 83.88 0.885 84.17 1.115 ;
      RECT 83.88 7.765 84.17 7.995 ;
      RECT 83.94 6.285 84.11 7.995 ;
      RECT 83.88 6.285 84.17 6.515 ;
      RECT 83.88 6.325 84.73 6.485 ;
      RECT 84.56 5.915 84.73 6.485 ;
      RECT 83.88 6.32 84.27 6.485 ;
      RECT 84.5 5.915 84.79 6.145 ;
      RECT 84.5 5.945 84.96 6.115 ;
      RECT 83.51 2.735 83.8 2.965 ;
      RECT 83.51 2.765 83.97 2.935 ;
      RECT 83.57 1.655 83.735 2.965 ;
      RECT 82.085 1.625 82.375 1.855 ;
      RECT 82.085 1.655 83.735 1.825 ;
      RECT 82.145 0.885 82.315 1.855 ;
      RECT 82.085 0.885 82.375 1.115 ;
      RECT 82.085 7.765 82.375 7.995 ;
      RECT 82.145 7.025 82.315 7.995 ;
      RECT 82.145 7.12 83.735 7.29 ;
      RECT 83.565 5.915 83.735 7.29 ;
      RECT 82.085 7.025 82.375 7.255 ;
      RECT 83.51 5.915 83.8 6.145 ;
      RECT 83.51 5.945 83.97 6.115 ;
      RECT 82.515 1.965 82.865 2.315 ;
      RECT 82.345 2.025 82.865 2.195 ;
      RECT 82.54 6.655 82.865 6.98 ;
      RECT 82.515 6.655 82.865 6.885 ;
      RECT 82.345 6.685 82.865 6.855 ;
      RECT 81.74 2.365 82.06 2.685 ;
      RECT 81.71 2.365 82.06 2.595 ;
      RECT 81.425 2.395 82.06 2.565 ;
      RECT 81.74 6.28 82.06 6.605 ;
      RECT 81.71 6.285 82.06 6.515 ;
      RECT 81.54 6.315 82.06 6.485 ;
      RECT 80.695 3.495 81.02 3.82 ;
      RECT 80.775 2.735 80.945 3.82 ;
      RECT 80.715 2.735 81.005 2.965 ;
      RECT 80.715 2.765 81.175 2.935 ;
      RECT 80.695 5.855 81.02 6.18 ;
      RECT 80.695 5.945 81.175 6.115 ;
      RECT 77.485 3.79 77.805 4.05 ;
      RECT 78.52 3.805 78.81 4.035 ;
      RECT 77.485 3.85 78.81 3.99 ;
      RECT 77.145 5.83 77.465 6.09 ;
      RECT 78.52 5.845 78.81 6.075 ;
      RECT 78.595 5.55 78.735 6.075 ;
      RECT 77.235 5.55 77.375 6.09 ;
      RECT 77.235 5.55 78.735 5.69 ;
      RECT 78.165 2.77 78.485 3.03 ;
      RECT 77.89 2.83 78.485 2.97 ;
      RECT 75.105 6.51 75.425 6.77 ;
      RECT 74.1 6.525 74.39 6.755 ;
      RECT 74.1 6.57 76.015 6.71 ;
      RECT 75.875 6.23 76.015 6.71 ;
      RECT 75.875 6.23 77.885 6.37 ;
      RECT 77.745 5.845 77.885 6.37 ;
      RECT 77.67 5.845 77.96 6.075 ;
      RECT 77.485 4.81 77.805 5.07 ;
      RECT 75.34 4.825 75.63 5.055 ;
      RECT 75.34 4.87 77.805 5.01 ;
      RECT 76.805 3.79 77.125 4.05 ;
      RECT 74.44 3.805 74.73 4.035 ;
      RECT 74.44 3.85 77.125 3.99 ;
      RECT 76.465 6.51 76.785 6.77 ;
      RECT 76.465 6.57 77.06 6.71 ;
      RECT 76.465 3.11 76.785 3.37 ;
      RECT 76.19 3.17 76.785 3.31 ;
      RECT 75.785 2.77 76.105 3.03 ;
      RECT 75.51 2.83 76.105 2.97 ;
      RECT 75.445 3.45 75.765 3.71 ;
      RECT 72.57 3.465 72.86 3.695 ;
      RECT 72.57 3.51 75.765 3.65 ;
      RECT 75.025 2.79 75.165 3.65 ;
      RECT 74.95 2.79 75.24 3.02 ;
      RECT 75.105 2.26 75.425 2.52 ;
      RECT 75.105 2.275 75.61 2.505 ;
      RECT 75.015 2.32 75.61 2.46 ;
      RECT 74.425 5.83 74.745 6.09 ;
      RECT 72.06 5.845 72.35 6.075 ;
      RECT 72.06 5.89 74.745 6.03 ;
      RECT 74.44 2.79 74.73 3.02 ;
      RECT 73.835 2.835 74.73 2.975 ;
      RECT 73.835 2.43 73.975 2.975 ;
      RECT 73.745 2.43 74.065 2.69 ;
      RECT 73.065 2.77 73.385 3.03 ;
      RECT 72.79 2.83 73.385 2.97 ;
      RECT 73.065 4.81 73.385 5.07 ;
      RECT 72.79 4.87 73.385 5.01 ;
      RECT 71.31 5.89 71.65 6.17 ;
      RECT 69.03 5.915 69.32 6.145 ;
      RECT 69.03 5.945 71.65 6.115 ;
      RECT 70.83 6.575 71.12 6.885 ;
      RECT 70.66 6.685 71.15 6.855 ;
      RECT 70.81 6.575 71.15 6.855 ;
      RECT 70.4 7.765 70.69 7.995 ;
      RECT 70.46 6.995 70.63 7.995 ;
      RECT 70.365 6.995 70.735 7.37 ;
      RECT 67.65 7.765 67.94 7.995 ;
      RECT 67.71 6.285 67.88 7.995 ;
      RECT 67.71 6.655 68.035 6.98 ;
      RECT 67.65 6.285 67.94 6.515 ;
      RECT 67.65 2.365 67.94 2.595 ;
      RECT 67.71 0.885 67.88 2.595 ;
      RECT 67.65 0.885 67.94 1.115 ;
      RECT 67.24 2.735 67.57 2.965 ;
      RECT 67.24 2.765 67.74 2.935 ;
      RECT 67.24 2.395 67.43 2.965 ;
      RECT 66.66 2.365 66.95 2.595 ;
      RECT 66.66 2.395 67.43 2.565 ;
      RECT 66.72 0.885 66.89 2.595 ;
      RECT 66.66 0.885 66.95 1.115 ;
      RECT 66.66 7.765 66.95 7.995 ;
      RECT 66.72 6.285 66.89 7.995 ;
      RECT 66.66 6.285 66.95 6.515 ;
      RECT 66.66 6.325 67.51 6.485 ;
      RECT 67.34 5.915 67.51 6.485 ;
      RECT 66.66 6.32 67.05 6.485 ;
      RECT 67.28 5.915 67.57 6.145 ;
      RECT 67.28 5.945 67.74 6.115 ;
      RECT 66.29 2.735 66.58 2.965 ;
      RECT 66.29 2.765 66.75 2.935 ;
      RECT 66.35 1.655 66.515 2.965 ;
      RECT 64.865 1.625 65.155 1.855 ;
      RECT 64.865 1.655 66.515 1.825 ;
      RECT 64.925 0.885 65.095 1.855 ;
      RECT 64.865 0.885 65.155 1.115 ;
      RECT 64.865 7.765 65.155 7.995 ;
      RECT 64.925 7.025 65.095 7.995 ;
      RECT 64.925 7.12 66.515 7.29 ;
      RECT 66.345 5.915 66.515 7.29 ;
      RECT 64.865 7.025 65.155 7.255 ;
      RECT 66.29 5.915 66.58 6.145 ;
      RECT 66.29 5.945 66.75 6.115 ;
      RECT 65.295 1.965 65.645 2.315 ;
      RECT 65.125 2.025 65.645 2.195 ;
      RECT 65.32 6.655 65.645 6.98 ;
      RECT 65.295 6.655 65.645 6.885 ;
      RECT 65.125 6.685 65.645 6.855 ;
      RECT 64.52 2.365 64.84 2.685 ;
      RECT 64.49 2.365 64.84 2.595 ;
      RECT 64.205 2.395 64.84 2.565 ;
      RECT 64.52 6.28 64.84 6.605 ;
      RECT 64.49 6.285 64.84 6.515 ;
      RECT 64.32 6.315 64.84 6.485 ;
      RECT 63.475 3.495 63.8 3.82 ;
      RECT 63.555 2.735 63.725 3.82 ;
      RECT 63.495 2.735 63.785 2.965 ;
      RECT 63.495 2.765 63.955 2.935 ;
      RECT 63.475 5.855 63.8 6.18 ;
      RECT 63.475 5.945 63.955 6.115 ;
      RECT 60.265 3.79 60.585 4.05 ;
      RECT 61.3 3.805 61.59 4.035 ;
      RECT 60.265 3.85 61.59 3.99 ;
      RECT 59.925 5.83 60.245 6.09 ;
      RECT 61.3 5.845 61.59 6.075 ;
      RECT 61.375 5.55 61.515 6.075 ;
      RECT 60.015 5.55 60.155 6.09 ;
      RECT 60.015 5.55 61.515 5.69 ;
      RECT 60.945 2.77 61.265 3.03 ;
      RECT 60.67 2.83 61.265 2.97 ;
      RECT 57.885 6.51 58.205 6.77 ;
      RECT 56.88 6.525 57.17 6.755 ;
      RECT 56.88 6.57 58.795 6.71 ;
      RECT 58.655 6.23 58.795 6.71 ;
      RECT 58.655 6.23 60.665 6.37 ;
      RECT 60.525 5.845 60.665 6.37 ;
      RECT 60.45 5.845 60.74 6.075 ;
      RECT 60.265 4.81 60.585 5.07 ;
      RECT 58.12 4.825 58.41 5.055 ;
      RECT 58.12 4.87 60.585 5.01 ;
      RECT 59.585 3.79 59.905 4.05 ;
      RECT 57.22 3.805 57.51 4.035 ;
      RECT 57.22 3.85 59.905 3.99 ;
      RECT 59.245 6.51 59.565 6.77 ;
      RECT 59.245 6.57 59.84 6.71 ;
      RECT 59.245 3.11 59.565 3.37 ;
      RECT 58.97 3.17 59.565 3.31 ;
      RECT 58.565 2.77 58.885 3.03 ;
      RECT 58.29 2.83 58.885 2.97 ;
      RECT 58.225 3.45 58.545 3.71 ;
      RECT 55.35 3.465 55.64 3.695 ;
      RECT 55.35 3.51 58.545 3.65 ;
      RECT 57.805 2.79 57.945 3.65 ;
      RECT 57.73 2.79 58.02 3.02 ;
      RECT 57.885 2.26 58.205 2.52 ;
      RECT 57.885 2.275 58.39 2.505 ;
      RECT 57.795 2.32 58.39 2.46 ;
      RECT 57.205 5.83 57.525 6.09 ;
      RECT 54.84 5.845 55.13 6.075 ;
      RECT 54.84 5.89 57.525 6.03 ;
      RECT 57.22 2.79 57.51 3.02 ;
      RECT 56.615 2.835 57.51 2.975 ;
      RECT 56.615 2.43 56.755 2.975 ;
      RECT 56.525 2.43 56.845 2.69 ;
      RECT 55.845 2.77 56.165 3.03 ;
      RECT 55.57 2.83 56.165 2.97 ;
      RECT 55.845 4.81 56.165 5.07 ;
      RECT 55.57 4.87 56.165 5.01 ;
      RECT 54.09 5.89 54.43 6.17 ;
      RECT 51.81 5.915 52.1 6.145 ;
      RECT 51.81 5.945 54.43 6.115 ;
      RECT 53.61 6.575 53.9 6.885 ;
      RECT 53.44 6.685 53.93 6.855 ;
      RECT 53.59 6.575 53.93 6.855 ;
      RECT 53.18 7.765 53.47 7.995 ;
      RECT 53.24 6.995 53.41 7.995 ;
      RECT 53.145 6.995 53.515 7.37 ;
      RECT 50.43 7.765 50.72 7.995 ;
      RECT 50.49 6.285 50.66 7.995 ;
      RECT 50.49 6.655 50.815 6.98 ;
      RECT 50.43 6.285 50.72 6.515 ;
      RECT 50.43 2.365 50.72 2.595 ;
      RECT 50.49 0.885 50.66 2.595 ;
      RECT 50.43 0.885 50.72 1.115 ;
      RECT 50.02 2.735 50.35 2.965 ;
      RECT 50.02 2.765 50.52 2.935 ;
      RECT 50.02 2.395 50.21 2.965 ;
      RECT 49.44 2.365 49.73 2.595 ;
      RECT 49.44 2.395 50.21 2.565 ;
      RECT 49.5 0.885 49.67 2.595 ;
      RECT 49.44 0.885 49.73 1.115 ;
      RECT 49.44 7.765 49.73 7.995 ;
      RECT 49.5 6.285 49.67 7.995 ;
      RECT 49.44 6.285 49.73 6.515 ;
      RECT 49.44 6.325 50.29 6.485 ;
      RECT 50.12 5.915 50.29 6.485 ;
      RECT 49.44 6.32 49.83 6.485 ;
      RECT 50.06 5.915 50.35 6.145 ;
      RECT 50.06 5.945 50.52 6.115 ;
      RECT 49.07 2.735 49.36 2.965 ;
      RECT 49.07 2.765 49.53 2.935 ;
      RECT 49.13 1.655 49.295 2.965 ;
      RECT 47.645 1.625 47.935 1.855 ;
      RECT 47.645 1.655 49.295 1.825 ;
      RECT 47.705 0.885 47.875 1.855 ;
      RECT 47.645 0.885 47.935 1.115 ;
      RECT 47.645 7.765 47.935 7.995 ;
      RECT 47.705 7.025 47.875 7.995 ;
      RECT 47.705 7.12 49.295 7.29 ;
      RECT 49.125 5.915 49.295 7.29 ;
      RECT 47.645 7.025 47.935 7.255 ;
      RECT 49.07 5.915 49.36 6.145 ;
      RECT 49.07 5.945 49.53 6.115 ;
      RECT 48.075 1.965 48.425 2.315 ;
      RECT 47.905 2.025 48.425 2.195 ;
      RECT 48.1 6.655 48.425 6.98 ;
      RECT 48.075 6.655 48.425 6.885 ;
      RECT 47.905 6.685 48.425 6.855 ;
      RECT 47.3 2.365 47.62 2.685 ;
      RECT 47.27 2.365 47.62 2.595 ;
      RECT 46.985 2.395 47.62 2.565 ;
      RECT 47.3 6.28 47.62 6.605 ;
      RECT 47.27 6.285 47.62 6.515 ;
      RECT 47.1 6.315 47.62 6.485 ;
      RECT 46.255 3.495 46.58 3.82 ;
      RECT 46.335 2.735 46.505 3.82 ;
      RECT 46.275 2.735 46.565 2.965 ;
      RECT 46.275 2.765 46.735 2.935 ;
      RECT 46.255 5.855 46.58 6.18 ;
      RECT 46.255 5.945 46.735 6.115 ;
      RECT 43.045 3.79 43.365 4.05 ;
      RECT 44.08 3.805 44.37 4.035 ;
      RECT 43.045 3.85 44.37 3.99 ;
      RECT 42.705 5.83 43.025 6.09 ;
      RECT 44.08 5.845 44.37 6.075 ;
      RECT 44.155 5.55 44.295 6.075 ;
      RECT 42.795 5.55 42.935 6.09 ;
      RECT 42.795 5.55 44.295 5.69 ;
      RECT 43.725 2.77 44.045 3.03 ;
      RECT 43.45 2.83 44.045 2.97 ;
      RECT 40.665 6.51 40.985 6.77 ;
      RECT 39.66 6.525 39.95 6.755 ;
      RECT 39.66 6.57 41.575 6.71 ;
      RECT 41.435 6.23 41.575 6.71 ;
      RECT 41.435 6.23 43.445 6.37 ;
      RECT 43.305 5.845 43.445 6.37 ;
      RECT 43.23 5.845 43.52 6.075 ;
      RECT 43.045 4.81 43.365 5.07 ;
      RECT 40.9 4.825 41.19 5.055 ;
      RECT 40.9 4.87 43.365 5.01 ;
      RECT 42.365 3.79 42.685 4.05 ;
      RECT 40 3.805 40.29 4.035 ;
      RECT 40 3.85 42.685 3.99 ;
      RECT 42.025 6.51 42.345 6.77 ;
      RECT 42.025 6.57 42.62 6.71 ;
      RECT 42.025 3.11 42.345 3.37 ;
      RECT 41.75 3.17 42.345 3.31 ;
      RECT 41.345 2.77 41.665 3.03 ;
      RECT 41.07 2.83 41.665 2.97 ;
      RECT 41.005 3.45 41.325 3.71 ;
      RECT 38.13 3.465 38.42 3.695 ;
      RECT 38.13 3.51 41.325 3.65 ;
      RECT 40.585 2.79 40.725 3.65 ;
      RECT 40.51 2.79 40.8 3.02 ;
      RECT 40.665 2.26 40.985 2.52 ;
      RECT 40.665 2.275 41.17 2.505 ;
      RECT 40.575 2.32 41.17 2.46 ;
      RECT 39.985 5.83 40.305 6.09 ;
      RECT 37.62 5.845 37.91 6.075 ;
      RECT 37.62 5.89 40.305 6.03 ;
      RECT 40 2.79 40.29 3.02 ;
      RECT 39.395 2.835 40.29 2.975 ;
      RECT 39.395 2.43 39.535 2.975 ;
      RECT 39.305 2.43 39.625 2.69 ;
      RECT 38.625 2.77 38.945 3.03 ;
      RECT 38.35 2.83 38.945 2.97 ;
      RECT 38.625 4.81 38.945 5.07 ;
      RECT 38.35 4.87 38.945 5.01 ;
      RECT 36.87 5.89 37.21 6.17 ;
      RECT 34.59 5.915 34.88 6.145 ;
      RECT 34.59 5.945 37.21 6.115 ;
      RECT 36.39 6.575 36.68 6.885 ;
      RECT 36.22 6.685 36.71 6.855 ;
      RECT 36.37 6.575 36.71 6.855 ;
      RECT 35.96 7.765 36.25 7.995 ;
      RECT 36.02 6.995 36.19 7.995 ;
      RECT 35.925 6.995 36.295 7.37 ;
      RECT 33.21 7.765 33.5 7.995 ;
      RECT 33.27 6.285 33.44 7.995 ;
      RECT 33.27 6.655 33.595 6.98 ;
      RECT 33.21 6.285 33.5 6.515 ;
      RECT 33.21 2.365 33.5 2.595 ;
      RECT 33.27 0.885 33.44 2.595 ;
      RECT 33.21 0.885 33.5 1.115 ;
      RECT 32.8 2.735 33.13 2.965 ;
      RECT 32.8 2.765 33.3 2.935 ;
      RECT 32.8 2.395 32.99 2.965 ;
      RECT 32.22 2.365 32.51 2.595 ;
      RECT 32.22 2.395 32.99 2.565 ;
      RECT 32.28 0.885 32.45 2.595 ;
      RECT 32.22 0.885 32.51 1.115 ;
      RECT 32.22 7.765 32.51 7.995 ;
      RECT 32.28 6.285 32.45 7.995 ;
      RECT 32.22 6.285 32.51 6.515 ;
      RECT 32.22 6.325 33.07 6.485 ;
      RECT 32.9 5.915 33.07 6.485 ;
      RECT 32.22 6.32 32.61 6.485 ;
      RECT 32.84 5.915 33.13 6.145 ;
      RECT 32.84 5.945 33.3 6.115 ;
      RECT 31.85 2.735 32.14 2.965 ;
      RECT 31.85 2.765 32.31 2.935 ;
      RECT 31.91 1.655 32.075 2.965 ;
      RECT 30.425 1.625 30.715 1.855 ;
      RECT 30.425 1.655 32.075 1.825 ;
      RECT 30.485 0.885 30.655 1.855 ;
      RECT 30.425 0.885 30.715 1.115 ;
      RECT 30.425 7.765 30.715 7.995 ;
      RECT 30.485 7.025 30.655 7.995 ;
      RECT 30.485 7.12 32.075 7.29 ;
      RECT 31.905 5.915 32.075 7.29 ;
      RECT 30.425 7.025 30.715 7.255 ;
      RECT 31.85 5.915 32.14 6.145 ;
      RECT 31.85 5.945 32.31 6.115 ;
      RECT 30.855 1.965 31.205 2.315 ;
      RECT 30.685 2.025 31.205 2.195 ;
      RECT 30.88 6.655 31.205 6.98 ;
      RECT 30.855 6.655 31.205 6.885 ;
      RECT 30.685 6.685 31.205 6.855 ;
      RECT 30.08 2.365 30.4 2.685 ;
      RECT 30.05 2.365 30.4 2.595 ;
      RECT 29.765 2.395 30.4 2.565 ;
      RECT 30.08 6.28 30.4 6.605 ;
      RECT 30.05 6.285 30.4 6.515 ;
      RECT 29.88 6.315 30.4 6.485 ;
      RECT 29.035 3.495 29.36 3.82 ;
      RECT 29.115 2.735 29.285 3.82 ;
      RECT 29.055 2.735 29.345 2.965 ;
      RECT 29.055 2.765 29.515 2.935 ;
      RECT 29.035 5.855 29.36 6.18 ;
      RECT 29.035 5.945 29.515 6.115 ;
      RECT 25.825 3.79 26.145 4.05 ;
      RECT 26.86 3.805 27.15 4.035 ;
      RECT 25.825 3.85 27.15 3.99 ;
      RECT 25.485 5.83 25.805 6.09 ;
      RECT 26.86 5.845 27.15 6.075 ;
      RECT 26.935 5.55 27.075 6.075 ;
      RECT 25.575 5.55 25.715 6.09 ;
      RECT 25.575 5.55 27.075 5.69 ;
      RECT 26.505 2.77 26.825 3.03 ;
      RECT 26.23 2.83 26.825 2.97 ;
      RECT 23.445 6.51 23.765 6.77 ;
      RECT 22.44 6.525 22.73 6.755 ;
      RECT 22.44 6.57 24.355 6.71 ;
      RECT 24.215 6.23 24.355 6.71 ;
      RECT 24.215 6.23 26.225 6.37 ;
      RECT 26.085 5.845 26.225 6.37 ;
      RECT 26.01 5.845 26.3 6.075 ;
      RECT 25.825 4.81 26.145 5.07 ;
      RECT 23.68 4.825 23.97 5.055 ;
      RECT 23.68 4.87 26.145 5.01 ;
      RECT 25.145 3.79 25.465 4.05 ;
      RECT 22.78 3.805 23.07 4.035 ;
      RECT 22.78 3.85 25.465 3.99 ;
      RECT 24.805 6.51 25.125 6.77 ;
      RECT 24.805 6.57 25.4 6.71 ;
      RECT 24.805 3.11 25.125 3.37 ;
      RECT 24.53 3.17 25.125 3.31 ;
      RECT 24.125 2.77 24.445 3.03 ;
      RECT 23.85 2.83 24.445 2.97 ;
      RECT 23.785 3.45 24.105 3.71 ;
      RECT 20.91 3.465 21.2 3.695 ;
      RECT 20.91 3.51 24.105 3.65 ;
      RECT 23.365 2.79 23.505 3.65 ;
      RECT 23.29 2.79 23.58 3.02 ;
      RECT 23.445 2.26 23.765 2.52 ;
      RECT 23.445 2.275 23.95 2.505 ;
      RECT 23.355 2.32 23.95 2.46 ;
      RECT 22.765 5.83 23.085 6.09 ;
      RECT 20.4 5.845 20.69 6.075 ;
      RECT 20.4 5.89 23.085 6.03 ;
      RECT 22.78 2.79 23.07 3.02 ;
      RECT 22.175 2.835 23.07 2.975 ;
      RECT 22.175 2.43 22.315 2.975 ;
      RECT 22.085 2.43 22.405 2.69 ;
      RECT 21.405 2.77 21.725 3.03 ;
      RECT 21.13 2.83 21.725 2.97 ;
      RECT 21.405 4.81 21.725 5.07 ;
      RECT 21.13 4.87 21.725 5.01 ;
      RECT 19.65 5.89 19.99 6.17 ;
      RECT 17.37 5.915 17.66 6.145 ;
      RECT 17.37 5.945 19.99 6.115 ;
      RECT 19.17 6.575 19.46 6.885 ;
      RECT 19 6.685 19.49 6.855 ;
      RECT 19.15 6.575 19.49 6.855 ;
      RECT 18.74 7.765 19.03 7.995 ;
      RECT 18.8 6.995 18.97 7.995 ;
      RECT 18.705 6.995 19.075 7.37 ;
      RECT 15.99 7.765 16.28 7.995 ;
      RECT 16.05 6.285 16.22 7.995 ;
      RECT 16.05 6.655 16.375 6.98 ;
      RECT 15.99 6.285 16.28 6.515 ;
      RECT 15.99 2.365 16.28 2.595 ;
      RECT 16.05 0.885 16.22 2.595 ;
      RECT 15.99 0.885 16.28 1.115 ;
      RECT 15.58 2.735 15.91 2.965 ;
      RECT 15.58 2.765 16.08 2.935 ;
      RECT 15.58 2.395 15.77 2.965 ;
      RECT 15 2.365 15.29 2.595 ;
      RECT 15 2.395 15.77 2.565 ;
      RECT 15.06 0.885 15.23 2.595 ;
      RECT 15 0.885 15.29 1.115 ;
      RECT 15 7.765 15.29 7.995 ;
      RECT 15.06 6.285 15.23 7.995 ;
      RECT 15 6.285 15.29 6.515 ;
      RECT 15 6.325 15.85 6.485 ;
      RECT 15.68 5.915 15.85 6.485 ;
      RECT 15 6.32 15.39 6.485 ;
      RECT 15.62 5.915 15.91 6.145 ;
      RECT 15.62 5.945 16.08 6.115 ;
      RECT 14.63 2.735 14.92 2.965 ;
      RECT 14.63 2.765 15.09 2.935 ;
      RECT 14.69 1.655 14.855 2.965 ;
      RECT 13.205 1.625 13.495 1.855 ;
      RECT 13.205 1.655 14.855 1.825 ;
      RECT 13.265 0.885 13.435 1.855 ;
      RECT 13.205 0.885 13.495 1.115 ;
      RECT 13.205 7.765 13.495 7.995 ;
      RECT 13.265 7.025 13.435 7.995 ;
      RECT 13.265 7.12 14.855 7.29 ;
      RECT 14.685 5.915 14.855 7.29 ;
      RECT 13.205 7.025 13.495 7.255 ;
      RECT 14.63 5.915 14.92 6.145 ;
      RECT 14.63 5.945 15.09 6.115 ;
      RECT 13.635 1.965 13.985 2.315 ;
      RECT 13.465 2.025 13.985 2.195 ;
      RECT 13.66 6.655 13.985 6.98 ;
      RECT 13.635 6.655 13.985 6.885 ;
      RECT 13.465 6.685 13.985 6.855 ;
      RECT 12.86 2.365 13.18 2.685 ;
      RECT 12.83 2.365 13.18 2.595 ;
      RECT 12.545 2.395 13.18 2.565 ;
      RECT 12.86 6.28 13.18 6.605 ;
      RECT 12.83 6.285 13.18 6.515 ;
      RECT 12.66 6.315 13.18 6.485 ;
      RECT 11.815 3.495 12.14 3.82 ;
      RECT 11.895 2.735 12.065 3.82 ;
      RECT 11.835 2.735 12.125 2.965 ;
      RECT 11.835 2.765 12.295 2.935 ;
      RECT 11.815 5.855 12.14 6.18 ;
      RECT 11.815 5.945 12.295 6.115 ;
      RECT 8.605 3.79 8.925 4.05 ;
      RECT 9.64 3.805 9.93 4.035 ;
      RECT 8.605 3.85 9.93 3.99 ;
      RECT 8.265 5.83 8.585 6.09 ;
      RECT 9.64 5.845 9.93 6.075 ;
      RECT 9.715 5.55 9.855 6.075 ;
      RECT 8.355 5.55 8.495 6.09 ;
      RECT 8.355 5.55 9.855 5.69 ;
      RECT 9.285 2.77 9.605 3.03 ;
      RECT 9.01 2.83 9.605 2.97 ;
      RECT 6.225 6.51 6.545 6.77 ;
      RECT 5.22 6.525 5.51 6.755 ;
      RECT 5.22 6.57 7.135 6.71 ;
      RECT 6.995 6.23 7.135 6.71 ;
      RECT 6.995 6.23 9.005 6.37 ;
      RECT 8.865 5.845 9.005 6.37 ;
      RECT 8.79 5.845 9.08 6.075 ;
      RECT 8.605 4.81 8.925 5.07 ;
      RECT 6.46 4.825 6.75 5.055 ;
      RECT 6.46 4.87 8.925 5.01 ;
      RECT 7.925 3.79 8.245 4.05 ;
      RECT 5.56 3.805 5.85 4.035 ;
      RECT 5.56 3.85 8.245 3.99 ;
      RECT 7.585 6.51 7.905 6.77 ;
      RECT 7.585 6.57 8.18 6.71 ;
      RECT 7.585 3.11 7.905 3.37 ;
      RECT 7.31 3.17 7.905 3.31 ;
      RECT 6.905 2.77 7.225 3.03 ;
      RECT 6.63 2.83 7.225 2.97 ;
      RECT 6.565 3.45 6.885 3.71 ;
      RECT 3.69 3.465 3.98 3.695 ;
      RECT 3.69 3.51 6.885 3.65 ;
      RECT 6.145 2.79 6.285 3.65 ;
      RECT 6.07 2.79 6.36 3.02 ;
      RECT 6.225 2.26 6.545 2.52 ;
      RECT 6.225 2.275 6.73 2.505 ;
      RECT 6.135 2.32 6.73 2.46 ;
      RECT 5.545 5.83 5.865 6.09 ;
      RECT 3.18 5.845 3.47 6.075 ;
      RECT 3.18 5.89 5.865 6.03 ;
      RECT 5.56 2.79 5.85 3.02 ;
      RECT 4.955 2.835 5.85 2.975 ;
      RECT 4.955 2.43 5.095 2.975 ;
      RECT 4.865 2.43 5.185 2.69 ;
      RECT 4.185 2.77 4.505 3.03 ;
      RECT 3.91 2.83 4.505 2.97 ;
      RECT 4.185 4.81 4.505 5.07 ;
      RECT 3.91 4.87 4.505 5.01 ;
      RECT 2.43 5.89 2.77 6.17 ;
      RECT 0.15 5.915 0.44 6.145 ;
      RECT 0.15 5.945 2.77 6.115 ;
      RECT 1.95 6.575 2.24 6.885 ;
      RECT 1.78 6.685 2.27 6.855 ;
      RECT 1.93 6.575 2.27 6.855 ;
      RECT 1.52 7.765 1.81 7.995 ;
      RECT 1.58 6.995 1.75 7.995 ;
      RECT 1.485 6.995 1.855 7.37 ;
      RECT -1.46 6.655 -1.17 6.885 ;
      RECT -1.63 6.685 -1.17 6.855 ;
      RECT -1.89 7.765 -1.6 7.995 ;
      RECT -1.83 7.025 -1.66 7.995 ;
      RECT -1.92 7.025 -1.58 7.305 ;
      RECT -2.295 6.285 -1.955 6.565 ;
      RECT -2.435 6.315 -1.955 6.485 ;
      RECT -3.26 5.915 -2.97 6.145 ;
      RECT -3.26 5.945 -2.8 6.115 ;
      RECT 80.07 1.995 80.395 2.32 ;
      RECT 77.84 6.51 78.485 6.77 ;
      RECT 75.79 5.83 76.435 6.09 ;
      RECT 62.85 1.995 63.175 2.32 ;
      RECT 60.62 6.51 61.265 6.77 ;
      RECT 58.57 5.83 59.215 6.09 ;
      RECT 45.63 1.995 45.955 2.32 ;
      RECT 43.4 6.51 44.045 6.77 ;
      RECT 41.35 5.83 41.995 6.09 ;
      RECT 28.41 1.995 28.735 2.32 ;
      RECT 26.18 6.51 26.825 6.77 ;
      RECT 24.13 5.83 24.775 6.09 ;
      RECT 11.19 1.995 11.515 2.32 ;
      RECT 8.96 6.51 9.605 6.77 ;
      RECT 6.91 5.83 7.555 6.09 ;
    LAYER mcon ;
      RECT 84.93 0.915 85.1 1.085 ;
      RECT 84.93 2.395 85.1 2.565 ;
      RECT 84.93 6.315 85.1 6.485 ;
      RECT 84.93 7.795 85.1 7.965 ;
      RECT 84.58 0.105 84.75 0.275 ;
      RECT 84.58 4.165 84.75 4.335 ;
      RECT 84.58 4.545 84.75 4.715 ;
      RECT 84.58 8.605 84.75 8.775 ;
      RECT 84.56 2.765 84.73 2.935 ;
      RECT 84.56 5.945 84.73 6.115 ;
      RECT 83.94 0.915 84.11 1.085 ;
      RECT 83.94 2.395 84.11 2.565 ;
      RECT 83.94 6.315 84.11 6.485 ;
      RECT 83.94 7.795 84.11 7.965 ;
      RECT 83.59 0.105 83.76 0.275 ;
      RECT 83.59 4.165 83.76 4.335 ;
      RECT 83.59 4.545 83.76 4.715 ;
      RECT 83.59 8.605 83.76 8.775 ;
      RECT 83.57 2.765 83.74 2.935 ;
      RECT 83.57 5.945 83.74 6.115 ;
      RECT 82.885 0.105 83.055 0.275 ;
      RECT 82.885 4.165 83.055 4.335 ;
      RECT 82.885 4.545 83.055 4.715 ;
      RECT 82.885 8.605 83.055 8.775 ;
      RECT 82.575 2.025 82.745 2.195 ;
      RECT 82.575 6.685 82.745 6.855 ;
      RECT 82.205 0.105 82.375 0.275 ;
      RECT 82.205 8.605 82.375 8.775 ;
      RECT 82.145 0.915 82.315 1.085 ;
      RECT 82.145 1.655 82.315 1.825 ;
      RECT 82.145 7.055 82.315 7.225 ;
      RECT 82.145 7.795 82.315 7.965 ;
      RECT 81.77 2.395 81.94 2.565 ;
      RECT 81.77 6.315 81.94 6.485 ;
      RECT 81.525 0.105 81.695 0.275 ;
      RECT 81.525 8.605 81.695 8.775 ;
      RECT 80.845 0.105 81.015 0.275 ;
      RECT 80.845 8.605 81.015 8.775 ;
      RECT 80.775 2.765 80.945 2.935 ;
      RECT 80.775 5.945 80.945 6.115 ;
      RECT 79.08 1.625 79.25 1.795 ;
      RECT 79.08 4.345 79.25 4.515 ;
      RECT 79.08 7.065 79.25 7.235 ;
      RECT 78.62 1.625 78.79 1.795 ;
      RECT 78.62 4.345 78.79 4.515 ;
      RECT 78.62 7.065 78.79 7.235 ;
      RECT 78.58 3.835 78.75 4.005 ;
      RECT 78.58 5.875 78.75 6.045 ;
      RECT 78.24 2.815 78.41 2.985 ;
      RECT 78.16 1.625 78.33 1.795 ;
      RECT 78.16 4.345 78.33 4.515 ;
      RECT 78.16 7.065 78.33 7.235 ;
      RECT 77.9 6.555 78.07 6.725 ;
      RECT 77.73 5.875 77.9 6.045 ;
      RECT 77.7 1.625 77.87 1.795 ;
      RECT 77.7 4.345 77.87 4.515 ;
      RECT 77.7 7.065 77.87 7.235 ;
      RECT 77.24 1.625 77.41 1.795 ;
      RECT 77.24 4.345 77.41 4.515 ;
      RECT 77.24 7.065 77.41 7.235 ;
      RECT 77.22 5.875 77.39 6.045 ;
      RECT 76.78 1.625 76.95 1.795 ;
      RECT 76.78 4.345 76.95 4.515 ;
      RECT 76.78 7.065 76.95 7.235 ;
      RECT 76.54 3.155 76.71 3.325 ;
      RECT 76.54 6.555 76.71 6.725 ;
      RECT 76.32 1.625 76.49 1.795 ;
      RECT 76.32 4.345 76.49 4.515 ;
      RECT 76.32 7.065 76.49 7.235 ;
      RECT 75.86 1.625 76.03 1.795 ;
      RECT 75.86 2.815 76.03 2.985 ;
      RECT 75.86 4.345 76.03 4.515 ;
      RECT 75.86 7.065 76.03 7.235 ;
      RECT 75.85 5.875 76.02 6.045 ;
      RECT 75.4 1.625 75.57 1.795 ;
      RECT 75.4 4.345 75.57 4.515 ;
      RECT 75.4 4.855 75.57 5.025 ;
      RECT 75.4 7.065 75.57 7.235 ;
      RECT 75.38 2.305 75.55 2.475 ;
      RECT 75.01 2.82 75.18 2.99 ;
      RECT 74.94 1.625 75.11 1.795 ;
      RECT 74.94 4.345 75.11 4.515 ;
      RECT 74.94 7.065 75.11 7.235 ;
      RECT 74.5 2.82 74.67 2.99 ;
      RECT 74.5 3.835 74.67 4.005 ;
      RECT 74.5 5.875 74.67 6.045 ;
      RECT 74.48 1.625 74.65 1.795 ;
      RECT 74.48 4.345 74.65 4.515 ;
      RECT 74.48 7.065 74.65 7.235 ;
      RECT 74.16 6.555 74.33 6.725 ;
      RECT 74.02 1.625 74.19 1.795 ;
      RECT 74.02 4.345 74.19 4.515 ;
      RECT 74.02 7.065 74.19 7.235 ;
      RECT 73.56 1.625 73.73 1.795 ;
      RECT 73.56 4.345 73.73 4.515 ;
      RECT 73.56 7.065 73.73 7.235 ;
      RECT 73.14 2.815 73.31 2.985 ;
      RECT 73.14 4.855 73.31 5.025 ;
      RECT 73.1 1.625 73.27 1.795 ;
      RECT 73.1 4.345 73.27 4.515 ;
      RECT 73.1 7.065 73.27 7.235 ;
      RECT 72.64 1.625 72.81 1.795 ;
      RECT 72.64 4.345 72.81 4.515 ;
      RECT 72.64 7.065 72.81 7.235 ;
      RECT 72.63 3.495 72.8 3.665 ;
      RECT 72.18 1.625 72.35 1.795 ;
      RECT 72.18 4.345 72.35 4.515 ;
      RECT 72.18 7.065 72.35 7.235 ;
      RECT 72.12 5.875 72.29 6.045 ;
      RECT 71.2 4.545 71.37 4.715 ;
      RECT 71.2 8.605 71.37 8.775 ;
      RECT 70.89 6.685 71.06 6.855 ;
      RECT 70.52 8.605 70.69 8.775 ;
      RECT 70.46 7.055 70.63 7.225 ;
      RECT 70.46 7.795 70.63 7.965 ;
      RECT 70.085 6.315 70.255 6.485 ;
      RECT 69.84 8.605 70.01 8.775 ;
      RECT 69.16 8.605 69.33 8.775 ;
      RECT 69.09 5.945 69.26 6.115 ;
      RECT 67.71 0.915 67.88 1.085 ;
      RECT 67.71 2.395 67.88 2.565 ;
      RECT 67.71 6.315 67.88 6.485 ;
      RECT 67.71 7.795 67.88 7.965 ;
      RECT 67.36 0.105 67.53 0.275 ;
      RECT 67.36 4.165 67.53 4.335 ;
      RECT 67.36 4.545 67.53 4.715 ;
      RECT 67.36 8.605 67.53 8.775 ;
      RECT 67.34 2.765 67.51 2.935 ;
      RECT 67.34 5.945 67.51 6.115 ;
      RECT 66.72 0.915 66.89 1.085 ;
      RECT 66.72 2.395 66.89 2.565 ;
      RECT 66.72 6.315 66.89 6.485 ;
      RECT 66.72 7.795 66.89 7.965 ;
      RECT 66.37 0.105 66.54 0.275 ;
      RECT 66.37 4.165 66.54 4.335 ;
      RECT 66.37 4.545 66.54 4.715 ;
      RECT 66.37 8.605 66.54 8.775 ;
      RECT 66.35 2.765 66.52 2.935 ;
      RECT 66.35 5.945 66.52 6.115 ;
      RECT 65.665 0.105 65.835 0.275 ;
      RECT 65.665 4.165 65.835 4.335 ;
      RECT 65.665 4.545 65.835 4.715 ;
      RECT 65.665 8.605 65.835 8.775 ;
      RECT 65.355 2.025 65.525 2.195 ;
      RECT 65.355 6.685 65.525 6.855 ;
      RECT 64.985 0.105 65.155 0.275 ;
      RECT 64.985 8.605 65.155 8.775 ;
      RECT 64.925 0.915 65.095 1.085 ;
      RECT 64.925 1.655 65.095 1.825 ;
      RECT 64.925 7.055 65.095 7.225 ;
      RECT 64.925 7.795 65.095 7.965 ;
      RECT 64.55 2.395 64.72 2.565 ;
      RECT 64.55 6.315 64.72 6.485 ;
      RECT 64.305 0.105 64.475 0.275 ;
      RECT 64.305 8.605 64.475 8.775 ;
      RECT 63.625 0.105 63.795 0.275 ;
      RECT 63.625 8.605 63.795 8.775 ;
      RECT 63.555 2.765 63.725 2.935 ;
      RECT 63.555 5.945 63.725 6.115 ;
      RECT 61.86 1.625 62.03 1.795 ;
      RECT 61.86 4.345 62.03 4.515 ;
      RECT 61.86 7.065 62.03 7.235 ;
      RECT 61.4 1.625 61.57 1.795 ;
      RECT 61.4 4.345 61.57 4.515 ;
      RECT 61.4 7.065 61.57 7.235 ;
      RECT 61.36 3.835 61.53 4.005 ;
      RECT 61.36 5.875 61.53 6.045 ;
      RECT 61.02 2.815 61.19 2.985 ;
      RECT 60.94 1.625 61.11 1.795 ;
      RECT 60.94 4.345 61.11 4.515 ;
      RECT 60.94 7.065 61.11 7.235 ;
      RECT 60.68 6.555 60.85 6.725 ;
      RECT 60.51 5.875 60.68 6.045 ;
      RECT 60.48 1.625 60.65 1.795 ;
      RECT 60.48 4.345 60.65 4.515 ;
      RECT 60.48 7.065 60.65 7.235 ;
      RECT 60.02 1.625 60.19 1.795 ;
      RECT 60.02 4.345 60.19 4.515 ;
      RECT 60.02 7.065 60.19 7.235 ;
      RECT 60 5.875 60.17 6.045 ;
      RECT 59.56 1.625 59.73 1.795 ;
      RECT 59.56 4.345 59.73 4.515 ;
      RECT 59.56 7.065 59.73 7.235 ;
      RECT 59.32 3.155 59.49 3.325 ;
      RECT 59.32 6.555 59.49 6.725 ;
      RECT 59.1 1.625 59.27 1.795 ;
      RECT 59.1 4.345 59.27 4.515 ;
      RECT 59.1 7.065 59.27 7.235 ;
      RECT 58.64 1.625 58.81 1.795 ;
      RECT 58.64 2.815 58.81 2.985 ;
      RECT 58.64 4.345 58.81 4.515 ;
      RECT 58.64 7.065 58.81 7.235 ;
      RECT 58.63 5.875 58.8 6.045 ;
      RECT 58.18 1.625 58.35 1.795 ;
      RECT 58.18 4.345 58.35 4.515 ;
      RECT 58.18 4.855 58.35 5.025 ;
      RECT 58.18 7.065 58.35 7.235 ;
      RECT 58.16 2.305 58.33 2.475 ;
      RECT 57.79 2.82 57.96 2.99 ;
      RECT 57.72 1.625 57.89 1.795 ;
      RECT 57.72 4.345 57.89 4.515 ;
      RECT 57.72 7.065 57.89 7.235 ;
      RECT 57.28 2.82 57.45 2.99 ;
      RECT 57.28 3.835 57.45 4.005 ;
      RECT 57.28 5.875 57.45 6.045 ;
      RECT 57.26 1.625 57.43 1.795 ;
      RECT 57.26 4.345 57.43 4.515 ;
      RECT 57.26 7.065 57.43 7.235 ;
      RECT 56.94 6.555 57.11 6.725 ;
      RECT 56.8 1.625 56.97 1.795 ;
      RECT 56.8 4.345 56.97 4.515 ;
      RECT 56.8 7.065 56.97 7.235 ;
      RECT 56.34 1.625 56.51 1.795 ;
      RECT 56.34 4.345 56.51 4.515 ;
      RECT 56.34 7.065 56.51 7.235 ;
      RECT 55.92 2.815 56.09 2.985 ;
      RECT 55.92 4.855 56.09 5.025 ;
      RECT 55.88 1.625 56.05 1.795 ;
      RECT 55.88 4.345 56.05 4.515 ;
      RECT 55.88 7.065 56.05 7.235 ;
      RECT 55.42 1.625 55.59 1.795 ;
      RECT 55.42 4.345 55.59 4.515 ;
      RECT 55.42 7.065 55.59 7.235 ;
      RECT 55.41 3.495 55.58 3.665 ;
      RECT 54.96 1.625 55.13 1.795 ;
      RECT 54.96 4.345 55.13 4.515 ;
      RECT 54.96 7.065 55.13 7.235 ;
      RECT 54.9 5.875 55.07 6.045 ;
      RECT 53.98 4.545 54.15 4.715 ;
      RECT 53.98 8.605 54.15 8.775 ;
      RECT 53.67 6.685 53.84 6.855 ;
      RECT 53.3 8.605 53.47 8.775 ;
      RECT 53.24 7.055 53.41 7.225 ;
      RECT 53.24 7.795 53.41 7.965 ;
      RECT 52.865 6.315 53.035 6.485 ;
      RECT 52.62 8.605 52.79 8.775 ;
      RECT 51.94 8.605 52.11 8.775 ;
      RECT 51.87 5.945 52.04 6.115 ;
      RECT 50.49 0.915 50.66 1.085 ;
      RECT 50.49 2.395 50.66 2.565 ;
      RECT 50.49 6.315 50.66 6.485 ;
      RECT 50.49 7.795 50.66 7.965 ;
      RECT 50.14 0.105 50.31 0.275 ;
      RECT 50.14 4.165 50.31 4.335 ;
      RECT 50.14 4.545 50.31 4.715 ;
      RECT 50.14 8.605 50.31 8.775 ;
      RECT 50.12 2.765 50.29 2.935 ;
      RECT 50.12 5.945 50.29 6.115 ;
      RECT 49.5 0.915 49.67 1.085 ;
      RECT 49.5 2.395 49.67 2.565 ;
      RECT 49.5 6.315 49.67 6.485 ;
      RECT 49.5 7.795 49.67 7.965 ;
      RECT 49.15 0.105 49.32 0.275 ;
      RECT 49.15 4.165 49.32 4.335 ;
      RECT 49.15 4.545 49.32 4.715 ;
      RECT 49.15 8.605 49.32 8.775 ;
      RECT 49.13 2.765 49.3 2.935 ;
      RECT 49.13 5.945 49.3 6.115 ;
      RECT 48.445 0.105 48.615 0.275 ;
      RECT 48.445 4.165 48.615 4.335 ;
      RECT 48.445 4.545 48.615 4.715 ;
      RECT 48.445 8.605 48.615 8.775 ;
      RECT 48.135 2.025 48.305 2.195 ;
      RECT 48.135 6.685 48.305 6.855 ;
      RECT 47.765 0.105 47.935 0.275 ;
      RECT 47.765 8.605 47.935 8.775 ;
      RECT 47.705 0.915 47.875 1.085 ;
      RECT 47.705 1.655 47.875 1.825 ;
      RECT 47.705 7.055 47.875 7.225 ;
      RECT 47.705 7.795 47.875 7.965 ;
      RECT 47.33 2.395 47.5 2.565 ;
      RECT 47.33 6.315 47.5 6.485 ;
      RECT 47.085 0.105 47.255 0.275 ;
      RECT 47.085 8.605 47.255 8.775 ;
      RECT 46.405 0.105 46.575 0.275 ;
      RECT 46.405 8.605 46.575 8.775 ;
      RECT 46.335 2.765 46.505 2.935 ;
      RECT 46.335 5.945 46.505 6.115 ;
      RECT 44.64 1.625 44.81 1.795 ;
      RECT 44.64 4.345 44.81 4.515 ;
      RECT 44.64 7.065 44.81 7.235 ;
      RECT 44.18 1.625 44.35 1.795 ;
      RECT 44.18 4.345 44.35 4.515 ;
      RECT 44.18 7.065 44.35 7.235 ;
      RECT 44.14 3.835 44.31 4.005 ;
      RECT 44.14 5.875 44.31 6.045 ;
      RECT 43.8 2.815 43.97 2.985 ;
      RECT 43.72 1.625 43.89 1.795 ;
      RECT 43.72 4.345 43.89 4.515 ;
      RECT 43.72 7.065 43.89 7.235 ;
      RECT 43.46 6.555 43.63 6.725 ;
      RECT 43.29 5.875 43.46 6.045 ;
      RECT 43.26 1.625 43.43 1.795 ;
      RECT 43.26 4.345 43.43 4.515 ;
      RECT 43.26 7.065 43.43 7.235 ;
      RECT 42.8 1.625 42.97 1.795 ;
      RECT 42.8 4.345 42.97 4.515 ;
      RECT 42.8 7.065 42.97 7.235 ;
      RECT 42.78 5.875 42.95 6.045 ;
      RECT 42.34 1.625 42.51 1.795 ;
      RECT 42.34 4.345 42.51 4.515 ;
      RECT 42.34 7.065 42.51 7.235 ;
      RECT 42.1 3.155 42.27 3.325 ;
      RECT 42.1 6.555 42.27 6.725 ;
      RECT 41.88 1.625 42.05 1.795 ;
      RECT 41.88 4.345 42.05 4.515 ;
      RECT 41.88 7.065 42.05 7.235 ;
      RECT 41.42 1.625 41.59 1.795 ;
      RECT 41.42 2.815 41.59 2.985 ;
      RECT 41.42 4.345 41.59 4.515 ;
      RECT 41.42 7.065 41.59 7.235 ;
      RECT 41.41 5.875 41.58 6.045 ;
      RECT 40.96 1.625 41.13 1.795 ;
      RECT 40.96 4.345 41.13 4.515 ;
      RECT 40.96 4.855 41.13 5.025 ;
      RECT 40.96 7.065 41.13 7.235 ;
      RECT 40.94 2.305 41.11 2.475 ;
      RECT 40.57 2.82 40.74 2.99 ;
      RECT 40.5 1.625 40.67 1.795 ;
      RECT 40.5 4.345 40.67 4.515 ;
      RECT 40.5 7.065 40.67 7.235 ;
      RECT 40.06 2.82 40.23 2.99 ;
      RECT 40.06 3.835 40.23 4.005 ;
      RECT 40.06 5.875 40.23 6.045 ;
      RECT 40.04 1.625 40.21 1.795 ;
      RECT 40.04 4.345 40.21 4.515 ;
      RECT 40.04 7.065 40.21 7.235 ;
      RECT 39.72 6.555 39.89 6.725 ;
      RECT 39.58 1.625 39.75 1.795 ;
      RECT 39.58 4.345 39.75 4.515 ;
      RECT 39.58 7.065 39.75 7.235 ;
      RECT 39.12 1.625 39.29 1.795 ;
      RECT 39.12 4.345 39.29 4.515 ;
      RECT 39.12 7.065 39.29 7.235 ;
      RECT 38.7 2.815 38.87 2.985 ;
      RECT 38.7 4.855 38.87 5.025 ;
      RECT 38.66 1.625 38.83 1.795 ;
      RECT 38.66 4.345 38.83 4.515 ;
      RECT 38.66 7.065 38.83 7.235 ;
      RECT 38.2 1.625 38.37 1.795 ;
      RECT 38.2 4.345 38.37 4.515 ;
      RECT 38.2 7.065 38.37 7.235 ;
      RECT 38.19 3.495 38.36 3.665 ;
      RECT 37.74 1.625 37.91 1.795 ;
      RECT 37.74 4.345 37.91 4.515 ;
      RECT 37.74 7.065 37.91 7.235 ;
      RECT 37.68 5.875 37.85 6.045 ;
      RECT 36.76 4.545 36.93 4.715 ;
      RECT 36.76 8.605 36.93 8.775 ;
      RECT 36.45 6.685 36.62 6.855 ;
      RECT 36.08 8.605 36.25 8.775 ;
      RECT 36.02 7.055 36.19 7.225 ;
      RECT 36.02 7.795 36.19 7.965 ;
      RECT 35.645 6.315 35.815 6.485 ;
      RECT 35.4 8.605 35.57 8.775 ;
      RECT 34.72 8.605 34.89 8.775 ;
      RECT 34.65 5.945 34.82 6.115 ;
      RECT 33.27 0.915 33.44 1.085 ;
      RECT 33.27 2.395 33.44 2.565 ;
      RECT 33.27 6.315 33.44 6.485 ;
      RECT 33.27 7.795 33.44 7.965 ;
      RECT 32.92 0.105 33.09 0.275 ;
      RECT 32.92 4.165 33.09 4.335 ;
      RECT 32.92 4.545 33.09 4.715 ;
      RECT 32.92 8.605 33.09 8.775 ;
      RECT 32.9 2.765 33.07 2.935 ;
      RECT 32.9 5.945 33.07 6.115 ;
      RECT 32.28 0.915 32.45 1.085 ;
      RECT 32.28 2.395 32.45 2.565 ;
      RECT 32.28 6.315 32.45 6.485 ;
      RECT 32.28 7.795 32.45 7.965 ;
      RECT 31.93 0.105 32.1 0.275 ;
      RECT 31.93 4.165 32.1 4.335 ;
      RECT 31.93 4.545 32.1 4.715 ;
      RECT 31.93 8.605 32.1 8.775 ;
      RECT 31.91 2.765 32.08 2.935 ;
      RECT 31.91 5.945 32.08 6.115 ;
      RECT 31.225 0.105 31.395 0.275 ;
      RECT 31.225 4.165 31.395 4.335 ;
      RECT 31.225 4.545 31.395 4.715 ;
      RECT 31.225 8.605 31.395 8.775 ;
      RECT 30.915 2.025 31.085 2.195 ;
      RECT 30.915 6.685 31.085 6.855 ;
      RECT 30.545 0.105 30.715 0.275 ;
      RECT 30.545 8.605 30.715 8.775 ;
      RECT 30.485 0.915 30.655 1.085 ;
      RECT 30.485 1.655 30.655 1.825 ;
      RECT 30.485 7.055 30.655 7.225 ;
      RECT 30.485 7.795 30.655 7.965 ;
      RECT 30.11 2.395 30.28 2.565 ;
      RECT 30.11 6.315 30.28 6.485 ;
      RECT 29.865 0.105 30.035 0.275 ;
      RECT 29.865 8.605 30.035 8.775 ;
      RECT 29.185 0.105 29.355 0.275 ;
      RECT 29.185 8.605 29.355 8.775 ;
      RECT 29.115 2.765 29.285 2.935 ;
      RECT 29.115 5.945 29.285 6.115 ;
      RECT 27.42 1.625 27.59 1.795 ;
      RECT 27.42 4.345 27.59 4.515 ;
      RECT 27.42 7.065 27.59 7.235 ;
      RECT 26.96 1.625 27.13 1.795 ;
      RECT 26.96 4.345 27.13 4.515 ;
      RECT 26.96 7.065 27.13 7.235 ;
      RECT 26.92 3.835 27.09 4.005 ;
      RECT 26.92 5.875 27.09 6.045 ;
      RECT 26.58 2.815 26.75 2.985 ;
      RECT 26.5 1.625 26.67 1.795 ;
      RECT 26.5 4.345 26.67 4.515 ;
      RECT 26.5 7.065 26.67 7.235 ;
      RECT 26.24 6.555 26.41 6.725 ;
      RECT 26.07 5.875 26.24 6.045 ;
      RECT 26.04 1.625 26.21 1.795 ;
      RECT 26.04 4.345 26.21 4.515 ;
      RECT 26.04 7.065 26.21 7.235 ;
      RECT 25.58 1.625 25.75 1.795 ;
      RECT 25.58 4.345 25.75 4.515 ;
      RECT 25.58 7.065 25.75 7.235 ;
      RECT 25.56 5.875 25.73 6.045 ;
      RECT 25.12 1.625 25.29 1.795 ;
      RECT 25.12 4.345 25.29 4.515 ;
      RECT 25.12 7.065 25.29 7.235 ;
      RECT 24.88 3.155 25.05 3.325 ;
      RECT 24.88 6.555 25.05 6.725 ;
      RECT 24.66 1.625 24.83 1.795 ;
      RECT 24.66 4.345 24.83 4.515 ;
      RECT 24.66 7.065 24.83 7.235 ;
      RECT 24.2 1.625 24.37 1.795 ;
      RECT 24.2 2.815 24.37 2.985 ;
      RECT 24.2 4.345 24.37 4.515 ;
      RECT 24.2 7.065 24.37 7.235 ;
      RECT 24.19 5.875 24.36 6.045 ;
      RECT 23.74 1.625 23.91 1.795 ;
      RECT 23.74 4.345 23.91 4.515 ;
      RECT 23.74 4.855 23.91 5.025 ;
      RECT 23.74 7.065 23.91 7.235 ;
      RECT 23.72 2.305 23.89 2.475 ;
      RECT 23.35 2.82 23.52 2.99 ;
      RECT 23.28 1.625 23.45 1.795 ;
      RECT 23.28 4.345 23.45 4.515 ;
      RECT 23.28 7.065 23.45 7.235 ;
      RECT 22.84 2.82 23.01 2.99 ;
      RECT 22.84 3.835 23.01 4.005 ;
      RECT 22.84 5.875 23.01 6.045 ;
      RECT 22.82 1.625 22.99 1.795 ;
      RECT 22.82 4.345 22.99 4.515 ;
      RECT 22.82 7.065 22.99 7.235 ;
      RECT 22.5 6.555 22.67 6.725 ;
      RECT 22.36 1.625 22.53 1.795 ;
      RECT 22.36 4.345 22.53 4.515 ;
      RECT 22.36 7.065 22.53 7.235 ;
      RECT 21.9 1.625 22.07 1.795 ;
      RECT 21.9 4.345 22.07 4.515 ;
      RECT 21.9 7.065 22.07 7.235 ;
      RECT 21.48 2.815 21.65 2.985 ;
      RECT 21.48 4.855 21.65 5.025 ;
      RECT 21.44 1.625 21.61 1.795 ;
      RECT 21.44 4.345 21.61 4.515 ;
      RECT 21.44 7.065 21.61 7.235 ;
      RECT 20.98 1.625 21.15 1.795 ;
      RECT 20.98 4.345 21.15 4.515 ;
      RECT 20.98 7.065 21.15 7.235 ;
      RECT 20.97 3.495 21.14 3.665 ;
      RECT 20.52 1.625 20.69 1.795 ;
      RECT 20.52 4.345 20.69 4.515 ;
      RECT 20.52 7.065 20.69 7.235 ;
      RECT 20.46 5.875 20.63 6.045 ;
      RECT 19.54 4.545 19.71 4.715 ;
      RECT 19.54 8.605 19.71 8.775 ;
      RECT 19.23 6.685 19.4 6.855 ;
      RECT 18.86 8.605 19.03 8.775 ;
      RECT 18.8 7.055 18.97 7.225 ;
      RECT 18.8 7.795 18.97 7.965 ;
      RECT 18.425 6.315 18.595 6.485 ;
      RECT 18.18 8.605 18.35 8.775 ;
      RECT 17.5 8.605 17.67 8.775 ;
      RECT 17.43 5.945 17.6 6.115 ;
      RECT 16.05 0.915 16.22 1.085 ;
      RECT 16.05 2.395 16.22 2.565 ;
      RECT 16.05 6.315 16.22 6.485 ;
      RECT 16.05 7.795 16.22 7.965 ;
      RECT 15.7 0.105 15.87 0.275 ;
      RECT 15.7 4.165 15.87 4.335 ;
      RECT 15.7 4.545 15.87 4.715 ;
      RECT 15.7 8.605 15.87 8.775 ;
      RECT 15.68 2.765 15.85 2.935 ;
      RECT 15.68 5.945 15.85 6.115 ;
      RECT 15.06 0.915 15.23 1.085 ;
      RECT 15.06 2.395 15.23 2.565 ;
      RECT 15.06 6.315 15.23 6.485 ;
      RECT 15.06 7.795 15.23 7.965 ;
      RECT 14.71 0.105 14.88 0.275 ;
      RECT 14.71 4.165 14.88 4.335 ;
      RECT 14.71 4.545 14.88 4.715 ;
      RECT 14.71 8.605 14.88 8.775 ;
      RECT 14.69 2.765 14.86 2.935 ;
      RECT 14.69 5.945 14.86 6.115 ;
      RECT 14.005 0.105 14.175 0.275 ;
      RECT 14.005 4.165 14.175 4.335 ;
      RECT 14.005 4.545 14.175 4.715 ;
      RECT 14.005 8.605 14.175 8.775 ;
      RECT 13.695 2.025 13.865 2.195 ;
      RECT 13.695 6.685 13.865 6.855 ;
      RECT 13.325 0.105 13.495 0.275 ;
      RECT 13.325 8.605 13.495 8.775 ;
      RECT 13.265 0.915 13.435 1.085 ;
      RECT 13.265 1.655 13.435 1.825 ;
      RECT 13.265 7.055 13.435 7.225 ;
      RECT 13.265 7.795 13.435 7.965 ;
      RECT 12.89 2.395 13.06 2.565 ;
      RECT 12.89 6.315 13.06 6.485 ;
      RECT 12.645 0.105 12.815 0.275 ;
      RECT 12.645 8.605 12.815 8.775 ;
      RECT 11.965 0.105 12.135 0.275 ;
      RECT 11.965 8.605 12.135 8.775 ;
      RECT 11.895 2.765 12.065 2.935 ;
      RECT 11.895 5.945 12.065 6.115 ;
      RECT 10.2 1.625 10.37 1.795 ;
      RECT 10.2 4.345 10.37 4.515 ;
      RECT 10.2 7.065 10.37 7.235 ;
      RECT 9.74 1.625 9.91 1.795 ;
      RECT 9.74 4.345 9.91 4.515 ;
      RECT 9.74 7.065 9.91 7.235 ;
      RECT 9.7 3.835 9.87 4.005 ;
      RECT 9.7 5.875 9.87 6.045 ;
      RECT 9.36 2.815 9.53 2.985 ;
      RECT 9.28 1.625 9.45 1.795 ;
      RECT 9.28 4.345 9.45 4.515 ;
      RECT 9.28 7.065 9.45 7.235 ;
      RECT 9.02 6.555 9.19 6.725 ;
      RECT 8.85 5.875 9.02 6.045 ;
      RECT 8.82 1.625 8.99 1.795 ;
      RECT 8.82 4.345 8.99 4.515 ;
      RECT 8.82 7.065 8.99 7.235 ;
      RECT 8.36 1.625 8.53 1.795 ;
      RECT 8.36 4.345 8.53 4.515 ;
      RECT 8.36 7.065 8.53 7.235 ;
      RECT 8.34 5.875 8.51 6.045 ;
      RECT 7.9 1.625 8.07 1.795 ;
      RECT 7.9 4.345 8.07 4.515 ;
      RECT 7.9 7.065 8.07 7.235 ;
      RECT 7.66 3.155 7.83 3.325 ;
      RECT 7.66 6.555 7.83 6.725 ;
      RECT 7.44 1.625 7.61 1.795 ;
      RECT 7.44 4.345 7.61 4.515 ;
      RECT 7.44 7.065 7.61 7.235 ;
      RECT 6.98 1.625 7.15 1.795 ;
      RECT 6.98 2.815 7.15 2.985 ;
      RECT 6.98 4.345 7.15 4.515 ;
      RECT 6.98 7.065 7.15 7.235 ;
      RECT 6.97 5.875 7.14 6.045 ;
      RECT 6.52 1.625 6.69 1.795 ;
      RECT 6.52 4.345 6.69 4.515 ;
      RECT 6.52 4.855 6.69 5.025 ;
      RECT 6.52 7.065 6.69 7.235 ;
      RECT 6.5 2.305 6.67 2.475 ;
      RECT 6.13 2.82 6.3 2.99 ;
      RECT 6.06 1.625 6.23 1.795 ;
      RECT 6.06 4.345 6.23 4.515 ;
      RECT 6.06 7.065 6.23 7.235 ;
      RECT 5.62 2.82 5.79 2.99 ;
      RECT 5.62 3.835 5.79 4.005 ;
      RECT 5.62 5.875 5.79 6.045 ;
      RECT 5.6 1.625 5.77 1.795 ;
      RECT 5.6 4.345 5.77 4.515 ;
      RECT 5.6 7.065 5.77 7.235 ;
      RECT 5.28 6.555 5.45 6.725 ;
      RECT 5.14 1.625 5.31 1.795 ;
      RECT 5.14 4.345 5.31 4.515 ;
      RECT 5.14 7.065 5.31 7.235 ;
      RECT 4.68 1.625 4.85 1.795 ;
      RECT 4.68 4.345 4.85 4.515 ;
      RECT 4.68 7.065 4.85 7.235 ;
      RECT 4.26 2.815 4.43 2.985 ;
      RECT 4.26 4.855 4.43 5.025 ;
      RECT 4.22 1.625 4.39 1.795 ;
      RECT 4.22 4.345 4.39 4.515 ;
      RECT 4.22 7.065 4.39 7.235 ;
      RECT 3.76 1.625 3.93 1.795 ;
      RECT 3.76 4.345 3.93 4.515 ;
      RECT 3.76 7.065 3.93 7.235 ;
      RECT 3.75 3.495 3.92 3.665 ;
      RECT 3.3 1.625 3.47 1.795 ;
      RECT 3.3 4.345 3.47 4.515 ;
      RECT 3.3 7.065 3.47 7.235 ;
      RECT 3.24 5.875 3.41 6.045 ;
      RECT 2.32 4.545 2.49 4.715 ;
      RECT 2.32 8.605 2.49 8.775 ;
      RECT 2.01 6.685 2.18 6.855 ;
      RECT 1.64 8.605 1.81 8.775 ;
      RECT 1.58 7.055 1.75 7.225 ;
      RECT 1.58 7.795 1.75 7.965 ;
      RECT 1.205 6.315 1.375 6.485 ;
      RECT 0.96 8.605 1.13 8.775 ;
      RECT 0.28 8.605 0.45 8.775 ;
      RECT 0.21 5.945 0.38 6.115 ;
      RECT -1.09 4.545 -0.92 4.715 ;
      RECT -1.09 8.605 -0.92 8.775 ;
      RECT -1.4 6.685 -1.23 6.855 ;
      RECT -1.77 8.605 -1.6 8.775 ;
      RECT -1.83 7.055 -1.66 7.225 ;
      RECT -1.83 7.795 -1.66 7.965 ;
      RECT -2.205 6.315 -2.035 6.485 ;
      RECT -2.45 8.605 -2.28 8.775 ;
      RECT -3.13 8.605 -2.96 8.775 ;
      RECT -3.2 5.945 -3.03 6.115 ;
    LAYER li ;
      RECT 76.26 0 76.55 2.63 ;
      RECT 59.04 0 59.33 2.63 ;
      RECT 41.82 0 42.11 2.63 ;
      RECT 24.6 0 24.89 2.63 ;
      RECT 7.38 0 7.67 2.63 ;
      RECT 73.06 0 73.29 2.615 ;
      RECT 72.18 0 72.39 2.615 ;
      RECT 55.84 0 56.07 2.615 ;
      RECT 54.96 0 55.17 2.615 ;
      RECT 38.62 0 38.85 2.615 ;
      RECT 37.74 0 37.95 2.615 ;
      RECT 21.4 0 21.63 2.615 ;
      RECT 20.52 0 20.73 2.615 ;
      RECT 4.18 0 4.41 2.615 ;
      RECT 3.3 0 3.51 2.615 ;
      RECT 75.81 0 76.08 2.605 ;
      RECT 74.9 0 75.14 2.605 ;
      RECT 74.45 0 74.69 2.605 ;
      RECT 73.51 0 73.78 2.605 ;
      RECT 58.59 0 58.86 2.605 ;
      RECT 57.68 0 57.92 2.605 ;
      RECT 57.23 0 57.47 2.605 ;
      RECT 56.29 0 56.56 2.605 ;
      RECT 41.37 0 41.64 2.605 ;
      RECT 40.46 0 40.7 2.605 ;
      RECT 40.01 0 40.25 2.605 ;
      RECT 39.07 0 39.34 2.605 ;
      RECT 24.15 0 24.42 2.605 ;
      RECT 23.24 0 23.48 2.605 ;
      RECT 22.79 0 23.03 2.605 ;
      RECT 21.85 0 22.12 2.605 ;
      RECT 6.93 0 7.2 2.605 ;
      RECT 6.02 0 6.26 2.605 ;
      RECT 5.57 0 5.81 2.605 ;
      RECT 4.63 0 4.9 2.605 ;
      RECT 78.93 0 79.26 2.185 ;
      RECT 78.09 0 78.42 2.185 ;
      RECT 61.71 0 62.04 2.185 ;
      RECT 60.87 0 61.2 2.185 ;
      RECT 44.49 0 44.82 2.185 ;
      RECT 43.65 0 43.98 2.185 ;
      RECT 27.27 0 27.6 2.185 ;
      RECT 26.43 0 26.76 2.185 ;
      RECT 10.05 0 10.38 2.185 ;
      RECT 9.21 0 9.54 2.185 ;
      RECT 72.035 0 79.69 1.795 ;
      RECT 54.815 0 62.47 1.795 ;
      RECT 37.595 0 45.25 1.795 ;
      RECT 20.375 0 28.03 1.795 ;
      RECT 3.155 0 10.81 1.795 ;
      RECT 72.03 0 79.69 1.635 ;
      RECT 54.81 0 62.47 1.635 ;
      RECT 37.59 0 45.25 1.635 ;
      RECT 20.37 0 28.03 1.635 ;
      RECT 3.15 0 10.81 1.635 ;
      RECT 84.5 0 84.67 0.935 ;
      RECT 83.51 0 83.68 0.935 ;
      RECT 80.765 0 80.935 0.935 ;
      RECT 67.28 0 67.45 0.935 ;
      RECT 66.29 0 66.46 0.935 ;
      RECT 63.545 0 63.715 0.935 ;
      RECT 50.06 0 50.23 0.935 ;
      RECT 49.07 0 49.24 0.935 ;
      RECT 46.325 0 46.495 0.935 ;
      RECT 32.84 0 33.01 0.935 ;
      RECT 31.85 0 32.02 0.935 ;
      RECT 29.105 0 29.275 0.935 ;
      RECT 15.62 0 15.79 0.935 ;
      RECT 14.63 0 14.8 0.935 ;
      RECT 11.885 0 12.055 0.935 ;
      RECT -3.385 0 85.47 0.305 ;
      RECT -1.4 4.13 -1.23 8.305 ;
      RECT 78.57 4.345 78.85 5.655 ;
      RECT 77.64 4.345 77.9 5.655 ;
      RECT 77.19 4.345 77.47 5.655 ;
      RECT 76.26 4.345 76.52 5.655 ;
      RECT 75.83 4.345 76.09 5.655 ;
      RECT 74.88 4.345 75.16 5.655 ;
      RECT 73.53 3.205 73.79 5.655 ;
      RECT 72.58 4.345 72.86 5.655 ;
      RECT 61.35 4.345 61.63 5.655 ;
      RECT 60.42 4.345 60.68 5.655 ;
      RECT 59.97 4.345 60.25 5.655 ;
      RECT 59.04 4.345 59.3 5.655 ;
      RECT 58.61 4.345 58.87 5.655 ;
      RECT 57.66 4.345 57.94 5.655 ;
      RECT 56.31 3.205 56.57 5.655 ;
      RECT 55.36 4.345 55.64 5.655 ;
      RECT 44.13 4.345 44.41 5.655 ;
      RECT 43.2 4.345 43.46 5.655 ;
      RECT 42.75 4.345 43.03 5.655 ;
      RECT 41.82 4.345 42.08 5.655 ;
      RECT 41.39 4.345 41.65 5.655 ;
      RECT 40.44 4.345 40.72 5.655 ;
      RECT 39.09 3.205 39.35 5.655 ;
      RECT 38.14 4.345 38.42 5.655 ;
      RECT 26.91 4.345 27.19 5.655 ;
      RECT 25.98 4.345 26.24 5.655 ;
      RECT 25.53 4.345 25.81 5.655 ;
      RECT 24.6 4.345 24.86 5.655 ;
      RECT 24.17 4.345 24.43 5.655 ;
      RECT 23.22 4.345 23.5 5.655 ;
      RECT 21.87 3.205 22.13 5.655 ;
      RECT 20.92 4.345 21.2 5.655 ;
      RECT 9.69 4.345 9.97 5.655 ;
      RECT 8.76 4.345 9.02 5.655 ;
      RECT 8.31 4.345 8.59 5.655 ;
      RECT 7.38 4.345 7.64 5.655 ;
      RECT 6.95 4.345 7.21 5.655 ;
      RECT 6 4.345 6.28 5.655 ;
      RECT 4.65 3.205 4.91 5.655 ;
      RECT 3.7 4.345 3.98 5.655 ;
      RECT 84.5 3.405 84.67 5.475 ;
      RECT 83.51 3.405 83.68 5.475 ;
      RECT 80.765 3.405 80.935 5.475 ;
      RECT 69.08 4.13 69.25 5.475 ;
      RECT 67.28 3.405 67.45 5.475 ;
      RECT 66.29 3.405 66.46 5.475 ;
      RECT 63.545 3.405 63.715 5.475 ;
      RECT 51.86 4.13 52.03 5.475 ;
      RECT 50.06 3.405 50.23 5.475 ;
      RECT 49.07 3.405 49.24 5.475 ;
      RECT 46.325 3.405 46.495 5.475 ;
      RECT 34.64 4.13 34.81 5.475 ;
      RECT 32.84 3.405 33.01 5.475 ;
      RECT 31.85 3.405 32.02 5.475 ;
      RECT 29.105 3.405 29.275 5.475 ;
      RECT 17.42 4.13 17.59 5.475 ;
      RECT 15.62 3.405 15.79 5.475 ;
      RECT 14.63 3.405 14.8 5.475 ;
      RECT 11.885 3.405 12.055 5.475 ;
      RECT 0.2 4.13 0.37 5.475 ;
      RECT -3.21 4.13 -3.04 5.475 ;
      RECT 79.485 4.135 85.47 4.745 ;
      RECT 68.905 4.13 71.655 4.745 ;
      RECT 62.265 4.135 68.25 4.745 ;
      RECT 51.685 4.13 54.435 4.745 ;
      RECT 45.045 4.135 51.03 4.745 ;
      RECT 34.465 4.13 37.215 4.745 ;
      RECT 27.825 4.135 33.81 4.745 ;
      RECT 17.245 4.13 19.995 4.745 ;
      RECT 10.605 4.135 16.59 4.745 ;
      RECT 0.025 4.13 2.775 4.745 ;
      RECT -3.385 4.13 -0.635 4.745 ;
      RECT 62.265 4.345 72.41 4.74 ;
      RECT 45.045 4.345 55.19 4.74 ;
      RECT 27.825 4.345 37.97 4.74 ;
      RECT 10.605 4.345 20.75 4.74 ;
      RECT -3.385 4.345 3.53 4.74 ;
      RECT -3.385 4.345 85.47 4.515 ;
      RECT 79.48 4.135 85.47 4.515 ;
      RECT 78.17 3.495 78.34 4.515 ;
      RECT 77.33 3.835 77.5 4.515 ;
      RECT 75.75 3.205 76.08 4.515 ;
      RECT 73.51 3.205 73.84 4.515 ;
      RECT 73.06 3.205 73.29 4.515 ;
      RECT 62.26 4.135 72.39 4.515 ;
      RECT 72.18 3.205 72.39 4.74 ;
      RECT 60.95 3.495 61.12 4.515 ;
      RECT 60.11 3.835 60.28 4.515 ;
      RECT 58.53 3.205 58.86 4.515 ;
      RECT 56.29 3.205 56.62 4.515 ;
      RECT 55.84 3.205 56.07 4.515 ;
      RECT 45.04 4.135 55.17 4.515 ;
      RECT 54.96 3.205 55.17 4.74 ;
      RECT 43.73 3.495 43.9 4.515 ;
      RECT 42.89 3.835 43.06 4.515 ;
      RECT 41.31 3.205 41.64 4.515 ;
      RECT 39.07 3.205 39.4 4.515 ;
      RECT 38.62 3.205 38.85 4.515 ;
      RECT 27.82 4.135 37.95 4.515 ;
      RECT 37.74 3.205 37.95 4.74 ;
      RECT 26.51 3.495 26.68 4.515 ;
      RECT 25.67 3.835 25.84 4.515 ;
      RECT 24.09 3.205 24.42 4.515 ;
      RECT 21.85 3.205 22.18 4.515 ;
      RECT 21.4 3.205 21.63 4.515 ;
      RECT 10.6 4.135 20.73 4.515 ;
      RECT 20.52 3.205 20.73 4.74 ;
      RECT 9.29 3.495 9.46 4.515 ;
      RECT 8.45 3.835 8.62 4.515 ;
      RECT 6.87 3.205 7.2 4.515 ;
      RECT 4.63 3.205 4.96 4.515 ;
      RECT 4.18 3.205 4.41 4.515 ;
      RECT -3.385 4.13 3.51 4.74 ;
      RECT 3.3 3.205 3.51 4.74 ;
      RECT 68.245 4.13 72.39 4.74 ;
      RECT 51.025 4.13 55.17 4.74 ;
      RECT 33.805 4.13 37.95 4.74 ;
      RECT 16.585 4.13 20.73 4.74 ;
      RECT -3.385 8.575 85.47 8.88 ;
      RECT 84.5 7.945 84.67 8.88 ;
      RECT 83.51 7.945 83.68 8.88 ;
      RECT 80.765 7.945 80.935 8.88 ;
      RECT 72.305 7.18 79.505 8.88 ;
      RECT 69.08 7.945 69.25 8.88 ;
      RECT 67.28 7.945 67.45 8.88 ;
      RECT 66.29 7.945 66.46 8.88 ;
      RECT 63.545 7.945 63.715 8.88 ;
      RECT 55.085 7.18 62.285 8.88 ;
      RECT 51.86 7.945 52.03 8.88 ;
      RECT 50.06 7.945 50.23 8.88 ;
      RECT 49.07 7.945 49.24 8.88 ;
      RECT 46.325 7.945 46.495 8.88 ;
      RECT 37.865 7.18 45.065 8.88 ;
      RECT 34.64 7.945 34.81 8.88 ;
      RECT 32.84 7.945 33.01 8.88 ;
      RECT 31.85 7.945 32.02 8.88 ;
      RECT 29.105 7.945 29.275 8.88 ;
      RECT 20.645 7.18 27.845 8.88 ;
      RECT 17.42 7.945 17.59 8.88 ;
      RECT 15.62 7.945 15.79 8.88 ;
      RECT 14.63 7.945 14.8 8.88 ;
      RECT 11.885 7.945 12.055 8.88 ;
      RECT 3.425 7.18 10.625 8.88 ;
      RECT 0.2 7.945 0.37 8.88 ;
      RECT -3.21 7.945 -3.04 8.88 ;
      RECT 72.035 7.065 79.395 7.235 ;
      RECT 54.815 7.065 62.175 7.235 ;
      RECT 37.595 7.065 44.955 7.235 ;
      RECT 20.375 7.065 27.735 7.235 ;
      RECT 3.155 7.065 10.515 7.235 ;
      RECT 78.54 6.265 78.85 8.88 ;
      RECT 77.16 6.265 77.47 8.88 ;
      RECT 74.88 6.265 75.19 8.88 ;
      RECT 74.51 5.875 74.68 8.88 ;
      RECT 72.58 6.265 72.89 8.88 ;
      RECT 61.32 6.265 61.63 8.88 ;
      RECT 59.94 6.265 60.25 8.88 ;
      RECT 57.66 6.265 57.97 8.88 ;
      RECT 57.29 5.875 57.46 8.88 ;
      RECT 55.36 6.265 55.67 8.88 ;
      RECT 44.1 6.265 44.41 8.88 ;
      RECT 42.72 6.265 43.03 8.88 ;
      RECT 40.44 6.265 40.75 8.88 ;
      RECT 40.07 5.875 40.24 8.88 ;
      RECT 38.14 6.265 38.45 8.88 ;
      RECT 26.88 6.265 27.19 8.88 ;
      RECT 25.5 6.265 25.81 8.88 ;
      RECT 23.22 6.265 23.53 8.88 ;
      RECT 22.85 5.875 23.02 8.88 ;
      RECT 20.92 6.265 21.23 8.88 ;
      RECT 9.66 6.265 9.97 8.88 ;
      RECT 8.28 6.265 8.59 8.88 ;
      RECT 6 6.265 6.31 8.88 ;
      RECT 5.63 5.875 5.8 8.88 ;
      RECT 3.7 6.265 4.01 8.88 ;
      RECT 74.89 5.825 75.225 6.095 ;
      RECT 57.67 5.825 58.005 6.095 ;
      RECT 40.45 5.825 40.785 6.095 ;
      RECT 23.23 5.825 23.565 6.095 ;
      RECT 6.01 5.825 6.345 6.095 ;
      RECT 74.5 5.875 75.225 6.045 ;
      RECT 57.28 5.875 58.005 6.045 ;
      RECT 40.06 5.875 40.785 6.045 ;
      RECT 22.84 5.875 23.565 6.045 ;
      RECT 5.62 5.875 6.345 6.045 ;
      RECT 84.56 1.74 84.73 2.935 ;
      RECT 84.56 1.74 85.025 1.91 ;
      RECT 84.56 6.97 85.025 7.14 ;
      RECT 84.56 5.945 84.73 7.14 ;
      RECT 83.57 1.74 83.74 2.935 ;
      RECT 83.57 1.74 84.035 1.91 ;
      RECT 83.57 6.97 84.035 7.14 ;
      RECT 83.57 5.945 83.74 7.14 ;
      RECT 81.715 2.635 81.885 3.865 ;
      RECT 81.77 0.855 81.94 2.805 ;
      RECT 81.715 0.575 81.885 1.025 ;
      RECT 81.715 7.855 81.885 8.305 ;
      RECT 81.77 6.075 81.94 8.025 ;
      RECT 81.715 5.015 81.885 6.245 ;
      RECT 81.195 0.575 81.365 3.865 ;
      RECT 81.195 2.075 81.6 2.405 ;
      RECT 81.195 1.235 81.6 1.565 ;
      RECT 81.195 5.015 81.365 8.305 ;
      RECT 81.195 7.315 81.6 7.645 ;
      RECT 81.195 6.475 81.6 6.805 ;
      RECT 80.775 5.94 80.945 7.22 ;
      RECT 80.765 5.94 80.945 6.18 ;
      RECT 78.93 3.495 79.31 4.175 ;
      RECT 79.14 2.365 79.31 4.175 ;
      RECT 77.06 2.365 77.29 3.035 ;
      RECT 77.06 2.365 79.31 2.535 ;
      RECT 78.59 2.045 78.76 2.535 ;
      RECT 78.58 3.155 78.75 4.005 ;
      RECT 77.665 3.155 78.97 3.325 ;
      RECT 78.725 2.705 78.97 3.325 ;
      RECT 77.665 2.785 77.835 3.325 ;
      RECT 77.46 2.785 77.835 2.955 ;
      RECT 77.64 6.265 78.335 6.895 ;
      RECT 78.165 4.685 78.335 6.895 ;
      RECT 78.07 4.685 78.4 5.665 ;
      RECT 77.67 3.495 78 4.175 ;
      RECT 76.76 3.495 77.16 4.175 ;
      RECT 76.76 3.495 78 3.665 ;
      RECT 76.26 3.075 76.58 4.175 ;
      RECT 76.26 3.075 76.71 3.325 ;
      RECT 76.26 3.075 76.89 3.245 ;
      RECT 76.72 2.025 76.89 3.245 ;
      RECT 76.72 2.025 77.675 2.195 ;
      RECT 76.26 6.265 76.955 6.895 ;
      RECT 76.785 4.685 76.955 6.895 ;
      RECT 76.69 4.685 77.02 5.665 ;
      RECT 76.28 5.825 76.615 6.075 ;
      RECT 75.735 5.825 76.07 6.075 ;
      RECT 75.735 5.875 76.615 6.045 ;
      RECT 75.395 6.265 76.09 6.895 ;
      RECT 75.395 4.685 75.565 6.895 ;
      RECT 75.33 4.685 75.66 5.665 ;
      RECT 74.89 3.205 75.22 4.16 ;
      RECT 74.89 3.205 75.57 3.375 ;
      RECT 75.4 1.965 75.57 3.375 ;
      RECT 75.31 1.965 75.64 2.605 ;
      RECT 74.37 3.205 74.7 4.16 ;
      RECT 74.02 3.205 74.7 3.375 ;
      RECT 74.02 1.965 74.19 3.375 ;
      RECT 73.95 1.965 74.28 2.605 ;
      RECT 74.16 5.875 74.33 6.725 ;
      RECT 73.435 5.825 73.77 6.075 ;
      RECT 73.435 5.875 74.33 6.045 ;
      RECT 73.5 2.785 73.85 3.035 ;
      RECT 72.98 2.785 73.31 3.035 ;
      RECT 72.98 2.815 73.85 2.985 ;
      RECT 73.095 6.265 73.79 6.895 ;
      RECT 73.095 4.685 73.265 6.895 ;
      RECT 73.03 4.685 73.36 5.665 ;
      RECT 72.59 5.825 72.925 6.095 ;
      RECT 72.12 5.875 72.925 6.045 ;
      RECT 72.56 3.195 72.89 4.175 ;
      RECT 72.56 1.965 72.81 4.175 ;
      RECT 72.56 1.965 72.89 2.595 ;
      RECT 70.03 7.855 70.2 8.305 ;
      RECT 70.085 6.075 70.255 8.025 ;
      RECT 70.03 5.015 70.2 6.245 ;
      RECT 69.51 5.015 69.68 8.305 ;
      RECT 69.51 7.315 69.915 7.645 ;
      RECT 69.51 6.475 69.915 6.805 ;
      RECT 67.34 1.74 67.51 2.935 ;
      RECT 67.34 1.74 67.805 1.91 ;
      RECT 67.34 6.97 67.805 7.14 ;
      RECT 67.34 5.945 67.51 7.14 ;
      RECT 66.35 1.74 66.52 2.935 ;
      RECT 66.35 1.74 66.815 1.91 ;
      RECT 66.35 6.97 66.815 7.14 ;
      RECT 66.35 5.945 66.52 7.14 ;
      RECT 64.495 2.635 64.665 3.865 ;
      RECT 64.55 0.855 64.72 2.805 ;
      RECT 64.495 0.575 64.665 1.025 ;
      RECT 64.495 7.855 64.665 8.305 ;
      RECT 64.55 6.075 64.72 8.025 ;
      RECT 64.495 5.015 64.665 6.245 ;
      RECT 63.975 0.575 64.145 3.865 ;
      RECT 63.975 2.075 64.38 2.405 ;
      RECT 63.975 1.235 64.38 1.565 ;
      RECT 63.975 5.015 64.145 8.305 ;
      RECT 63.975 7.315 64.38 7.645 ;
      RECT 63.975 6.475 64.38 6.805 ;
      RECT 63.555 5.94 63.725 7.22 ;
      RECT 63.545 5.94 63.725 6.18 ;
      RECT 61.71 3.495 62.09 4.175 ;
      RECT 61.92 2.365 62.09 4.175 ;
      RECT 59.84 2.365 60.07 3.035 ;
      RECT 59.84 2.365 62.09 2.535 ;
      RECT 61.37 2.045 61.54 2.535 ;
      RECT 61.36 3.155 61.53 4.005 ;
      RECT 60.445 3.155 61.75 3.325 ;
      RECT 61.505 2.705 61.75 3.325 ;
      RECT 60.445 2.785 60.615 3.325 ;
      RECT 60.24 2.785 60.615 2.955 ;
      RECT 60.42 6.265 61.115 6.895 ;
      RECT 60.945 4.685 61.115 6.895 ;
      RECT 60.85 4.685 61.18 5.665 ;
      RECT 60.45 3.495 60.78 4.175 ;
      RECT 59.54 3.495 59.94 4.175 ;
      RECT 59.54 3.495 60.78 3.665 ;
      RECT 59.04 3.075 59.36 4.175 ;
      RECT 59.04 3.075 59.49 3.325 ;
      RECT 59.04 3.075 59.67 3.245 ;
      RECT 59.5 2.025 59.67 3.245 ;
      RECT 59.5 2.025 60.455 2.195 ;
      RECT 59.04 6.265 59.735 6.895 ;
      RECT 59.565 4.685 59.735 6.895 ;
      RECT 59.47 4.685 59.8 5.665 ;
      RECT 59.06 5.825 59.395 6.075 ;
      RECT 58.515 5.825 58.85 6.075 ;
      RECT 58.515 5.875 59.395 6.045 ;
      RECT 58.175 6.265 58.87 6.895 ;
      RECT 58.175 4.685 58.345 6.895 ;
      RECT 58.11 4.685 58.44 5.665 ;
      RECT 57.67 3.205 58 4.16 ;
      RECT 57.67 3.205 58.35 3.375 ;
      RECT 58.18 1.965 58.35 3.375 ;
      RECT 58.09 1.965 58.42 2.605 ;
      RECT 57.15 3.205 57.48 4.16 ;
      RECT 56.8 3.205 57.48 3.375 ;
      RECT 56.8 1.965 56.97 3.375 ;
      RECT 56.73 1.965 57.06 2.605 ;
      RECT 56.94 5.875 57.11 6.725 ;
      RECT 56.215 5.825 56.55 6.075 ;
      RECT 56.215 5.875 57.11 6.045 ;
      RECT 56.28 2.785 56.63 3.035 ;
      RECT 55.76 2.785 56.09 3.035 ;
      RECT 55.76 2.815 56.63 2.985 ;
      RECT 55.875 6.265 56.57 6.895 ;
      RECT 55.875 4.685 56.045 6.895 ;
      RECT 55.81 4.685 56.14 5.665 ;
      RECT 55.37 5.825 55.705 6.095 ;
      RECT 54.9 5.875 55.705 6.045 ;
      RECT 55.34 3.195 55.67 4.175 ;
      RECT 55.34 1.965 55.59 4.175 ;
      RECT 55.34 1.965 55.67 2.595 ;
      RECT 52.81 7.855 52.98 8.305 ;
      RECT 52.865 6.075 53.035 8.025 ;
      RECT 52.81 5.015 52.98 6.245 ;
      RECT 52.29 5.015 52.46 8.305 ;
      RECT 52.29 7.315 52.695 7.645 ;
      RECT 52.29 6.475 52.695 6.805 ;
      RECT 50.12 1.74 50.29 2.935 ;
      RECT 50.12 1.74 50.585 1.91 ;
      RECT 50.12 6.97 50.585 7.14 ;
      RECT 50.12 5.945 50.29 7.14 ;
      RECT 49.13 1.74 49.3 2.935 ;
      RECT 49.13 1.74 49.595 1.91 ;
      RECT 49.13 6.97 49.595 7.14 ;
      RECT 49.13 5.945 49.3 7.14 ;
      RECT 47.275 2.635 47.445 3.865 ;
      RECT 47.33 0.855 47.5 2.805 ;
      RECT 47.275 0.575 47.445 1.025 ;
      RECT 47.275 7.855 47.445 8.305 ;
      RECT 47.33 6.075 47.5 8.025 ;
      RECT 47.275 5.015 47.445 6.245 ;
      RECT 46.755 0.575 46.925 3.865 ;
      RECT 46.755 2.075 47.16 2.405 ;
      RECT 46.755 1.235 47.16 1.565 ;
      RECT 46.755 5.015 46.925 8.305 ;
      RECT 46.755 7.315 47.16 7.645 ;
      RECT 46.755 6.475 47.16 6.805 ;
      RECT 46.335 5.94 46.505 7.22 ;
      RECT 46.325 5.94 46.505 6.18 ;
      RECT 44.49 3.495 44.87 4.175 ;
      RECT 44.7 2.365 44.87 4.175 ;
      RECT 42.62 2.365 42.85 3.035 ;
      RECT 42.62 2.365 44.87 2.535 ;
      RECT 44.15 2.045 44.32 2.535 ;
      RECT 44.14 3.155 44.31 4.005 ;
      RECT 43.225 3.155 44.53 3.325 ;
      RECT 44.285 2.705 44.53 3.325 ;
      RECT 43.225 2.785 43.395 3.325 ;
      RECT 43.02 2.785 43.395 2.955 ;
      RECT 43.2 6.265 43.895 6.895 ;
      RECT 43.725 4.685 43.895 6.895 ;
      RECT 43.63 4.685 43.96 5.665 ;
      RECT 43.23 3.495 43.56 4.175 ;
      RECT 42.32 3.495 42.72 4.175 ;
      RECT 42.32 3.495 43.56 3.665 ;
      RECT 41.82 3.075 42.14 4.175 ;
      RECT 41.82 3.075 42.27 3.325 ;
      RECT 41.82 3.075 42.45 3.245 ;
      RECT 42.28 2.025 42.45 3.245 ;
      RECT 42.28 2.025 43.235 2.195 ;
      RECT 41.82 6.265 42.515 6.895 ;
      RECT 42.345 4.685 42.515 6.895 ;
      RECT 42.25 4.685 42.58 5.665 ;
      RECT 41.84 5.825 42.175 6.075 ;
      RECT 41.295 5.825 41.63 6.075 ;
      RECT 41.295 5.875 42.175 6.045 ;
      RECT 40.955 6.265 41.65 6.895 ;
      RECT 40.955 4.685 41.125 6.895 ;
      RECT 40.89 4.685 41.22 5.665 ;
      RECT 40.45 3.205 40.78 4.16 ;
      RECT 40.45 3.205 41.13 3.375 ;
      RECT 40.96 1.965 41.13 3.375 ;
      RECT 40.87 1.965 41.2 2.605 ;
      RECT 39.93 3.205 40.26 4.16 ;
      RECT 39.58 3.205 40.26 3.375 ;
      RECT 39.58 1.965 39.75 3.375 ;
      RECT 39.51 1.965 39.84 2.605 ;
      RECT 39.72 5.875 39.89 6.725 ;
      RECT 38.995 5.825 39.33 6.075 ;
      RECT 38.995 5.875 39.89 6.045 ;
      RECT 39.06 2.785 39.41 3.035 ;
      RECT 38.54 2.785 38.87 3.035 ;
      RECT 38.54 2.815 39.41 2.985 ;
      RECT 38.655 6.265 39.35 6.895 ;
      RECT 38.655 4.685 38.825 6.895 ;
      RECT 38.59 4.685 38.92 5.665 ;
      RECT 38.15 5.825 38.485 6.095 ;
      RECT 37.68 5.875 38.485 6.045 ;
      RECT 38.12 3.195 38.45 4.175 ;
      RECT 38.12 1.965 38.37 4.175 ;
      RECT 38.12 1.965 38.45 2.595 ;
      RECT 35.59 7.855 35.76 8.305 ;
      RECT 35.645 6.075 35.815 8.025 ;
      RECT 35.59 5.015 35.76 6.245 ;
      RECT 35.07 5.015 35.24 8.305 ;
      RECT 35.07 7.315 35.475 7.645 ;
      RECT 35.07 6.475 35.475 6.805 ;
      RECT 32.9 1.74 33.07 2.935 ;
      RECT 32.9 1.74 33.365 1.91 ;
      RECT 32.9 6.97 33.365 7.14 ;
      RECT 32.9 5.945 33.07 7.14 ;
      RECT 31.91 1.74 32.08 2.935 ;
      RECT 31.91 1.74 32.375 1.91 ;
      RECT 31.91 6.97 32.375 7.14 ;
      RECT 31.91 5.945 32.08 7.14 ;
      RECT 30.055 2.635 30.225 3.865 ;
      RECT 30.11 0.855 30.28 2.805 ;
      RECT 30.055 0.575 30.225 1.025 ;
      RECT 30.055 7.855 30.225 8.305 ;
      RECT 30.11 6.075 30.28 8.025 ;
      RECT 30.055 5.015 30.225 6.245 ;
      RECT 29.535 0.575 29.705 3.865 ;
      RECT 29.535 2.075 29.94 2.405 ;
      RECT 29.535 1.235 29.94 1.565 ;
      RECT 29.535 5.015 29.705 8.305 ;
      RECT 29.535 7.315 29.94 7.645 ;
      RECT 29.535 6.475 29.94 6.805 ;
      RECT 29.115 5.94 29.285 7.22 ;
      RECT 29.105 5.94 29.285 6.18 ;
      RECT 27.27 3.495 27.65 4.175 ;
      RECT 27.48 2.365 27.65 4.175 ;
      RECT 25.4 2.365 25.63 3.035 ;
      RECT 25.4 2.365 27.65 2.535 ;
      RECT 26.93 2.045 27.1 2.535 ;
      RECT 26.92 3.155 27.09 4.005 ;
      RECT 26.005 3.155 27.31 3.325 ;
      RECT 27.065 2.705 27.31 3.325 ;
      RECT 26.005 2.785 26.175 3.325 ;
      RECT 25.8 2.785 26.175 2.955 ;
      RECT 25.98 6.265 26.675 6.895 ;
      RECT 26.505 4.685 26.675 6.895 ;
      RECT 26.41 4.685 26.74 5.665 ;
      RECT 26.01 3.495 26.34 4.175 ;
      RECT 25.1 3.495 25.5 4.175 ;
      RECT 25.1 3.495 26.34 3.665 ;
      RECT 24.6 3.075 24.92 4.175 ;
      RECT 24.6 3.075 25.05 3.325 ;
      RECT 24.6 3.075 25.23 3.245 ;
      RECT 25.06 2.025 25.23 3.245 ;
      RECT 25.06 2.025 26.015 2.195 ;
      RECT 24.6 6.265 25.295 6.895 ;
      RECT 25.125 4.685 25.295 6.895 ;
      RECT 25.03 4.685 25.36 5.665 ;
      RECT 24.62 5.825 24.955 6.075 ;
      RECT 24.075 5.825 24.41 6.075 ;
      RECT 24.075 5.875 24.955 6.045 ;
      RECT 23.735 6.265 24.43 6.895 ;
      RECT 23.735 4.685 23.905 6.895 ;
      RECT 23.67 4.685 24 5.665 ;
      RECT 23.23 3.205 23.56 4.16 ;
      RECT 23.23 3.205 23.91 3.375 ;
      RECT 23.74 1.965 23.91 3.375 ;
      RECT 23.65 1.965 23.98 2.605 ;
      RECT 22.71 3.205 23.04 4.16 ;
      RECT 22.36 3.205 23.04 3.375 ;
      RECT 22.36 1.965 22.53 3.375 ;
      RECT 22.29 1.965 22.62 2.605 ;
      RECT 22.5 5.875 22.67 6.725 ;
      RECT 21.775 5.825 22.11 6.075 ;
      RECT 21.775 5.875 22.67 6.045 ;
      RECT 21.84 2.785 22.19 3.035 ;
      RECT 21.32 2.785 21.65 3.035 ;
      RECT 21.32 2.815 22.19 2.985 ;
      RECT 21.435 6.265 22.13 6.895 ;
      RECT 21.435 4.685 21.605 6.895 ;
      RECT 21.37 4.685 21.7 5.665 ;
      RECT 20.93 5.825 21.265 6.095 ;
      RECT 20.46 5.875 21.265 6.045 ;
      RECT 20.9 3.195 21.23 4.175 ;
      RECT 20.9 1.965 21.15 4.175 ;
      RECT 20.9 1.965 21.23 2.595 ;
      RECT 18.37 7.855 18.54 8.305 ;
      RECT 18.425 6.075 18.595 8.025 ;
      RECT 18.37 5.015 18.54 6.245 ;
      RECT 17.85 5.015 18.02 8.305 ;
      RECT 17.85 7.315 18.255 7.645 ;
      RECT 17.85 6.475 18.255 6.805 ;
      RECT 15.68 1.74 15.85 2.935 ;
      RECT 15.68 1.74 16.145 1.91 ;
      RECT 15.68 6.97 16.145 7.14 ;
      RECT 15.68 5.945 15.85 7.14 ;
      RECT 14.69 1.74 14.86 2.935 ;
      RECT 14.69 1.74 15.155 1.91 ;
      RECT 14.69 6.97 15.155 7.14 ;
      RECT 14.69 5.945 14.86 7.14 ;
      RECT 12.835 2.635 13.005 3.865 ;
      RECT 12.89 0.855 13.06 2.805 ;
      RECT 12.835 0.575 13.005 1.025 ;
      RECT 12.835 7.855 13.005 8.305 ;
      RECT 12.89 6.075 13.06 8.025 ;
      RECT 12.835 5.015 13.005 6.245 ;
      RECT 12.315 0.575 12.485 3.865 ;
      RECT 12.315 2.075 12.72 2.405 ;
      RECT 12.315 1.235 12.72 1.565 ;
      RECT 12.315 5.015 12.485 8.305 ;
      RECT 12.315 7.315 12.72 7.645 ;
      RECT 12.315 6.475 12.72 6.805 ;
      RECT 11.895 5.94 12.065 7.22 ;
      RECT 11.885 5.94 12.065 6.18 ;
      RECT 10.05 3.495 10.43 4.175 ;
      RECT 10.26 2.365 10.43 4.175 ;
      RECT 8.18 2.365 8.41 3.035 ;
      RECT 8.18 2.365 10.43 2.535 ;
      RECT 9.71 2.045 9.88 2.535 ;
      RECT 9.7 3.155 9.87 4.005 ;
      RECT 8.785 3.155 10.09 3.325 ;
      RECT 9.845 2.705 10.09 3.325 ;
      RECT 8.785 2.785 8.955 3.325 ;
      RECT 8.58 2.785 8.955 2.955 ;
      RECT 8.76 6.265 9.455 6.895 ;
      RECT 9.285 4.685 9.455 6.895 ;
      RECT 9.19 4.685 9.52 5.665 ;
      RECT 8.79 3.495 9.12 4.175 ;
      RECT 7.88 3.495 8.28 4.175 ;
      RECT 7.88 3.495 9.12 3.665 ;
      RECT 7.38 3.075 7.7 4.175 ;
      RECT 7.38 3.075 7.83 3.325 ;
      RECT 7.38 3.075 8.01 3.245 ;
      RECT 7.84 2.025 8.01 3.245 ;
      RECT 7.84 2.025 8.795 2.195 ;
      RECT 7.38 6.265 8.075 6.895 ;
      RECT 7.905 4.685 8.075 6.895 ;
      RECT 7.81 4.685 8.14 5.665 ;
      RECT 7.4 5.825 7.735 6.075 ;
      RECT 6.855 5.825 7.19 6.075 ;
      RECT 6.855 5.875 7.735 6.045 ;
      RECT 6.515 6.265 7.21 6.895 ;
      RECT 6.515 4.685 6.685 6.895 ;
      RECT 6.45 4.685 6.78 5.665 ;
      RECT 6.01 3.205 6.34 4.16 ;
      RECT 6.01 3.205 6.69 3.375 ;
      RECT 6.52 1.965 6.69 3.375 ;
      RECT 6.43 1.965 6.76 2.605 ;
      RECT 5.49 3.205 5.82 4.16 ;
      RECT 5.14 3.205 5.82 3.375 ;
      RECT 5.14 1.965 5.31 3.375 ;
      RECT 5.07 1.965 5.4 2.605 ;
      RECT 5.28 5.875 5.45 6.725 ;
      RECT 4.555 5.825 4.89 6.075 ;
      RECT 4.555 5.875 5.45 6.045 ;
      RECT 4.62 2.785 4.97 3.035 ;
      RECT 4.1 2.785 4.43 3.035 ;
      RECT 4.1 2.815 4.97 2.985 ;
      RECT 4.215 6.265 4.91 6.895 ;
      RECT 4.215 4.685 4.385 6.895 ;
      RECT 4.15 4.685 4.48 5.665 ;
      RECT 3.71 5.825 4.045 6.095 ;
      RECT 3.24 5.875 4.045 6.045 ;
      RECT 3.68 3.195 4.01 4.175 ;
      RECT 3.68 1.965 3.93 4.175 ;
      RECT 3.68 1.965 4.01 2.595 ;
      RECT 1.15 7.855 1.32 8.305 ;
      RECT 1.205 6.075 1.375 8.025 ;
      RECT 1.15 5.015 1.32 6.245 ;
      RECT 0.63 5.015 0.8 8.305 ;
      RECT 0.63 7.315 1.035 7.645 ;
      RECT 0.63 6.475 1.035 6.805 ;
      RECT -2.26 7.855 -2.09 8.305 ;
      RECT -2.205 6.075 -2.035 8.025 ;
      RECT -2.26 5.015 -2.09 6.245 ;
      RECT -2.78 5.015 -2.61 8.305 ;
      RECT -2.78 7.315 -2.375 7.645 ;
      RECT -2.78 6.475 -2.375 6.805 ;
      RECT 84.93 0.575 85.1 1.085 ;
      RECT 84.93 2.395 85.1 3.865 ;
      RECT 84.93 5.015 85.1 6.485 ;
      RECT 84.93 7.795 85.1 8.305 ;
      RECT 83.94 0.575 84.11 1.085 ;
      RECT 83.94 2.395 84.11 3.865 ;
      RECT 83.94 5.015 84.11 6.485 ;
      RECT 83.94 7.795 84.11 8.305 ;
      RECT 82.575 0.575 82.745 3.865 ;
      RECT 82.575 5.015 82.745 8.305 ;
      RECT 82.145 0.575 82.315 1.085 ;
      RECT 82.145 1.655 82.315 3.865 ;
      RECT 82.145 5.015 82.315 7.225 ;
      RECT 82.145 7.795 82.315 8.305 ;
      RECT 80.775 1.66 80.945 2.935 ;
      RECT 78.505 5.825 78.84 6.095 ;
      RECT 78.005 2.785 78.555 2.985 ;
      RECT 77.66 5.825 77.995 6.075 ;
      RECT 77.125 5.825 77.46 6.095 ;
      RECT 75.74 2.785 76.09 3.035 ;
      RECT 74.88 2.785 75.23 3.035 ;
      RECT 74.36 2.785 74.71 3.035 ;
      RECT 70.89 5.015 71.06 8.305 ;
      RECT 70.46 5.015 70.63 7.225 ;
      RECT 70.46 7.795 70.63 8.305 ;
      RECT 69.09 5.945 69.26 7.22 ;
      RECT 67.71 0.575 67.88 1.085 ;
      RECT 67.71 2.395 67.88 3.865 ;
      RECT 67.71 5.015 67.88 6.485 ;
      RECT 67.71 7.795 67.88 8.305 ;
      RECT 66.72 0.575 66.89 1.085 ;
      RECT 66.72 2.395 66.89 3.865 ;
      RECT 66.72 5.015 66.89 6.485 ;
      RECT 66.72 7.795 66.89 8.305 ;
      RECT 65.355 0.575 65.525 3.865 ;
      RECT 65.355 5.015 65.525 8.305 ;
      RECT 64.925 0.575 65.095 1.085 ;
      RECT 64.925 1.655 65.095 3.865 ;
      RECT 64.925 5.015 65.095 7.225 ;
      RECT 64.925 7.795 65.095 8.305 ;
      RECT 63.555 1.66 63.725 2.935 ;
      RECT 61.285 5.825 61.62 6.095 ;
      RECT 60.785 2.785 61.335 2.985 ;
      RECT 60.44 5.825 60.775 6.075 ;
      RECT 59.905 5.825 60.24 6.095 ;
      RECT 58.52 2.785 58.87 3.035 ;
      RECT 57.66 2.785 58.01 3.035 ;
      RECT 57.14 2.785 57.49 3.035 ;
      RECT 53.67 5.015 53.84 8.305 ;
      RECT 53.24 5.015 53.41 7.225 ;
      RECT 53.24 7.795 53.41 8.305 ;
      RECT 51.87 5.945 52.04 7.22 ;
      RECT 50.49 0.575 50.66 1.085 ;
      RECT 50.49 2.395 50.66 3.865 ;
      RECT 50.49 5.015 50.66 6.485 ;
      RECT 50.49 7.795 50.66 8.305 ;
      RECT 49.5 0.575 49.67 1.085 ;
      RECT 49.5 2.395 49.67 3.865 ;
      RECT 49.5 5.015 49.67 6.485 ;
      RECT 49.5 7.795 49.67 8.305 ;
      RECT 48.135 0.575 48.305 3.865 ;
      RECT 48.135 5.015 48.305 8.305 ;
      RECT 47.705 0.575 47.875 1.085 ;
      RECT 47.705 1.655 47.875 3.865 ;
      RECT 47.705 5.015 47.875 7.225 ;
      RECT 47.705 7.795 47.875 8.305 ;
      RECT 46.335 1.66 46.505 2.935 ;
      RECT 44.065 5.825 44.4 6.095 ;
      RECT 43.565 2.785 44.115 2.985 ;
      RECT 43.22 5.825 43.555 6.075 ;
      RECT 42.685 5.825 43.02 6.095 ;
      RECT 41.3 2.785 41.65 3.035 ;
      RECT 40.44 2.785 40.79 3.035 ;
      RECT 39.92 2.785 40.27 3.035 ;
      RECT 36.45 5.015 36.62 8.305 ;
      RECT 36.02 5.015 36.19 7.225 ;
      RECT 36.02 7.795 36.19 8.305 ;
      RECT 34.65 5.945 34.82 7.22 ;
      RECT 33.27 0.575 33.44 1.085 ;
      RECT 33.27 2.395 33.44 3.865 ;
      RECT 33.27 5.015 33.44 6.485 ;
      RECT 33.27 7.795 33.44 8.305 ;
      RECT 32.28 0.575 32.45 1.085 ;
      RECT 32.28 2.395 32.45 3.865 ;
      RECT 32.28 5.015 32.45 6.485 ;
      RECT 32.28 7.795 32.45 8.305 ;
      RECT 30.915 0.575 31.085 3.865 ;
      RECT 30.915 5.015 31.085 8.305 ;
      RECT 30.485 0.575 30.655 1.085 ;
      RECT 30.485 1.655 30.655 3.865 ;
      RECT 30.485 5.015 30.655 7.225 ;
      RECT 30.485 7.795 30.655 8.305 ;
      RECT 29.115 1.66 29.285 2.935 ;
      RECT 26.845 5.825 27.18 6.095 ;
      RECT 26.345 2.785 26.895 2.985 ;
      RECT 26 5.825 26.335 6.075 ;
      RECT 25.465 5.825 25.8 6.095 ;
      RECT 24.08 2.785 24.43 3.035 ;
      RECT 23.22 2.785 23.57 3.035 ;
      RECT 22.7 2.785 23.05 3.035 ;
      RECT 19.23 5.015 19.4 8.305 ;
      RECT 18.8 5.015 18.97 7.225 ;
      RECT 18.8 7.795 18.97 8.305 ;
      RECT 17.43 5.945 17.6 7.22 ;
      RECT 16.05 0.575 16.22 1.085 ;
      RECT 16.05 2.395 16.22 3.865 ;
      RECT 16.05 5.015 16.22 6.485 ;
      RECT 16.05 7.795 16.22 8.305 ;
      RECT 15.06 0.575 15.23 1.085 ;
      RECT 15.06 2.395 15.23 3.865 ;
      RECT 15.06 5.015 15.23 6.485 ;
      RECT 15.06 7.795 15.23 8.305 ;
      RECT 13.695 0.575 13.865 3.865 ;
      RECT 13.695 5.015 13.865 8.305 ;
      RECT 13.265 0.575 13.435 1.085 ;
      RECT 13.265 1.655 13.435 3.865 ;
      RECT 13.265 5.015 13.435 7.225 ;
      RECT 13.265 7.795 13.435 8.305 ;
      RECT 11.895 1.66 12.065 2.935 ;
      RECT 9.625 5.825 9.96 6.095 ;
      RECT 9.125 2.785 9.675 2.985 ;
      RECT 8.78 5.825 9.115 6.075 ;
      RECT 8.245 5.825 8.58 6.095 ;
      RECT 6.86 2.785 7.21 3.035 ;
      RECT 6 2.785 6.35 3.035 ;
      RECT 5.48 2.785 5.83 3.035 ;
      RECT 2.01 5.015 2.18 8.305 ;
      RECT 1.58 5.015 1.75 7.225 ;
      RECT 1.58 7.795 1.75 8.305 ;
      RECT 0.21 5.945 0.38 7.22 ;
      RECT -1.83 5.015 -1.66 7.225 ;
      RECT -1.83 7.795 -1.66 8.305 ;
      RECT -3.2 5.945 -3.03 7.22 ;
  END
END sky130_osu_ring_oscillator_mpr2ct_8_b0r1

MACRO sky130_osu_ring_oscillator_mpr2ct_8_b0r2
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 3.43 0 ;
  SIZE 88.9 BY 8.88 ;
  SYMMETRY X Y R90 ;
  SITE CoreSite ;
  OBS
    LAYER met3 ;
      RECT 71.5 7.435 77.515 7.735 ;
      RECT 77.215 5.805 77.515 7.735 ;
      RECT 76.16 5.785 76.46 7.735 ;
      RECT 75.13 6.48 75.43 7.735 ;
      RECT 71.5 7.035 71.8 7.735 ;
      RECT 70.365 7 70.735 7.37 ;
      RECT 70.365 7.035 71.8 7.335 ;
      RECT 75.1 6.48 75.43 6.81 ;
      RECT 74.63 6.495 75.43 6.795 ;
      RECT 75.01 6.455 75.31 6.795 ;
      RECT 77.14 5.805 77.515 6.17 ;
      RECT 77.205 5.765 77.505 6.17 ;
      RECT 76.12 5.785 76.46 6.135 ;
      RECT 76.135 5.745 76.435 6.135 ;
      RECT 76.11 5.79 76.46 6.12 ;
      RECT 77.14 5.805 77.95 6.105 ;
      RECT 75.64 5.805 76.46 6.105 ;
      RECT 77.15 5.79 77.505 6.17 ;
      RECT 76.8 3.755 77.13 4.085 ;
      RECT 76.8 3.77 77.6 4.07 ;
      RECT 76.815 3.725 77.115 4.085 ;
      RECT 76.46 3.075 76.79 3.405 ;
      RECT 76.46 3.09 77.26 3.39 ;
      RECT 76.545 3.065 76.845 3.39 ;
      RECT 75.78 4.155 76.11 4.485 ;
      RECT 73.74 4.155 74.07 4.485 ;
      RECT 73.74 4.17 76.11 4.47 ;
      RECT 75.43 3.415 75.76 3.745 ;
      RECT 74.97 3.43 75.77 3.73 ;
      RECT 75.1 2.225 75.43 2.555 ;
      RECT 74.63 2.24 75.43 2.54 ;
      RECT 75.09 2.235 75.43 2.54 ;
      RECT 74.42 5.79 74.75 6.12 ;
      RECT 73.95 5.805 74.75 6.105 ;
      RECT 54.28 7.435 60.295 7.735 ;
      RECT 59.995 5.805 60.295 7.735 ;
      RECT 58.94 5.785 59.24 7.735 ;
      RECT 57.91 6.48 58.21 7.735 ;
      RECT 54.28 7.035 54.58 7.735 ;
      RECT 53.145 7 53.515 7.37 ;
      RECT 53.145 7.035 54.58 7.335 ;
      RECT 57.88 6.48 58.21 6.81 ;
      RECT 57.41 6.495 58.21 6.795 ;
      RECT 57.79 6.455 58.09 6.795 ;
      RECT 59.92 5.805 60.295 6.17 ;
      RECT 59.985 5.765 60.285 6.17 ;
      RECT 58.9 5.785 59.24 6.135 ;
      RECT 58.915 5.745 59.215 6.135 ;
      RECT 58.89 5.79 59.24 6.12 ;
      RECT 59.92 5.805 60.73 6.105 ;
      RECT 58.42 5.805 59.24 6.105 ;
      RECT 59.93 5.79 60.285 6.17 ;
      RECT 59.58 3.755 59.91 4.085 ;
      RECT 59.58 3.77 60.38 4.07 ;
      RECT 59.595 3.725 59.895 4.085 ;
      RECT 59.24 3.075 59.57 3.405 ;
      RECT 59.24 3.09 60.04 3.39 ;
      RECT 59.325 3.065 59.625 3.39 ;
      RECT 58.56 4.155 58.89 4.485 ;
      RECT 56.52 4.155 56.85 4.485 ;
      RECT 56.52 4.17 58.89 4.47 ;
      RECT 58.21 3.415 58.54 3.745 ;
      RECT 57.75 3.43 58.55 3.73 ;
      RECT 57.88 2.225 58.21 2.555 ;
      RECT 57.41 2.24 58.21 2.54 ;
      RECT 57.87 2.235 58.21 2.54 ;
      RECT 57.2 5.79 57.53 6.12 ;
      RECT 56.73 5.805 57.53 6.105 ;
      RECT 37.06 7.435 43.075 7.735 ;
      RECT 42.775 5.805 43.075 7.735 ;
      RECT 41.72 5.785 42.02 7.735 ;
      RECT 40.69 6.48 40.99 7.735 ;
      RECT 37.06 7.035 37.36 7.735 ;
      RECT 35.925 7 36.295 7.37 ;
      RECT 35.925 7.035 37.36 7.335 ;
      RECT 40.66 6.48 40.99 6.81 ;
      RECT 40.19 6.495 40.99 6.795 ;
      RECT 40.57 6.455 40.87 6.795 ;
      RECT 42.7 5.805 43.075 6.17 ;
      RECT 42.765 5.765 43.065 6.17 ;
      RECT 41.68 5.785 42.02 6.135 ;
      RECT 41.695 5.745 41.995 6.135 ;
      RECT 41.67 5.79 42.02 6.12 ;
      RECT 42.7 5.805 43.51 6.105 ;
      RECT 41.2 5.805 42.02 6.105 ;
      RECT 42.71 5.79 43.065 6.17 ;
      RECT 42.36 3.755 42.69 4.085 ;
      RECT 42.36 3.77 43.16 4.07 ;
      RECT 42.375 3.725 42.675 4.085 ;
      RECT 42.02 3.075 42.35 3.405 ;
      RECT 42.02 3.09 42.82 3.39 ;
      RECT 42.105 3.065 42.405 3.39 ;
      RECT 41.34 4.155 41.67 4.485 ;
      RECT 39.3 4.155 39.63 4.485 ;
      RECT 39.3 4.17 41.67 4.47 ;
      RECT 40.99 3.415 41.32 3.745 ;
      RECT 40.53 3.43 41.33 3.73 ;
      RECT 40.66 2.225 40.99 2.555 ;
      RECT 40.19 2.24 40.99 2.54 ;
      RECT 40.65 2.235 40.99 2.54 ;
      RECT 39.98 5.79 40.31 6.12 ;
      RECT 39.51 5.805 40.31 6.105 ;
      RECT 19.84 7.435 25.855 7.735 ;
      RECT 25.555 5.805 25.855 7.735 ;
      RECT 24.5 5.785 24.8 7.735 ;
      RECT 23.47 6.48 23.77 7.735 ;
      RECT 19.84 7.035 20.14 7.735 ;
      RECT 18.705 7 19.075 7.37 ;
      RECT 18.705 7.035 20.14 7.335 ;
      RECT 23.44 6.48 23.77 6.81 ;
      RECT 22.97 6.495 23.77 6.795 ;
      RECT 23.35 6.455 23.65 6.795 ;
      RECT 25.48 5.805 25.855 6.17 ;
      RECT 25.545 5.765 25.845 6.17 ;
      RECT 24.46 5.785 24.8 6.135 ;
      RECT 24.475 5.745 24.775 6.135 ;
      RECT 24.45 5.79 24.8 6.12 ;
      RECT 25.48 5.805 26.29 6.105 ;
      RECT 23.98 5.805 24.8 6.105 ;
      RECT 25.49 5.79 25.845 6.17 ;
      RECT 25.14 3.755 25.47 4.085 ;
      RECT 25.14 3.77 25.94 4.07 ;
      RECT 25.155 3.725 25.455 4.085 ;
      RECT 24.8 3.075 25.13 3.405 ;
      RECT 24.8 3.09 25.6 3.39 ;
      RECT 24.885 3.065 25.185 3.39 ;
      RECT 24.12 4.155 24.45 4.485 ;
      RECT 22.08 4.155 22.41 4.485 ;
      RECT 22.08 4.17 24.45 4.47 ;
      RECT 23.77 3.415 24.1 3.745 ;
      RECT 23.31 3.43 24.11 3.73 ;
      RECT 23.44 2.225 23.77 2.555 ;
      RECT 22.97 2.24 23.77 2.54 ;
      RECT 23.43 2.235 23.77 2.54 ;
      RECT 22.76 5.79 23.09 6.12 ;
      RECT 22.29 5.805 23.09 6.105 ;
      RECT 2.62 7.435 8.635 7.735 ;
      RECT 8.335 5.805 8.635 7.735 ;
      RECT 7.28 5.785 7.58 7.735 ;
      RECT 6.25 6.48 6.55 7.735 ;
      RECT 2.62 7.035 2.92 7.735 ;
      RECT 1.485 7 1.855 7.37 ;
      RECT 1.485 7.035 2.92 7.335 ;
      RECT 6.22 6.48 6.55 6.81 ;
      RECT 5.75 6.495 6.55 6.795 ;
      RECT 6.13 6.455 6.43 6.795 ;
      RECT 8.26 5.805 8.635 6.17 ;
      RECT 8.325 5.765 8.625 6.17 ;
      RECT 7.24 5.785 7.58 6.135 ;
      RECT 7.255 5.745 7.555 6.135 ;
      RECT 7.23 5.79 7.58 6.12 ;
      RECT 8.26 5.805 9.07 6.105 ;
      RECT 6.76 5.805 7.58 6.105 ;
      RECT 8.27 5.79 8.625 6.17 ;
      RECT 7.92 3.755 8.25 4.085 ;
      RECT 7.92 3.77 8.72 4.07 ;
      RECT 7.935 3.725 8.235 4.085 ;
      RECT 7.58 3.075 7.91 3.405 ;
      RECT 7.58 3.09 8.38 3.39 ;
      RECT 7.665 3.065 7.965 3.39 ;
      RECT 6.9 4.155 7.23 4.485 ;
      RECT 4.86 4.155 5.19 4.485 ;
      RECT 4.86 4.17 7.23 4.47 ;
      RECT 6.55 3.415 6.88 3.745 ;
      RECT 6.09 3.43 6.89 3.73 ;
      RECT 6.22 2.225 6.55 2.555 ;
      RECT 5.75 2.24 6.55 2.54 ;
      RECT 6.21 2.235 6.55 2.54 ;
      RECT 5.54 5.79 5.87 6.12 ;
      RECT 5.07 5.805 5.87 6.105 ;
    LAYER via2 ;
      RECT 77.215 5.855 77.415 6.055 ;
      RECT 76.865 3.82 77.065 4.02 ;
      RECT 76.525 3.14 76.725 3.34 ;
      RECT 76.175 5.855 76.375 6.055 ;
      RECT 75.845 4.22 76.045 4.42 ;
      RECT 75.495 3.48 75.695 3.68 ;
      RECT 75.165 2.29 75.365 2.49 ;
      RECT 75.165 6.545 75.365 6.745 ;
      RECT 74.485 5.855 74.685 6.055 ;
      RECT 73.805 4.22 74.005 4.42 ;
      RECT 70.45 7.085 70.65 7.285 ;
      RECT 59.995 5.855 60.195 6.055 ;
      RECT 59.645 3.82 59.845 4.02 ;
      RECT 59.305 3.14 59.505 3.34 ;
      RECT 58.955 5.855 59.155 6.055 ;
      RECT 58.625 4.22 58.825 4.42 ;
      RECT 58.275 3.48 58.475 3.68 ;
      RECT 57.945 2.29 58.145 2.49 ;
      RECT 57.945 6.545 58.145 6.745 ;
      RECT 57.265 5.855 57.465 6.055 ;
      RECT 56.585 4.22 56.785 4.42 ;
      RECT 53.23 7.085 53.43 7.285 ;
      RECT 42.775 5.855 42.975 6.055 ;
      RECT 42.425 3.82 42.625 4.02 ;
      RECT 42.085 3.14 42.285 3.34 ;
      RECT 41.735 5.855 41.935 6.055 ;
      RECT 41.405 4.22 41.605 4.42 ;
      RECT 41.055 3.48 41.255 3.68 ;
      RECT 40.725 2.29 40.925 2.49 ;
      RECT 40.725 6.545 40.925 6.745 ;
      RECT 40.045 5.855 40.245 6.055 ;
      RECT 39.365 4.22 39.565 4.42 ;
      RECT 36.01 7.085 36.21 7.285 ;
      RECT 25.555 5.855 25.755 6.055 ;
      RECT 25.205 3.82 25.405 4.02 ;
      RECT 24.865 3.14 25.065 3.34 ;
      RECT 24.515 5.855 24.715 6.055 ;
      RECT 24.185 4.22 24.385 4.42 ;
      RECT 23.835 3.48 24.035 3.68 ;
      RECT 23.505 2.29 23.705 2.49 ;
      RECT 23.505 6.545 23.705 6.745 ;
      RECT 22.825 5.855 23.025 6.055 ;
      RECT 22.145 4.22 22.345 4.42 ;
      RECT 18.79 7.085 18.99 7.285 ;
      RECT 8.335 5.855 8.535 6.055 ;
      RECT 7.985 3.82 8.185 4.02 ;
      RECT 7.645 3.14 7.845 3.34 ;
      RECT 7.295 5.855 7.495 6.055 ;
      RECT 6.965 4.22 7.165 4.42 ;
      RECT 6.615 3.48 6.815 3.68 ;
      RECT 6.285 2.29 6.485 2.49 ;
      RECT 6.285 6.545 6.485 6.745 ;
      RECT 5.605 5.855 5.805 6.055 ;
      RECT 4.925 4.22 5.125 4.42 ;
      RECT 1.57 7.085 1.77 7.285 ;
    LAYER met2 ;
      RECT -2.22 8.6 85.1 8.77 ;
      RECT 84.93 7.3 85.1 8.77 ;
      RECT -2.22 6.255 -2.05 8.77 ;
      RECT 84.895 7.3 85.22 7.625 ;
      RECT -2.265 6.255 -1.985 6.595 ;
      RECT 81.74 6.28 82.06 6.605 ;
      RECT 81.77 5.695 81.94 6.605 ;
      RECT 81.77 5.695 81.945 6.045 ;
      RECT 81.77 5.695 82.745 5.87 ;
      RECT 82.57 1.965 82.745 5.87 ;
      RECT 75.125 2.205 75.405 2.575 ;
      RECT 75.125 2.345 79.775 2.52 ;
      RECT 79.6 2.025 79.775 2.52 ;
      RECT 80.07 1.995 80.395 2.32 ;
      RECT 82.515 1.965 82.865 2.315 ;
      RECT 79.6 2.025 82.865 2.195 ;
      RECT 70.89 8.29 81.585 8.46 ;
      RECT 81.425 2.395 81.585 8.46 ;
      RECT 70.89 6.545 71.06 8.46 ;
      RECT 82.54 6.655 82.865 6.98 ;
      RECT 67.71 6.655 68.035 6.98 ;
      RECT 81.425 6.745 82.865 6.915 ;
      RECT 70.84 6.545 71.12 6.885 ;
      RECT 67.71 6.685 71.12 6.855 ;
      RECT 81.74 2.365 82.06 2.685 ;
      RECT 81.425 2.395 82.06 2.565 ;
      RECT 71.395 7.55 80.945 7.72 ;
      RECT 80.775 5.855 80.945 7.72 ;
      RECT 71.395 5.86 71.565 7.72 ;
      RECT 71.34 5.86 71.62 6.2 ;
      RECT 80.695 5.855 81.02 6.18 ;
      RECT 80.765 3.495 80.935 6.18 ;
      RECT 80.695 3.495 81.02 3.82 ;
      RECT 78.195 6.48 78.455 6.8 ;
      RECT 78.255 2.74 78.395 6.8 ;
      RECT 78.195 2.74 78.455 3.06 ;
      RECT 77.515 4.78 77.775 5.1 ;
      RECT 77.575 3.76 77.715 5.1 ;
      RECT 77.515 3.76 77.775 4.08 ;
      RECT 76.495 6.48 76.755 6.8 ;
      RECT 76.555 5.21 76.695 6.8 ;
      RECT 75.875 5.21 76.695 5.35 ;
      RECT 75.875 2.74 76.015 5.35 ;
      RECT 75.805 4.135 76.085 4.505 ;
      RECT 75.815 2.74 76.075 3.06 ;
      RECT 73.765 4.135 74.045 4.505 ;
      RECT 73.835 2.4 73.975 4.505 ;
      RECT 73.775 2.4 74.035 2.72 ;
      RECT 73.095 4.78 73.355 5.1 ;
      RECT 73.155 2.74 73.295 5.1 ;
      RECT 73.095 2.74 73.355 3.06 ;
      RECT 64.52 6.28 64.84 6.605 ;
      RECT 64.55 5.695 64.72 6.605 ;
      RECT 64.55 5.695 64.725 6.045 ;
      RECT 64.55 5.695 65.525 5.87 ;
      RECT 65.35 1.965 65.525 5.87 ;
      RECT 57.905 2.205 58.185 2.575 ;
      RECT 57.905 2.345 62.555 2.52 ;
      RECT 62.38 2.025 62.555 2.52 ;
      RECT 62.85 1.995 63.175 2.32 ;
      RECT 65.295 1.965 65.645 2.315 ;
      RECT 62.38 2.025 65.645 2.195 ;
      RECT 53.67 8.29 64.365 8.46 ;
      RECT 64.205 2.395 64.365 8.46 ;
      RECT 53.67 6.545 53.84 8.46 ;
      RECT 65.32 6.655 65.645 6.98 ;
      RECT 50.49 6.655 50.815 6.98 ;
      RECT 64.205 6.745 65.645 6.915 ;
      RECT 53.62 6.545 53.9 6.885 ;
      RECT 50.49 6.685 53.9 6.855 ;
      RECT 64.52 2.365 64.84 2.685 ;
      RECT 64.205 2.395 64.84 2.565 ;
      RECT 54.175 7.55 63.725 7.72 ;
      RECT 63.555 5.855 63.725 7.72 ;
      RECT 54.175 5.86 54.345 7.72 ;
      RECT 54.12 5.86 54.4 6.2 ;
      RECT 63.475 5.855 63.8 6.18 ;
      RECT 63.545 3.495 63.715 6.18 ;
      RECT 63.475 3.495 63.8 3.82 ;
      RECT 60.975 6.48 61.235 6.8 ;
      RECT 61.035 2.74 61.175 6.8 ;
      RECT 60.975 2.74 61.235 3.06 ;
      RECT 60.295 4.78 60.555 5.1 ;
      RECT 60.355 3.76 60.495 5.1 ;
      RECT 60.295 3.76 60.555 4.08 ;
      RECT 59.275 6.48 59.535 6.8 ;
      RECT 59.335 5.21 59.475 6.8 ;
      RECT 58.655 5.21 59.475 5.35 ;
      RECT 58.655 2.74 58.795 5.35 ;
      RECT 58.585 4.135 58.865 4.505 ;
      RECT 58.595 2.74 58.855 3.06 ;
      RECT 56.545 4.135 56.825 4.505 ;
      RECT 56.615 2.4 56.755 4.505 ;
      RECT 56.555 2.4 56.815 2.72 ;
      RECT 55.875 4.78 56.135 5.1 ;
      RECT 55.935 2.74 56.075 5.1 ;
      RECT 55.875 2.74 56.135 3.06 ;
      RECT 47.3 6.28 47.62 6.605 ;
      RECT 47.33 5.695 47.5 6.605 ;
      RECT 47.33 5.695 47.505 6.045 ;
      RECT 47.33 5.695 48.305 5.87 ;
      RECT 48.13 1.965 48.305 5.87 ;
      RECT 40.685 2.205 40.965 2.575 ;
      RECT 40.685 2.345 45.335 2.52 ;
      RECT 45.16 2.025 45.335 2.52 ;
      RECT 45.63 1.995 45.955 2.32 ;
      RECT 48.075 1.965 48.425 2.315 ;
      RECT 45.16 2.025 48.425 2.195 ;
      RECT 36.45 8.29 47.145 8.46 ;
      RECT 46.985 2.395 47.145 8.46 ;
      RECT 36.45 6.545 36.62 8.46 ;
      RECT 48.1 6.655 48.425 6.98 ;
      RECT 33.27 6.655 33.595 6.98 ;
      RECT 46.985 6.745 48.425 6.915 ;
      RECT 36.4 6.545 36.68 6.885 ;
      RECT 33.27 6.685 36.69 6.855 ;
      RECT 47.3 2.365 47.62 2.685 ;
      RECT 46.985 2.395 47.62 2.565 ;
      RECT 36.955 7.55 46.505 7.72 ;
      RECT 46.335 5.855 46.505 7.72 ;
      RECT 36.955 5.86 37.125 7.72 ;
      RECT 36.9 5.86 37.18 6.2 ;
      RECT 46.255 5.855 46.58 6.18 ;
      RECT 46.325 3.495 46.495 6.18 ;
      RECT 46.255 3.495 46.58 3.82 ;
      RECT 43.755 6.48 44.015 6.8 ;
      RECT 43.815 2.74 43.955 6.8 ;
      RECT 43.755 2.74 44.015 3.06 ;
      RECT 43.075 4.78 43.335 5.1 ;
      RECT 43.135 3.76 43.275 5.1 ;
      RECT 43.075 3.76 43.335 4.08 ;
      RECT 42.055 6.48 42.315 6.8 ;
      RECT 42.115 5.21 42.255 6.8 ;
      RECT 41.435 5.21 42.255 5.35 ;
      RECT 41.435 2.74 41.575 5.35 ;
      RECT 41.365 4.135 41.645 4.505 ;
      RECT 41.375 2.74 41.635 3.06 ;
      RECT 39.325 4.135 39.605 4.505 ;
      RECT 39.395 2.4 39.535 4.505 ;
      RECT 39.335 2.4 39.595 2.72 ;
      RECT 38.655 4.78 38.915 5.1 ;
      RECT 38.715 2.74 38.855 5.1 ;
      RECT 38.655 2.74 38.915 3.06 ;
      RECT 30.08 6.28 30.4 6.605 ;
      RECT 30.11 5.695 30.28 6.605 ;
      RECT 30.11 5.695 30.285 6.045 ;
      RECT 30.11 5.695 31.085 5.87 ;
      RECT 30.91 1.965 31.085 5.87 ;
      RECT 23.465 2.205 23.745 2.575 ;
      RECT 23.465 2.345 28.115 2.52 ;
      RECT 27.94 2.025 28.115 2.52 ;
      RECT 28.41 1.995 28.735 2.32 ;
      RECT 30.855 1.965 31.205 2.315 ;
      RECT 27.94 2.025 31.205 2.195 ;
      RECT 19.23 8.29 29.925 8.46 ;
      RECT 29.765 2.395 29.925 8.46 ;
      RECT 19.23 6.545 19.4 8.46 ;
      RECT 30.88 6.655 31.205 6.98 ;
      RECT 16.05 6.655 16.375 6.98 ;
      RECT 29.765 6.745 31.205 6.915 ;
      RECT 19.18 6.545 19.46 6.885 ;
      RECT 16.05 6.685 19.46 6.855 ;
      RECT 30.08 2.365 30.4 2.685 ;
      RECT 29.765 2.395 30.4 2.565 ;
      RECT 19.735 7.55 29.285 7.72 ;
      RECT 29.115 5.855 29.285 7.72 ;
      RECT 19.735 5.86 19.905 7.72 ;
      RECT 19.68 5.86 19.96 6.2 ;
      RECT 29.035 5.855 29.36 6.18 ;
      RECT 29.105 3.495 29.275 6.18 ;
      RECT 29.035 3.495 29.36 3.82 ;
      RECT 26.535 6.48 26.795 6.8 ;
      RECT 26.595 2.74 26.735 6.8 ;
      RECT 26.535 2.74 26.795 3.06 ;
      RECT 25.855 4.78 26.115 5.1 ;
      RECT 25.915 3.76 26.055 5.1 ;
      RECT 25.855 3.76 26.115 4.08 ;
      RECT 24.835 6.48 25.095 6.8 ;
      RECT 24.895 5.21 25.035 6.8 ;
      RECT 24.215 5.21 25.035 5.35 ;
      RECT 24.215 2.74 24.355 5.35 ;
      RECT 24.145 4.135 24.425 4.505 ;
      RECT 24.155 2.74 24.415 3.06 ;
      RECT 22.105 4.135 22.385 4.505 ;
      RECT 22.175 2.4 22.315 4.505 ;
      RECT 22.115 2.4 22.375 2.72 ;
      RECT 21.435 4.78 21.695 5.1 ;
      RECT 21.495 2.74 21.635 5.1 ;
      RECT 21.435 2.74 21.695 3.06 ;
      RECT 12.86 6.28 13.18 6.605 ;
      RECT 12.89 5.695 13.06 6.605 ;
      RECT 12.89 5.695 13.065 6.045 ;
      RECT 12.89 5.695 13.865 5.87 ;
      RECT 13.69 1.965 13.865 5.87 ;
      RECT 6.245 2.205 6.525 2.575 ;
      RECT 6.245 2.345 10.895 2.52 ;
      RECT 10.72 2.025 10.895 2.52 ;
      RECT 11.19 1.995 11.515 2.32 ;
      RECT 13.635 1.965 13.985 2.315 ;
      RECT 10.72 2.025 13.985 2.195 ;
      RECT 2.01 8.29 12.705 8.46 ;
      RECT 12.545 2.395 12.705 8.46 ;
      RECT 2.01 6.545 2.18 8.46 ;
      RECT -1.89 6.995 -1.61 7.335 ;
      RECT -1.89 7.06 -0.685 7.23 ;
      RECT -0.855 6.685 -0.685 7.23 ;
      RECT 13.66 6.655 13.985 6.98 ;
      RECT 12.545 6.745 13.985 6.915 ;
      RECT 1.96 6.545 2.24 6.885 ;
      RECT -0.855 6.685 2.24 6.855 ;
      RECT 12.86 2.365 13.18 2.685 ;
      RECT 12.545 2.395 13.18 2.565 ;
      RECT 2.515 7.55 12.065 7.72 ;
      RECT 11.895 5.855 12.065 7.72 ;
      RECT 2.515 5.86 2.685 7.72 ;
      RECT 2.46 5.86 2.74 6.2 ;
      RECT 11.815 5.855 12.14 6.18 ;
      RECT 11.885 3.495 12.055 6.18 ;
      RECT 11.815 3.495 12.14 3.82 ;
      RECT 9.315 6.48 9.575 6.8 ;
      RECT 9.375 2.74 9.515 6.8 ;
      RECT 9.315 2.74 9.575 3.06 ;
      RECT 8.635 4.78 8.895 5.1 ;
      RECT 8.695 3.76 8.835 5.1 ;
      RECT 8.635 3.76 8.895 4.08 ;
      RECT 7.615 6.48 7.875 6.8 ;
      RECT 7.675 5.21 7.815 6.8 ;
      RECT 6.995 5.21 7.815 5.35 ;
      RECT 6.995 2.74 7.135 5.35 ;
      RECT 6.925 4.135 7.205 4.505 ;
      RECT 6.935 2.74 7.195 3.06 ;
      RECT 4.885 4.135 5.165 4.505 ;
      RECT 4.955 2.4 5.095 4.505 ;
      RECT 4.895 2.4 5.155 2.72 ;
      RECT 4.215 4.78 4.475 5.1 ;
      RECT 4.275 2.74 4.415 5.1 ;
      RECT 4.215 2.74 4.475 3.06 ;
      RECT 77.175 5.77 77.455 6.14 ;
      RECT 76.825 3.735 77.105 4.105 ;
      RECT 76.485 3.055 76.765 3.425 ;
      RECT 76.135 5.77 76.415 6.14 ;
      RECT 75.455 3.395 75.735 3.765 ;
      RECT 75.125 6.46 75.405 6.83 ;
      RECT 74.445 5.77 74.725 6.14 ;
      RECT 70.365 7 70.735 7.37 ;
      RECT 59.955 5.77 60.235 6.14 ;
      RECT 59.605 3.735 59.885 4.105 ;
      RECT 59.265 3.055 59.545 3.425 ;
      RECT 58.915 5.77 59.195 6.14 ;
      RECT 58.235 3.395 58.515 3.765 ;
      RECT 57.905 6.46 58.185 6.83 ;
      RECT 57.225 5.77 57.505 6.14 ;
      RECT 53.145 7 53.515 7.37 ;
      RECT 42.735 5.77 43.015 6.14 ;
      RECT 42.385 3.735 42.665 4.105 ;
      RECT 42.045 3.055 42.325 3.425 ;
      RECT 41.695 5.77 41.975 6.14 ;
      RECT 41.015 3.395 41.295 3.765 ;
      RECT 40.685 6.46 40.965 6.83 ;
      RECT 40.005 5.77 40.285 6.14 ;
      RECT 35.925 7 36.295 7.37 ;
      RECT 25.515 5.77 25.795 6.14 ;
      RECT 25.165 3.735 25.445 4.105 ;
      RECT 24.825 3.055 25.105 3.425 ;
      RECT 24.475 5.77 24.755 6.14 ;
      RECT 23.795 3.395 24.075 3.765 ;
      RECT 23.465 6.46 23.745 6.83 ;
      RECT 22.785 5.77 23.065 6.14 ;
      RECT 18.705 7 19.075 7.37 ;
      RECT 8.295 5.77 8.575 6.14 ;
      RECT 7.945 3.735 8.225 4.105 ;
      RECT 7.605 3.055 7.885 3.425 ;
      RECT 7.255 5.77 7.535 6.14 ;
      RECT 6.575 3.395 6.855 3.765 ;
      RECT 6.245 6.46 6.525 6.83 ;
      RECT 5.565 5.77 5.845 6.14 ;
      RECT 1.485 7 1.855 7.37 ;
    LAYER via1 ;
      RECT 84.985 7.385 85.135 7.535 ;
      RECT 82.63 6.74 82.78 6.89 ;
      RECT 82.615 2.065 82.765 2.215 ;
      RECT 81.825 2.45 81.975 2.6 ;
      RECT 81.825 6.37 81.975 6.52 ;
      RECT 80.785 3.58 80.935 3.73 ;
      RECT 80.785 5.94 80.935 6.09 ;
      RECT 80.16 2.08 80.31 2.23 ;
      RECT 78.25 2.825 78.4 2.975 ;
      RECT 78.25 6.565 78.4 6.715 ;
      RECT 77.57 3.845 77.72 3.995 ;
      RECT 77.57 4.865 77.72 5.015 ;
      RECT 77.23 5.885 77.38 6.035 ;
      RECT 76.89 3.845 77.04 3.995 ;
      RECT 76.55 3.165 76.7 3.315 ;
      RECT 76.55 6.565 76.7 6.715 ;
      RECT 76.2 5.885 76.35 6.035 ;
      RECT 75.87 2.825 76.02 2.975 ;
      RECT 75.53 3.505 75.68 3.655 ;
      RECT 75.19 2.315 75.34 2.465 ;
      RECT 75.19 6.565 75.34 6.715 ;
      RECT 74.51 5.885 74.66 6.035 ;
      RECT 73.83 2.485 73.98 2.635 ;
      RECT 73.15 2.825 73.3 2.975 ;
      RECT 73.15 4.865 73.3 5.015 ;
      RECT 71.405 5.955 71.555 6.105 ;
      RECT 70.905 6.64 71.055 6.79 ;
      RECT 70.475 7.11 70.625 7.26 ;
      RECT 67.8 6.74 67.95 6.89 ;
      RECT 65.41 6.74 65.56 6.89 ;
      RECT 65.395 2.065 65.545 2.215 ;
      RECT 64.605 2.45 64.755 2.6 ;
      RECT 64.605 6.37 64.755 6.52 ;
      RECT 63.565 3.58 63.715 3.73 ;
      RECT 63.565 5.94 63.715 6.09 ;
      RECT 62.94 2.08 63.09 2.23 ;
      RECT 61.03 2.825 61.18 2.975 ;
      RECT 61.03 6.565 61.18 6.715 ;
      RECT 60.35 3.845 60.5 3.995 ;
      RECT 60.35 4.865 60.5 5.015 ;
      RECT 60.01 5.885 60.16 6.035 ;
      RECT 59.67 3.845 59.82 3.995 ;
      RECT 59.33 3.165 59.48 3.315 ;
      RECT 59.33 6.565 59.48 6.715 ;
      RECT 58.98 5.885 59.13 6.035 ;
      RECT 58.65 2.825 58.8 2.975 ;
      RECT 58.31 3.505 58.46 3.655 ;
      RECT 57.97 2.315 58.12 2.465 ;
      RECT 57.97 6.565 58.12 6.715 ;
      RECT 57.29 5.885 57.44 6.035 ;
      RECT 56.61 2.485 56.76 2.635 ;
      RECT 55.93 2.825 56.08 2.975 ;
      RECT 55.93 4.865 56.08 5.015 ;
      RECT 54.185 5.955 54.335 6.105 ;
      RECT 53.685 6.64 53.835 6.79 ;
      RECT 53.255 7.11 53.405 7.26 ;
      RECT 50.58 6.74 50.73 6.89 ;
      RECT 48.19 6.74 48.34 6.89 ;
      RECT 48.175 2.065 48.325 2.215 ;
      RECT 47.385 2.45 47.535 2.6 ;
      RECT 47.385 6.37 47.535 6.52 ;
      RECT 46.345 3.58 46.495 3.73 ;
      RECT 46.345 5.94 46.495 6.09 ;
      RECT 45.72 2.08 45.87 2.23 ;
      RECT 43.81 2.825 43.96 2.975 ;
      RECT 43.81 6.565 43.96 6.715 ;
      RECT 43.13 3.845 43.28 3.995 ;
      RECT 43.13 4.865 43.28 5.015 ;
      RECT 42.79 5.885 42.94 6.035 ;
      RECT 42.45 3.845 42.6 3.995 ;
      RECT 42.11 3.165 42.26 3.315 ;
      RECT 42.11 6.565 42.26 6.715 ;
      RECT 41.76 5.885 41.91 6.035 ;
      RECT 41.43 2.825 41.58 2.975 ;
      RECT 41.09 3.505 41.24 3.655 ;
      RECT 40.75 2.315 40.9 2.465 ;
      RECT 40.75 6.565 40.9 6.715 ;
      RECT 40.07 5.885 40.22 6.035 ;
      RECT 39.39 2.485 39.54 2.635 ;
      RECT 38.71 2.825 38.86 2.975 ;
      RECT 38.71 4.865 38.86 5.015 ;
      RECT 36.965 5.955 37.115 6.105 ;
      RECT 36.465 6.64 36.615 6.79 ;
      RECT 36.035 7.11 36.185 7.26 ;
      RECT 33.36 6.74 33.51 6.89 ;
      RECT 30.97 6.74 31.12 6.89 ;
      RECT 30.955 2.065 31.105 2.215 ;
      RECT 30.165 2.45 30.315 2.6 ;
      RECT 30.165 6.37 30.315 6.52 ;
      RECT 29.125 3.58 29.275 3.73 ;
      RECT 29.125 5.94 29.275 6.09 ;
      RECT 28.5 2.08 28.65 2.23 ;
      RECT 26.59 2.825 26.74 2.975 ;
      RECT 26.59 6.565 26.74 6.715 ;
      RECT 25.91 3.845 26.06 3.995 ;
      RECT 25.91 4.865 26.06 5.015 ;
      RECT 25.57 5.885 25.72 6.035 ;
      RECT 25.23 3.845 25.38 3.995 ;
      RECT 24.89 3.165 25.04 3.315 ;
      RECT 24.89 6.565 25.04 6.715 ;
      RECT 24.54 5.885 24.69 6.035 ;
      RECT 24.21 2.825 24.36 2.975 ;
      RECT 23.87 3.505 24.02 3.655 ;
      RECT 23.53 2.315 23.68 2.465 ;
      RECT 23.53 6.565 23.68 6.715 ;
      RECT 22.85 5.885 23 6.035 ;
      RECT 22.17 2.485 22.32 2.635 ;
      RECT 21.49 2.825 21.64 2.975 ;
      RECT 21.49 4.865 21.64 5.015 ;
      RECT 19.745 5.955 19.895 6.105 ;
      RECT 19.245 6.64 19.395 6.79 ;
      RECT 18.815 7.11 18.965 7.26 ;
      RECT 16.14 6.74 16.29 6.89 ;
      RECT 13.75 6.74 13.9 6.89 ;
      RECT 13.735 2.065 13.885 2.215 ;
      RECT 12.945 2.45 13.095 2.6 ;
      RECT 12.945 6.37 13.095 6.52 ;
      RECT 11.905 3.58 12.055 3.73 ;
      RECT 11.905 5.94 12.055 6.09 ;
      RECT 11.28 2.08 11.43 2.23 ;
      RECT 9.37 2.825 9.52 2.975 ;
      RECT 9.37 6.565 9.52 6.715 ;
      RECT 8.69 3.845 8.84 3.995 ;
      RECT 8.69 4.865 8.84 5.015 ;
      RECT 8.35 5.885 8.5 6.035 ;
      RECT 8.01 3.845 8.16 3.995 ;
      RECT 7.67 3.165 7.82 3.315 ;
      RECT 7.67 6.565 7.82 6.715 ;
      RECT 7.32 5.885 7.47 6.035 ;
      RECT 6.99 2.825 7.14 2.975 ;
      RECT 6.65 3.505 6.8 3.655 ;
      RECT 6.31 2.315 6.46 2.465 ;
      RECT 6.31 6.565 6.46 6.715 ;
      RECT 5.63 5.885 5.78 6.035 ;
      RECT 4.95 2.485 5.1 2.635 ;
      RECT 4.27 2.825 4.42 2.975 ;
      RECT 4.27 4.865 4.42 5.015 ;
      RECT 2.525 5.955 2.675 6.105 ;
      RECT 2.025 6.64 2.175 6.79 ;
      RECT 1.595 7.11 1.745 7.26 ;
      RECT -1.825 7.09 -1.675 7.24 ;
      RECT -2.2 6.35 -2.05 6.5 ;
    LAYER met1 ;
      RECT 72.035 0 79.395 1.95 ;
      RECT 54.815 0 62.175 1.95 ;
      RECT 37.595 0 44.955 1.95 ;
      RECT 20.375 0 27.735 1.95 ;
      RECT 3.155 0 10.515 1.95 ;
      RECT 72.035 0 79.69 1.795 ;
      RECT 54.815 0 62.47 1.795 ;
      RECT 37.595 0 45.25 1.795 ;
      RECT 20.375 0 28.03 1.795 ;
      RECT 3.155 0 10.81 1.795 ;
      RECT 72.03 0 79.69 1.635 ;
      RECT 54.81 0 62.47 1.635 ;
      RECT 37.59 0 45.25 1.635 ;
      RECT 20.37 0 28.03 1.635 ;
      RECT 3.15 0 10.81 1.635 ;
      RECT -3.385 0 85.47 0.305 ;
      RECT 79.485 4.135 85.47 4.745 ;
      RECT 68.905 4.13 71.655 4.745 ;
      RECT 62.265 4.135 68.25 4.745 ;
      RECT 51.685 4.13 54.435 4.745 ;
      RECT 45.045 4.135 51.03 4.745 ;
      RECT 34.465 4.13 37.215 4.745 ;
      RECT 27.825 4.135 33.81 4.745 ;
      RECT 17.245 4.13 19.995 4.745 ;
      RECT 10.605 4.135 16.59 4.745 ;
      RECT 0.025 4.13 2.775 4.745 ;
      RECT -3.385 4.13 -0.635 4.745 ;
      RECT 62.265 4.19 72.41 4.74 ;
      RECT 45.045 4.19 55.19 4.74 ;
      RECT 27.825 4.19 37.97 4.74 ;
      RECT 10.605 4.19 20.75 4.74 ;
      RECT -3.385 4.19 3.53 4.74 ;
      RECT -3.385 4.19 85.47 4.67 ;
      RECT 79.48 4.135 85.47 4.67 ;
      RECT 62.26 4.135 72.39 4.67 ;
      RECT 68.245 4.13 72.39 4.74 ;
      RECT 45.04 4.135 55.17 4.67 ;
      RECT 51.025 4.13 55.17 4.74 ;
      RECT 27.82 4.135 37.95 4.67 ;
      RECT 33.805 4.13 37.95 4.74 ;
      RECT 10.6 4.135 20.73 4.67 ;
      RECT 16.585 4.13 20.73 4.74 ;
      RECT -3.385 4.13 3.51 4.74 ;
      RECT -3.385 8.575 85.47 8.88 ;
      RECT 72.305 7.18 79.505 8.88 ;
      RECT 69.625 6.315 69.795 8.88 ;
      RECT 55.085 7.18 62.285 8.88 ;
      RECT 52.405 6.315 52.575 8.88 ;
      RECT 37.865 7.18 45.065 8.88 ;
      RECT 35.185 6.315 35.355 8.88 ;
      RECT 20.645 7.18 27.845 8.88 ;
      RECT 17.965 6.315 18.135 8.88 ;
      RECT 3.425 7.18 10.625 8.88 ;
      RECT 0.745 6.315 0.915 8.88 ;
      RECT 72.035 6.91 79.395 7.39 ;
      RECT 54.815 6.91 62.175 7.39 ;
      RECT 37.595 6.91 44.955 7.39 ;
      RECT 20.375 6.91 27.735 7.39 ;
      RECT 3.155 6.91 10.515 7.39 ;
      RECT 70.025 6.285 70.315 6.515 ;
      RECT 52.805 6.285 53.095 6.515 ;
      RECT 35.585 6.285 35.875 6.515 ;
      RECT 18.365 6.285 18.655 6.515 ;
      RECT 1.145 6.285 1.435 6.515 ;
      RECT 69.625 6.315 70.315 6.485 ;
      RECT 52.405 6.315 53.095 6.485 ;
      RECT 35.185 6.315 35.875 6.485 ;
      RECT 17.965 6.315 18.655 6.485 ;
      RECT 0.745 6.315 1.435 6.485 ;
      RECT 84.87 7.765 85.16 7.995 ;
      RECT 84.93 6.285 85.1 7.995 ;
      RECT 84.895 7.3 85.22 7.625 ;
      RECT 84.87 6.285 85.16 6.515 ;
      RECT 84.87 2.365 85.16 2.595 ;
      RECT 84.93 0.885 85.1 2.595 ;
      RECT 84.87 0.885 85.16 1.115 ;
      RECT 84.46 2.735 84.79 2.965 ;
      RECT 84.46 2.765 84.96 2.935 ;
      RECT 84.46 2.395 84.65 2.965 ;
      RECT 83.88 2.365 84.17 2.595 ;
      RECT 83.88 2.395 84.65 2.565 ;
      RECT 83.94 0.885 84.11 2.595 ;
      RECT 83.88 0.885 84.17 1.115 ;
      RECT 83.88 7.765 84.17 7.995 ;
      RECT 83.94 6.285 84.11 7.995 ;
      RECT 83.88 6.285 84.17 6.515 ;
      RECT 83.88 6.325 84.73 6.485 ;
      RECT 84.56 5.915 84.73 6.485 ;
      RECT 83.88 6.32 84.27 6.485 ;
      RECT 84.5 5.915 84.79 6.145 ;
      RECT 84.5 5.945 84.96 6.115 ;
      RECT 83.51 2.735 83.8 2.965 ;
      RECT 83.51 2.765 83.97 2.935 ;
      RECT 83.57 1.655 83.735 2.965 ;
      RECT 82.085 1.625 82.375 1.855 ;
      RECT 82.085 1.655 83.735 1.825 ;
      RECT 82.145 0.885 82.315 1.855 ;
      RECT 82.085 0.885 82.375 1.115 ;
      RECT 82.085 7.765 82.375 7.995 ;
      RECT 82.145 7.025 82.315 7.995 ;
      RECT 82.145 7.12 83.735 7.29 ;
      RECT 83.565 5.915 83.735 7.29 ;
      RECT 82.085 7.025 82.375 7.255 ;
      RECT 83.51 5.915 83.8 6.145 ;
      RECT 83.51 5.945 83.97 6.115 ;
      RECT 82.515 1.965 82.865 2.315 ;
      RECT 82.345 2.025 82.865 2.195 ;
      RECT 82.54 6.655 82.865 6.98 ;
      RECT 82.515 6.655 82.865 6.885 ;
      RECT 82.345 6.685 82.865 6.855 ;
      RECT 81.74 2.365 82.06 2.685 ;
      RECT 81.71 2.365 82.06 2.595 ;
      RECT 81.425 2.395 82.06 2.565 ;
      RECT 81.74 6.28 82.06 6.605 ;
      RECT 81.71 6.285 82.06 6.515 ;
      RECT 81.54 6.315 82.06 6.485 ;
      RECT 80.695 3.495 81.02 3.82 ;
      RECT 80.775 2.735 80.945 3.82 ;
      RECT 80.715 2.735 81.005 2.965 ;
      RECT 80.715 2.765 81.175 2.935 ;
      RECT 80.695 5.855 81.02 6.18 ;
      RECT 80.695 5.945 81.175 6.115 ;
      RECT 77.485 3.79 77.805 4.05 ;
      RECT 78.52 3.805 78.81 4.035 ;
      RECT 77.485 3.85 78.81 3.99 ;
      RECT 77.145 5.83 77.465 6.09 ;
      RECT 78.52 5.845 78.81 6.075 ;
      RECT 78.595 5.55 78.735 6.075 ;
      RECT 77.235 5.55 77.375 6.09 ;
      RECT 77.235 5.55 78.735 5.69 ;
      RECT 78.165 2.77 78.485 3.03 ;
      RECT 77.89 2.83 78.485 2.97 ;
      RECT 75.105 6.51 75.425 6.77 ;
      RECT 74.1 6.525 74.39 6.755 ;
      RECT 74.1 6.57 76.015 6.71 ;
      RECT 75.875 6.23 76.015 6.71 ;
      RECT 75.875 6.23 77.885 6.37 ;
      RECT 77.745 5.845 77.885 6.37 ;
      RECT 77.67 5.845 77.96 6.075 ;
      RECT 77.485 4.81 77.805 5.07 ;
      RECT 75.34 4.825 75.63 5.055 ;
      RECT 75.34 4.87 77.805 5.01 ;
      RECT 76.805 3.79 77.125 4.05 ;
      RECT 74.44 3.805 74.73 4.035 ;
      RECT 74.44 3.85 77.125 3.99 ;
      RECT 76.465 6.51 76.785 6.77 ;
      RECT 76.465 6.57 77.06 6.71 ;
      RECT 76.465 3.11 76.785 3.37 ;
      RECT 76.19 3.17 76.785 3.31 ;
      RECT 75.785 2.77 76.105 3.03 ;
      RECT 75.51 2.83 76.105 2.97 ;
      RECT 75.445 3.45 75.765 3.71 ;
      RECT 72.57 3.465 72.86 3.695 ;
      RECT 72.57 3.51 75.765 3.65 ;
      RECT 75.025 2.79 75.165 3.65 ;
      RECT 74.95 2.79 75.24 3.02 ;
      RECT 75.105 2.26 75.425 2.52 ;
      RECT 75.105 2.275 75.61 2.505 ;
      RECT 75.015 2.32 75.61 2.46 ;
      RECT 74.425 5.83 74.745 6.09 ;
      RECT 72.06 5.845 72.35 6.075 ;
      RECT 72.06 5.89 74.745 6.03 ;
      RECT 74.44 2.79 74.73 3.02 ;
      RECT 73.835 2.835 74.73 2.975 ;
      RECT 73.835 2.43 73.975 2.975 ;
      RECT 73.745 2.43 74.065 2.69 ;
      RECT 73.065 2.77 73.385 3.03 ;
      RECT 72.79 2.83 73.385 2.97 ;
      RECT 73.065 4.81 73.385 5.07 ;
      RECT 72.79 4.87 73.385 5.01 ;
      RECT 71.31 5.89 71.65 6.17 ;
      RECT 69.03 5.915 69.32 6.145 ;
      RECT 69.03 5.945 71.65 6.115 ;
      RECT 70.83 6.575 71.12 6.885 ;
      RECT 70.66 6.685 71.15 6.855 ;
      RECT 70.81 6.575 71.15 6.855 ;
      RECT 70.4 7.765 70.69 7.995 ;
      RECT 70.46 6.995 70.63 7.995 ;
      RECT 70.365 6.995 70.735 7.37 ;
      RECT 67.65 7.765 67.94 7.995 ;
      RECT 67.71 6.285 67.88 7.995 ;
      RECT 67.71 6.655 68.035 6.98 ;
      RECT 67.65 6.285 67.94 6.515 ;
      RECT 67.65 2.365 67.94 2.595 ;
      RECT 67.71 0.885 67.88 2.595 ;
      RECT 67.65 0.885 67.94 1.115 ;
      RECT 67.24 2.735 67.57 2.965 ;
      RECT 67.24 2.765 67.74 2.935 ;
      RECT 67.24 2.395 67.43 2.965 ;
      RECT 66.66 2.365 66.95 2.595 ;
      RECT 66.66 2.395 67.43 2.565 ;
      RECT 66.72 0.885 66.89 2.595 ;
      RECT 66.66 0.885 66.95 1.115 ;
      RECT 66.66 7.765 66.95 7.995 ;
      RECT 66.72 6.285 66.89 7.995 ;
      RECT 66.66 6.285 66.95 6.515 ;
      RECT 66.66 6.325 67.51 6.485 ;
      RECT 67.34 5.915 67.51 6.485 ;
      RECT 66.66 6.32 67.05 6.485 ;
      RECT 67.28 5.915 67.57 6.145 ;
      RECT 67.28 5.945 67.74 6.115 ;
      RECT 66.29 2.735 66.58 2.965 ;
      RECT 66.29 2.765 66.75 2.935 ;
      RECT 66.35 1.655 66.515 2.965 ;
      RECT 64.865 1.625 65.155 1.855 ;
      RECT 64.865 1.655 66.515 1.825 ;
      RECT 64.925 0.885 65.095 1.855 ;
      RECT 64.865 0.885 65.155 1.115 ;
      RECT 64.865 7.765 65.155 7.995 ;
      RECT 64.925 7.025 65.095 7.995 ;
      RECT 64.925 7.12 66.515 7.29 ;
      RECT 66.345 5.915 66.515 7.29 ;
      RECT 64.865 7.025 65.155 7.255 ;
      RECT 66.29 5.915 66.58 6.145 ;
      RECT 66.29 5.945 66.75 6.115 ;
      RECT 65.295 1.965 65.645 2.315 ;
      RECT 65.125 2.025 65.645 2.195 ;
      RECT 65.32 6.655 65.645 6.98 ;
      RECT 65.295 6.655 65.645 6.885 ;
      RECT 65.125 6.685 65.645 6.855 ;
      RECT 64.52 2.365 64.84 2.685 ;
      RECT 64.49 2.365 64.84 2.595 ;
      RECT 64.205 2.395 64.84 2.565 ;
      RECT 64.52 6.28 64.84 6.605 ;
      RECT 64.49 6.285 64.84 6.515 ;
      RECT 64.32 6.315 64.84 6.485 ;
      RECT 63.475 3.495 63.8 3.82 ;
      RECT 63.555 2.735 63.725 3.82 ;
      RECT 63.495 2.735 63.785 2.965 ;
      RECT 63.495 2.765 63.955 2.935 ;
      RECT 63.475 5.855 63.8 6.18 ;
      RECT 63.475 5.945 63.955 6.115 ;
      RECT 60.265 3.79 60.585 4.05 ;
      RECT 61.3 3.805 61.59 4.035 ;
      RECT 60.265 3.85 61.59 3.99 ;
      RECT 59.925 5.83 60.245 6.09 ;
      RECT 61.3 5.845 61.59 6.075 ;
      RECT 61.375 5.55 61.515 6.075 ;
      RECT 60.015 5.55 60.155 6.09 ;
      RECT 60.015 5.55 61.515 5.69 ;
      RECT 60.945 2.77 61.265 3.03 ;
      RECT 60.67 2.83 61.265 2.97 ;
      RECT 57.885 6.51 58.205 6.77 ;
      RECT 56.88 6.525 57.17 6.755 ;
      RECT 56.88 6.57 58.795 6.71 ;
      RECT 58.655 6.23 58.795 6.71 ;
      RECT 58.655 6.23 60.665 6.37 ;
      RECT 60.525 5.845 60.665 6.37 ;
      RECT 60.45 5.845 60.74 6.075 ;
      RECT 60.265 4.81 60.585 5.07 ;
      RECT 58.12 4.825 58.41 5.055 ;
      RECT 58.12 4.87 60.585 5.01 ;
      RECT 59.585 3.79 59.905 4.05 ;
      RECT 57.22 3.805 57.51 4.035 ;
      RECT 57.22 3.85 59.905 3.99 ;
      RECT 59.245 6.51 59.565 6.77 ;
      RECT 59.245 6.57 59.84 6.71 ;
      RECT 59.245 3.11 59.565 3.37 ;
      RECT 58.97 3.17 59.565 3.31 ;
      RECT 58.565 2.77 58.885 3.03 ;
      RECT 58.29 2.83 58.885 2.97 ;
      RECT 58.225 3.45 58.545 3.71 ;
      RECT 55.35 3.465 55.64 3.695 ;
      RECT 55.35 3.51 58.545 3.65 ;
      RECT 57.805 2.79 57.945 3.65 ;
      RECT 57.73 2.79 58.02 3.02 ;
      RECT 57.885 2.26 58.205 2.52 ;
      RECT 57.885 2.275 58.39 2.505 ;
      RECT 57.795 2.32 58.39 2.46 ;
      RECT 57.205 5.83 57.525 6.09 ;
      RECT 54.84 5.845 55.13 6.075 ;
      RECT 54.84 5.89 57.525 6.03 ;
      RECT 57.22 2.79 57.51 3.02 ;
      RECT 56.615 2.835 57.51 2.975 ;
      RECT 56.615 2.43 56.755 2.975 ;
      RECT 56.525 2.43 56.845 2.69 ;
      RECT 55.845 2.77 56.165 3.03 ;
      RECT 55.57 2.83 56.165 2.97 ;
      RECT 55.845 4.81 56.165 5.07 ;
      RECT 55.57 4.87 56.165 5.01 ;
      RECT 54.09 5.89 54.43 6.17 ;
      RECT 51.81 5.915 52.1 6.145 ;
      RECT 51.81 5.945 54.43 6.115 ;
      RECT 53.61 6.575 53.9 6.885 ;
      RECT 53.44 6.685 53.93 6.855 ;
      RECT 53.59 6.575 53.93 6.855 ;
      RECT 53.18 7.765 53.47 7.995 ;
      RECT 53.24 6.995 53.41 7.995 ;
      RECT 53.145 6.995 53.515 7.37 ;
      RECT 50.43 7.765 50.72 7.995 ;
      RECT 50.49 6.285 50.66 7.995 ;
      RECT 50.49 6.655 50.815 6.98 ;
      RECT 50.43 6.285 50.72 6.515 ;
      RECT 50.43 2.365 50.72 2.595 ;
      RECT 50.49 0.885 50.66 2.595 ;
      RECT 50.43 0.885 50.72 1.115 ;
      RECT 50.02 2.735 50.35 2.965 ;
      RECT 50.02 2.765 50.52 2.935 ;
      RECT 50.02 2.395 50.21 2.965 ;
      RECT 49.44 2.365 49.73 2.595 ;
      RECT 49.44 2.395 50.21 2.565 ;
      RECT 49.5 0.885 49.67 2.595 ;
      RECT 49.44 0.885 49.73 1.115 ;
      RECT 49.44 7.765 49.73 7.995 ;
      RECT 49.5 6.285 49.67 7.995 ;
      RECT 49.44 6.285 49.73 6.515 ;
      RECT 49.44 6.325 50.29 6.485 ;
      RECT 50.12 5.915 50.29 6.485 ;
      RECT 49.44 6.32 49.83 6.485 ;
      RECT 50.06 5.915 50.35 6.145 ;
      RECT 50.06 5.945 50.52 6.115 ;
      RECT 49.07 2.735 49.36 2.965 ;
      RECT 49.07 2.765 49.53 2.935 ;
      RECT 49.13 1.655 49.295 2.965 ;
      RECT 47.645 1.625 47.935 1.855 ;
      RECT 47.645 1.655 49.295 1.825 ;
      RECT 47.705 0.885 47.875 1.855 ;
      RECT 47.645 0.885 47.935 1.115 ;
      RECT 47.645 7.765 47.935 7.995 ;
      RECT 47.705 7.025 47.875 7.995 ;
      RECT 47.705 7.12 49.295 7.29 ;
      RECT 49.125 5.915 49.295 7.29 ;
      RECT 47.645 7.025 47.935 7.255 ;
      RECT 49.07 5.915 49.36 6.145 ;
      RECT 49.07 5.945 49.53 6.115 ;
      RECT 48.075 1.965 48.425 2.315 ;
      RECT 47.905 2.025 48.425 2.195 ;
      RECT 48.1 6.655 48.425 6.98 ;
      RECT 48.075 6.655 48.425 6.885 ;
      RECT 47.905 6.685 48.425 6.855 ;
      RECT 47.3 2.365 47.62 2.685 ;
      RECT 47.27 2.365 47.62 2.595 ;
      RECT 46.985 2.395 47.62 2.565 ;
      RECT 47.3 6.28 47.62 6.605 ;
      RECT 47.27 6.285 47.62 6.515 ;
      RECT 47.1 6.315 47.62 6.485 ;
      RECT 46.255 3.495 46.58 3.82 ;
      RECT 46.335 2.735 46.505 3.82 ;
      RECT 46.275 2.735 46.565 2.965 ;
      RECT 46.275 2.765 46.735 2.935 ;
      RECT 46.255 5.855 46.58 6.18 ;
      RECT 46.255 5.945 46.735 6.115 ;
      RECT 43.045 3.79 43.365 4.05 ;
      RECT 44.08 3.805 44.37 4.035 ;
      RECT 43.045 3.85 44.37 3.99 ;
      RECT 42.705 5.83 43.025 6.09 ;
      RECT 44.08 5.845 44.37 6.075 ;
      RECT 44.155 5.55 44.295 6.075 ;
      RECT 42.795 5.55 42.935 6.09 ;
      RECT 42.795 5.55 44.295 5.69 ;
      RECT 43.725 2.77 44.045 3.03 ;
      RECT 43.45 2.83 44.045 2.97 ;
      RECT 40.665 6.51 40.985 6.77 ;
      RECT 39.66 6.525 39.95 6.755 ;
      RECT 39.66 6.57 41.575 6.71 ;
      RECT 41.435 6.23 41.575 6.71 ;
      RECT 41.435 6.23 43.445 6.37 ;
      RECT 43.305 5.845 43.445 6.37 ;
      RECT 43.23 5.845 43.52 6.075 ;
      RECT 43.045 4.81 43.365 5.07 ;
      RECT 40.9 4.825 41.19 5.055 ;
      RECT 40.9 4.87 43.365 5.01 ;
      RECT 42.365 3.79 42.685 4.05 ;
      RECT 40 3.805 40.29 4.035 ;
      RECT 40 3.85 42.685 3.99 ;
      RECT 42.025 6.51 42.345 6.77 ;
      RECT 42.025 6.57 42.62 6.71 ;
      RECT 42.025 3.11 42.345 3.37 ;
      RECT 41.75 3.17 42.345 3.31 ;
      RECT 41.345 2.77 41.665 3.03 ;
      RECT 41.07 2.83 41.665 2.97 ;
      RECT 41.005 3.45 41.325 3.71 ;
      RECT 38.13 3.465 38.42 3.695 ;
      RECT 38.13 3.51 41.325 3.65 ;
      RECT 40.585 2.79 40.725 3.65 ;
      RECT 40.51 2.79 40.8 3.02 ;
      RECT 40.665 2.26 40.985 2.52 ;
      RECT 40.665 2.275 41.17 2.505 ;
      RECT 40.575 2.32 41.17 2.46 ;
      RECT 39.985 5.83 40.305 6.09 ;
      RECT 37.62 5.845 37.91 6.075 ;
      RECT 37.62 5.89 40.305 6.03 ;
      RECT 40 2.79 40.29 3.02 ;
      RECT 39.395 2.835 40.29 2.975 ;
      RECT 39.395 2.43 39.535 2.975 ;
      RECT 39.305 2.43 39.625 2.69 ;
      RECT 38.625 2.77 38.945 3.03 ;
      RECT 38.35 2.83 38.945 2.97 ;
      RECT 38.625 4.81 38.945 5.07 ;
      RECT 38.35 4.87 38.945 5.01 ;
      RECT 36.87 5.89 37.21 6.17 ;
      RECT 34.59 5.915 34.88 6.145 ;
      RECT 34.59 5.945 37.21 6.115 ;
      RECT 36.39 6.575 36.68 6.885 ;
      RECT 36.22 6.685 36.71 6.855 ;
      RECT 36.37 6.575 36.71 6.855 ;
      RECT 35.96 7.765 36.25 7.995 ;
      RECT 36.02 6.995 36.19 7.995 ;
      RECT 35.925 6.995 36.295 7.37 ;
      RECT 33.21 7.765 33.5 7.995 ;
      RECT 33.27 6.285 33.44 7.995 ;
      RECT 33.27 6.655 33.595 6.98 ;
      RECT 33.21 6.285 33.5 6.515 ;
      RECT 33.21 2.365 33.5 2.595 ;
      RECT 33.27 0.885 33.44 2.595 ;
      RECT 33.21 0.885 33.5 1.115 ;
      RECT 32.8 2.735 33.13 2.965 ;
      RECT 32.8 2.765 33.3 2.935 ;
      RECT 32.8 2.395 32.99 2.965 ;
      RECT 32.22 2.365 32.51 2.595 ;
      RECT 32.22 2.395 32.99 2.565 ;
      RECT 32.28 0.885 32.45 2.595 ;
      RECT 32.22 0.885 32.51 1.115 ;
      RECT 32.22 7.765 32.51 7.995 ;
      RECT 32.28 6.285 32.45 7.995 ;
      RECT 32.22 6.285 32.51 6.515 ;
      RECT 32.22 6.325 33.07 6.485 ;
      RECT 32.9 5.915 33.07 6.485 ;
      RECT 32.22 6.32 32.61 6.485 ;
      RECT 32.84 5.915 33.13 6.145 ;
      RECT 32.84 5.945 33.3 6.115 ;
      RECT 31.85 2.735 32.14 2.965 ;
      RECT 31.85 2.765 32.31 2.935 ;
      RECT 31.91 1.655 32.075 2.965 ;
      RECT 30.425 1.625 30.715 1.855 ;
      RECT 30.425 1.655 32.075 1.825 ;
      RECT 30.485 0.885 30.655 1.855 ;
      RECT 30.425 0.885 30.715 1.115 ;
      RECT 30.425 7.765 30.715 7.995 ;
      RECT 30.485 7.025 30.655 7.995 ;
      RECT 30.485 7.12 32.075 7.29 ;
      RECT 31.905 5.915 32.075 7.29 ;
      RECT 30.425 7.025 30.715 7.255 ;
      RECT 31.85 5.915 32.14 6.145 ;
      RECT 31.85 5.945 32.31 6.115 ;
      RECT 30.855 1.965 31.205 2.315 ;
      RECT 30.685 2.025 31.205 2.195 ;
      RECT 30.88 6.655 31.205 6.98 ;
      RECT 30.855 6.655 31.205 6.885 ;
      RECT 30.685 6.685 31.205 6.855 ;
      RECT 30.08 2.365 30.4 2.685 ;
      RECT 30.05 2.365 30.4 2.595 ;
      RECT 29.765 2.395 30.4 2.565 ;
      RECT 30.08 6.28 30.4 6.605 ;
      RECT 30.05 6.285 30.4 6.515 ;
      RECT 29.88 6.315 30.4 6.485 ;
      RECT 29.035 3.495 29.36 3.82 ;
      RECT 29.115 2.735 29.285 3.82 ;
      RECT 29.055 2.735 29.345 2.965 ;
      RECT 29.055 2.765 29.515 2.935 ;
      RECT 29.035 5.855 29.36 6.18 ;
      RECT 29.035 5.945 29.515 6.115 ;
      RECT 25.825 3.79 26.145 4.05 ;
      RECT 26.86 3.805 27.15 4.035 ;
      RECT 25.825 3.85 27.15 3.99 ;
      RECT 25.485 5.83 25.805 6.09 ;
      RECT 26.86 5.845 27.15 6.075 ;
      RECT 26.935 5.55 27.075 6.075 ;
      RECT 25.575 5.55 25.715 6.09 ;
      RECT 25.575 5.55 27.075 5.69 ;
      RECT 26.505 2.77 26.825 3.03 ;
      RECT 26.23 2.83 26.825 2.97 ;
      RECT 23.445 6.51 23.765 6.77 ;
      RECT 22.44 6.525 22.73 6.755 ;
      RECT 22.44 6.57 24.355 6.71 ;
      RECT 24.215 6.23 24.355 6.71 ;
      RECT 24.215 6.23 26.225 6.37 ;
      RECT 26.085 5.845 26.225 6.37 ;
      RECT 26.01 5.845 26.3 6.075 ;
      RECT 25.825 4.81 26.145 5.07 ;
      RECT 23.68 4.825 23.97 5.055 ;
      RECT 23.68 4.87 26.145 5.01 ;
      RECT 25.145 3.79 25.465 4.05 ;
      RECT 22.78 3.805 23.07 4.035 ;
      RECT 22.78 3.85 25.465 3.99 ;
      RECT 24.805 6.51 25.125 6.77 ;
      RECT 24.805 6.57 25.4 6.71 ;
      RECT 24.805 3.11 25.125 3.37 ;
      RECT 24.53 3.17 25.125 3.31 ;
      RECT 24.125 2.77 24.445 3.03 ;
      RECT 23.85 2.83 24.445 2.97 ;
      RECT 23.785 3.45 24.105 3.71 ;
      RECT 20.91 3.465 21.2 3.695 ;
      RECT 20.91 3.51 24.105 3.65 ;
      RECT 23.365 2.79 23.505 3.65 ;
      RECT 23.29 2.79 23.58 3.02 ;
      RECT 23.445 2.26 23.765 2.52 ;
      RECT 23.445 2.275 23.95 2.505 ;
      RECT 23.355 2.32 23.95 2.46 ;
      RECT 22.765 5.83 23.085 6.09 ;
      RECT 20.4 5.845 20.69 6.075 ;
      RECT 20.4 5.89 23.085 6.03 ;
      RECT 22.78 2.79 23.07 3.02 ;
      RECT 22.175 2.835 23.07 2.975 ;
      RECT 22.175 2.43 22.315 2.975 ;
      RECT 22.085 2.43 22.405 2.69 ;
      RECT 21.405 2.77 21.725 3.03 ;
      RECT 21.13 2.83 21.725 2.97 ;
      RECT 21.405 4.81 21.725 5.07 ;
      RECT 21.13 4.87 21.725 5.01 ;
      RECT 19.65 5.89 19.99 6.17 ;
      RECT 17.37 5.915 17.66 6.145 ;
      RECT 17.37 5.945 19.99 6.115 ;
      RECT 19.17 6.575 19.46 6.885 ;
      RECT 19 6.685 19.49 6.855 ;
      RECT 19.15 6.575 19.49 6.855 ;
      RECT 18.74 7.765 19.03 7.995 ;
      RECT 18.8 6.995 18.97 7.995 ;
      RECT 18.705 6.995 19.075 7.37 ;
      RECT 15.99 7.765 16.28 7.995 ;
      RECT 16.05 6.285 16.22 7.995 ;
      RECT 16.05 6.655 16.375 6.98 ;
      RECT 15.99 6.285 16.28 6.515 ;
      RECT 15.99 2.365 16.28 2.595 ;
      RECT 16.05 0.885 16.22 2.595 ;
      RECT 15.99 0.885 16.28 1.115 ;
      RECT 15.58 2.735 15.91 2.965 ;
      RECT 15.58 2.765 16.08 2.935 ;
      RECT 15.58 2.395 15.77 2.965 ;
      RECT 15 2.365 15.29 2.595 ;
      RECT 15 2.395 15.77 2.565 ;
      RECT 15.06 0.885 15.23 2.595 ;
      RECT 15 0.885 15.29 1.115 ;
      RECT 15 7.765 15.29 7.995 ;
      RECT 15.06 6.285 15.23 7.995 ;
      RECT 15 6.285 15.29 6.515 ;
      RECT 15 6.325 15.85 6.485 ;
      RECT 15.68 5.915 15.85 6.485 ;
      RECT 15 6.32 15.39 6.485 ;
      RECT 15.62 5.915 15.91 6.145 ;
      RECT 15.62 5.945 16.08 6.115 ;
      RECT 14.63 2.735 14.92 2.965 ;
      RECT 14.63 2.765 15.09 2.935 ;
      RECT 14.69 1.655 14.855 2.965 ;
      RECT 13.205 1.625 13.495 1.855 ;
      RECT 13.205 1.655 14.855 1.825 ;
      RECT 13.265 0.885 13.435 1.855 ;
      RECT 13.205 0.885 13.495 1.115 ;
      RECT 13.205 7.765 13.495 7.995 ;
      RECT 13.265 7.025 13.435 7.995 ;
      RECT 13.265 7.12 14.855 7.29 ;
      RECT 14.685 5.915 14.855 7.29 ;
      RECT 13.205 7.025 13.495 7.255 ;
      RECT 14.63 5.915 14.92 6.145 ;
      RECT 14.63 5.945 15.09 6.115 ;
      RECT 13.635 1.965 13.985 2.315 ;
      RECT 13.465 2.025 13.985 2.195 ;
      RECT 13.66 6.655 13.985 6.98 ;
      RECT 13.635 6.655 13.985 6.885 ;
      RECT 13.465 6.685 13.985 6.855 ;
      RECT 12.86 2.365 13.18 2.685 ;
      RECT 12.83 2.365 13.18 2.595 ;
      RECT 12.545 2.395 13.18 2.565 ;
      RECT 12.86 6.28 13.18 6.605 ;
      RECT 12.83 6.285 13.18 6.515 ;
      RECT 12.66 6.315 13.18 6.485 ;
      RECT 11.815 3.495 12.14 3.82 ;
      RECT 11.895 2.735 12.065 3.82 ;
      RECT 11.835 2.735 12.125 2.965 ;
      RECT 11.835 2.765 12.295 2.935 ;
      RECT 11.815 5.855 12.14 6.18 ;
      RECT 11.815 5.945 12.295 6.115 ;
      RECT 8.605 3.79 8.925 4.05 ;
      RECT 9.64 3.805 9.93 4.035 ;
      RECT 8.605 3.85 9.93 3.99 ;
      RECT 8.265 5.83 8.585 6.09 ;
      RECT 9.64 5.845 9.93 6.075 ;
      RECT 9.715 5.55 9.855 6.075 ;
      RECT 8.355 5.55 8.495 6.09 ;
      RECT 8.355 5.55 9.855 5.69 ;
      RECT 9.285 2.77 9.605 3.03 ;
      RECT 9.01 2.83 9.605 2.97 ;
      RECT 6.225 6.51 6.545 6.77 ;
      RECT 5.22 6.525 5.51 6.755 ;
      RECT 5.22 6.57 7.135 6.71 ;
      RECT 6.995 6.23 7.135 6.71 ;
      RECT 6.995 6.23 9.005 6.37 ;
      RECT 8.865 5.845 9.005 6.37 ;
      RECT 8.79 5.845 9.08 6.075 ;
      RECT 8.605 4.81 8.925 5.07 ;
      RECT 6.46 4.825 6.75 5.055 ;
      RECT 6.46 4.87 8.925 5.01 ;
      RECT 7.925 3.79 8.245 4.05 ;
      RECT 5.56 3.805 5.85 4.035 ;
      RECT 5.56 3.85 8.245 3.99 ;
      RECT 7.585 6.51 7.905 6.77 ;
      RECT 7.585 6.57 8.18 6.71 ;
      RECT 7.585 3.11 7.905 3.37 ;
      RECT 7.31 3.17 7.905 3.31 ;
      RECT 6.905 2.77 7.225 3.03 ;
      RECT 6.63 2.83 7.225 2.97 ;
      RECT 6.565 3.45 6.885 3.71 ;
      RECT 3.69 3.465 3.98 3.695 ;
      RECT 3.69 3.51 6.885 3.65 ;
      RECT 6.145 2.79 6.285 3.65 ;
      RECT 6.07 2.79 6.36 3.02 ;
      RECT 6.225 2.26 6.545 2.52 ;
      RECT 6.225 2.275 6.73 2.505 ;
      RECT 6.135 2.32 6.73 2.46 ;
      RECT 5.545 5.83 5.865 6.09 ;
      RECT 3.18 5.845 3.47 6.075 ;
      RECT 3.18 5.89 5.865 6.03 ;
      RECT 5.56 2.79 5.85 3.02 ;
      RECT 4.955 2.835 5.85 2.975 ;
      RECT 4.955 2.43 5.095 2.975 ;
      RECT 4.865 2.43 5.185 2.69 ;
      RECT 4.185 2.77 4.505 3.03 ;
      RECT 3.91 2.83 4.505 2.97 ;
      RECT 4.185 4.81 4.505 5.07 ;
      RECT 3.91 4.87 4.505 5.01 ;
      RECT 2.43 5.89 2.77 6.17 ;
      RECT 0.15 5.915 0.44 6.145 ;
      RECT 0.15 5.945 2.77 6.115 ;
      RECT 1.95 6.575 2.24 6.885 ;
      RECT 1.78 6.685 2.27 6.855 ;
      RECT 1.93 6.575 2.27 6.855 ;
      RECT 1.52 7.765 1.81 7.995 ;
      RECT 1.58 6.995 1.75 7.995 ;
      RECT 1.485 6.995 1.855 7.37 ;
      RECT -1.46 6.655 -1.17 6.885 ;
      RECT -1.63 6.685 -1.17 6.855 ;
      RECT -1.89 7.765 -1.6 7.995 ;
      RECT -1.83 7.025 -1.66 7.995 ;
      RECT -1.92 7.025 -1.58 7.305 ;
      RECT -2.295 6.285 -1.955 6.565 ;
      RECT -2.435 6.315 -1.955 6.485 ;
      RECT -3.26 5.915 -2.97 6.145 ;
      RECT -3.26 5.945 -2.8 6.115 ;
      RECT 80.07 1.995 80.395 2.32 ;
      RECT 77.84 6.51 78.485 6.77 ;
      RECT 75.79 5.83 76.435 6.09 ;
      RECT 62.85 1.995 63.175 2.32 ;
      RECT 60.62 6.51 61.265 6.77 ;
      RECT 58.57 5.83 59.215 6.09 ;
      RECT 45.63 1.995 45.955 2.32 ;
      RECT 43.4 6.51 44.045 6.77 ;
      RECT 41.35 5.83 41.995 6.09 ;
      RECT 28.41 1.995 28.735 2.32 ;
      RECT 26.18 6.51 26.825 6.77 ;
      RECT 24.13 5.83 24.775 6.09 ;
      RECT 11.19 1.995 11.515 2.32 ;
      RECT 8.96 6.51 9.605 6.77 ;
      RECT 6.91 5.83 7.555 6.09 ;
    LAYER mcon ;
      RECT 84.93 0.915 85.1 1.085 ;
      RECT 84.93 2.395 85.1 2.565 ;
      RECT 84.93 6.315 85.1 6.485 ;
      RECT 84.93 7.795 85.1 7.965 ;
      RECT 84.58 0.105 84.75 0.275 ;
      RECT 84.58 4.165 84.75 4.335 ;
      RECT 84.58 4.545 84.75 4.715 ;
      RECT 84.58 8.605 84.75 8.775 ;
      RECT 84.56 2.765 84.73 2.935 ;
      RECT 84.56 5.945 84.73 6.115 ;
      RECT 83.94 0.915 84.11 1.085 ;
      RECT 83.94 2.395 84.11 2.565 ;
      RECT 83.94 6.315 84.11 6.485 ;
      RECT 83.94 7.795 84.11 7.965 ;
      RECT 83.59 0.105 83.76 0.275 ;
      RECT 83.59 4.165 83.76 4.335 ;
      RECT 83.59 4.545 83.76 4.715 ;
      RECT 83.59 8.605 83.76 8.775 ;
      RECT 83.57 2.765 83.74 2.935 ;
      RECT 83.57 5.945 83.74 6.115 ;
      RECT 82.885 0.105 83.055 0.275 ;
      RECT 82.885 4.165 83.055 4.335 ;
      RECT 82.885 4.545 83.055 4.715 ;
      RECT 82.885 8.605 83.055 8.775 ;
      RECT 82.575 2.025 82.745 2.195 ;
      RECT 82.575 6.685 82.745 6.855 ;
      RECT 82.205 0.105 82.375 0.275 ;
      RECT 82.205 8.605 82.375 8.775 ;
      RECT 82.145 0.915 82.315 1.085 ;
      RECT 82.145 1.655 82.315 1.825 ;
      RECT 82.145 7.055 82.315 7.225 ;
      RECT 82.145 7.795 82.315 7.965 ;
      RECT 81.77 2.395 81.94 2.565 ;
      RECT 81.77 6.315 81.94 6.485 ;
      RECT 81.525 0.105 81.695 0.275 ;
      RECT 81.525 8.605 81.695 8.775 ;
      RECT 80.845 0.105 81.015 0.275 ;
      RECT 80.845 8.605 81.015 8.775 ;
      RECT 80.775 2.765 80.945 2.935 ;
      RECT 80.775 5.945 80.945 6.115 ;
      RECT 79.08 1.625 79.25 1.795 ;
      RECT 79.08 4.345 79.25 4.515 ;
      RECT 79.08 7.065 79.25 7.235 ;
      RECT 78.62 1.625 78.79 1.795 ;
      RECT 78.62 4.345 78.79 4.515 ;
      RECT 78.62 7.065 78.79 7.235 ;
      RECT 78.58 3.835 78.75 4.005 ;
      RECT 78.58 5.875 78.75 6.045 ;
      RECT 78.24 2.815 78.41 2.985 ;
      RECT 78.16 1.625 78.33 1.795 ;
      RECT 78.16 4.345 78.33 4.515 ;
      RECT 78.16 7.065 78.33 7.235 ;
      RECT 77.9 6.555 78.07 6.725 ;
      RECT 77.73 5.875 77.9 6.045 ;
      RECT 77.7 1.625 77.87 1.795 ;
      RECT 77.7 4.345 77.87 4.515 ;
      RECT 77.7 7.065 77.87 7.235 ;
      RECT 77.24 1.625 77.41 1.795 ;
      RECT 77.24 4.345 77.41 4.515 ;
      RECT 77.24 7.065 77.41 7.235 ;
      RECT 77.22 5.875 77.39 6.045 ;
      RECT 76.78 1.625 76.95 1.795 ;
      RECT 76.78 4.345 76.95 4.515 ;
      RECT 76.78 7.065 76.95 7.235 ;
      RECT 76.54 3.155 76.71 3.325 ;
      RECT 76.54 6.555 76.71 6.725 ;
      RECT 76.32 1.625 76.49 1.795 ;
      RECT 76.32 4.345 76.49 4.515 ;
      RECT 76.32 7.065 76.49 7.235 ;
      RECT 75.86 1.625 76.03 1.795 ;
      RECT 75.86 2.815 76.03 2.985 ;
      RECT 75.86 4.345 76.03 4.515 ;
      RECT 75.86 7.065 76.03 7.235 ;
      RECT 75.85 5.875 76.02 6.045 ;
      RECT 75.4 1.625 75.57 1.795 ;
      RECT 75.4 4.345 75.57 4.515 ;
      RECT 75.4 4.855 75.57 5.025 ;
      RECT 75.4 7.065 75.57 7.235 ;
      RECT 75.38 2.305 75.55 2.475 ;
      RECT 75.01 2.82 75.18 2.99 ;
      RECT 74.94 1.625 75.11 1.795 ;
      RECT 74.94 4.345 75.11 4.515 ;
      RECT 74.94 7.065 75.11 7.235 ;
      RECT 74.5 2.82 74.67 2.99 ;
      RECT 74.5 3.835 74.67 4.005 ;
      RECT 74.5 5.875 74.67 6.045 ;
      RECT 74.48 1.625 74.65 1.795 ;
      RECT 74.48 4.345 74.65 4.515 ;
      RECT 74.48 7.065 74.65 7.235 ;
      RECT 74.16 6.555 74.33 6.725 ;
      RECT 74.02 1.625 74.19 1.795 ;
      RECT 74.02 4.345 74.19 4.515 ;
      RECT 74.02 7.065 74.19 7.235 ;
      RECT 73.56 1.625 73.73 1.795 ;
      RECT 73.56 4.345 73.73 4.515 ;
      RECT 73.56 7.065 73.73 7.235 ;
      RECT 73.14 2.815 73.31 2.985 ;
      RECT 73.14 4.855 73.31 5.025 ;
      RECT 73.1 1.625 73.27 1.795 ;
      RECT 73.1 4.345 73.27 4.515 ;
      RECT 73.1 7.065 73.27 7.235 ;
      RECT 72.64 1.625 72.81 1.795 ;
      RECT 72.64 4.345 72.81 4.515 ;
      RECT 72.64 7.065 72.81 7.235 ;
      RECT 72.63 3.495 72.8 3.665 ;
      RECT 72.18 1.625 72.35 1.795 ;
      RECT 72.18 4.345 72.35 4.515 ;
      RECT 72.18 7.065 72.35 7.235 ;
      RECT 72.12 5.875 72.29 6.045 ;
      RECT 71.2 4.545 71.37 4.715 ;
      RECT 71.2 8.605 71.37 8.775 ;
      RECT 70.89 6.685 71.06 6.855 ;
      RECT 70.52 8.605 70.69 8.775 ;
      RECT 70.46 7.055 70.63 7.225 ;
      RECT 70.46 7.795 70.63 7.965 ;
      RECT 70.085 6.315 70.255 6.485 ;
      RECT 69.84 8.605 70.01 8.775 ;
      RECT 69.16 8.605 69.33 8.775 ;
      RECT 69.09 5.945 69.26 6.115 ;
      RECT 67.71 0.915 67.88 1.085 ;
      RECT 67.71 2.395 67.88 2.565 ;
      RECT 67.71 6.315 67.88 6.485 ;
      RECT 67.71 7.795 67.88 7.965 ;
      RECT 67.36 0.105 67.53 0.275 ;
      RECT 67.36 4.165 67.53 4.335 ;
      RECT 67.36 4.545 67.53 4.715 ;
      RECT 67.36 8.605 67.53 8.775 ;
      RECT 67.34 2.765 67.51 2.935 ;
      RECT 67.34 5.945 67.51 6.115 ;
      RECT 66.72 0.915 66.89 1.085 ;
      RECT 66.72 2.395 66.89 2.565 ;
      RECT 66.72 6.315 66.89 6.485 ;
      RECT 66.72 7.795 66.89 7.965 ;
      RECT 66.37 0.105 66.54 0.275 ;
      RECT 66.37 4.165 66.54 4.335 ;
      RECT 66.37 4.545 66.54 4.715 ;
      RECT 66.37 8.605 66.54 8.775 ;
      RECT 66.35 2.765 66.52 2.935 ;
      RECT 66.35 5.945 66.52 6.115 ;
      RECT 65.665 0.105 65.835 0.275 ;
      RECT 65.665 4.165 65.835 4.335 ;
      RECT 65.665 4.545 65.835 4.715 ;
      RECT 65.665 8.605 65.835 8.775 ;
      RECT 65.355 2.025 65.525 2.195 ;
      RECT 65.355 6.685 65.525 6.855 ;
      RECT 64.985 0.105 65.155 0.275 ;
      RECT 64.985 8.605 65.155 8.775 ;
      RECT 64.925 0.915 65.095 1.085 ;
      RECT 64.925 1.655 65.095 1.825 ;
      RECT 64.925 7.055 65.095 7.225 ;
      RECT 64.925 7.795 65.095 7.965 ;
      RECT 64.55 2.395 64.72 2.565 ;
      RECT 64.55 6.315 64.72 6.485 ;
      RECT 64.305 0.105 64.475 0.275 ;
      RECT 64.305 8.605 64.475 8.775 ;
      RECT 63.625 0.105 63.795 0.275 ;
      RECT 63.625 8.605 63.795 8.775 ;
      RECT 63.555 2.765 63.725 2.935 ;
      RECT 63.555 5.945 63.725 6.115 ;
      RECT 61.86 1.625 62.03 1.795 ;
      RECT 61.86 4.345 62.03 4.515 ;
      RECT 61.86 7.065 62.03 7.235 ;
      RECT 61.4 1.625 61.57 1.795 ;
      RECT 61.4 4.345 61.57 4.515 ;
      RECT 61.4 7.065 61.57 7.235 ;
      RECT 61.36 3.835 61.53 4.005 ;
      RECT 61.36 5.875 61.53 6.045 ;
      RECT 61.02 2.815 61.19 2.985 ;
      RECT 60.94 1.625 61.11 1.795 ;
      RECT 60.94 4.345 61.11 4.515 ;
      RECT 60.94 7.065 61.11 7.235 ;
      RECT 60.68 6.555 60.85 6.725 ;
      RECT 60.51 5.875 60.68 6.045 ;
      RECT 60.48 1.625 60.65 1.795 ;
      RECT 60.48 4.345 60.65 4.515 ;
      RECT 60.48 7.065 60.65 7.235 ;
      RECT 60.02 1.625 60.19 1.795 ;
      RECT 60.02 4.345 60.19 4.515 ;
      RECT 60.02 7.065 60.19 7.235 ;
      RECT 60 5.875 60.17 6.045 ;
      RECT 59.56 1.625 59.73 1.795 ;
      RECT 59.56 4.345 59.73 4.515 ;
      RECT 59.56 7.065 59.73 7.235 ;
      RECT 59.32 3.155 59.49 3.325 ;
      RECT 59.32 6.555 59.49 6.725 ;
      RECT 59.1 1.625 59.27 1.795 ;
      RECT 59.1 4.345 59.27 4.515 ;
      RECT 59.1 7.065 59.27 7.235 ;
      RECT 58.64 1.625 58.81 1.795 ;
      RECT 58.64 2.815 58.81 2.985 ;
      RECT 58.64 4.345 58.81 4.515 ;
      RECT 58.64 7.065 58.81 7.235 ;
      RECT 58.63 5.875 58.8 6.045 ;
      RECT 58.18 1.625 58.35 1.795 ;
      RECT 58.18 4.345 58.35 4.515 ;
      RECT 58.18 4.855 58.35 5.025 ;
      RECT 58.18 7.065 58.35 7.235 ;
      RECT 58.16 2.305 58.33 2.475 ;
      RECT 57.79 2.82 57.96 2.99 ;
      RECT 57.72 1.625 57.89 1.795 ;
      RECT 57.72 4.345 57.89 4.515 ;
      RECT 57.72 7.065 57.89 7.235 ;
      RECT 57.28 2.82 57.45 2.99 ;
      RECT 57.28 3.835 57.45 4.005 ;
      RECT 57.28 5.875 57.45 6.045 ;
      RECT 57.26 1.625 57.43 1.795 ;
      RECT 57.26 4.345 57.43 4.515 ;
      RECT 57.26 7.065 57.43 7.235 ;
      RECT 56.94 6.555 57.11 6.725 ;
      RECT 56.8 1.625 56.97 1.795 ;
      RECT 56.8 4.345 56.97 4.515 ;
      RECT 56.8 7.065 56.97 7.235 ;
      RECT 56.34 1.625 56.51 1.795 ;
      RECT 56.34 4.345 56.51 4.515 ;
      RECT 56.34 7.065 56.51 7.235 ;
      RECT 55.92 2.815 56.09 2.985 ;
      RECT 55.92 4.855 56.09 5.025 ;
      RECT 55.88 1.625 56.05 1.795 ;
      RECT 55.88 4.345 56.05 4.515 ;
      RECT 55.88 7.065 56.05 7.235 ;
      RECT 55.42 1.625 55.59 1.795 ;
      RECT 55.42 4.345 55.59 4.515 ;
      RECT 55.42 7.065 55.59 7.235 ;
      RECT 55.41 3.495 55.58 3.665 ;
      RECT 54.96 1.625 55.13 1.795 ;
      RECT 54.96 4.345 55.13 4.515 ;
      RECT 54.96 7.065 55.13 7.235 ;
      RECT 54.9 5.875 55.07 6.045 ;
      RECT 53.98 4.545 54.15 4.715 ;
      RECT 53.98 8.605 54.15 8.775 ;
      RECT 53.67 6.685 53.84 6.855 ;
      RECT 53.3 8.605 53.47 8.775 ;
      RECT 53.24 7.055 53.41 7.225 ;
      RECT 53.24 7.795 53.41 7.965 ;
      RECT 52.865 6.315 53.035 6.485 ;
      RECT 52.62 8.605 52.79 8.775 ;
      RECT 51.94 8.605 52.11 8.775 ;
      RECT 51.87 5.945 52.04 6.115 ;
      RECT 50.49 0.915 50.66 1.085 ;
      RECT 50.49 2.395 50.66 2.565 ;
      RECT 50.49 6.315 50.66 6.485 ;
      RECT 50.49 7.795 50.66 7.965 ;
      RECT 50.14 0.105 50.31 0.275 ;
      RECT 50.14 4.165 50.31 4.335 ;
      RECT 50.14 4.545 50.31 4.715 ;
      RECT 50.14 8.605 50.31 8.775 ;
      RECT 50.12 2.765 50.29 2.935 ;
      RECT 50.12 5.945 50.29 6.115 ;
      RECT 49.5 0.915 49.67 1.085 ;
      RECT 49.5 2.395 49.67 2.565 ;
      RECT 49.5 6.315 49.67 6.485 ;
      RECT 49.5 7.795 49.67 7.965 ;
      RECT 49.15 0.105 49.32 0.275 ;
      RECT 49.15 4.165 49.32 4.335 ;
      RECT 49.15 4.545 49.32 4.715 ;
      RECT 49.15 8.605 49.32 8.775 ;
      RECT 49.13 2.765 49.3 2.935 ;
      RECT 49.13 5.945 49.3 6.115 ;
      RECT 48.445 0.105 48.615 0.275 ;
      RECT 48.445 4.165 48.615 4.335 ;
      RECT 48.445 4.545 48.615 4.715 ;
      RECT 48.445 8.605 48.615 8.775 ;
      RECT 48.135 2.025 48.305 2.195 ;
      RECT 48.135 6.685 48.305 6.855 ;
      RECT 47.765 0.105 47.935 0.275 ;
      RECT 47.765 8.605 47.935 8.775 ;
      RECT 47.705 0.915 47.875 1.085 ;
      RECT 47.705 1.655 47.875 1.825 ;
      RECT 47.705 7.055 47.875 7.225 ;
      RECT 47.705 7.795 47.875 7.965 ;
      RECT 47.33 2.395 47.5 2.565 ;
      RECT 47.33 6.315 47.5 6.485 ;
      RECT 47.085 0.105 47.255 0.275 ;
      RECT 47.085 8.605 47.255 8.775 ;
      RECT 46.405 0.105 46.575 0.275 ;
      RECT 46.405 8.605 46.575 8.775 ;
      RECT 46.335 2.765 46.505 2.935 ;
      RECT 46.335 5.945 46.505 6.115 ;
      RECT 44.64 1.625 44.81 1.795 ;
      RECT 44.64 4.345 44.81 4.515 ;
      RECT 44.64 7.065 44.81 7.235 ;
      RECT 44.18 1.625 44.35 1.795 ;
      RECT 44.18 4.345 44.35 4.515 ;
      RECT 44.18 7.065 44.35 7.235 ;
      RECT 44.14 3.835 44.31 4.005 ;
      RECT 44.14 5.875 44.31 6.045 ;
      RECT 43.8 2.815 43.97 2.985 ;
      RECT 43.72 1.625 43.89 1.795 ;
      RECT 43.72 4.345 43.89 4.515 ;
      RECT 43.72 7.065 43.89 7.235 ;
      RECT 43.46 6.555 43.63 6.725 ;
      RECT 43.29 5.875 43.46 6.045 ;
      RECT 43.26 1.625 43.43 1.795 ;
      RECT 43.26 4.345 43.43 4.515 ;
      RECT 43.26 7.065 43.43 7.235 ;
      RECT 42.8 1.625 42.97 1.795 ;
      RECT 42.8 4.345 42.97 4.515 ;
      RECT 42.8 7.065 42.97 7.235 ;
      RECT 42.78 5.875 42.95 6.045 ;
      RECT 42.34 1.625 42.51 1.795 ;
      RECT 42.34 4.345 42.51 4.515 ;
      RECT 42.34 7.065 42.51 7.235 ;
      RECT 42.1 3.155 42.27 3.325 ;
      RECT 42.1 6.555 42.27 6.725 ;
      RECT 41.88 1.625 42.05 1.795 ;
      RECT 41.88 4.345 42.05 4.515 ;
      RECT 41.88 7.065 42.05 7.235 ;
      RECT 41.42 1.625 41.59 1.795 ;
      RECT 41.42 2.815 41.59 2.985 ;
      RECT 41.42 4.345 41.59 4.515 ;
      RECT 41.42 7.065 41.59 7.235 ;
      RECT 41.41 5.875 41.58 6.045 ;
      RECT 40.96 1.625 41.13 1.795 ;
      RECT 40.96 4.345 41.13 4.515 ;
      RECT 40.96 4.855 41.13 5.025 ;
      RECT 40.96 7.065 41.13 7.235 ;
      RECT 40.94 2.305 41.11 2.475 ;
      RECT 40.57 2.82 40.74 2.99 ;
      RECT 40.5 1.625 40.67 1.795 ;
      RECT 40.5 4.345 40.67 4.515 ;
      RECT 40.5 7.065 40.67 7.235 ;
      RECT 40.06 2.82 40.23 2.99 ;
      RECT 40.06 3.835 40.23 4.005 ;
      RECT 40.06 5.875 40.23 6.045 ;
      RECT 40.04 1.625 40.21 1.795 ;
      RECT 40.04 4.345 40.21 4.515 ;
      RECT 40.04 7.065 40.21 7.235 ;
      RECT 39.72 6.555 39.89 6.725 ;
      RECT 39.58 1.625 39.75 1.795 ;
      RECT 39.58 4.345 39.75 4.515 ;
      RECT 39.58 7.065 39.75 7.235 ;
      RECT 39.12 1.625 39.29 1.795 ;
      RECT 39.12 4.345 39.29 4.515 ;
      RECT 39.12 7.065 39.29 7.235 ;
      RECT 38.7 2.815 38.87 2.985 ;
      RECT 38.7 4.855 38.87 5.025 ;
      RECT 38.66 1.625 38.83 1.795 ;
      RECT 38.66 4.345 38.83 4.515 ;
      RECT 38.66 7.065 38.83 7.235 ;
      RECT 38.2 1.625 38.37 1.795 ;
      RECT 38.2 4.345 38.37 4.515 ;
      RECT 38.2 7.065 38.37 7.235 ;
      RECT 38.19 3.495 38.36 3.665 ;
      RECT 37.74 1.625 37.91 1.795 ;
      RECT 37.74 4.345 37.91 4.515 ;
      RECT 37.74 7.065 37.91 7.235 ;
      RECT 37.68 5.875 37.85 6.045 ;
      RECT 36.76 4.545 36.93 4.715 ;
      RECT 36.76 8.605 36.93 8.775 ;
      RECT 36.45 6.685 36.62 6.855 ;
      RECT 36.08 8.605 36.25 8.775 ;
      RECT 36.02 7.055 36.19 7.225 ;
      RECT 36.02 7.795 36.19 7.965 ;
      RECT 35.645 6.315 35.815 6.485 ;
      RECT 35.4 8.605 35.57 8.775 ;
      RECT 34.72 8.605 34.89 8.775 ;
      RECT 34.65 5.945 34.82 6.115 ;
      RECT 33.27 0.915 33.44 1.085 ;
      RECT 33.27 2.395 33.44 2.565 ;
      RECT 33.27 6.315 33.44 6.485 ;
      RECT 33.27 7.795 33.44 7.965 ;
      RECT 32.92 0.105 33.09 0.275 ;
      RECT 32.92 4.165 33.09 4.335 ;
      RECT 32.92 4.545 33.09 4.715 ;
      RECT 32.92 8.605 33.09 8.775 ;
      RECT 32.9 2.765 33.07 2.935 ;
      RECT 32.9 5.945 33.07 6.115 ;
      RECT 32.28 0.915 32.45 1.085 ;
      RECT 32.28 2.395 32.45 2.565 ;
      RECT 32.28 6.315 32.45 6.485 ;
      RECT 32.28 7.795 32.45 7.965 ;
      RECT 31.93 0.105 32.1 0.275 ;
      RECT 31.93 4.165 32.1 4.335 ;
      RECT 31.93 4.545 32.1 4.715 ;
      RECT 31.93 8.605 32.1 8.775 ;
      RECT 31.91 2.765 32.08 2.935 ;
      RECT 31.91 5.945 32.08 6.115 ;
      RECT 31.225 0.105 31.395 0.275 ;
      RECT 31.225 4.165 31.395 4.335 ;
      RECT 31.225 4.545 31.395 4.715 ;
      RECT 31.225 8.605 31.395 8.775 ;
      RECT 30.915 2.025 31.085 2.195 ;
      RECT 30.915 6.685 31.085 6.855 ;
      RECT 30.545 0.105 30.715 0.275 ;
      RECT 30.545 8.605 30.715 8.775 ;
      RECT 30.485 0.915 30.655 1.085 ;
      RECT 30.485 1.655 30.655 1.825 ;
      RECT 30.485 7.055 30.655 7.225 ;
      RECT 30.485 7.795 30.655 7.965 ;
      RECT 30.11 2.395 30.28 2.565 ;
      RECT 30.11 6.315 30.28 6.485 ;
      RECT 29.865 0.105 30.035 0.275 ;
      RECT 29.865 8.605 30.035 8.775 ;
      RECT 29.185 0.105 29.355 0.275 ;
      RECT 29.185 8.605 29.355 8.775 ;
      RECT 29.115 2.765 29.285 2.935 ;
      RECT 29.115 5.945 29.285 6.115 ;
      RECT 27.42 1.625 27.59 1.795 ;
      RECT 27.42 4.345 27.59 4.515 ;
      RECT 27.42 7.065 27.59 7.235 ;
      RECT 26.96 1.625 27.13 1.795 ;
      RECT 26.96 4.345 27.13 4.515 ;
      RECT 26.96 7.065 27.13 7.235 ;
      RECT 26.92 3.835 27.09 4.005 ;
      RECT 26.92 5.875 27.09 6.045 ;
      RECT 26.58 2.815 26.75 2.985 ;
      RECT 26.5 1.625 26.67 1.795 ;
      RECT 26.5 4.345 26.67 4.515 ;
      RECT 26.5 7.065 26.67 7.235 ;
      RECT 26.24 6.555 26.41 6.725 ;
      RECT 26.07 5.875 26.24 6.045 ;
      RECT 26.04 1.625 26.21 1.795 ;
      RECT 26.04 4.345 26.21 4.515 ;
      RECT 26.04 7.065 26.21 7.235 ;
      RECT 25.58 1.625 25.75 1.795 ;
      RECT 25.58 4.345 25.75 4.515 ;
      RECT 25.58 7.065 25.75 7.235 ;
      RECT 25.56 5.875 25.73 6.045 ;
      RECT 25.12 1.625 25.29 1.795 ;
      RECT 25.12 4.345 25.29 4.515 ;
      RECT 25.12 7.065 25.29 7.235 ;
      RECT 24.88 3.155 25.05 3.325 ;
      RECT 24.88 6.555 25.05 6.725 ;
      RECT 24.66 1.625 24.83 1.795 ;
      RECT 24.66 4.345 24.83 4.515 ;
      RECT 24.66 7.065 24.83 7.235 ;
      RECT 24.2 1.625 24.37 1.795 ;
      RECT 24.2 2.815 24.37 2.985 ;
      RECT 24.2 4.345 24.37 4.515 ;
      RECT 24.2 7.065 24.37 7.235 ;
      RECT 24.19 5.875 24.36 6.045 ;
      RECT 23.74 1.625 23.91 1.795 ;
      RECT 23.74 4.345 23.91 4.515 ;
      RECT 23.74 4.855 23.91 5.025 ;
      RECT 23.74 7.065 23.91 7.235 ;
      RECT 23.72 2.305 23.89 2.475 ;
      RECT 23.35 2.82 23.52 2.99 ;
      RECT 23.28 1.625 23.45 1.795 ;
      RECT 23.28 4.345 23.45 4.515 ;
      RECT 23.28 7.065 23.45 7.235 ;
      RECT 22.84 2.82 23.01 2.99 ;
      RECT 22.84 3.835 23.01 4.005 ;
      RECT 22.84 5.875 23.01 6.045 ;
      RECT 22.82 1.625 22.99 1.795 ;
      RECT 22.82 4.345 22.99 4.515 ;
      RECT 22.82 7.065 22.99 7.235 ;
      RECT 22.5 6.555 22.67 6.725 ;
      RECT 22.36 1.625 22.53 1.795 ;
      RECT 22.36 4.345 22.53 4.515 ;
      RECT 22.36 7.065 22.53 7.235 ;
      RECT 21.9 1.625 22.07 1.795 ;
      RECT 21.9 4.345 22.07 4.515 ;
      RECT 21.9 7.065 22.07 7.235 ;
      RECT 21.48 2.815 21.65 2.985 ;
      RECT 21.48 4.855 21.65 5.025 ;
      RECT 21.44 1.625 21.61 1.795 ;
      RECT 21.44 4.345 21.61 4.515 ;
      RECT 21.44 7.065 21.61 7.235 ;
      RECT 20.98 1.625 21.15 1.795 ;
      RECT 20.98 4.345 21.15 4.515 ;
      RECT 20.98 7.065 21.15 7.235 ;
      RECT 20.97 3.495 21.14 3.665 ;
      RECT 20.52 1.625 20.69 1.795 ;
      RECT 20.52 4.345 20.69 4.515 ;
      RECT 20.52 7.065 20.69 7.235 ;
      RECT 20.46 5.875 20.63 6.045 ;
      RECT 19.54 4.545 19.71 4.715 ;
      RECT 19.54 8.605 19.71 8.775 ;
      RECT 19.23 6.685 19.4 6.855 ;
      RECT 18.86 8.605 19.03 8.775 ;
      RECT 18.8 7.055 18.97 7.225 ;
      RECT 18.8 7.795 18.97 7.965 ;
      RECT 18.425 6.315 18.595 6.485 ;
      RECT 18.18 8.605 18.35 8.775 ;
      RECT 17.5 8.605 17.67 8.775 ;
      RECT 17.43 5.945 17.6 6.115 ;
      RECT 16.05 0.915 16.22 1.085 ;
      RECT 16.05 2.395 16.22 2.565 ;
      RECT 16.05 6.315 16.22 6.485 ;
      RECT 16.05 7.795 16.22 7.965 ;
      RECT 15.7 0.105 15.87 0.275 ;
      RECT 15.7 4.165 15.87 4.335 ;
      RECT 15.7 4.545 15.87 4.715 ;
      RECT 15.7 8.605 15.87 8.775 ;
      RECT 15.68 2.765 15.85 2.935 ;
      RECT 15.68 5.945 15.85 6.115 ;
      RECT 15.06 0.915 15.23 1.085 ;
      RECT 15.06 2.395 15.23 2.565 ;
      RECT 15.06 6.315 15.23 6.485 ;
      RECT 15.06 7.795 15.23 7.965 ;
      RECT 14.71 0.105 14.88 0.275 ;
      RECT 14.71 4.165 14.88 4.335 ;
      RECT 14.71 4.545 14.88 4.715 ;
      RECT 14.71 8.605 14.88 8.775 ;
      RECT 14.69 2.765 14.86 2.935 ;
      RECT 14.69 5.945 14.86 6.115 ;
      RECT 14.005 0.105 14.175 0.275 ;
      RECT 14.005 4.165 14.175 4.335 ;
      RECT 14.005 4.545 14.175 4.715 ;
      RECT 14.005 8.605 14.175 8.775 ;
      RECT 13.695 2.025 13.865 2.195 ;
      RECT 13.695 6.685 13.865 6.855 ;
      RECT 13.325 0.105 13.495 0.275 ;
      RECT 13.325 8.605 13.495 8.775 ;
      RECT 13.265 0.915 13.435 1.085 ;
      RECT 13.265 1.655 13.435 1.825 ;
      RECT 13.265 7.055 13.435 7.225 ;
      RECT 13.265 7.795 13.435 7.965 ;
      RECT 12.89 2.395 13.06 2.565 ;
      RECT 12.89 6.315 13.06 6.485 ;
      RECT 12.645 0.105 12.815 0.275 ;
      RECT 12.645 8.605 12.815 8.775 ;
      RECT 11.965 0.105 12.135 0.275 ;
      RECT 11.965 8.605 12.135 8.775 ;
      RECT 11.895 2.765 12.065 2.935 ;
      RECT 11.895 5.945 12.065 6.115 ;
      RECT 10.2 1.625 10.37 1.795 ;
      RECT 10.2 4.345 10.37 4.515 ;
      RECT 10.2 7.065 10.37 7.235 ;
      RECT 9.74 1.625 9.91 1.795 ;
      RECT 9.74 4.345 9.91 4.515 ;
      RECT 9.74 7.065 9.91 7.235 ;
      RECT 9.7 3.835 9.87 4.005 ;
      RECT 9.7 5.875 9.87 6.045 ;
      RECT 9.36 2.815 9.53 2.985 ;
      RECT 9.28 1.625 9.45 1.795 ;
      RECT 9.28 4.345 9.45 4.515 ;
      RECT 9.28 7.065 9.45 7.235 ;
      RECT 9.02 6.555 9.19 6.725 ;
      RECT 8.85 5.875 9.02 6.045 ;
      RECT 8.82 1.625 8.99 1.795 ;
      RECT 8.82 4.345 8.99 4.515 ;
      RECT 8.82 7.065 8.99 7.235 ;
      RECT 8.36 1.625 8.53 1.795 ;
      RECT 8.36 4.345 8.53 4.515 ;
      RECT 8.36 7.065 8.53 7.235 ;
      RECT 8.34 5.875 8.51 6.045 ;
      RECT 7.9 1.625 8.07 1.795 ;
      RECT 7.9 4.345 8.07 4.515 ;
      RECT 7.9 7.065 8.07 7.235 ;
      RECT 7.66 3.155 7.83 3.325 ;
      RECT 7.66 6.555 7.83 6.725 ;
      RECT 7.44 1.625 7.61 1.795 ;
      RECT 7.44 4.345 7.61 4.515 ;
      RECT 7.44 7.065 7.61 7.235 ;
      RECT 6.98 1.625 7.15 1.795 ;
      RECT 6.98 2.815 7.15 2.985 ;
      RECT 6.98 4.345 7.15 4.515 ;
      RECT 6.98 7.065 7.15 7.235 ;
      RECT 6.97 5.875 7.14 6.045 ;
      RECT 6.52 1.625 6.69 1.795 ;
      RECT 6.52 4.345 6.69 4.515 ;
      RECT 6.52 4.855 6.69 5.025 ;
      RECT 6.52 7.065 6.69 7.235 ;
      RECT 6.5 2.305 6.67 2.475 ;
      RECT 6.13 2.82 6.3 2.99 ;
      RECT 6.06 1.625 6.23 1.795 ;
      RECT 6.06 4.345 6.23 4.515 ;
      RECT 6.06 7.065 6.23 7.235 ;
      RECT 5.62 2.82 5.79 2.99 ;
      RECT 5.62 3.835 5.79 4.005 ;
      RECT 5.62 5.875 5.79 6.045 ;
      RECT 5.6 1.625 5.77 1.795 ;
      RECT 5.6 4.345 5.77 4.515 ;
      RECT 5.6 7.065 5.77 7.235 ;
      RECT 5.28 6.555 5.45 6.725 ;
      RECT 5.14 1.625 5.31 1.795 ;
      RECT 5.14 4.345 5.31 4.515 ;
      RECT 5.14 7.065 5.31 7.235 ;
      RECT 4.68 1.625 4.85 1.795 ;
      RECT 4.68 4.345 4.85 4.515 ;
      RECT 4.68 7.065 4.85 7.235 ;
      RECT 4.26 2.815 4.43 2.985 ;
      RECT 4.26 4.855 4.43 5.025 ;
      RECT 4.22 1.625 4.39 1.795 ;
      RECT 4.22 4.345 4.39 4.515 ;
      RECT 4.22 7.065 4.39 7.235 ;
      RECT 3.76 1.625 3.93 1.795 ;
      RECT 3.76 4.345 3.93 4.515 ;
      RECT 3.76 7.065 3.93 7.235 ;
      RECT 3.75 3.495 3.92 3.665 ;
      RECT 3.3 1.625 3.47 1.795 ;
      RECT 3.3 4.345 3.47 4.515 ;
      RECT 3.3 7.065 3.47 7.235 ;
      RECT 3.24 5.875 3.41 6.045 ;
      RECT 2.32 4.545 2.49 4.715 ;
      RECT 2.32 8.605 2.49 8.775 ;
      RECT 2.01 6.685 2.18 6.855 ;
      RECT 1.64 8.605 1.81 8.775 ;
      RECT 1.58 7.055 1.75 7.225 ;
      RECT 1.58 7.795 1.75 7.965 ;
      RECT 1.205 6.315 1.375 6.485 ;
      RECT 0.96 8.605 1.13 8.775 ;
      RECT 0.28 8.605 0.45 8.775 ;
      RECT 0.21 5.945 0.38 6.115 ;
      RECT -1.09 4.545 -0.92 4.715 ;
      RECT -1.09 8.605 -0.92 8.775 ;
      RECT -1.4 6.685 -1.23 6.855 ;
      RECT -1.77 8.605 -1.6 8.775 ;
      RECT -1.83 7.055 -1.66 7.225 ;
      RECT -1.83 7.795 -1.66 7.965 ;
      RECT -2.205 6.315 -2.035 6.485 ;
      RECT -2.45 8.605 -2.28 8.775 ;
      RECT -3.13 8.605 -2.96 8.775 ;
      RECT -3.2 5.945 -3.03 6.115 ;
    LAYER li ;
      RECT 76.26 0 76.55 2.63 ;
      RECT 59.04 0 59.33 2.63 ;
      RECT 41.82 0 42.11 2.63 ;
      RECT 24.6 0 24.89 2.63 ;
      RECT 7.38 0 7.67 2.63 ;
      RECT 73.06 0 73.29 2.615 ;
      RECT 72.18 0 72.39 2.615 ;
      RECT 55.84 0 56.07 2.615 ;
      RECT 54.96 0 55.17 2.615 ;
      RECT 38.62 0 38.85 2.615 ;
      RECT 37.74 0 37.95 2.615 ;
      RECT 21.4 0 21.63 2.615 ;
      RECT 20.52 0 20.73 2.615 ;
      RECT 4.18 0 4.41 2.615 ;
      RECT 3.3 0 3.51 2.615 ;
      RECT 75.81 0 76.08 2.605 ;
      RECT 74.9 0 75.14 2.605 ;
      RECT 74.45 0 74.69 2.605 ;
      RECT 73.51 0 73.78 2.605 ;
      RECT 58.59 0 58.86 2.605 ;
      RECT 57.68 0 57.92 2.605 ;
      RECT 57.23 0 57.47 2.605 ;
      RECT 56.29 0 56.56 2.605 ;
      RECT 41.37 0 41.64 2.605 ;
      RECT 40.46 0 40.7 2.605 ;
      RECT 40.01 0 40.25 2.605 ;
      RECT 39.07 0 39.34 2.605 ;
      RECT 24.15 0 24.42 2.605 ;
      RECT 23.24 0 23.48 2.605 ;
      RECT 22.79 0 23.03 2.605 ;
      RECT 21.85 0 22.12 2.605 ;
      RECT 6.93 0 7.2 2.605 ;
      RECT 6.02 0 6.26 2.605 ;
      RECT 5.57 0 5.81 2.605 ;
      RECT 4.63 0 4.9 2.605 ;
      RECT 78.93 0 79.26 2.185 ;
      RECT 78.09 0 78.42 2.185 ;
      RECT 61.71 0 62.04 2.185 ;
      RECT 60.87 0 61.2 2.185 ;
      RECT 44.49 0 44.82 2.185 ;
      RECT 43.65 0 43.98 2.185 ;
      RECT 27.27 0 27.6 2.185 ;
      RECT 26.43 0 26.76 2.185 ;
      RECT 10.05 0 10.38 2.185 ;
      RECT 9.21 0 9.54 2.185 ;
      RECT 72.035 0 79.69 1.795 ;
      RECT 54.815 0 62.47 1.795 ;
      RECT 37.595 0 45.25 1.795 ;
      RECT 20.375 0 28.03 1.795 ;
      RECT 3.155 0 10.81 1.795 ;
      RECT 72.03 0 79.69 1.635 ;
      RECT 54.81 0 62.47 1.635 ;
      RECT 37.59 0 45.25 1.635 ;
      RECT 20.37 0 28.03 1.635 ;
      RECT 3.15 0 10.81 1.635 ;
      RECT 84.5 0 84.67 0.935 ;
      RECT 83.51 0 83.68 0.935 ;
      RECT 80.765 0 80.935 0.935 ;
      RECT 67.28 0 67.45 0.935 ;
      RECT 66.29 0 66.46 0.935 ;
      RECT 63.545 0 63.715 0.935 ;
      RECT 50.06 0 50.23 0.935 ;
      RECT 49.07 0 49.24 0.935 ;
      RECT 46.325 0 46.495 0.935 ;
      RECT 32.84 0 33.01 0.935 ;
      RECT 31.85 0 32.02 0.935 ;
      RECT 29.105 0 29.275 0.935 ;
      RECT 15.62 0 15.79 0.935 ;
      RECT 14.63 0 14.8 0.935 ;
      RECT 11.885 0 12.055 0.935 ;
      RECT -3.385 0 85.47 0.305 ;
      RECT -1.4 4.13 -1.23 8.305 ;
      RECT 78.57 4.345 78.85 5.655 ;
      RECT 77.64 4.345 77.9 5.655 ;
      RECT 77.19 4.345 77.47 5.655 ;
      RECT 76.26 4.345 76.52 5.655 ;
      RECT 75.83 4.345 76.09 5.655 ;
      RECT 74.88 4.345 75.16 5.655 ;
      RECT 73.53 3.205 73.79 5.655 ;
      RECT 72.58 4.345 72.86 5.655 ;
      RECT 61.35 4.345 61.63 5.655 ;
      RECT 60.42 4.345 60.68 5.655 ;
      RECT 59.97 4.345 60.25 5.655 ;
      RECT 59.04 4.345 59.3 5.655 ;
      RECT 58.61 4.345 58.87 5.655 ;
      RECT 57.66 4.345 57.94 5.655 ;
      RECT 56.31 3.205 56.57 5.655 ;
      RECT 55.36 4.345 55.64 5.655 ;
      RECT 44.13 4.345 44.41 5.655 ;
      RECT 43.2 4.345 43.46 5.655 ;
      RECT 42.75 4.345 43.03 5.655 ;
      RECT 41.82 4.345 42.08 5.655 ;
      RECT 41.39 4.345 41.65 5.655 ;
      RECT 40.44 4.345 40.72 5.655 ;
      RECT 39.09 3.205 39.35 5.655 ;
      RECT 38.14 4.345 38.42 5.655 ;
      RECT 26.91 4.345 27.19 5.655 ;
      RECT 25.98 4.345 26.24 5.655 ;
      RECT 25.53 4.345 25.81 5.655 ;
      RECT 24.6 4.345 24.86 5.655 ;
      RECT 24.17 4.345 24.43 5.655 ;
      RECT 23.22 4.345 23.5 5.655 ;
      RECT 21.87 3.205 22.13 5.655 ;
      RECT 20.92 4.345 21.2 5.655 ;
      RECT 9.69 4.345 9.97 5.655 ;
      RECT 8.76 4.345 9.02 5.655 ;
      RECT 8.31 4.345 8.59 5.655 ;
      RECT 7.38 4.345 7.64 5.655 ;
      RECT 6.95 4.345 7.21 5.655 ;
      RECT 6 4.345 6.28 5.655 ;
      RECT 4.65 3.205 4.91 5.655 ;
      RECT 3.7 4.345 3.98 5.655 ;
      RECT 84.5 3.405 84.67 5.475 ;
      RECT 83.51 3.405 83.68 5.475 ;
      RECT 80.765 3.405 80.935 5.475 ;
      RECT 69.08 4.13 69.25 5.475 ;
      RECT 67.28 3.405 67.45 5.475 ;
      RECT 66.29 3.405 66.46 5.475 ;
      RECT 63.545 3.405 63.715 5.475 ;
      RECT 51.86 4.13 52.03 5.475 ;
      RECT 50.06 3.405 50.23 5.475 ;
      RECT 49.07 3.405 49.24 5.475 ;
      RECT 46.325 3.405 46.495 5.475 ;
      RECT 34.64 4.13 34.81 5.475 ;
      RECT 32.84 3.405 33.01 5.475 ;
      RECT 31.85 3.405 32.02 5.475 ;
      RECT 29.105 3.405 29.275 5.475 ;
      RECT 17.42 4.13 17.59 5.475 ;
      RECT 15.62 3.405 15.79 5.475 ;
      RECT 14.63 3.405 14.8 5.475 ;
      RECT 11.885 3.405 12.055 5.475 ;
      RECT 0.2 4.13 0.37 5.475 ;
      RECT -3.21 4.13 -3.04 5.475 ;
      RECT 79.485 4.135 85.47 4.745 ;
      RECT 68.905 4.13 71.655 4.745 ;
      RECT 62.265 4.135 68.25 4.745 ;
      RECT 51.685 4.13 54.435 4.745 ;
      RECT 45.045 4.135 51.03 4.745 ;
      RECT 34.465 4.13 37.215 4.745 ;
      RECT 27.825 4.135 33.81 4.745 ;
      RECT 17.245 4.13 19.995 4.745 ;
      RECT 10.605 4.135 16.59 4.745 ;
      RECT 0.025 4.13 2.775 4.745 ;
      RECT -3.385 4.13 -0.635 4.745 ;
      RECT 62.265 4.345 72.41 4.74 ;
      RECT 45.045 4.345 55.19 4.74 ;
      RECT 27.825 4.345 37.97 4.74 ;
      RECT 10.605 4.345 20.75 4.74 ;
      RECT -3.385 4.345 3.53 4.74 ;
      RECT -3.385 4.345 85.47 4.515 ;
      RECT 79.48 4.135 85.47 4.515 ;
      RECT 78.17 3.495 78.34 4.515 ;
      RECT 77.33 3.835 77.5 4.515 ;
      RECT 75.75 3.205 76.08 4.515 ;
      RECT 73.51 3.205 73.84 4.515 ;
      RECT 73.06 3.205 73.29 4.515 ;
      RECT 62.26 4.135 72.39 4.515 ;
      RECT 72.18 3.205 72.39 4.74 ;
      RECT 60.95 3.495 61.12 4.515 ;
      RECT 60.11 3.835 60.28 4.515 ;
      RECT 58.53 3.205 58.86 4.515 ;
      RECT 56.29 3.205 56.62 4.515 ;
      RECT 55.84 3.205 56.07 4.515 ;
      RECT 45.04 4.135 55.17 4.515 ;
      RECT 54.96 3.205 55.17 4.74 ;
      RECT 43.73 3.495 43.9 4.515 ;
      RECT 42.89 3.835 43.06 4.515 ;
      RECT 41.31 3.205 41.64 4.515 ;
      RECT 39.07 3.205 39.4 4.515 ;
      RECT 38.62 3.205 38.85 4.515 ;
      RECT 27.82 4.135 37.95 4.515 ;
      RECT 37.74 3.205 37.95 4.74 ;
      RECT 26.51 3.495 26.68 4.515 ;
      RECT 25.67 3.835 25.84 4.515 ;
      RECT 24.09 3.205 24.42 4.515 ;
      RECT 21.85 3.205 22.18 4.515 ;
      RECT 21.4 3.205 21.63 4.515 ;
      RECT 10.6 4.135 20.73 4.515 ;
      RECT 20.52 3.205 20.73 4.74 ;
      RECT 9.29 3.495 9.46 4.515 ;
      RECT 8.45 3.835 8.62 4.515 ;
      RECT 6.87 3.205 7.2 4.515 ;
      RECT 4.63 3.205 4.96 4.515 ;
      RECT 4.18 3.205 4.41 4.515 ;
      RECT -3.385 4.13 3.51 4.74 ;
      RECT 3.3 3.205 3.51 4.74 ;
      RECT 68.245 4.13 72.39 4.74 ;
      RECT 51.025 4.13 55.17 4.74 ;
      RECT 33.805 4.13 37.95 4.74 ;
      RECT 16.585 4.13 20.73 4.74 ;
      RECT -3.385 8.575 85.47 8.88 ;
      RECT 84.5 7.945 84.67 8.88 ;
      RECT 83.51 7.945 83.68 8.88 ;
      RECT 80.765 7.945 80.935 8.88 ;
      RECT 72.305 7.18 79.505 8.88 ;
      RECT 69.08 7.945 69.25 8.88 ;
      RECT 67.28 7.945 67.45 8.88 ;
      RECT 66.29 7.945 66.46 8.88 ;
      RECT 63.545 7.945 63.715 8.88 ;
      RECT 55.085 7.18 62.285 8.88 ;
      RECT 51.86 7.945 52.03 8.88 ;
      RECT 50.06 7.945 50.23 8.88 ;
      RECT 49.07 7.945 49.24 8.88 ;
      RECT 46.325 7.945 46.495 8.88 ;
      RECT 37.865 7.18 45.065 8.88 ;
      RECT 34.64 7.945 34.81 8.88 ;
      RECT 32.84 7.945 33.01 8.88 ;
      RECT 31.85 7.945 32.02 8.88 ;
      RECT 29.105 7.945 29.275 8.88 ;
      RECT 20.645 7.18 27.845 8.88 ;
      RECT 17.42 7.945 17.59 8.88 ;
      RECT 15.62 7.945 15.79 8.88 ;
      RECT 14.63 7.945 14.8 8.88 ;
      RECT 11.885 7.945 12.055 8.88 ;
      RECT 3.425 7.18 10.625 8.88 ;
      RECT 0.2 7.945 0.37 8.88 ;
      RECT -3.21 7.945 -3.04 8.88 ;
      RECT 72.035 7.065 79.395 7.235 ;
      RECT 54.815 7.065 62.175 7.235 ;
      RECT 37.595 7.065 44.955 7.235 ;
      RECT 20.375 7.065 27.735 7.235 ;
      RECT 3.155 7.065 10.515 7.235 ;
      RECT 78.54 6.265 78.85 8.88 ;
      RECT 77.16 6.265 77.47 8.88 ;
      RECT 74.88 6.265 75.19 8.88 ;
      RECT 74.51 5.875 74.68 8.88 ;
      RECT 72.58 6.265 72.89 8.88 ;
      RECT 61.32 6.265 61.63 8.88 ;
      RECT 59.94 6.265 60.25 8.88 ;
      RECT 57.66 6.265 57.97 8.88 ;
      RECT 57.29 5.875 57.46 8.88 ;
      RECT 55.36 6.265 55.67 8.88 ;
      RECT 44.1 6.265 44.41 8.88 ;
      RECT 42.72 6.265 43.03 8.88 ;
      RECT 40.44 6.265 40.75 8.88 ;
      RECT 40.07 5.875 40.24 8.88 ;
      RECT 38.14 6.265 38.45 8.88 ;
      RECT 26.88 6.265 27.19 8.88 ;
      RECT 25.5 6.265 25.81 8.88 ;
      RECT 23.22 6.265 23.53 8.88 ;
      RECT 22.85 5.875 23.02 8.88 ;
      RECT 20.92 6.265 21.23 8.88 ;
      RECT 9.66 6.265 9.97 8.88 ;
      RECT 8.28 6.265 8.59 8.88 ;
      RECT 6 6.265 6.31 8.88 ;
      RECT 5.63 5.875 5.8 8.88 ;
      RECT 3.7 6.265 4.01 8.88 ;
      RECT 74.89 5.825 75.225 6.095 ;
      RECT 57.67 5.825 58.005 6.095 ;
      RECT 40.45 5.825 40.785 6.095 ;
      RECT 23.23 5.825 23.565 6.095 ;
      RECT 6.01 5.825 6.345 6.095 ;
      RECT 74.5 5.875 75.225 6.045 ;
      RECT 57.28 5.875 58.005 6.045 ;
      RECT 40.06 5.875 40.785 6.045 ;
      RECT 22.84 5.875 23.565 6.045 ;
      RECT 5.62 5.875 6.345 6.045 ;
      RECT 84.56 1.74 84.73 2.935 ;
      RECT 84.56 1.74 85.025 1.91 ;
      RECT 84.56 6.97 85.025 7.14 ;
      RECT 84.56 5.945 84.73 7.14 ;
      RECT 83.57 1.74 83.74 2.935 ;
      RECT 83.57 1.74 84.035 1.91 ;
      RECT 83.57 6.97 84.035 7.14 ;
      RECT 83.57 5.945 83.74 7.14 ;
      RECT 81.715 2.635 81.885 3.865 ;
      RECT 81.77 0.855 81.94 2.805 ;
      RECT 81.715 0.575 81.885 1.025 ;
      RECT 81.715 7.855 81.885 8.305 ;
      RECT 81.77 6.075 81.94 8.025 ;
      RECT 81.715 5.015 81.885 6.245 ;
      RECT 81.195 0.575 81.365 3.865 ;
      RECT 81.195 2.075 81.6 2.405 ;
      RECT 81.195 1.235 81.6 1.565 ;
      RECT 81.195 5.015 81.365 8.305 ;
      RECT 81.195 7.315 81.6 7.645 ;
      RECT 81.195 6.475 81.6 6.805 ;
      RECT 80.775 5.94 80.945 7.22 ;
      RECT 80.765 5.94 80.945 6.18 ;
      RECT 78.93 3.495 79.31 4.175 ;
      RECT 79.14 2.365 79.31 4.175 ;
      RECT 77.06 2.365 77.29 3.035 ;
      RECT 77.06 2.365 79.31 2.535 ;
      RECT 78.59 2.045 78.76 2.535 ;
      RECT 78.58 3.155 78.75 4.005 ;
      RECT 77.665 3.155 78.97 3.325 ;
      RECT 78.725 2.705 78.97 3.325 ;
      RECT 77.665 2.785 77.835 3.325 ;
      RECT 77.46 2.785 77.835 2.955 ;
      RECT 77.64 6.265 78.335 6.895 ;
      RECT 78.165 4.685 78.335 6.895 ;
      RECT 78.07 4.685 78.4 5.665 ;
      RECT 77.67 3.495 78 4.175 ;
      RECT 76.76 3.495 77.16 4.175 ;
      RECT 76.76 3.495 78 3.665 ;
      RECT 76.26 3.075 76.58 4.175 ;
      RECT 76.26 3.075 76.71 3.325 ;
      RECT 76.26 3.075 76.89 3.245 ;
      RECT 76.72 2.025 76.89 3.245 ;
      RECT 76.72 2.025 77.675 2.195 ;
      RECT 76.26 6.265 76.955 6.895 ;
      RECT 76.785 4.685 76.955 6.895 ;
      RECT 76.69 4.685 77.02 5.665 ;
      RECT 76.28 5.825 76.615 6.075 ;
      RECT 75.735 5.825 76.07 6.075 ;
      RECT 75.735 5.875 76.615 6.045 ;
      RECT 75.395 6.265 76.09 6.895 ;
      RECT 75.395 4.685 75.565 6.895 ;
      RECT 75.33 4.685 75.66 5.665 ;
      RECT 74.89 3.205 75.22 4.16 ;
      RECT 74.89 3.205 75.57 3.375 ;
      RECT 75.4 1.965 75.57 3.375 ;
      RECT 75.31 1.965 75.64 2.605 ;
      RECT 74.37 3.205 74.7 4.16 ;
      RECT 74.02 3.205 74.7 3.375 ;
      RECT 74.02 1.965 74.19 3.375 ;
      RECT 73.95 1.965 74.28 2.605 ;
      RECT 74.16 5.875 74.33 6.725 ;
      RECT 73.435 5.825 73.77 6.075 ;
      RECT 73.435 5.875 74.33 6.045 ;
      RECT 73.5 2.785 73.85 3.035 ;
      RECT 72.98 2.785 73.31 3.035 ;
      RECT 72.98 2.815 73.85 2.985 ;
      RECT 73.095 6.265 73.79 6.895 ;
      RECT 73.095 4.685 73.265 6.895 ;
      RECT 73.03 4.685 73.36 5.665 ;
      RECT 72.59 5.825 72.925 6.095 ;
      RECT 72.12 5.875 72.925 6.045 ;
      RECT 72.56 3.195 72.89 4.175 ;
      RECT 72.56 1.965 72.81 4.175 ;
      RECT 72.56 1.965 72.89 2.595 ;
      RECT 70.03 7.855 70.2 8.305 ;
      RECT 70.085 6.075 70.255 8.025 ;
      RECT 70.03 5.015 70.2 6.245 ;
      RECT 69.51 5.015 69.68 8.305 ;
      RECT 69.51 7.315 69.915 7.645 ;
      RECT 69.51 6.475 69.915 6.805 ;
      RECT 67.34 1.74 67.51 2.935 ;
      RECT 67.34 1.74 67.805 1.91 ;
      RECT 67.34 6.97 67.805 7.14 ;
      RECT 67.34 5.945 67.51 7.14 ;
      RECT 66.35 1.74 66.52 2.935 ;
      RECT 66.35 1.74 66.815 1.91 ;
      RECT 66.35 6.97 66.815 7.14 ;
      RECT 66.35 5.945 66.52 7.14 ;
      RECT 64.495 2.635 64.665 3.865 ;
      RECT 64.55 0.855 64.72 2.805 ;
      RECT 64.495 0.575 64.665 1.025 ;
      RECT 64.495 7.855 64.665 8.305 ;
      RECT 64.55 6.075 64.72 8.025 ;
      RECT 64.495 5.015 64.665 6.245 ;
      RECT 63.975 0.575 64.145 3.865 ;
      RECT 63.975 2.075 64.38 2.405 ;
      RECT 63.975 1.235 64.38 1.565 ;
      RECT 63.975 5.015 64.145 8.305 ;
      RECT 63.975 7.315 64.38 7.645 ;
      RECT 63.975 6.475 64.38 6.805 ;
      RECT 63.555 5.94 63.725 7.22 ;
      RECT 63.545 5.94 63.725 6.18 ;
      RECT 61.71 3.495 62.09 4.175 ;
      RECT 61.92 2.365 62.09 4.175 ;
      RECT 59.84 2.365 60.07 3.035 ;
      RECT 59.84 2.365 62.09 2.535 ;
      RECT 61.37 2.045 61.54 2.535 ;
      RECT 61.36 3.155 61.53 4.005 ;
      RECT 60.445 3.155 61.75 3.325 ;
      RECT 61.505 2.705 61.75 3.325 ;
      RECT 60.445 2.785 60.615 3.325 ;
      RECT 60.24 2.785 60.615 2.955 ;
      RECT 60.42 6.265 61.115 6.895 ;
      RECT 60.945 4.685 61.115 6.895 ;
      RECT 60.85 4.685 61.18 5.665 ;
      RECT 60.45 3.495 60.78 4.175 ;
      RECT 59.54 3.495 59.94 4.175 ;
      RECT 59.54 3.495 60.78 3.665 ;
      RECT 59.04 3.075 59.36 4.175 ;
      RECT 59.04 3.075 59.49 3.325 ;
      RECT 59.04 3.075 59.67 3.245 ;
      RECT 59.5 2.025 59.67 3.245 ;
      RECT 59.5 2.025 60.455 2.195 ;
      RECT 59.04 6.265 59.735 6.895 ;
      RECT 59.565 4.685 59.735 6.895 ;
      RECT 59.47 4.685 59.8 5.665 ;
      RECT 59.06 5.825 59.395 6.075 ;
      RECT 58.515 5.825 58.85 6.075 ;
      RECT 58.515 5.875 59.395 6.045 ;
      RECT 58.175 6.265 58.87 6.895 ;
      RECT 58.175 4.685 58.345 6.895 ;
      RECT 58.11 4.685 58.44 5.665 ;
      RECT 57.67 3.205 58 4.16 ;
      RECT 57.67 3.205 58.35 3.375 ;
      RECT 58.18 1.965 58.35 3.375 ;
      RECT 58.09 1.965 58.42 2.605 ;
      RECT 57.15 3.205 57.48 4.16 ;
      RECT 56.8 3.205 57.48 3.375 ;
      RECT 56.8 1.965 56.97 3.375 ;
      RECT 56.73 1.965 57.06 2.605 ;
      RECT 56.94 5.875 57.11 6.725 ;
      RECT 56.215 5.825 56.55 6.075 ;
      RECT 56.215 5.875 57.11 6.045 ;
      RECT 56.28 2.785 56.63 3.035 ;
      RECT 55.76 2.785 56.09 3.035 ;
      RECT 55.76 2.815 56.63 2.985 ;
      RECT 55.875 6.265 56.57 6.895 ;
      RECT 55.875 4.685 56.045 6.895 ;
      RECT 55.81 4.685 56.14 5.665 ;
      RECT 55.37 5.825 55.705 6.095 ;
      RECT 54.9 5.875 55.705 6.045 ;
      RECT 55.34 3.195 55.67 4.175 ;
      RECT 55.34 1.965 55.59 4.175 ;
      RECT 55.34 1.965 55.67 2.595 ;
      RECT 52.81 7.855 52.98 8.305 ;
      RECT 52.865 6.075 53.035 8.025 ;
      RECT 52.81 5.015 52.98 6.245 ;
      RECT 52.29 5.015 52.46 8.305 ;
      RECT 52.29 7.315 52.695 7.645 ;
      RECT 52.29 6.475 52.695 6.805 ;
      RECT 50.12 1.74 50.29 2.935 ;
      RECT 50.12 1.74 50.585 1.91 ;
      RECT 50.12 6.97 50.585 7.14 ;
      RECT 50.12 5.945 50.29 7.14 ;
      RECT 49.13 1.74 49.3 2.935 ;
      RECT 49.13 1.74 49.595 1.91 ;
      RECT 49.13 6.97 49.595 7.14 ;
      RECT 49.13 5.945 49.3 7.14 ;
      RECT 47.275 2.635 47.445 3.865 ;
      RECT 47.33 0.855 47.5 2.805 ;
      RECT 47.275 0.575 47.445 1.025 ;
      RECT 47.275 7.855 47.445 8.305 ;
      RECT 47.33 6.075 47.5 8.025 ;
      RECT 47.275 5.015 47.445 6.245 ;
      RECT 46.755 0.575 46.925 3.865 ;
      RECT 46.755 2.075 47.16 2.405 ;
      RECT 46.755 1.235 47.16 1.565 ;
      RECT 46.755 5.015 46.925 8.305 ;
      RECT 46.755 7.315 47.16 7.645 ;
      RECT 46.755 6.475 47.16 6.805 ;
      RECT 46.335 5.94 46.505 7.22 ;
      RECT 46.325 5.94 46.505 6.18 ;
      RECT 44.49 3.495 44.87 4.175 ;
      RECT 44.7 2.365 44.87 4.175 ;
      RECT 42.62 2.365 42.85 3.035 ;
      RECT 42.62 2.365 44.87 2.535 ;
      RECT 44.15 2.045 44.32 2.535 ;
      RECT 44.14 3.155 44.31 4.005 ;
      RECT 43.225 3.155 44.53 3.325 ;
      RECT 44.285 2.705 44.53 3.325 ;
      RECT 43.225 2.785 43.395 3.325 ;
      RECT 43.02 2.785 43.395 2.955 ;
      RECT 43.2 6.265 43.895 6.895 ;
      RECT 43.725 4.685 43.895 6.895 ;
      RECT 43.63 4.685 43.96 5.665 ;
      RECT 43.23 3.495 43.56 4.175 ;
      RECT 42.32 3.495 42.72 4.175 ;
      RECT 42.32 3.495 43.56 3.665 ;
      RECT 41.82 3.075 42.14 4.175 ;
      RECT 41.82 3.075 42.27 3.325 ;
      RECT 41.82 3.075 42.45 3.245 ;
      RECT 42.28 2.025 42.45 3.245 ;
      RECT 42.28 2.025 43.235 2.195 ;
      RECT 41.82 6.265 42.515 6.895 ;
      RECT 42.345 4.685 42.515 6.895 ;
      RECT 42.25 4.685 42.58 5.665 ;
      RECT 41.84 5.825 42.175 6.075 ;
      RECT 41.295 5.825 41.63 6.075 ;
      RECT 41.295 5.875 42.175 6.045 ;
      RECT 40.955 6.265 41.65 6.895 ;
      RECT 40.955 4.685 41.125 6.895 ;
      RECT 40.89 4.685 41.22 5.665 ;
      RECT 40.45 3.205 40.78 4.16 ;
      RECT 40.45 3.205 41.13 3.375 ;
      RECT 40.96 1.965 41.13 3.375 ;
      RECT 40.87 1.965 41.2 2.605 ;
      RECT 39.93 3.205 40.26 4.16 ;
      RECT 39.58 3.205 40.26 3.375 ;
      RECT 39.58 1.965 39.75 3.375 ;
      RECT 39.51 1.965 39.84 2.605 ;
      RECT 39.72 5.875 39.89 6.725 ;
      RECT 38.995 5.825 39.33 6.075 ;
      RECT 38.995 5.875 39.89 6.045 ;
      RECT 39.06 2.785 39.41 3.035 ;
      RECT 38.54 2.785 38.87 3.035 ;
      RECT 38.54 2.815 39.41 2.985 ;
      RECT 38.655 6.265 39.35 6.895 ;
      RECT 38.655 4.685 38.825 6.895 ;
      RECT 38.59 4.685 38.92 5.665 ;
      RECT 38.15 5.825 38.485 6.095 ;
      RECT 37.68 5.875 38.485 6.045 ;
      RECT 38.12 3.195 38.45 4.175 ;
      RECT 38.12 1.965 38.37 4.175 ;
      RECT 38.12 1.965 38.45 2.595 ;
      RECT 35.59 7.855 35.76 8.305 ;
      RECT 35.645 6.075 35.815 8.025 ;
      RECT 35.59 5.015 35.76 6.245 ;
      RECT 35.07 5.015 35.24 8.305 ;
      RECT 35.07 7.315 35.475 7.645 ;
      RECT 35.07 6.475 35.475 6.805 ;
      RECT 32.9 1.74 33.07 2.935 ;
      RECT 32.9 1.74 33.365 1.91 ;
      RECT 32.9 6.97 33.365 7.14 ;
      RECT 32.9 5.945 33.07 7.14 ;
      RECT 31.91 1.74 32.08 2.935 ;
      RECT 31.91 1.74 32.375 1.91 ;
      RECT 31.91 6.97 32.375 7.14 ;
      RECT 31.91 5.945 32.08 7.14 ;
      RECT 30.055 2.635 30.225 3.865 ;
      RECT 30.11 0.855 30.28 2.805 ;
      RECT 30.055 0.575 30.225 1.025 ;
      RECT 30.055 7.855 30.225 8.305 ;
      RECT 30.11 6.075 30.28 8.025 ;
      RECT 30.055 5.015 30.225 6.245 ;
      RECT 29.535 0.575 29.705 3.865 ;
      RECT 29.535 2.075 29.94 2.405 ;
      RECT 29.535 1.235 29.94 1.565 ;
      RECT 29.535 5.015 29.705 8.305 ;
      RECT 29.535 7.315 29.94 7.645 ;
      RECT 29.535 6.475 29.94 6.805 ;
      RECT 29.115 5.94 29.285 7.22 ;
      RECT 29.105 5.94 29.285 6.18 ;
      RECT 27.27 3.495 27.65 4.175 ;
      RECT 27.48 2.365 27.65 4.175 ;
      RECT 25.4 2.365 25.63 3.035 ;
      RECT 25.4 2.365 27.65 2.535 ;
      RECT 26.93 2.045 27.1 2.535 ;
      RECT 26.92 3.155 27.09 4.005 ;
      RECT 26.005 3.155 27.31 3.325 ;
      RECT 27.065 2.705 27.31 3.325 ;
      RECT 26.005 2.785 26.175 3.325 ;
      RECT 25.8 2.785 26.175 2.955 ;
      RECT 25.98 6.265 26.675 6.895 ;
      RECT 26.505 4.685 26.675 6.895 ;
      RECT 26.41 4.685 26.74 5.665 ;
      RECT 26.01 3.495 26.34 4.175 ;
      RECT 25.1 3.495 25.5 4.175 ;
      RECT 25.1 3.495 26.34 3.665 ;
      RECT 24.6 3.075 24.92 4.175 ;
      RECT 24.6 3.075 25.05 3.325 ;
      RECT 24.6 3.075 25.23 3.245 ;
      RECT 25.06 2.025 25.23 3.245 ;
      RECT 25.06 2.025 26.015 2.195 ;
      RECT 24.6 6.265 25.295 6.895 ;
      RECT 25.125 4.685 25.295 6.895 ;
      RECT 25.03 4.685 25.36 5.665 ;
      RECT 24.62 5.825 24.955 6.075 ;
      RECT 24.075 5.825 24.41 6.075 ;
      RECT 24.075 5.875 24.955 6.045 ;
      RECT 23.735 6.265 24.43 6.895 ;
      RECT 23.735 4.685 23.905 6.895 ;
      RECT 23.67 4.685 24 5.665 ;
      RECT 23.23 3.205 23.56 4.16 ;
      RECT 23.23 3.205 23.91 3.375 ;
      RECT 23.74 1.965 23.91 3.375 ;
      RECT 23.65 1.965 23.98 2.605 ;
      RECT 22.71 3.205 23.04 4.16 ;
      RECT 22.36 3.205 23.04 3.375 ;
      RECT 22.36 1.965 22.53 3.375 ;
      RECT 22.29 1.965 22.62 2.605 ;
      RECT 22.5 5.875 22.67 6.725 ;
      RECT 21.775 5.825 22.11 6.075 ;
      RECT 21.775 5.875 22.67 6.045 ;
      RECT 21.84 2.785 22.19 3.035 ;
      RECT 21.32 2.785 21.65 3.035 ;
      RECT 21.32 2.815 22.19 2.985 ;
      RECT 21.435 6.265 22.13 6.895 ;
      RECT 21.435 4.685 21.605 6.895 ;
      RECT 21.37 4.685 21.7 5.665 ;
      RECT 20.93 5.825 21.265 6.095 ;
      RECT 20.46 5.875 21.265 6.045 ;
      RECT 20.9 3.195 21.23 4.175 ;
      RECT 20.9 1.965 21.15 4.175 ;
      RECT 20.9 1.965 21.23 2.595 ;
      RECT 18.37 7.855 18.54 8.305 ;
      RECT 18.425 6.075 18.595 8.025 ;
      RECT 18.37 5.015 18.54 6.245 ;
      RECT 17.85 5.015 18.02 8.305 ;
      RECT 17.85 7.315 18.255 7.645 ;
      RECT 17.85 6.475 18.255 6.805 ;
      RECT 15.68 1.74 15.85 2.935 ;
      RECT 15.68 1.74 16.145 1.91 ;
      RECT 15.68 6.97 16.145 7.14 ;
      RECT 15.68 5.945 15.85 7.14 ;
      RECT 14.69 1.74 14.86 2.935 ;
      RECT 14.69 1.74 15.155 1.91 ;
      RECT 14.69 6.97 15.155 7.14 ;
      RECT 14.69 5.945 14.86 7.14 ;
      RECT 12.835 2.635 13.005 3.865 ;
      RECT 12.89 0.855 13.06 2.805 ;
      RECT 12.835 0.575 13.005 1.025 ;
      RECT 12.835 7.855 13.005 8.305 ;
      RECT 12.89 6.075 13.06 8.025 ;
      RECT 12.835 5.015 13.005 6.245 ;
      RECT 12.315 0.575 12.485 3.865 ;
      RECT 12.315 2.075 12.72 2.405 ;
      RECT 12.315 1.235 12.72 1.565 ;
      RECT 12.315 5.015 12.485 8.305 ;
      RECT 12.315 7.315 12.72 7.645 ;
      RECT 12.315 6.475 12.72 6.805 ;
      RECT 11.895 5.94 12.065 7.22 ;
      RECT 11.885 5.94 12.065 6.18 ;
      RECT 10.05 3.495 10.43 4.175 ;
      RECT 10.26 2.365 10.43 4.175 ;
      RECT 8.18 2.365 8.41 3.035 ;
      RECT 8.18 2.365 10.43 2.535 ;
      RECT 9.71 2.045 9.88 2.535 ;
      RECT 9.7 3.155 9.87 4.005 ;
      RECT 8.785 3.155 10.09 3.325 ;
      RECT 9.845 2.705 10.09 3.325 ;
      RECT 8.785 2.785 8.955 3.325 ;
      RECT 8.58 2.785 8.955 2.955 ;
      RECT 8.76 6.265 9.455 6.895 ;
      RECT 9.285 4.685 9.455 6.895 ;
      RECT 9.19 4.685 9.52 5.665 ;
      RECT 8.79 3.495 9.12 4.175 ;
      RECT 7.88 3.495 8.28 4.175 ;
      RECT 7.88 3.495 9.12 3.665 ;
      RECT 7.38 3.075 7.7 4.175 ;
      RECT 7.38 3.075 7.83 3.325 ;
      RECT 7.38 3.075 8.01 3.245 ;
      RECT 7.84 2.025 8.01 3.245 ;
      RECT 7.84 2.025 8.795 2.195 ;
      RECT 7.38 6.265 8.075 6.895 ;
      RECT 7.905 4.685 8.075 6.895 ;
      RECT 7.81 4.685 8.14 5.665 ;
      RECT 7.4 5.825 7.735 6.075 ;
      RECT 6.855 5.825 7.19 6.075 ;
      RECT 6.855 5.875 7.735 6.045 ;
      RECT 6.515 6.265 7.21 6.895 ;
      RECT 6.515 4.685 6.685 6.895 ;
      RECT 6.45 4.685 6.78 5.665 ;
      RECT 6.01 3.205 6.34 4.16 ;
      RECT 6.01 3.205 6.69 3.375 ;
      RECT 6.52 1.965 6.69 3.375 ;
      RECT 6.43 1.965 6.76 2.605 ;
      RECT 5.49 3.205 5.82 4.16 ;
      RECT 5.14 3.205 5.82 3.375 ;
      RECT 5.14 1.965 5.31 3.375 ;
      RECT 5.07 1.965 5.4 2.605 ;
      RECT 5.28 5.875 5.45 6.725 ;
      RECT 4.555 5.825 4.89 6.075 ;
      RECT 4.555 5.875 5.45 6.045 ;
      RECT 4.62 2.785 4.97 3.035 ;
      RECT 4.1 2.785 4.43 3.035 ;
      RECT 4.1 2.815 4.97 2.985 ;
      RECT 4.215 6.265 4.91 6.895 ;
      RECT 4.215 4.685 4.385 6.895 ;
      RECT 4.15 4.685 4.48 5.665 ;
      RECT 3.71 5.825 4.045 6.095 ;
      RECT 3.24 5.875 4.045 6.045 ;
      RECT 3.68 3.195 4.01 4.175 ;
      RECT 3.68 1.965 3.93 4.175 ;
      RECT 3.68 1.965 4.01 2.595 ;
      RECT 1.15 7.855 1.32 8.305 ;
      RECT 1.205 6.075 1.375 8.025 ;
      RECT 1.15 5.015 1.32 6.245 ;
      RECT 0.63 5.015 0.8 8.305 ;
      RECT 0.63 7.315 1.035 7.645 ;
      RECT 0.63 6.475 1.035 6.805 ;
      RECT -2.26 7.855 -2.09 8.305 ;
      RECT -2.205 6.075 -2.035 8.025 ;
      RECT -2.26 5.015 -2.09 6.245 ;
      RECT -2.78 5.015 -2.61 8.305 ;
      RECT -2.78 7.315 -2.375 7.645 ;
      RECT -2.78 6.475 -2.375 6.805 ;
      RECT 84.93 0.575 85.1 1.085 ;
      RECT 84.93 2.395 85.1 3.865 ;
      RECT 84.93 5.015 85.1 6.485 ;
      RECT 84.93 7.795 85.1 8.305 ;
      RECT 83.94 0.575 84.11 1.085 ;
      RECT 83.94 2.395 84.11 3.865 ;
      RECT 83.94 5.015 84.11 6.485 ;
      RECT 83.94 7.795 84.11 8.305 ;
      RECT 82.575 0.575 82.745 3.865 ;
      RECT 82.575 5.015 82.745 8.305 ;
      RECT 82.145 0.575 82.315 1.085 ;
      RECT 82.145 1.655 82.315 3.865 ;
      RECT 82.145 5.015 82.315 7.225 ;
      RECT 82.145 7.795 82.315 8.305 ;
      RECT 80.775 1.66 80.945 2.935 ;
      RECT 78.505 5.825 78.84 6.095 ;
      RECT 78.005 2.785 78.555 2.985 ;
      RECT 77.66 5.825 77.995 6.075 ;
      RECT 77.125 5.825 77.46 6.095 ;
      RECT 75.74 2.785 76.09 3.035 ;
      RECT 74.88 2.785 75.23 3.035 ;
      RECT 74.36 2.785 74.71 3.035 ;
      RECT 70.89 5.015 71.06 8.305 ;
      RECT 70.46 5.015 70.63 7.225 ;
      RECT 70.46 7.795 70.63 8.305 ;
      RECT 69.09 5.945 69.26 7.22 ;
      RECT 67.71 0.575 67.88 1.085 ;
      RECT 67.71 2.395 67.88 3.865 ;
      RECT 67.71 5.015 67.88 6.485 ;
      RECT 67.71 7.795 67.88 8.305 ;
      RECT 66.72 0.575 66.89 1.085 ;
      RECT 66.72 2.395 66.89 3.865 ;
      RECT 66.72 5.015 66.89 6.485 ;
      RECT 66.72 7.795 66.89 8.305 ;
      RECT 65.355 0.575 65.525 3.865 ;
      RECT 65.355 5.015 65.525 8.305 ;
      RECT 64.925 0.575 65.095 1.085 ;
      RECT 64.925 1.655 65.095 3.865 ;
      RECT 64.925 5.015 65.095 7.225 ;
      RECT 64.925 7.795 65.095 8.305 ;
      RECT 63.555 1.66 63.725 2.935 ;
      RECT 61.285 5.825 61.62 6.095 ;
      RECT 60.785 2.785 61.335 2.985 ;
      RECT 60.44 5.825 60.775 6.075 ;
      RECT 59.905 5.825 60.24 6.095 ;
      RECT 58.52 2.785 58.87 3.035 ;
      RECT 57.66 2.785 58.01 3.035 ;
      RECT 57.14 2.785 57.49 3.035 ;
      RECT 53.67 5.015 53.84 8.305 ;
      RECT 53.24 5.015 53.41 7.225 ;
      RECT 53.24 7.795 53.41 8.305 ;
      RECT 51.87 5.945 52.04 7.22 ;
      RECT 50.49 0.575 50.66 1.085 ;
      RECT 50.49 2.395 50.66 3.865 ;
      RECT 50.49 5.015 50.66 6.485 ;
      RECT 50.49 7.795 50.66 8.305 ;
      RECT 49.5 0.575 49.67 1.085 ;
      RECT 49.5 2.395 49.67 3.865 ;
      RECT 49.5 5.015 49.67 6.485 ;
      RECT 49.5 7.795 49.67 8.305 ;
      RECT 48.135 0.575 48.305 3.865 ;
      RECT 48.135 5.015 48.305 8.305 ;
      RECT 47.705 0.575 47.875 1.085 ;
      RECT 47.705 1.655 47.875 3.865 ;
      RECT 47.705 5.015 47.875 7.225 ;
      RECT 47.705 7.795 47.875 8.305 ;
      RECT 46.335 1.66 46.505 2.935 ;
      RECT 44.065 5.825 44.4 6.095 ;
      RECT 43.565 2.785 44.115 2.985 ;
      RECT 43.22 5.825 43.555 6.075 ;
      RECT 42.685 5.825 43.02 6.095 ;
      RECT 41.3 2.785 41.65 3.035 ;
      RECT 40.44 2.785 40.79 3.035 ;
      RECT 39.92 2.785 40.27 3.035 ;
      RECT 36.45 5.015 36.62 8.305 ;
      RECT 36.02 5.015 36.19 7.225 ;
      RECT 36.02 7.795 36.19 8.305 ;
      RECT 34.65 5.945 34.82 7.22 ;
      RECT 33.27 0.575 33.44 1.085 ;
      RECT 33.27 2.395 33.44 3.865 ;
      RECT 33.27 5.015 33.44 6.485 ;
      RECT 33.27 7.795 33.44 8.305 ;
      RECT 32.28 0.575 32.45 1.085 ;
      RECT 32.28 2.395 32.45 3.865 ;
      RECT 32.28 5.015 32.45 6.485 ;
      RECT 32.28 7.795 32.45 8.305 ;
      RECT 30.915 0.575 31.085 3.865 ;
      RECT 30.915 5.015 31.085 8.305 ;
      RECT 30.485 0.575 30.655 1.085 ;
      RECT 30.485 1.655 30.655 3.865 ;
      RECT 30.485 5.015 30.655 7.225 ;
      RECT 30.485 7.795 30.655 8.305 ;
      RECT 29.115 1.66 29.285 2.935 ;
      RECT 26.845 5.825 27.18 6.095 ;
      RECT 26.345 2.785 26.895 2.985 ;
      RECT 26 5.825 26.335 6.075 ;
      RECT 25.465 5.825 25.8 6.095 ;
      RECT 24.08 2.785 24.43 3.035 ;
      RECT 23.22 2.785 23.57 3.035 ;
      RECT 22.7 2.785 23.05 3.035 ;
      RECT 19.23 5.015 19.4 8.305 ;
      RECT 18.8 5.015 18.97 7.225 ;
      RECT 18.8 7.795 18.97 8.305 ;
      RECT 17.43 5.945 17.6 7.22 ;
      RECT 16.05 0.575 16.22 1.085 ;
      RECT 16.05 2.395 16.22 3.865 ;
      RECT 16.05 5.015 16.22 6.485 ;
      RECT 16.05 7.795 16.22 8.305 ;
      RECT 15.06 0.575 15.23 1.085 ;
      RECT 15.06 2.395 15.23 3.865 ;
      RECT 15.06 5.015 15.23 6.485 ;
      RECT 15.06 7.795 15.23 8.305 ;
      RECT 13.695 0.575 13.865 3.865 ;
      RECT 13.695 5.015 13.865 8.305 ;
      RECT 13.265 0.575 13.435 1.085 ;
      RECT 13.265 1.655 13.435 3.865 ;
      RECT 13.265 5.015 13.435 7.225 ;
      RECT 13.265 7.795 13.435 8.305 ;
      RECT 11.895 1.66 12.065 2.935 ;
      RECT 9.625 5.825 9.96 6.095 ;
      RECT 9.125 2.785 9.675 2.985 ;
      RECT 8.78 5.825 9.115 6.075 ;
      RECT 8.245 5.825 8.58 6.095 ;
      RECT 6.86 2.785 7.21 3.035 ;
      RECT 6 2.785 6.35 3.035 ;
      RECT 5.48 2.785 5.83 3.035 ;
      RECT 2.01 5.015 2.18 8.305 ;
      RECT 1.58 5.015 1.75 7.225 ;
      RECT 1.58 7.795 1.75 8.305 ;
      RECT 0.21 5.945 0.38 7.22 ;
      RECT -1.83 5.015 -1.66 7.225 ;
      RECT -1.83 7.795 -1.66 8.305 ;
      RECT -3.2 5.945 -3.03 7.22 ;
  END
END sky130_osu_ring_oscillator_mpr2ct_8_b0r2

MACRO sky130_osu_ring_oscillator_mpr2ea_8_b0r1
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 3.275 0 ;
  SIZE 84.425 BY 8.88 ;
  SYMMETRY X Y R90 ;
  SITE CoreSite ;
  OBS
    LAYER met3 ;
      RECT 72.13 7.055 72.5 7.425 ;
      RECT 72.13 7.09 74.115 7.39 ;
      RECT 73.815 2.28 74.115 7.39 ;
      RECT 70.815 2.015 71.145 2.745 ;
      RECT 69.935 2.015 70.265 2.745 ;
      RECT 73.015 2.28 74.305 2.58 ;
      RECT 73.975 1.85 74.305 2.58 ;
      RECT 69.935 2.28 72.075 2.58 ;
      RECT 71.775 1.965 72.075 2.58 ;
      RECT 73.015 1.98 73.32 2.58 ;
      RECT 71.775 1.965 73.135 2.275 ;
      RECT 70.435 3.535 70.765 3.865 ;
      RECT 69.23 3.55 70.765 3.85 ;
      RECT 69.23 2.43 69.53 3.85 ;
      RECT 68.975 2.415 69.305 2.745 ;
      RECT 55.805 7.055 56.175 7.425 ;
      RECT 55.805 7.09 57.79 7.39 ;
      RECT 57.49 2.28 57.79 7.39 ;
      RECT 54.49 2.015 54.82 2.745 ;
      RECT 53.61 2.015 53.94 2.745 ;
      RECT 56.69 2.28 57.98 2.58 ;
      RECT 57.65 1.85 57.98 2.58 ;
      RECT 53.61 2.28 55.75 2.58 ;
      RECT 55.45 1.965 55.75 2.58 ;
      RECT 56.69 1.98 56.995 2.58 ;
      RECT 55.45 1.965 56.81 2.275 ;
      RECT 54.11 3.535 54.44 3.865 ;
      RECT 52.905 3.55 54.44 3.85 ;
      RECT 52.905 2.43 53.205 3.85 ;
      RECT 52.65 2.415 52.98 2.745 ;
      RECT 39.48 7.055 39.85 7.425 ;
      RECT 39.48 7.09 41.465 7.39 ;
      RECT 41.165 2.28 41.465 7.39 ;
      RECT 38.165 2.015 38.495 2.745 ;
      RECT 37.285 2.015 37.615 2.745 ;
      RECT 40.365 2.28 41.655 2.58 ;
      RECT 41.325 1.85 41.655 2.58 ;
      RECT 37.285 2.28 39.425 2.58 ;
      RECT 39.125 1.965 39.425 2.58 ;
      RECT 40.365 1.98 40.67 2.58 ;
      RECT 39.125 1.965 40.485 2.275 ;
      RECT 37.785 3.535 38.115 3.865 ;
      RECT 36.58 3.55 38.115 3.85 ;
      RECT 36.58 2.43 36.88 3.85 ;
      RECT 36.325 2.415 36.655 2.745 ;
      RECT 23.155 7.055 23.525 7.425 ;
      RECT 23.155 7.09 25.14 7.39 ;
      RECT 24.84 2.28 25.14 7.39 ;
      RECT 21.84 2.015 22.17 2.745 ;
      RECT 20.96 2.015 21.29 2.745 ;
      RECT 24.04 2.28 25.33 2.58 ;
      RECT 25 1.85 25.33 2.58 ;
      RECT 20.96 2.28 23.1 2.58 ;
      RECT 22.8 1.965 23.1 2.58 ;
      RECT 24.04 1.98 24.345 2.58 ;
      RECT 22.8 1.965 24.16 2.275 ;
      RECT 21.46 3.535 21.79 3.865 ;
      RECT 20.255 3.55 21.79 3.85 ;
      RECT 20.255 2.43 20.555 3.85 ;
      RECT 20 2.415 20.33 2.745 ;
      RECT 6.83 7.055 7.2 7.425 ;
      RECT 6.83 7.09 8.815 7.39 ;
      RECT 8.515 2.28 8.815 7.39 ;
      RECT 5.515 2.015 5.845 2.745 ;
      RECT 4.635 2.015 4.965 2.745 ;
      RECT 7.715 2.28 9.005 2.58 ;
      RECT 8.675 1.85 9.005 2.58 ;
      RECT 4.635 2.28 6.775 2.58 ;
      RECT 6.475 1.965 6.775 2.58 ;
      RECT 7.715 1.98 8.02 2.58 ;
      RECT 6.475 1.965 7.835 2.275 ;
      RECT 5.135 3.535 5.465 3.865 ;
      RECT 3.93 3.55 5.465 3.85 ;
      RECT 3.93 2.43 4.23 3.85 ;
      RECT 3.675 2.415 4.005 2.745 ;
      RECT 74.455 2.975 74.785 3.705 ;
      RECT 72.375 2.575 72.705 3.305 ;
      RECT 68.255 2.415 68.585 3.145 ;
      RECT 67.255 1.855 67.585 2.585 ;
      RECT 65.815 2.575 66.145 3.305 ;
      RECT 58.13 2.975 58.46 3.705 ;
      RECT 56.05 2.575 56.38 3.305 ;
      RECT 51.93 2.415 52.26 3.145 ;
      RECT 50.93 1.855 51.26 2.585 ;
      RECT 49.49 2.575 49.82 3.305 ;
      RECT 41.805 2.975 42.135 3.705 ;
      RECT 39.725 2.575 40.055 3.305 ;
      RECT 35.605 2.415 35.935 3.145 ;
      RECT 34.605 1.855 34.935 2.585 ;
      RECT 33.165 2.575 33.495 3.305 ;
      RECT 25.48 2.975 25.81 3.705 ;
      RECT 23.4 2.575 23.73 3.305 ;
      RECT 19.28 2.415 19.61 3.145 ;
      RECT 18.28 1.855 18.61 2.585 ;
      RECT 16.84 2.575 17.17 3.305 ;
      RECT 9.155 2.975 9.485 3.705 ;
      RECT 7.075 2.575 7.405 3.305 ;
      RECT 2.955 2.415 3.285 3.145 ;
      RECT 1.955 1.855 2.285 2.585 ;
      RECT 0.515 2.575 0.845 3.305 ;
    LAYER via2 ;
      RECT 74.52 3.04 74.72 3.24 ;
      RECT 74.04 2.315 74.24 2.515 ;
      RECT 72.44 3.04 72.64 3.24 ;
      RECT 72.215 7.14 72.415 7.34 ;
      RECT 70.88 2.48 71.08 2.68 ;
      RECT 70.5 3.6 70.7 3.8 ;
      RECT 70 2.48 70.2 2.68 ;
      RECT 69.04 2.48 69.24 2.68 ;
      RECT 68.32 2.48 68.52 2.68 ;
      RECT 67.32 1.92 67.52 2.12 ;
      RECT 65.88 3.04 66.08 3.24 ;
      RECT 58.195 3.04 58.395 3.24 ;
      RECT 57.715 2.315 57.915 2.515 ;
      RECT 56.115 3.04 56.315 3.24 ;
      RECT 55.89 7.14 56.09 7.34 ;
      RECT 54.555 2.48 54.755 2.68 ;
      RECT 54.175 3.6 54.375 3.8 ;
      RECT 53.675 2.48 53.875 2.68 ;
      RECT 52.715 2.48 52.915 2.68 ;
      RECT 51.995 2.48 52.195 2.68 ;
      RECT 50.995 1.92 51.195 2.12 ;
      RECT 49.555 3.04 49.755 3.24 ;
      RECT 41.87 3.04 42.07 3.24 ;
      RECT 41.39 2.315 41.59 2.515 ;
      RECT 39.79 3.04 39.99 3.24 ;
      RECT 39.565 7.14 39.765 7.34 ;
      RECT 38.23 2.48 38.43 2.68 ;
      RECT 37.85 3.6 38.05 3.8 ;
      RECT 37.35 2.48 37.55 2.68 ;
      RECT 36.39 2.48 36.59 2.68 ;
      RECT 35.67 2.48 35.87 2.68 ;
      RECT 34.67 1.92 34.87 2.12 ;
      RECT 33.23 3.04 33.43 3.24 ;
      RECT 25.545 3.04 25.745 3.24 ;
      RECT 25.065 2.315 25.265 2.515 ;
      RECT 23.465 3.04 23.665 3.24 ;
      RECT 23.24 7.14 23.44 7.34 ;
      RECT 21.905 2.48 22.105 2.68 ;
      RECT 21.525 3.6 21.725 3.8 ;
      RECT 21.025 2.48 21.225 2.68 ;
      RECT 20.065 2.48 20.265 2.68 ;
      RECT 19.345 2.48 19.545 2.68 ;
      RECT 18.345 1.92 18.545 2.12 ;
      RECT 16.905 3.04 17.105 3.24 ;
      RECT 9.22 3.04 9.42 3.24 ;
      RECT 8.74 2.315 8.94 2.515 ;
      RECT 7.14 3.04 7.34 3.24 ;
      RECT 6.915 7.14 7.115 7.34 ;
      RECT 5.58 2.48 5.78 2.68 ;
      RECT 5.2 3.6 5.4 3.8 ;
      RECT 4.7 2.48 4.9 2.68 ;
      RECT 3.74 2.48 3.94 2.68 ;
      RECT 3.02 2.48 3.22 2.68 ;
      RECT 2.02 1.92 2.22 2.12 ;
      RECT 0.58 3.04 0.78 3.24 ;
    LAYER met2 ;
      RECT -2.045 8.4 80.78 8.57 ;
      RECT 80.61 7.275 80.78 8.57 ;
      RECT -2.045 6.255 -1.875 8.57 ;
      RECT 80.58 7.275 80.93 7.625 ;
      RECT -2.105 6.255 -1.815 6.605 ;
      RECT 77.42 6.22 77.74 6.545 ;
      RECT 77.45 5.695 77.62 6.545 ;
      RECT 77.45 5.695 77.625 6.045 ;
      RECT 77.45 5.695 78.425 5.87 ;
      RECT 78.25 1.965 78.425 5.87 ;
      RECT 78.195 1.965 78.545 2.315 ;
      RECT 78.22 6.655 78.545 6.98 ;
      RECT 77.105 6.745 78.545 6.915 ;
      RECT 77.105 2.395 77.265 6.915 ;
      RECT 77.42 2.365 77.74 2.685 ;
      RECT 77.105 2.395 77.74 2.565 ;
      RECT 76.37 5.84 76.71 6.19 ;
      RECT 76.455 2.705 76.625 6.19 ;
      RECT 76.38 2.705 76.72 3.055 ;
      RECT 67.28 1.835 67.56 2.205 ;
      RECT 67.315 1.29 67.485 2.205 ;
      RECT 75.89 1.29 76.06 1.815 ;
      RECT 75.8 1.46 76.14 1.81 ;
      RECT 67.315 1.29 76.06 1.46 ;
      RECT 72.52 2.395 72.8 2.765 ;
      RECT 71.45 2.42 71.71 2.74 ;
      RECT 74 2.23 74.28 2.6 ;
      RECT 74.61 2.14 74.87 2.46 ;
      RECT 71.51 1.58 71.65 2.74 ;
      RECT 72.59 1.58 72.73 2.765 ;
      RECT 73.71 2.23 74.87 2.37 ;
      RECT 73.71 1.58 73.85 2.37 ;
      RECT 71.51 1.58 73.85 1.72 ;
      RECT 74.48 2.955 74.76 3.325 ;
      RECT 74.49 2.7 74.75 3.325 ;
      RECT 71.54 3.72 73.715 3.885 ;
      RECT 73.57 2.6 73.715 3.885 ;
      RECT 70.46 3.515 70.74 3.885 ;
      RECT 70.46 3.63 71.68 3.77 ;
      RECT 73.29 2.6 73.715 2.74 ;
      RECT 73.29 2.42 73.55 2.74 ;
      RECT 66.63 4 70.29 4.14 ;
      RECT 70.15 3.185 70.29 4.14 ;
      RECT 66.63 3.07 66.77 4.14 ;
      RECT 73.17 3.26 73.43 3.58 ;
      RECT 70.15 3.185 72.68 3.325 ;
      RECT 72.4 2.955 72.68 3.325 ;
      RECT 66.63 3.07 67.08 3.325 ;
      RECT 66.8 2.955 67.08 3.325 ;
      RECT 73.17 3.07 73.37 3.58 ;
      RECT 72.4 3.07 73.37 3.21 ;
      RECT 72.97 1.86 73.11 3.21 ;
      RECT 72.91 1.86 73.17 2.18 ;
      RECT 64.23 6.655 64.58 7.005 ;
      RECT 72.785 6.61 73.135 6.96 ;
      RECT 64.23 6.685 73.135 6.885 ;
      RECT 66.81 2.42 67.07 2.74 ;
      RECT 66.81 2.51 67.85 2.65 ;
      RECT 67.71 1.72 67.85 2.65 ;
      RECT 70.47 1.86 70.73 2.18 ;
      RECT 67.71 1.72 70.67 1.86 ;
      RECT 69.85 2.7 70.11 3.02 ;
      RECT 69.85 2.7 70.17 2.93 ;
      RECT 69.96 2.395 70.24 2.765 ;
      RECT 69.55 3.26 69.87 3.58 ;
      RECT 69.55 2.14 69.69 3.58 ;
      RECT 69.49 2.14 69.75 2.46 ;
      RECT 67.05 3.54 67.31 3.86 ;
      RECT 67.05 3.63 68.73 3.77 ;
      RECT 68.59 3.35 68.73 3.77 ;
      RECT 68.59 3.35 69.03 3.58 ;
      RECT 68.77 3.26 69.03 3.58 ;
      RECT 68.09 2.42 68.49 2.93 ;
      RECT 68.28 2.395 68.56 2.765 ;
      RECT 68.03 2.42 68.56 2.74 ;
      RECT 61.095 6.22 61.415 6.545 ;
      RECT 61.125 5.695 61.295 6.545 ;
      RECT 61.125 5.695 61.3 6.045 ;
      RECT 61.125 5.695 62.1 5.87 ;
      RECT 61.925 1.965 62.1 5.87 ;
      RECT 61.87 1.965 62.22 2.315 ;
      RECT 61.895 6.655 62.22 6.98 ;
      RECT 60.78 6.745 62.22 6.915 ;
      RECT 60.78 2.395 60.94 6.915 ;
      RECT 61.095 2.365 61.415 2.685 ;
      RECT 60.78 2.395 61.415 2.565 ;
      RECT 60.045 5.84 60.385 6.19 ;
      RECT 60.13 2.705 60.3 6.19 ;
      RECT 60.055 2.705 60.395 3.055 ;
      RECT 50.955 1.835 51.235 2.205 ;
      RECT 50.99 1.29 51.16 2.205 ;
      RECT 59.565 1.29 59.735 1.815 ;
      RECT 59.475 1.46 59.815 1.81 ;
      RECT 50.99 1.29 59.735 1.46 ;
      RECT 56.195 2.395 56.475 2.765 ;
      RECT 55.125 2.42 55.385 2.74 ;
      RECT 57.675 2.23 57.955 2.6 ;
      RECT 58.285 2.14 58.545 2.46 ;
      RECT 55.185 1.58 55.325 2.74 ;
      RECT 56.265 1.58 56.405 2.765 ;
      RECT 57.385 2.23 58.545 2.37 ;
      RECT 57.385 1.58 57.525 2.37 ;
      RECT 55.185 1.58 57.525 1.72 ;
      RECT 58.155 2.955 58.435 3.325 ;
      RECT 58.165 2.7 58.425 3.325 ;
      RECT 55.215 3.72 57.39 3.885 ;
      RECT 57.245 2.6 57.39 3.885 ;
      RECT 54.135 3.515 54.415 3.885 ;
      RECT 54.135 3.63 55.355 3.77 ;
      RECT 56.965 2.6 57.39 2.74 ;
      RECT 56.965 2.42 57.225 2.74 ;
      RECT 50.305 4 53.965 4.14 ;
      RECT 53.825 3.185 53.965 4.14 ;
      RECT 50.305 3.07 50.445 4.14 ;
      RECT 56.845 3.26 57.105 3.58 ;
      RECT 53.825 3.185 56.355 3.325 ;
      RECT 56.075 2.955 56.355 3.325 ;
      RECT 50.305 3.07 50.755 3.325 ;
      RECT 50.475 2.955 50.755 3.325 ;
      RECT 56.845 3.07 57.045 3.58 ;
      RECT 56.075 3.07 57.045 3.21 ;
      RECT 56.645 1.86 56.785 3.21 ;
      RECT 56.585 1.86 56.845 2.18 ;
      RECT 47.905 6.655 48.255 7.005 ;
      RECT 56.455 6.61 56.805 6.96 ;
      RECT 47.905 6.685 56.805 6.885 ;
      RECT 50.485 2.42 50.745 2.74 ;
      RECT 50.485 2.51 51.525 2.65 ;
      RECT 51.385 1.72 51.525 2.65 ;
      RECT 54.145 1.86 54.405 2.18 ;
      RECT 51.385 1.72 54.345 1.86 ;
      RECT 53.525 2.7 53.785 3.02 ;
      RECT 53.525 2.7 53.845 2.93 ;
      RECT 53.635 2.395 53.915 2.765 ;
      RECT 53.225 3.26 53.545 3.58 ;
      RECT 53.225 2.14 53.365 3.58 ;
      RECT 53.165 2.14 53.425 2.46 ;
      RECT 50.725 3.54 50.985 3.86 ;
      RECT 50.725 3.63 52.405 3.77 ;
      RECT 52.265 3.35 52.405 3.77 ;
      RECT 52.265 3.35 52.705 3.58 ;
      RECT 52.445 3.26 52.705 3.58 ;
      RECT 51.765 2.42 52.165 2.93 ;
      RECT 51.955 2.395 52.235 2.765 ;
      RECT 51.705 2.42 52.235 2.74 ;
      RECT 44.77 6.22 45.09 6.545 ;
      RECT 44.8 5.695 44.97 6.545 ;
      RECT 44.8 5.695 44.975 6.045 ;
      RECT 44.8 5.695 45.775 5.87 ;
      RECT 45.6 1.965 45.775 5.87 ;
      RECT 45.545 1.965 45.895 2.315 ;
      RECT 45.57 6.655 45.895 6.98 ;
      RECT 44.455 6.745 45.895 6.915 ;
      RECT 44.455 2.395 44.615 6.915 ;
      RECT 44.77 2.365 45.09 2.685 ;
      RECT 44.455 2.395 45.09 2.565 ;
      RECT 43.72 5.84 44.06 6.19 ;
      RECT 43.805 2.705 43.975 6.19 ;
      RECT 43.73 2.705 44.07 3.055 ;
      RECT 34.63 1.835 34.91 2.205 ;
      RECT 34.665 1.29 34.835 2.205 ;
      RECT 43.24 1.29 43.41 1.815 ;
      RECT 43.15 1.46 43.49 1.81 ;
      RECT 34.665 1.29 43.41 1.46 ;
      RECT 39.87 2.395 40.15 2.765 ;
      RECT 38.8 2.42 39.06 2.74 ;
      RECT 41.35 2.23 41.63 2.6 ;
      RECT 41.96 2.14 42.22 2.46 ;
      RECT 38.86 1.58 39 2.74 ;
      RECT 39.94 1.58 40.08 2.765 ;
      RECT 41.06 2.23 42.22 2.37 ;
      RECT 41.06 1.58 41.2 2.37 ;
      RECT 38.86 1.58 41.2 1.72 ;
      RECT 41.83 2.955 42.11 3.325 ;
      RECT 41.84 2.7 42.1 3.325 ;
      RECT 38.89 3.72 41.065 3.885 ;
      RECT 40.92 2.6 41.065 3.885 ;
      RECT 37.81 3.515 38.09 3.885 ;
      RECT 37.81 3.63 39.03 3.77 ;
      RECT 40.64 2.6 41.065 2.74 ;
      RECT 40.64 2.42 40.9 2.74 ;
      RECT 33.98 4 37.64 4.14 ;
      RECT 37.5 3.185 37.64 4.14 ;
      RECT 33.98 3.07 34.12 4.14 ;
      RECT 40.52 3.26 40.78 3.58 ;
      RECT 37.5 3.185 40.03 3.325 ;
      RECT 39.75 2.955 40.03 3.325 ;
      RECT 33.98 3.07 34.43 3.325 ;
      RECT 34.15 2.955 34.43 3.325 ;
      RECT 40.52 3.07 40.72 3.58 ;
      RECT 39.75 3.07 40.72 3.21 ;
      RECT 40.32 1.86 40.46 3.21 ;
      RECT 40.26 1.86 40.52 2.18 ;
      RECT 31.625 6.66 31.975 7.01 ;
      RECT 40.13 6.615 40.48 6.965 ;
      RECT 31.625 6.69 40.48 6.89 ;
      RECT 34.16 2.42 34.42 2.74 ;
      RECT 34.16 2.51 35.2 2.65 ;
      RECT 35.06 1.72 35.2 2.65 ;
      RECT 37.82 1.86 38.08 2.18 ;
      RECT 35.06 1.72 38.02 1.86 ;
      RECT 37.2 2.7 37.46 3.02 ;
      RECT 37.2 2.7 37.52 2.93 ;
      RECT 37.31 2.395 37.59 2.765 ;
      RECT 36.9 3.26 37.22 3.58 ;
      RECT 36.9 2.14 37.04 3.58 ;
      RECT 36.84 2.14 37.1 2.46 ;
      RECT 34.4 3.54 34.66 3.86 ;
      RECT 34.4 3.63 36.08 3.77 ;
      RECT 35.94 3.35 36.08 3.77 ;
      RECT 35.94 3.35 36.38 3.58 ;
      RECT 36.12 3.26 36.38 3.58 ;
      RECT 35.44 2.42 35.84 2.93 ;
      RECT 35.63 2.395 35.91 2.765 ;
      RECT 35.38 2.42 35.91 2.74 ;
      RECT 28.445 6.22 28.765 6.545 ;
      RECT 28.475 5.695 28.645 6.545 ;
      RECT 28.475 5.695 28.65 6.045 ;
      RECT 28.475 5.695 29.45 5.87 ;
      RECT 29.275 1.965 29.45 5.87 ;
      RECT 29.22 1.965 29.57 2.315 ;
      RECT 29.245 6.655 29.57 6.98 ;
      RECT 28.13 6.745 29.57 6.915 ;
      RECT 28.13 2.395 28.29 6.915 ;
      RECT 28.445 2.365 28.765 2.685 ;
      RECT 28.13 2.395 28.765 2.565 ;
      RECT 27.395 5.84 27.735 6.19 ;
      RECT 27.48 2.705 27.65 6.19 ;
      RECT 27.405 2.705 27.745 3.055 ;
      RECT 18.305 1.835 18.585 2.205 ;
      RECT 18.34 1.29 18.51 2.205 ;
      RECT 26.915 1.29 27.085 1.815 ;
      RECT 26.825 1.46 27.165 1.81 ;
      RECT 18.34 1.29 27.085 1.46 ;
      RECT 23.545 2.395 23.825 2.765 ;
      RECT 22.475 2.42 22.735 2.74 ;
      RECT 25.025 2.23 25.305 2.6 ;
      RECT 25.635 2.14 25.895 2.46 ;
      RECT 22.535 1.58 22.675 2.74 ;
      RECT 23.615 1.58 23.755 2.765 ;
      RECT 24.735 2.23 25.895 2.37 ;
      RECT 24.735 1.58 24.875 2.37 ;
      RECT 22.535 1.58 24.875 1.72 ;
      RECT 25.505 2.955 25.785 3.325 ;
      RECT 25.515 2.7 25.775 3.325 ;
      RECT 22.565 3.72 24.74 3.885 ;
      RECT 24.595 2.6 24.74 3.885 ;
      RECT 21.485 3.515 21.765 3.885 ;
      RECT 21.485 3.63 22.705 3.77 ;
      RECT 24.315 2.6 24.74 2.74 ;
      RECT 24.315 2.42 24.575 2.74 ;
      RECT 17.655 4 21.315 4.14 ;
      RECT 21.175 3.185 21.315 4.14 ;
      RECT 17.655 3.07 17.795 4.14 ;
      RECT 24.195 3.26 24.455 3.58 ;
      RECT 21.175 3.185 23.705 3.325 ;
      RECT 23.425 2.955 23.705 3.325 ;
      RECT 17.655 3.07 18.105 3.325 ;
      RECT 17.825 2.955 18.105 3.325 ;
      RECT 24.195 3.07 24.395 3.58 ;
      RECT 23.425 3.07 24.395 3.21 ;
      RECT 23.995 1.86 24.135 3.21 ;
      RECT 23.935 1.86 24.195 2.18 ;
      RECT 15.3 6.655 15.65 7.005 ;
      RECT 23.805 6.61 24.155 6.96 ;
      RECT 15.3 6.685 24.155 6.885 ;
      RECT 17.835 2.42 18.095 2.74 ;
      RECT 17.835 2.51 18.875 2.65 ;
      RECT 18.735 1.72 18.875 2.65 ;
      RECT 21.495 1.86 21.755 2.18 ;
      RECT 18.735 1.72 21.695 1.86 ;
      RECT 20.875 2.7 21.135 3.02 ;
      RECT 20.875 2.7 21.195 2.93 ;
      RECT 20.985 2.395 21.265 2.765 ;
      RECT 20.575 3.26 20.895 3.58 ;
      RECT 20.575 2.14 20.715 3.58 ;
      RECT 20.515 2.14 20.775 2.46 ;
      RECT 18.075 3.54 18.335 3.86 ;
      RECT 18.075 3.63 19.755 3.77 ;
      RECT 19.615 3.35 19.755 3.77 ;
      RECT 19.615 3.35 20.055 3.58 ;
      RECT 19.795 3.26 20.055 3.58 ;
      RECT 19.115 2.42 19.515 2.93 ;
      RECT 19.305 2.395 19.585 2.765 ;
      RECT 19.055 2.42 19.585 2.74 ;
      RECT 12.12 6.22 12.44 6.545 ;
      RECT 12.15 5.695 12.32 6.545 ;
      RECT 12.15 5.695 12.325 6.045 ;
      RECT 12.15 5.695 13.125 5.87 ;
      RECT 12.95 1.965 13.125 5.87 ;
      RECT 12.895 1.965 13.245 2.315 ;
      RECT 12.92 6.655 13.245 6.98 ;
      RECT 11.805 6.745 13.245 6.915 ;
      RECT 11.805 2.395 11.965 6.915 ;
      RECT 12.12 2.365 12.44 2.685 ;
      RECT 11.805 2.395 12.44 2.565 ;
      RECT 11.07 5.84 11.41 6.19 ;
      RECT 11.155 2.705 11.325 6.19 ;
      RECT 11.08 2.705 11.42 3.055 ;
      RECT 1.98 1.835 2.26 2.205 ;
      RECT 2.015 1.29 2.185 2.205 ;
      RECT 10.59 1.29 10.76 1.815 ;
      RECT 10.5 1.46 10.84 1.81 ;
      RECT 2.015 1.29 10.76 1.46 ;
      RECT 7.22 2.395 7.5 2.765 ;
      RECT 6.15 2.42 6.41 2.74 ;
      RECT 8.7 2.23 8.98 2.6 ;
      RECT 9.31 2.14 9.57 2.46 ;
      RECT 6.21 1.58 6.35 2.74 ;
      RECT 7.29 1.58 7.43 2.765 ;
      RECT 8.41 2.23 9.57 2.37 ;
      RECT 8.41 1.58 8.55 2.37 ;
      RECT 6.21 1.58 8.55 1.72 ;
      RECT 9.18 2.955 9.46 3.325 ;
      RECT 9.19 2.7 9.45 3.325 ;
      RECT -1.73 6.995 -1.44 7.345 ;
      RECT -1.73 7.05 -0.445 7.225 ;
      RECT -0.62 6.685 -0.445 7.225 ;
      RECT 8.315 6.605 8.665 6.955 ;
      RECT -0.62 6.685 8.665 6.86 ;
      RECT 6.24 3.72 8.415 3.885 ;
      RECT 8.27 2.6 8.415 3.885 ;
      RECT 5.16 3.515 5.44 3.885 ;
      RECT 5.16 3.63 6.38 3.77 ;
      RECT 7.99 2.6 8.415 2.74 ;
      RECT 7.99 2.42 8.25 2.74 ;
      RECT 1.33 4 4.99 4.14 ;
      RECT 4.85 3.185 4.99 4.14 ;
      RECT 1.33 3.07 1.47 4.14 ;
      RECT 7.87 3.26 8.13 3.58 ;
      RECT 4.85 3.185 7.38 3.325 ;
      RECT 7.1 2.955 7.38 3.325 ;
      RECT 1.33 3.07 1.78 3.325 ;
      RECT 1.5 2.955 1.78 3.325 ;
      RECT 7.87 3.07 8.07 3.58 ;
      RECT 7.1 3.07 8.07 3.21 ;
      RECT 7.67 1.86 7.81 3.21 ;
      RECT 7.61 1.86 7.87 2.18 ;
      RECT 1.51 2.42 1.77 2.74 ;
      RECT 1.51 2.51 2.55 2.65 ;
      RECT 2.41 1.72 2.55 2.65 ;
      RECT 5.17 1.86 5.43 2.18 ;
      RECT 2.41 1.72 5.37 1.86 ;
      RECT 4.55 2.7 4.81 3.02 ;
      RECT 4.55 2.7 4.87 2.93 ;
      RECT 4.66 2.395 4.94 2.765 ;
      RECT 4.25 3.26 4.57 3.58 ;
      RECT 4.25 2.14 4.39 3.58 ;
      RECT 4.19 2.14 4.45 2.46 ;
      RECT 1.75 3.54 2.01 3.86 ;
      RECT 1.75 3.63 3.43 3.77 ;
      RECT 3.29 3.35 3.43 3.77 ;
      RECT 3.29 3.35 3.73 3.58 ;
      RECT 3.47 3.26 3.73 3.58 ;
      RECT 2.79 2.42 3.19 2.93 ;
      RECT 2.98 2.395 3.26 2.765 ;
      RECT 2.73 2.42 3.26 2.74 ;
      RECT 72.13 7.055 72.5 7.425 ;
      RECT 70.84 2.395 71.12 2.765 ;
      RECT 69 2.395 69.28 2.765 ;
      RECT 65.84 2.955 66.12 3.325 ;
      RECT 55.805 7.055 56.175 7.425 ;
      RECT 54.515 2.395 54.795 2.765 ;
      RECT 52.675 2.395 52.955 2.765 ;
      RECT 49.515 2.955 49.795 3.325 ;
      RECT 39.48 7.055 39.85 7.425 ;
      RECT 38.19 2.395 38.47 2.765 ;
      RECT 36.35 2.395 36.63 2.765 ;
      RECT 33.19 2.955 33.47 3.325 ;
      RECT 23.155 7.055 23.525 7.425 ;
      RECT 21.865 2.395 22.145 2.765 ;
      RECT 20.025 2.395 20.305 2.765 ;
      RECT 16.865 2.955 17.145 3.325 ;
      RECT 6.83 7.055 7.2 7.425 ;
      RECT 5.54 2.395 5.82 2.765 ;
      RECT 3.7 2.395 3.98 2.765 ;
      RECT 0.54 2.955 0.82 3.325 ;
    LAYER via1 ;
      RECT 80.68 7.375 80.83 7.525 ;
      RECT 78.31 6.74 78.46 6.89 ;
      RECT 78.295 2.065 78.445 2.215 ;
      RECT 77.505 2.45 77.655 2.6 ;
      RECT 77.505 6.325 77.655 6.475 ;
      RECT 76.48 2.805 76.63 2.955 ;
      RECT 76.47 5.94 76.62 6.09 ;
      RECT 75.9 1.56 76.05 1.71 ;
      RECT 74.665 2.225 74.815 2.375 ;
      RECT 74.545 2.785 74.695 2.935 ;
      RECT 73.345 2.505 73.495 2.655 ;
      RECT 73.225 3.345 73.375 3.495 ;
      RECT 72.965 1.945 73.115 2.095 ;
      RECT 72.885 6.71 73.035 6.86 ;
      RECT 72.24 7.165 72.39 7.315 ;
      RECT 71.505 2.505 71.655 2.655 ;
      RECT 70.905 2.505 71.055 2.655 ;
      RECT 70.525 1.945 70.675 2.095 ;
      RECT 69.905 2.785 70.055 2.935 ;
      RECT 69.665 3.345 69.815 3.495 ;
      RECT 69.545 2.225 69.695 2.375 ;
      RECT 69.065 2.505 69.215 2.655 ;
      RECT 68.825 3.345 68.975 3.495 ;
      RECT 68.085 2.505 68.235 2.655 ;
      RECT 67.345 1.945 67.495 2.095 ;
      RECT 67.105 3.625 67.255 3.775 ;
      RECT 66.865 2.505 67.015 2.655 ;
      RECT 66.865 3.065 67.015 3.215 ;
      RECT 65.905 3.065 66.055 3.215 ;
      RECT 64.33 6.755 64.48 6.905 ;
      RECT 61.985 6.74 62.135 6.89 ;
      RECT 61.97 2.065 62.12 2.215 ;
      RECT 61.18 2.45 61.33 2.6 ;
      RECT 61.18 6.325 61.33 6.475 ;
      RECT 60.155 2.805 60.305 2.955 ;
      RECT 60.145 5.94 60.295 6.09 ;
      RECT 59.575 1.56 59.725 1.71 ;
      RECT 58.34 2.225 58.49 2.375 ;
      RECT 58.22 2.785 58.37 2.935 ;
      RECT 57.02 2.505 57.17 2.655 ;
      RECT 56.9 3.345 57.05 3.495 ;
      RECT 56.64 1.945 56.79 2.095 ;
      RECT 56.555 6.71 56.705 6.86 ;
      RECT 55.915 7.165 56.065 7.315 ;
      RECT 55.18 2.505 55.33 2.655 ;
      RECT 54.58 2.505 54.73 2.655 ;
      RECT 54.2 1.945 54.35 2.095 ;
      RECT 53.58 2.785 53.73 2.935 ;
      RECT 53.34 3.345 53.49 3.495 ;
      RECT 53.22 2.225 53.37 2.375 ;
      RECT 52.74 2.505 52.89 2.655 ;
      RECT 52.5 3.345 52.65 3.495 ;
      RECT 51.76 2.505 51.91 2.655 ;
      RECT 51.02 1.945 51.17 2.095 ;
      RECT 50.78 3.625 50.93 3.775 ;
      RECT 50.54 2.505 50.69 2.655 ;
      RECT 50.54 3.065 50.69 3.215 ;
      RECT 49.58 3.065 49.73 3.215 ;
      RECT 48.005 6.755 48.155 6.905 ;
      RECT 45.66 6.74 45.81 6.89 ;
      RECT 45.645 2.065 45.795 2.215 ;
      RECT 44.855 2.45 45.005 2.6 ;
      RECT 44.855 6.325 45.005 6.475 ;
      RECT 43.83 2.805 43.98 2.955 ;
      RECT 43.82 5.94 43.97 6.09 ;
      RECT 43.25 1.56 43.4 1.71 ;
      RECT 42.015 2.225 42.165 2.375 ;
      RECT 41.895 2.785 42.045 2.935 ;
      RECT 40.695 2.505 40.845 2.655 ;
      RECT 40.575 3.345 40.725 3.495 ;
      RECT 40.315 1.945 40.465 2.095 ;
      RECT 40.23 6.715 40.38 6.865 ;
      RECT 39.59 7.165 39.74 7.315 ;
      RECT 38.855 2.505 39.005 2.655 ;
      RECT 38.255 2.505 38.405 2.655 ;
      RECT 37.875 1.945 38.025 2.095 ;
      RECT 37.255 2.785 37.405 2.935 ;
      RECT 37.015 3.345 37.165 3.495 ;
      RECT 36.895 2.225 37.045 2.375 ;
      RECT 36.415 2.505 36.565 2.655 ;
      RECT 36.175 3.345 36.325 3.495 ;
      RECT 35.435 2.505 35.585 2.655 ;
      RECT 34.695 1.945 34.845 2.095 ;
      RECT 34.455 3.625 34.605 3.775 ;
      RECT 34.215 2.505 34.365 2.655 ;
      RECT 34.215 3.065 34.365 3.215 ;
      RECT 33.255 3.065 33.405 3.215 ;
      RECT 31.725 6.76 31.875 6.91 ;
      RECT 29.335 6.74 29.485 6.89 ;
      RECT 29.32 2.065 29.47 2.215 ;
      RECT 28.53 2.45 28.68 2.6 ;
      RECT 28.53 6.325 28.68 6.475 ;
      RECT 27.505 2.805 27.655 2.955 ;
      RECT 27.495 5.94 27.645 6.09 ;
      RECT 26.925 1.56 27.075 1.71 ;
      RECT 25.69 2.225 25.84 2.375 ;
      RECT 25.57 2.785 25.72 2.935 ;
      RECT 24.37 2.505 24.52 2.655 ;
      RECT 24.25 3.345 24.4 3.495 ;
      RECT 23.99 1.945 24.14 2.095 ;
      RECT 23.905 6.71 24.055 6.86 ;
      RECT 23.265 7.165 23.415 7.315 ;
      RECT 22.53 2.505 22.68 2.655 ;
      RECT 21.93 2.505 22.08 2.655 ;
      RECT 21.55 1.945 21.7 2.095 ;
      RECT 20.93 2.785 21.08 2.935 ;
      RECT 20.69 3.345 20.84 3.495 ;
      RECT 20.57 2.225 20.72 2.375 ;
      RECT 20.09 2.505 20.24 2.655 ;
      RECT 19.85 3.345 20 3.495 ;
      RECT 19.11 2.505 19.26 2.655 ;
      RECT 18.37 1.945 18.52 2.095 ;
      RECT 18.13 3.625 18.28 3.775 ;
      RECT 17.89 2.505 18.04 2.655 ;
      RECT 17.89 3.065 18.04 3.215 ;
      RECT 16.93 3.065 17.08 3.215 ;
      RECT 15.4 6.755 15.55 6.905 ;
      RECT 13.01 6.74 13.16 6.89 ;
      RECT 12.995 2.065 13.145 2.215 ;
      RECT 12.205 2.45 12.355 2.6 ;
      RECT 12.205 6.325 12.355 6.475 ;
      RECT 11.18 2.805 11.33 2.955 ;
      RECT 11.17 5.94 11.32 6.09 ;
      RECT 10.6 1.56 10.75 1.71 ;
      RECT 9.365 2.225 9.515 2.375 ;
      RECT 9.245 2.785 9.395 2.935 ;
      RECT 8.415 6.705 8.565 6.855 ;
      RECT 8.045 2.505 8.195 2.655 ;
      RECT 7.925 3.345 8.075 3.495 ;
      RECT 7.665 1.945 7.815 2.095 ;
      RECT 6.94 7.165 7.09 7.315 ;
      RECT 6.205 2.505 6.355 2.655 ;
      RECT 5.605 2.505 5.755 2.655 ;
      RECT 5.225 1.945 5.375 2.095 ;
      RECT 4.605 2.785 4.755 2.935 ;
      RECT 4.365 3.345 4.515 3.495 ;
      RECT 4.245 2.225 4.395 2.375 ;
      RECT 3.765 2.505 3.915 2.655 ;
      RECT 3.525 3.345 3.675 3.495 ;
      RECT 2.785 2.505 2.935 2.655 ;
      RECT 2.045 1.945 2.195 2.095 ;
      RECT 1.805 3.625 1.955 3.775 ;
      RECT 1.565 2.505 1.715 2.655 ;
      RECT 1.565 3.065 1.715 3.215 ;
      RECT 0.605 3.065 0.755 3.215 ;
      RECT -1.66 7.095 -1.51 7.245 ;
      RECT -2.035 6.355 -1.885 6.505 ;
    LAYER met1 ;
      RECT 72.97 2.93 74.57 3.07 ;
      RECT 56.645 2.93 58.245 3.07 ;
      RECT 40.32 2.93 41.92 3.07 ;
      RECT 23.995 2.93 25.595 3.07 ;
      RECT 7.67 2.93 9.27 3.07 ;
      RECT 72.97 2.93 74.735 3.055 ;
      RECT 56.645 2.93 58.41 3.055 ;
      RECT 40.32 2.93 42.085 3.055 ;
      RECT 23.995 2.93 25.76 3.055 ;
      RECT 7.67 2.93 9.435 3.055 ;
      RECT 74.46 2.73 74.78 2.99 ;
      RECT 58.135 2.73 58.455 2.99 ;
      RECT 41.81 2.73 42.13 2.99 ;
      RECT 25.485 2.73 25.805 2.99 ;
      RECT 9.16 2.73 9.48 2.99 ;
      RECT 74.46 2.745 74.885 2.975 ;
      RECT 58.135 2.745 58.56 2.975 ;
      RECT 41.81 2.745 42.235 2.975 ;
      RECT 25.485 2.745 25.91 2.975 ;
      RECT 9.16 2.745 9.585 2.975 ;
      RECT 75.195 0 75.38 2.945 ;
      RECT 58.87 0 59.055 2.945 ;
      RECT 42.545 0 42.73 2.945 ;
      RECT 26.22 0 26.405 2.945 ;
      RECT 9.895 0 10.08 2.945 ;
      RECT 74.43 2.79 75.38 2.945 ;
      RECT 74.46 2.76 75.38 2.945 ;
      RECT 72.635 2.79 73.11 2.975 ;
      RECT 58.105 2.79 59.055 2.945 ;
      RECT 58.135 2.76 59.055 2.945 ;
      RECT 56.31 2.79 56.785 2.975 ;
      RECT 41.78 2.79 42.73 2.945 ;
      RECT 41.81 2.76 42.73 2.945 ;
      RECT 39.985 2.79 40.46 2.975 ;
      RECT 25.455 2.79 26.405 2.945 ;
      RECT 25.485 2.76 26.405 2.945 ;
      RECT 23.66 2.79 24.135 2.975 ;
      RECT 9.13 2.79 10.08 2.945 ;
      RECT 9.16 2.76 10.08 2.945 ;
      RECT 7.335 2.79 7.81 2.975 ;
      RECT 72.635 2.745 72.925 2.975 ;
      RECT 56.31 2.745 56.6 2.975 ;
      RECT 39.985 2.745 40.275 2.975 ;
      RECT 23.66 2.745 23.95 2.975 ;
      RECT 7.335 2.745 7.625 2.975 ;
      RECT 65.565 0 75.38 1.74 ;
      RECT 49.24 0 59.055 1.74 ;
      RECT 32.915 0 42.73 1.74 ;
      RECT 16.59 0 26.405 1.74 ;
      RECT 0.265 0 10.08 1.74 ;
      RECT -3.225 0 81.15 0.305 ;
      RECT -3.225 4.135 81.15 4.745 ;
      RECT 65.565 3.98 75.225 4.745 ;
      RECT 49.24 3.98 58.9 4.745 ;
      RECT 32.915 3.98 42.575 4.745 ;
      RECT 16.59 3.98 26.25 4.745 ;
      RECT 0.265 3.98 9.925 4.745 ;
      RECT -3.225 8.575 81.15 8.88 ;
      RECT 71.4 6.315 71.575 8.88 ;
      RECT 55.075 6.315 55.25 8.88 ;
      RECT 38.75 6.315 38.925 8.88 ;
      RECT 22.425 6.315 22.6 8.88 ;
      RECT 6.1 6.315 6.275 8.88 ;
      RECT 71.775 6.285 72.065 6.515 ;
      RECT 55.45 6.285 55.74 6.515 ;
      RECT 39.125 6.285 39.415 6.515 ;
      RECT 22.8 6.285 23.09 6.515 ;
      RECT 6.475 6.285 6.765 6.515 ;
      RECT 71.4 6.315 72.065 6.485 ;
      RECT 55.075 6.315 55.74 6.485 ;
      RECT 38.75 6.315 39.415 6.485 ;
      RECT 22.425 6.315 23.09 6.485 ;
      RECT 6.1 6.315 6.765 6.485 ;
      RECT 80.55 7.765 80.84 7.995 ;
      RECT 80.61 6.285 80.78 7.995 ;
      RECT 80.58 7.275 80.93 7.625 ;
      RECT 80.55 6.285 80.84 6.515 ;
      RECT 80.55 2.365 80.84 2.595 ;
      RECT 80.61 0.885 80.78 2.595 ;
      RECT 80.55 0.885 80.84 1.115 ;
      RECT 80.14 2.735 80.47 2.965 ;
      RECT 80.14 2.765 80.64 2.935 ;
      RECT 80.14 2.395 80.33 2.965 ;
      RECT 79.56 2.365 79.85 2.595 ;
      RECT 79.56 2.395 80.33 2.565 ;
      RECT 79.62 0.885 79.79 2.595 ;
      RECT 79.56 0.885 79.85 1.115 ;
      RECT 79.56 7.765 79.85 7.995 ;
      RECT 79.62 6.285 79.79 7.995 ;
      RECT 79.56 6.285 79.85 6.515 ;
      RECT 79.56 6.325 80.41 6.485 ;
      RECT 80.24 5.915 80.41 6.485 ;
      RECT 79.56 6.32 79.95 6.485 ;
      RECT 80.18 5.915 80.47 6.145 ;
      RECT 80.18 5.945 80.64 6.115 ;
      RECT 79.19 2.735 79.48 2.965 ;
      RECT 79.19 2.765 79.65 2.935 ;
      RECT 79.25 1.655 79.415 2.965 ;
      RECT 77.765 1.625 78.055 1.855 ;
      RECT 77.765 1.655 79.415 1.825 ;
      RECT 77.825 0.885 77.995 1.855 ;
      RECT 77.765 0.885 78.055 1.115 ;
      RECT 77.765 7.765 78.055 7.995 ;
      RECT 77.825 7.025 77.995 7.995 ;
      RECT 77.825 7.12 79.415 7.29 ;
      RECT 79.245 5.915 79.415 7.29 ;
      RECT 77.765 7.025 78.055 7.255 ;
      RECT 79.19 5.915 79.48 6.145 ;
      RECT 79.19 5.945 79.65 6.115 ;
      RECT 78.195 1.965 78.545 2.315 ;
      RECT 75.89 2.025 78.545 2.195 ;
      RECT 75.89 1.46 76.06 2.195 ;
      RECT 75.8 1.46 76.14 1.81 ;
      RECT 78.22 6.655 78.545 6.98 ;
      RECT 72.785 6.61 73.135 6.96 ;
      RECT 78.195 6.655 78.545 6.885 ;
      RECT 72.58 6.655 73.135 6.885 ;
      RECT 72.41 6.685 78.545 6.855 ;
      RECT 77.42 2.365 77.74 2.685 ;
      RECT 77.39 2.365 77.74 2.595 ;
      RECT 77.22 2.395 77.74 2.565 ;
      RECT 77.42 6.255 77.74 6.545 ;
      RECT 77.39 6.285 77.74 6.515 ;
      RECT 77.22 6.315 77.74 6.485 ;
      RECT 76.38 2.705 76.72 3.055 ;
      RECT 76.38 2.765 76.855 2.935 ;
      RECT 76.37 5.84 76.71 6.19 ;
      RECT 70.78 5.915 71.07 6.145 ;
      RECT 70.78 5.945 76.855 6.115 ;
      RECT 73.875 2.465 74.165 2.695 ;
      RECT 73.875 2.465 74.33 2.65 ;
      RECT 74.19 2.37 74.81 2.51 ;
      RECT 74.58 2.17 74.9 2.43 ;
      RECT 73.26 2.45 73.58 2.71 ;
      RECT 73.26 2.45 73.725 2.695 ;
      RECT 73.585 2.07 73.725 2.695 ;
      RECT 73.585 2.07 73.85 2.21 ;
      RECT 74.115 1.905 74.405 2.135 ;
      RECT 73.71 1.95 74.405 2.09 ;
      RECT 73.155 3.29 73.445 3.815 ;
      RECT 73.14 3.29 73.46 3.55 ;
      RECT 72.88 1.89 73.2 2.15 ;
      RECT 72.88 1.905 73.445 2.135 ;
      RECT 72.155 3.585 72.445 3.815 ;
      RECT 72.35 2.23 72.49 3.77 ;
      RECT 72.395 2.185 72.685 2.415 ;
      RECT 71.99 2.23 72.685 2.37 ;
      RECT 71.99 2.07 72.13 2.37 ;
      RECT 70.53 2.07 72.13 2.21 ;
      RECT 70.44 1.89 70.76 2.15 ;
      RECT 70.44 1.905 71.005 2.15 ;
      RECT 72.15 7.765 72.44 7.995 ;
      RECT 72.21 7.025 72.38 7.995 ;
      RECT 72.13 7.075 72.5 7.425 ;
      RECT 72.13 7.055 72.44 7.425 ;
      RECT 72.15 7.025 72.44 7.425 ;
      RECT 69.55 2.93 72.13 3.07 ;
      RECT 71.915 2.745 72.205 2.975 ;
      RECT 69.475 2.745 70.14 2.975 ;
      RECT 69.82 2.73 70.14 3.07 ;
      RECT 70.82 2.45 71.14 2.71 ;
      RECT 70.82 2.465 71.245 2.695 ;
      RECT 69.46 2.17 69.78 2.43 ;
      RECT 69.955 2.185 70.245 2.415 ;
      RECT 69.46 2.23 70.245 2.37 ;
      RECT 69.58 3.29 69.9 3.55 ;
      RECT 68.74 3.29 69.06 3.55 ;
      RECT 69.58 3.305 70.005 3.535 ;
      RECT 68.74 3.35 70.005 3.49 ;
      RECT 68.275 3.025 68.565 3.255 ;
      RECT 68.35 1.95 68.49 3.255 ;
      RECT 68 2.45 68.49 2.71 ;
      RECT 67.755 2.465 68.49 2.695 ;
      RECT 68.755 1.905 69.045 2.135 ;
      RECT 68.35 1.95 69.045 2.09 ;
      RECT 67.515 3.305 67.805 3.535 ;
      RECT 67.515 3.305 67.97 3.49 ;
      RECT 67.83 2.93 67.97 3.49 ;
      RECT 67.47 2.93 67.97 3.07 ;
      RECT 67.47 1.95 67.61 3.07 ;
      RECT 67.26 1.89 67.58 2.15 ;
      RECT 67.02 3.57 67.34 3.83 ;
      RECT 66.315 3.585 66.605 3.815 ;
      RECT 66.315 3.63 67.34 3.77 ;
      RECT 66.39 3.58 66.65 3.77 ;
      RECT 66.78 2.45 67.1 2.71 ;
      RECT 66.78 2.465 67.325 2.695 ;
      RECT 66.78 3.01 67.1 3.27 ;
      RECT 66.78 3.025 67.325 3.255 ;
      RECT 65.82 3.01 66.14 3.27 ;
      RECT 65.91 1.95 66.05 3.27 ;
      RECT 66.315 1.905 66.605 2.135 ;
      RECT 65.91 1.95 66.605 2.09 ;
      RECT 64.225 7.765 64.515 7.995 ;
      RECT 64.285 6.285 64.455 7.995 ;
      RECT 64.23 6.655 64.58 7.005 ;
      RECT 64.225 6.285 64.515 6.515 ;
      RECT 64.225 2.365 64.515 2.595 ;
      RECT 64.285 0.885 64.455 2.595 ;
      RECT 64.225 0.885 64.515 1.115 ;
      RECT 63.815 2.735 64.145 2.965 ;
      RECT 63.815 2.765 64.315 2.935 ;
      RECT 63.815 2.395 64.005 2.965 ;
      RECT 63.235 2.365 63.525 2.595 ;
      RECT 63.235 2.395 64.005 2.565 ;
      RECT 63.295 0.885 63.465 2.595 ;
      RECT 63.235 0.885 63.525 1.115 ;
      RECT 63.235 7.765 63.525 7.995 ;
      RECT 63.295 6.285 63.465 7.995 ;
      RECT 63.235 6.285 63.525 6.515 ;
      RECT 63.235 6.325 64.085 6.485 ;
      RECT 63.915 5.915 64.085 6.485 ;
      RECT 63.235 6.32 63.625 6.485 ;
      RECT 63.855 5.915 64.145 6.145 ;
      RECT 63.855 5.945 64.315 6.115 ;
      RECT 62.865 2.735 63.155 2.965 ;
      RECT 62.865 2.765 63.325 2.935 ;
      RECT 62.925 1.655 63.09 2.965 ;
      RECT 61.44 1.625 61.73 1.855 ;
      RECT 61.44 1.655 63.09 1.825 ;
      RECT 61.5 0.885 61.67 1.855 ;
      RECT 61.44 0.885 61.73 1.115 ;
      RECT 61.44 7.765 61.73 7.995 ;
      RECT 61.5 7.025 61.67 7.995 ;
      RECT 61.5 7.12 63.09 7.29 ;
      RECT 62.92 5.915 63.09 7.29 ;
      RECT 61.44 7.025 61.73 7.255 ;
      RECT 62.865 5.915 63.155 6.145 ;
      RECT 62.865 5.945 63.325 6.115 ;
      RECT 61.87 1.965 62.22 2.315 ;
      RECT 59.565 2.025 62.22 2.195 ;
      RECT 59.565 1.46 59.735 2.195 ;
      RECT 59.475 1.46 59.815 1.81 ;
      RECT 61.895 6.655 62.22 6.98 ;
      RECT 56.455 6.61 56.805 6.96 ;
      RECT 61.87 6.655 62.22 6.885 ;
      RECT 56.255 6.655 56.805 6.885 ;
      RECT 56.085 6.685 62.22 6.855 ;
      RECT 61.095 2.365 61.415 2.685 ;
      RECT 61.065 2.365 61.415 2.595 ;
      RECT 60.895 2.395 61.415 2.565 ;
      RECT 61.095 6.255 61.415 6.545 ;
      RECT 61.065 6.285 61.415 6.515 ;
      RECT 60.895 6.315 61.415 6.485 ;
      RECT 60.055 2.705 60.395 3.055 ;
      RECT 60.055 2.765 60.53 2.935 ;
      RECT 60.045 5.84 60.385 6.19 ;
      RECT 54.455 5.915 54.745 6.145 ;
      RECT 54.455 5.945 60.53 6.115 ;
      RECT 57.55 2.465 57.84 2.695 ;
      RECT 57.55 2.465 58.005 2.65 ;
      RECT 57.865 2.37 58.485 2.51 ;
      RECT 58.255 2.17 58.575 2.43 ;
      RECT 56.935 2.45 57.255 2.71 ;
      RECT 56.935 2.45 57.4 2.695 ;
      RECT 57.26 2.07 57.4 2.695 ;
      RECT 57.26 2.07 57.525 2.21 ;
      RECT 57.79 1.905 58.08 2.135 ;
      RECT 57.385 1.95 58.08 2.09 ;
      RECT 56.83 3.29 57.12 3.815 ;
      RECT 56.815 3.29 57.135 3.55 ;
      RECT 56.555 1.89 56.875 2.15 ;
      RECT 56.555 1.905 57.12 2.135 ;
      RECT 55.83 3.585 56.12 3.815 ;
      RECT 56.025 2.23 56.165 3.77 ;
      RECT 56.07 2.185 56.36 2.415 ;
      RECT 55.665 2.23 56.36 2.37 ;
      RECT 55.665 2.07 55.805 2.37 ;
      RECT 54.205 2.07 55.805 2.21 ;
      RECT 54.115 1.89 54.435 2.15 ;
      RECT 54.115 1.905 54.68 2.15 ;
      RECT 55.825 7.765 56.115 7.995 ;
      RECT 55.885 7.025 56.055 7.995 ;
      RECT 55.805 7.075 56.175 7.425 ;
      RECT 55.805 7.055 56.115 7.425 ;
      RECT 55.825 7.025 56.115 7.425 ;
      RECT 53.225 2.93 55.805 3.07 ;
      RECT 55.59 2.745 55.88 2.975 ;
      RECT 53.15 2.745 53.815 2.975 ;
      RECT 53.495 2.73 53.815 3.07 ;
      RECT 54.495 2.45 54.815 2.71 ;
      RECT 54.495 2.465 54.92 2.695 ;
      RECT 53.135 2.17 53.455 2.43 ;
      RECT 53.63 2.185 53.92 2.415 ;
      RECT 53.135 2.23 53.92 2.37 ;
      RECT 53.255 3.29 53.575 3.55 ;
      RECT 52.415 3.29 52.735 3.55 ;
      RECT 53.255 3.305 53.68 3.535 ;
      RECT 52.415 3.35 53.68 3.49 ;
      RECT 51.95 3.025 52.24 3.255 ;
      RECT 52.025 1.95 52.165 3.255 ;
      RECT 51.675 2.45 52.165 2.71 ;
      RECT 51.43 2.465 52.165 2.695 ;
      RECT 52.43 1.905 52.72 2.135 ;
      RECT 52.025 1.95 52.72 2.09 ;
      RECT 51.19 3.305 51.48 3.535 ;
      RECT 51.19 3.305 51.645 3.49 ;
      RECT 51.505 2.93 51.645 3.49 ;
      RECT 51.145 2.93 51.645 3.07 ;
      RECT 51.145 1.95 51.285 3.07 ;
      RECT 50.935 1.89 51.255 2.15 ;
      RECT 50.695 3.57 51.015 3.83 ;
      RECT 49.99 3.585 50.28 3.815 ;
      RECT 49.99 3.63 51.015 3.77 ;
      RECT 50.065 3.58 50.325 3.77 ;
      RECT 50.455 2.45 50.775 2.71 ;
      RECT 50.455 2.465 51 2.695 ;
      RECT 50.455 3.01 50.775 3.27 ;
      RECT 50.455 3.025 51 3.255 ;
      RECT 49.495 3.01 49.815 3.27 ;
      RECT 49.585 1.95 49.725 3.27 ;
      RECT 49.99 1.905 50.28 2.135 ;
      RECT 49.585 1.95 50.28 2.09 ;
      RECT 47.9 7.765 48.19 7.995 ;
      RECT 47.96 6.285 48.13 7.995 ;
      RECT 47.905 6.655 48.255 7.005 ;
      RECT 47.9 6.285 48.19 6.515 ;
      RECT 47.9 2.365 48.19 2.595 ;
      RECT 47.96 0.885 48.13 2.595 ;
      RECT 47.9 0.885 48.19 1.115 ;
      RECT 47.49 2.735 47.82 2.965 ;
      RECT 47.49 2.765 47.99 2.935 ;
      RECT 47.49 2.395 47.68 2.965 ;
      RECT 46.91 2.365 47.2 2.595 ;
      RECT 46.91 2.395 47.68 2.565 ;
      RECT 46.97 0.885 47.14 2.595 ;
      RECT 46.91 0.885 47.2 1.115 ;
      RECT 46.91 7.765 47.2 7.995 ;
      RECT 46.97 6.285 47.14 7.995 ;
      RECT 46.91 6.285 47.2 6.515 ;
      RECT 46.91 6.325 47.76 6.485 ;
      RECT 47.59 5.915 47.76 6.485 ;
      RECT 46.91 6.32 47.3 6.485 ;
      RECT 47.53 5.915 47.82 6.145 ;
      RECT 47.53 5.945 47.99 6.115 ;
      RECT 46.54 2.735 46.83 2.965 ;
      RECT 46.54 2.765 47 2.935 ;
      RECT 46.6 1.655 46.765 2.965 ;
      RECT 45.115 1.625 45.405 1.855 ;
      RECT 45.115 1.655 46.765 1.825 ;
      RECT 45.175 0.885 45.345 1.855 ;
      RECT 45.115 0.885 45.405 1.115 ;
      RECT 45.115 7.765 45.405 7.995 ;
      RECT 45.175 7.025 45.345 7.995 ;
      RECT 45.175 7.12 46.765 7.29 ;
      RECT 46.595 5.915 46.765 7.29 ;
      RECT 45.115 7.025 45.405 7.255 ;
      RECT 46.54 5.915 46.83 6.145 ;
      RECT 46.54 5.945 47 6.115 ;
      RECT 45.545 1.965 45.895 2.315 ;
      RECT 43.24 2.025 45.895 2.195 ;
      RECT 43.24 1.46 43.41 2.195 ;
      RECT 43.15 1.46 43.49 1.81 ;
      RECT 45.57 6.655 45.895 6.98 ;
      RECT 40.13 6.615 40.48 6.965 ;
      RECT 45.545 6.655 45.895 6.885 ;
      RECT 39.93 6.655 40.48 6.885 ;
      RECT 39.76 6.685 45.895 6.855 ;
      RECT 44.77 2.365 45.09 2.685 ;
      RECT 44.74 2.365 45.09 2.595 ;
      RECT 44.57 2.395 45.09 2.565 ;
      RECT 44.77 6.255 45.09 6.545 ;
      RECT 44.74 6.285 45.09 6.515 ;
      RECT 44.57 6.315 45.09 6.485 ;
      RECT 43.73 2.705 44.07 3.055 ;
      RECT 43.73 2.765 44.205 2.935 ;
      RECT 43.72 5.84 44.06 6.19 ;
      RECT 38.13 5.915 38.42 6.145 ;
      RECT 38.13 5.945 44.205 6.115 ;
      RECT 41.225 2.465 41.515 2.695 ;
      RECT 41.225 2.465 41.68 2.65 ;
      RECT 41.54 2.37 42.16 2.51 ;
      RECT 41.93 2.17 42.25 2.43 ;
      RECT 40.61 2.45 40.93 2.71 ;
      RECT 40.61 2.45 41.075 2.695 ;
      RECT 40.935 2.07 41.075 2.695 ;
      RECT 40.935 2.07 41.2 2.21 ;
      RECT 41.465 1.905 41.755 2.135 ;
      RECT 41.06 1.95 41.755 2.09 ;
      RECT 40.505 3.29 40.795 3.815 ;
      RECT 40.49 3.29 40.81 3.55 ;
      RECT 40.23 1.89 40.55 2.15 ;
      RECT 40.23 1.905 40.795 2.135 ;
      RECT 39.505 3.585 39.795 3.815 ;
      RECT 39.7 2.23 39.84 3.77 ;
      RECT 39.745 2.185 40.035 2.415 ;
      RECT 39.34 2.23 40.035 2.37 ;
      RECT 39.34 2.07 39.48 2.37 ;
      RECT 37.88 2.07 39.48 2.21 ;
      RECT 37.79 1.89 38.11 2.15 ;
      RECT 37.79 1.905 38.355 2.15 ;
      RECT 39.5 7.765 39.79 7.995 ;
      RECT 39.56 7.025 39.73 7.995 ;
      RECT 39.48 7.075 39.85 7.425 ;
      RECT 39.48 7.055 39.79 7.425 ;
      RECT 39.5 7.025 39.79 7.425 ;
      RECT 36.9 2.93 39.48 3.07 ;
      RECT 39.265 2.745 39.555 2.975 ;
      RECT 36.825 2.745 37.49 2.975 ;
      RECT 37.17 2.73 37.49 3.07 ;
      RECT 38.17 2.45 38.49 2.71 ;
      RECT 38.17 2.465 38.595 2.695 ;
      RECT 36.81 2.17 37.13 2.43 ;
      RECT 37.305 2.185 37.595 2.415 ;
      RECT 36.81 2.23 37.595 2.37 ;
      RECT 36.93 3.29 37.25 3.55 ;
      RECT 36.09 3.29 36.41 3.55 ;
      RECT 36.93 3.305 37.355 3.535 ;
      RECT 36.09 3.35 37.355 3.49 ;
      RECT 35.625 3.025 35.915 3.255 ;
      RECT 35.7 1.95 35.84 3.255 ;
      RECT 35.35 2.45 35.84 2.71 ;
      RECT 35.105 2.465 35.84 2.695 ;
      RECT 36.105 1.905 36.395 2.135 ;
      RECT 35.7 1.95 36.395 2.09 ;
      RECT 34.865 3.305 35.155 3.535 ;
      RECT 34.865 3.305 35.32 3.49 ;
      RECT 35.18 2.93 35.32 3.49 ;
      RECT 34.82 2.93 35.32 3.07 ;
      RECT 34.82 1.95 34.96 3.07 ;
      RECT 34.61 1.89 34.93 2.15 ;
      RECT 34.37 3.57 34.69 3.83 ;
      RECT 33.665 3.585 33.955 3.815 ;
      RECT 33.665 3.63 34.69 3.77 ;
      RECT 33.74 3.58 34 3.77 ;
      RECT 34.13 2.45 34.45 2.71 ;
      RECT 34.13 2.465 34.675 2.695 ;
      RECT 34.13 3.01 34.45 3.27 ;
      RECT 34.13 3.025 34.675 3.255 ;
      RECT 33.17 3.01 33.49 3.27 ;
      RECT 33.26 1.95 33.4 3.27 ;
      RECT 33.665 1.905 33.955 2.135 ;
      RECT 33.26 1.95 33.955 2.09 ;
      RECT 31.575 7.765 31.865 7.995 ;
      RECT 31.635 6.285 31.805 7.995 ;
      RECT 31.62 6.66 31.975 7.015 ;
      RECT 31.575 6.285 31.865 6.515 ;
      RECT 31.575 2.365 31.865 2.595 ;
      RECT 31.635 0.885 31.805 2.595 ;
      RECT 31.575 0.885 31.865 1.115 ;
      RECT 31.165 2.735 31.495 2.965 ;
      RECT 31.165 2.765 31.665 2.935 ;
      RECT 31.165 2.395 31.355 2.965 ;
      RECT 30.585 2.365 30.875 2.595 ;
      RECT 30.585 2.395 31.355 2.565 ;
      RECT 30.645 0.885 30.815 2.595 ;
      RECT 30.585 0.885 30.875 1.115 ;
      RECT 30.585 7.765 30.875 7.995 ;
      RECT 30.645 6.285 30.815 7.995 ;
      RECT 30.585 6.285 30.875 6.515 ;
      RECT 30.585 6.325 31.435 6.485 ;
      RECT 31.265 5.915 31.435 6.485 ;
      RECT 30.585 6.32 30.975 6.485 ;
      RECT 31.205 5.915 31.495 6.145 ;
      RECT 31.205 5.945 31.665 6.115 ;
      RECT 30.215 2.735 30.505 2.965 ;
      RECT 30.215 2.765 30.675 2.935 ;
      RECT 30.275 1.655 30.44 2.965 ;
      RECT 28.79 1.625 29.08 1.855 ;
      RECT 28.79 1.655 30.44 1.825 ;
      RECT 28.85 0.885 29.02 1.855 ;
      RECT 28.79 0.885 29.08 1.115 ;
      RECT 28.79 7.765 29.08 7.995 ;
      RECT 28.85 7.025 29.02 7.995 ;
      RECT 28.85 7.12 30.44 7.29 ;
      RECT 30.27 5.915 30.44 7.29 ;
      RECT 28.79 7.025 29.08 7.255 ;
      RECT 30.215 5.915 30.505 6.145 ;
      RECT 30.215 5.945 30.675 6.115 ;
      RECT 29.22 1.965 29.57 2.315 ;
      RECT 26.915 2.025 29.57 2.195 ;
      RECT 26.915 1.46 27.085 2.195 ;
      RECT 26.825 1.46 27.165 1.81 ;
      RECT 29.245 6.655 29.57 6.98 ;
      RECT 23.805 6.61 24.155 6.96 ;
      RECT 29.22 6.655 29.57 6.885 ;
      RECT 23.605 6.655 24.155 6.885 ;
      RECT 23.435 6.685 29.57 6.855 ;
      RECT 28.445 2.365 28.765 2.685 ;
      RECT 28.415 2.365 28.765 2.595 ;
      RECT 28.245 2.395 28.765 2.565 ;
      RECT 28.445 6.255 28.765 6.545 ;
      RECT 28.415 6.285 28.765 6.515 ;
      RECT 28.245 6.315 28.765 6.485 ;
      RECT 27.405 2.705 27.745 3.055 ;
      RECT 27.405 2.765 27.88 2.935 ;
      RECT 27.395 5.84 27.735 6.19 ;
      RECT 21.805 5.915 22.095 6.145 ;
      RECT 21.805 5.945 27.88 6.115 ;
      RECT 24.9 2.465 25.19 2.695 ;
      RECT 24.9 2.465 25.355 2.65 ;
      RECT 25.215 2.37 25.835 2.51 ;
      RECT 25.605 2.17 25.925 2.43 ;
      RECT 24.285 2.45 24.605 2.71 ;
      RECT 24.285 2.45 24.75 2.695 ;
      RECT 24.61 2.07 24.75 2.695 ;
      RECT 24.61 2.07 24.875 2.21 ;
      RECT 25.14 1.905 25.43 2.135 ;
      RECT 24.735 1.95 25.43 2.09 ;
      RECT 24.18 3.29 24.47 3.815 ;
      RECT 24.165 3.29 24.485 3.55 ;
      RECT 23.905 1.89 24.225 2.15 ;
      RECT 23.905 1.905 24.47 2.135 ;
      RECT 23.18 3.585 23.47 3.815 ;
      RECT 23.375 2.23 23.515 3.77 ;
      RECT 23.42 2.185 23.71 2.415 ;
      RECT 23.015 2.23 23.71 2.37 ;
      RECT 23.015 2.07 23.155 2.37 ;
      RECT 21.555 2.07 23.155 2.21 ;
      RECT 21.465 1.89 21.785 2.15 ;
      RECT 21.465 1.905 22.03 2.15 ;
      RECT 23.175 7.765 23.465 7.995 ;
      RECT 23.235 7.025 23.405 7.995 ;
      RECT 23.155 7.075 23.525 7.425 ;
      RECT 23.155 7.055 23.465 7.425 ;
      RECT 23.175 7.025 23.465 7.425 ;
      RECT 20.575 2.93 23.155 3.07 ;
      RECT 22.94 2.745 23.23 2.975 ;
      RECT 20.5 2.745 21.165 2.975 ;
      RECT 20.845 2.73 21.165 3.07 ;
      RECT 21.845 2.45 22.165 2.71 ;
      RECT 21.845 2.465 22.27 2.695 ;
      RECT 20.485 2.17 20.805 2.43 ;
      RECT 20.98 2.185 21.27 2.415 ;
      RECT 20.485 2.23 21.27 2.37 ;
      RECT 20.605 3.29 20.925 3.55 ;
      RECT 19.765 3.29 20.085 3.55 ;
      RECT 20.605 3.305 21.03 3.535 ;
      RECT 19.765 3.35 21.03 3.49 ;
      RECT 19.3 3.025 19.59 3.255 ;
      RECT 19.375 1.95 19.515 3.255 ;
      RECT 19.025 2.45 19.515 2.71 ;
      RECT 18.78 2.465 19.515 2.695 ;
      RECT 19.78 1.905 20.07 2.135 ;
      RECT 19.375 1.95 20.07 2.09 ;
      RECT 18.54 3.305 18.83 3.535 ;
      RECT 18.54 3.305 18.995 3.49 ;
      RECT 18.855 2.93 18.995 3.49 ;
      RECT 18.495 2.93 18.995 3.07 ;
      RECT 18.495 1.95 18.635 3.07 ;
      RECT 18.285 1.89 18.605 2.15 ;
      RECT 18.045 3.57 18.365 3.83 ;
      RECT 17.34 3.585 17.63 3.815 ;
      RECT 17.34 3.63 18.365 3.77 ;
      RECT 17.415 3.58 17.675 3.77 ;
      RECT 17.805 2.45 18.125 2.71 ;
      RECT 17.805 2.465 18.35 2.695 ;
      RECT 17.805 3.01 18.125 3.27 ;
      RECT 17.805 3.025 18.35 3.255 ;
      RECT 16.845 3.01 17.165 3.27 ;
      RECT 16.935 1.95 17.075 3.27 ;
      RECT 17.34 1.905 17.63 2.135 ;
      RECT 16.935 1.95 17.63 2.09 ;
      RECT 15.25 7.765 15.54 7.995 ;
      RECT 15.31 6.285 15.48 7.995 ;
      RECT 15.3 6.655 15.65 7.005 ;
      RECT 15.25 6.285 15.54 6.515 ;
      RECT 15.25 2.365 15.54 2.595 ;
      RECT 15.31 0.885 15.48 2.595 ;
      RECT 15.25 0.885 15.54 1.115 ;
      RECT 14.84 2.735 15.17 2.965 ;
      RECT 14.84 2.765 15.34 2.935 ;
      RECT 14.84 2.395 15.03 2.965 ;
      RECT 14.26 2.365 14.55 2.595 ;
      RECT 14.26 2.395 15.03 2.565 ;
      RECT 14.32 0.885 14.49 2.595 ;
      RECT 14.26 0.885 14.55 1.115 ;
      RECT 14.26 7.765 14.55 7.995 ;
      RECT 14.32 6.285 14.49 7.995 ;
      RECT 14.26 6.285 14.55 6.515 ;
      RECT 14.26 6.325 15.11 6.485 ;
      RECT 14.94 5.915 15.11 6.485 ;
      RECT 14.26 6.32 14.65 6.485 ;
      RECT 14.88 5.915 15.17 6.145 ;
      RECT 14.88 5.945 15.34 6.115 ;
      RECT 13.89 2.735 14.18 2.965 ;
      RECT 13.89 2.765 14.35 2.935 ;
      RECT 13.95 1.655 14.115 2.965 ;
      RECT 12.465 1.625 12.755 1.855 ;
      RECT 12.465 1.655 14.115 1.825 ;
      RECT 12.525 0.885 12.695 1.855 ;
      RECT 12.465 0.885 12.755 1.115 ;
      RECT 12.465 7.765 12.755 7.995 ;
      RECT 12.525 7.025 12.695 7.995 ;
      RECT 12.525 7.12 14.115 7.29 ;
      RECT 13.945 5.915 14.115 7.29 ;
      RECT 12.465 7.025 12.755 7.255 ;
      RECT 13.89 5.915 14.18 6.145 ;
      RECT 13.89 5.945 14.35 6.115 ;
      RECT 12.895 1.965 13.245 2.315 ;
      RECT 10.59 2.025 13.245 2.195 ;
      RECT 10.59 1.46 10.76 2.195 ;
      RECT 10.5 1.46 10.84 1.81 ;
      RECT 12.92 6.655 13.245 6.98 ;
      RECT 8.315 6.605 8.665 6.955 ;
      RECT 12.895 6.655 13.245 6.885 ;
      RECT 7.28 6.655 7.57 6.885 ;
      RECT 7.11 6.685 13.245 6.855 ;
      RECT 12.12 2.365 12.44 2.685 ;
      RECT 12.09 2.365 12.44 2.595 ;
      RECT 11.92 2.395 12.44 2.565 ;
      RECT 12.12 6.255 12.44 6.545 ;
      RECT 12.09 6.285 12.44 6.515 ;
      RECT 11.92 6.315 12.44 6.485 ;
      RECT 11.08 2.705 11.42 3.055 ;
      RECT 11.08 2.765 11.555 2.935 ;
      RECT 11.07 5.84 11.41 6.19 ;
      RECT 5.48 5.915 5.77 6.145 ;
      RECT 5.48 5.945 11.555 6.115 ;
      RECT 8.575 2.465 8.865 2.695 ;
      RECT 8.575 2.465 9.03 2.65 ;
      RECT 8.89 2.37 9.51 2.51 ;
      RECT 9.28 2.17 9.6 2.43 ;
      RECT 7.96 2.45 8.28 2.71 ;
      RECT 7.96 2.45 8.425 2.695 ;
      RECT 8.285 2.07 8.425 2.695 ;
      RECT 8.285 2.07 8.55 2.21 ;
      RECT 8.815 1.905 9.105 2.135 ;
      RECT 8.41 1.95 9.105 2.09 ;
      RECT 7.855 3.29 8.145 3.815 ;
      RECT 7.84 3.29 8.16 3.55 ;
      RECT 7.58 1.89 7.9 2.15 ;
      RECT 7.58 1.905 8.145 2.135 ;
      RECT 6.855 3.585 7.145 3.815 ;
      RECT 7.05 2.23 7.19 3.77 ;
      RECT 7.095 2.185 7.385 2.415 ;
      RECT 6.69 2.23 7.385 2.37 ;
      RECT 6.69 2.07 6.83 2.37 ;
      RECT 5.23 2.07 6.83 2.21 ;
      RECT 5.14 1.89 5.46 2.15 ;
      RECT 5.14 1.905 5.705 2.15 ;
      RECT 6.85 7.765 7.14 7.995 ;
      RECT 6.91 7.025 7.08 7.995 ;
      RECT 6.83 7.075 7.2 7.425 ;
      RECT 6.83 7.055 7.14 7.425 ;
      RECT 6.85 7.025 7.14 7.425 ;
      RECT 4.25 2.93 6.83 3.07 ;
      RECT 6.615 2.745 6.905 2.975 ;
      RECT 4.175 2.745 4.84 2.975 ;
      RECT 4.52 2.73 4.84 3.07 ;
      RECT 5.52 2.45 5.84 2.71 ;
      RECT 5.52 2.465 5.945 2.695 ;
      RECT 4.16 2.17 4.48 2.43 ;
      RECT 4.655 2.185 4.945 2.415 ;
      RECT 4.16 2.23 4.945 2.37 ;
      RECT 4.28 3.29 4.6 3.55 ;
      RECT 3.44 3.29 3.76 3.55 ;
      RECT 4.28 3.305 4.705 3.535 ;
      RECT 3.44 3.35 4.705 3.49 ;
      RECT 2.975 3.025 3.265 3.255 ;
      RECT 3.05 1.95 3.19 3.255 ;
      RECT 2.7 2.45 3.19 2.71 ;
      RECT 2.455 2.465 3.19 2.695 ;
      RECT 3.455 1.905 3.745 2.135 ;
      RECT 3.05 1.95 3.745 2.09 ;
      RECT 2.215 3.305 2.505 3.535 ;
      RECT 2.215 3.305 2.67 3.49 ;
      RECT 2.53 2.93 2.67 3.49 ;
      RECT 2.17 2.93 2.67 3.07 ;
      RECT 2.17 1.95 2.31 3.07 ;
      RECT 1.96 1.89 2.28 2.15 ;
      RECT 1.72 3.57 2.04 3.83 ;
      RECT 1.015 3.585 1.305 3.815 ;
      RECT 1.015 3.63 2.04 3.77 ;
      RECT 1.09 3.58 1.35 3.77 ;
      RECT 1.48 2.45 1.8 2.71 ;
      RECT 1.48 2.465 2.025 2.695 ;
      RECT 1.48 3.01 1.8 3.27 ;
      RECT 1.48 3.025 2.025 3.255 ;
      RECT 0.52 3.01 0.84 3.27 ;
      RECT 0.61 1.95 0.75 3.27 ;
      RECT 1.015 1.905 1.305 2.135 ;
      RECT 0.61 1.95 1.305 2.09 ;
      RECT -1.3 6.655 -1.01 6.885 ;
      RECT -1.47 6.685 -1.01 6.855 ;
      RECT -1.73 7.765 -1.44 7.995 ;
      RECT -1.67 7.025 -1.5 7.995 ;
      RECT -1.76 7.025 -1.41 7.315 ;
      RECT -2.135 6.285 -1.785 6.575 ;
      RECT -2.275 6.315 -1.785 6.485 ;
      RECT -3.1 5.915 -2.81 6.145 ;
      RECT -3.1 5.945 -2.64 6.115 ;
      RECT 71.42 2.45 71.74 2.71 ;
      RECT 68.98 2.45 69.3 2.71 ;
      RECT 55.095 2.45 55.415 2.71 ;
      RECT 52.655 2.45 52.975 2.71 ;
      RECT 38.77 2.45 39.09 2.71 ;
      RECT 36.33 2.45 36.65 2.71 ;
      RECT 22.445 2.45 22.765 2.71 ;
      RECT 20.005 2.45 20.325 2.71 ;
      RECT 6.12 2.45 6.44 2.71 ;
      RECT 3.68 2.45 4 2.71 ;
    LAYER mcon ;
      RECT 80.61 0.915 80.78 1.085 ;
      RECT 80.61 2.395 80.78 2.565 ;
      RECT 80.61 6.315 80.78 6.485 ;
      RECT 80.61 7.795 80.78 7.965 ;
      RECT 80.26 0.105 80.43 0.275 ;
      RECT 80.26 4.165 80.43 4.335 ;
      RECT 80.26 4.545 80.43 4.715 ;
      RECT 80.26 8.605 80.43 8.775 ;
      RECT 80.24 2.765 80.41 2.935 ;
      RECT 80.24 5.945 80.41 6.115 ;
      RECT 79.62 0.915 79.79 1.085 ;
      RECT 79.62 2.395 79.79 2.565 ;
      RECT 79.62 6.315 79.79 6.485 ;
      RECT 79.62 7.795 79.79 7.965 ;
      RECT 79.27 0.105 79.44 0.275 ;
      RECT 79.27 4.165 79.44 4.335 ;
      RECT 79.27 4.545 79.44 4.715 ;
      RECT 79.27 8.605 79.44 8.775 ;
      RECT 79.25 2.765 79.42 2.935 ;
      RECT 79.25 5.945 79.42 6.115 ;
      RECT 78.565 0.105 78.735 0.275 ;
      RECT 78.565 4.165 78.735 4.335 ;
      RECT 78.565 4.545 78.735 4.715 ;
      RECT 78.565 8.605 78.735 8.775 ;
      RECT 78.255 2.025 78.425 2.195 ;
      RECT 78.255 6.685 78.425 6.855 ;
      RECT 77.885 0.105 78.055 0.275 ;
      RECT 77.885 8.605 78.055 8.775 ;
      RECT 77.825 0.915 77.995 1.085 ;
      RECT 77.825 1.655 77.995 1.825 ;
      RECT 77.825 7.055 77.995 7.225 ;
      RECT 77.825 7.795 77.995 7.965 ;
      RECT 77.45 2.395 77.62 2.565 ;
      RECT 77.45 6.315 77.62 6.485 ;
      RECT 77.205 0.105 77.375 0.275 ;
      RECT 77.205 8.605 77.375 8.775 ;
      RECT 76.525 0.105 76.695 0.275 ;
      RECT 76.525 8.605 76.695 8.775 ;
      RECT 76.455 2.765 76.625 2.935 ;
      RECT 76.455 5.945 76.625 6.115 ;
      RECT 74.91 1.415 75.08 1.585 ;
      RECT 74.91 4.135 75.08 4.305 ;
      RECT 74.655 2.775 74.825 2.945 ;
      RECT 74.45 1.415 74.62 1.585 ;
      RECT 74.45 4.135 74.62 4.305 ;
      RECT 74.175 1.935 74.345 2.105 ;
      RECT 73.99 1.415 74.16 1.585 ;
      RECT 73.99 4.135 74.16 4.305 ;
      RECT 73.935 2.495 74.105 2.665 ;
      RECT 73.53 1.415 73.7 1.585 ;
      RECT 73.53 4.135 73.7 4.305 ;
      RECT 73.455 2.495 73.625 2.665 ;
      RECT 73.215 1.935 73.385 2.105 ;
      RECT 73.215 3.615 73.385 3.785 ;
      RECT 73.07 1.415 73.24 1.585 ;
      RECT 73.07 4.135 73.24 4.305 ;
      RECT 72.95 4.545 73.12 4.715 ;
      RECT 72.95 8.605 73.12 8.775 ;
      RECT 72.695 2.775 72.865 2.945 ;
      RECT 72.64 6.685 72.81 6.855 ;
      RECT 72.61 1.415 72.78 1.585 ;
      RECT 72.61 4.135 72.78 4.305 ;
      RECT 72.455 2.215 72.625 2.385 ;
      RECT 72.27 8.605 72.44 8.775 ;
      RECT 72.215 3.615 72.385 3.785 ;
      RECT 72.21 7.055 72.38 7.225 ;
      RECT 72.21 7.795 72.38 7.965 ;
      RECT 72.15 1.415 72.32 1.585 ;
      RECT 72.15 4.135 72.32 4.305 ;
      RECT 71.975 2.775 72.145 2.945 ;
      RECT 71.835 6.315 72.005 6.485 ;
      RECT 71.69 1.415 71.86 1.585 ;
      RECT 71.69 4.135 71.86 4.305 ;
      RECT 71.59 8.605 71.76 8.775 ;
      RECT 71.495 2.495 71.665 2.665 ;
      RECT 71.23 1.415 71.4 1.585 ;
      RECT 71.23 4.135 71.4 4.305 ;
      RECT 71.015 2.495 71.185 2.665 ;
      RECT 70.91 8.605 71.08 8.775 ;
      RECT 70.84 5.945 71.01 6.115 ;
      RECT 70.775 1.935 70.945 2.105 ;
      RECT 70.77 1.415 70.94 1.585 ;
      RECT 70.77 4.135 70.94 4.305 ;
      RECT 70.31 1.415 70.48 1.585 ;
      RECT 70.31 4.135 70.48 4.305 ;
      RECT 70.015 2.215 70.185 2.385 ;
      RECT 69.85 1.415 70.02 1.585 ;
      RECT 69.85 4.135 70.02 4.305 ;
      RECT 69.775 3.335 69.945 3.505 ;
      RECT 69.535 2.775 69.705 2.945 ;
      RECT 69.39 1.415 69.56 1.585 ;
      RECT 69.39 4.135 69.56 4.305 ;
      RECT 69.055 2.495 69.225 2.665 ;
      RECT 68.93 1.415 69.1 1.585 ;
      RECT 68.93 4.135 69.1 4.305 ;
      RECT 68.815 1.935 68.985 2.105 ;
      RECT 68.815 3.335 68.985 3.505 ;
      RECT 68.47 1.415 68.64 1.585 ;
      RECT 68.47 4.135 68.64 4.305 ;
      RECT 68.335 3.055 68.505 3.225 ;
      RECT 68.01 1.415 68.18 1.585 ;
      RECT 68.01 4.135 68.18 4.305 ;
      RECT 67.815 2.495 67.985 2.665 ;
      RECT 67.575 3.335 67.745 3.505 ;
      RECT 67.55 1.415 67.72 1.585 ;
      RECT 67.55 4.135 67.72 4.305 ;
      RECT 67.335 1.935 67.505 2.105 ;
      RECT 67.095 2.495 67.265 2.665 ;
      RECT 67.095 3.055 67.265 3.225 ;
      RECT 67.09 1.415 67.26 1.585 ;
      RECT 67.09 4.135 67.26 4.305 ;
      RECT 66.63 1.415 66.8 1.585 ;
      RECT 66.63 4.135 66.8 4.305 ;
      RECT 66.375 1.935 66.545 2.105 ;
      RECT 66.375 3.615 66.545 3.785 ;
      RECT 66.17 1.415 66.34 1.585 ;
      RECT 66.17 4.135 66.34 4.305 ;
      RECT 65.895 3.055 66.065 3.225 ;
      RECT 65.71 1.415 65.88 1.585 ;
      RECT 65.71 4.135 65.88 4.305 ;
      RECT 64.285 0.915 64.455 1.085 ;
      RECT 64.285 2.395 64.455 2.565 ;
      RECT 64.285 6.315 64.455 6.485 ;
      RECT 64.285 7.795 64.455 7.965 ;
      RECT 63.935 0.105 64.105 0.275 ;
      RECT 63.935 4.165 64.105 4.335 ;
      RECT 63.935 4.545 64.105 4.715 ;
      RECT 63.935 8.605 64.105 8.775 ;
      RECT 63.915 2.765 64.085 2.935 ;
      RECT 63.915 5.945 64.085 6.115 ;
      RECT 63.295 0.915 63.465 1.085 ;
      RECT 63.295 2.395 63.465 2.565 ;
      RECT 63.295 6.315 63.465 6.485 ;
      RECT 63.295 7.795 63.465 7.965 ;
      RECT 62.945 0.105 63.115 0.275 ;
      RECT 62.945 4.165 63.115 4.335 ;
      RECT 62.945 4.545 63.115 4.715 ;
      RECT 62.945 8.605 63.115 8.775 ;
      RECT 62.925 2.765 63.095 2.935 ;
      RECT 62.925 5.945 63.095 6.115 ;
      RECT 62.24 0.105 62.41 0.275 ;
      RECT 62.24 4.165 62.41 4.335 ;
      RECT 62.24 4.545 62.41 4.715 ;
      RECT 62.24 8.605 62.41 8.775 ;
      RECT 61.93 2.025 62.1 2.195 ;
      RECT 61.93 6.685 62.1 6.855 ;
      RECT 61.56 0.105 61.73 0.275 ;
      RECT 61.56 8.605 61.73 8.775 ;
      RECT 61.5 0.915 61.67 1.085 ;
      RECT 61.5 1.655 61.67 1.825 ;
      RECT 61.5 7.055 61.67 7.225 ;
      RECT 61.5 7.795 61.67 7.965 ;
      RECT 61.125 2.395 61.295 2.565 ;
      RECT 61.125 6.315 61.295 6.485 ;
      RECT 60.88 0.105 61.05 0.275 ;
      RECT 60.88 8.605 61.05 8.775 ;
      RECT 60.2 0.105 60.37 0.275 ;
      RECT 60.2 8.605 60.37 8.775 ;
      RECT 60.13 2.765 60.3 2.935 ;
      RECT 60.13 5.945 60.3 6.115 ;
      RECT 58.585 1.415 58.755 1.585 ;
      RECT 58.585 4.135 58.755 4.305 ;
      RECT 58.33 2.775 58.5 2.945 ;
      RECT 58.125 1.415 58.295 1.585 ;
      RECT 58.125 4.135 58.295 4.305 ;
      RECT 57.85 1.935 58.02 2.105 ;
      RECT 57.665 1.415 57.835 1.585 ;
      RECT 57.665 4.135 57.835 4.305 ;
      RECT 57.61 2.495 57.78 2.665 ;
      RECT 57.205 1.415 57.375 1.585 ;
      RECT 57.205 4.135 57.375 4.305 ;
      RECT 57.13 2.495 57.3 2.665 ;
      RECT 56.89 1.935 57.06 2.105 ;
      RECT 56.89 3.615 57.06 3.785 ;
      RECT 56.745 1.415 56.915 1.585 ;
      RECT 56.745 4.135 56.915 4.305 ;
      RECT 56.625 4.545 56.795 4.715 ;
      RECT 56.625 8.605 56.795 8.775 ;
      RECT 56.37 2.775 56.54 2.945 ;
      RECT 56.315 6.685 56.485 6.855 ;
      RECT 56.285 1.415 56.455 1.585 ;
      RECT 56.285 4.135 56.455 4.305 ;
      RECT 56.13 2.215 56.3 2.385 ;
      RECT 55.945 8.605 56.115 8.775 ;
      RECT 55.89 3.615 56.06 3.785 ;
      RECT 55.885 7.055 56.055 7.225 ;
      RECT 55.885 7.795 56.055 7.965 ;
      RECT 55.825 1.415 55.995 1.585 ;
      RECT 55.825 4.135 55.995 4.305 ;
      RECT 55.65 2.775 55.82 2.945 ;
      RECT 55.51 6.315 55.68 6.485 ;
      RECT 55.365 1.415 55.535 1.585 ;
      RECT 55.365 4.135 55.535 4.305 ;
      RECT 55.265 8.605 55.435 8.775 ;
      RECT 55.17 2.495 55.34 2.665 ;
      RECT 54.905 1.415 55.075 1.585 ;
      RECT 54.905 4.135 55.075 4.305 ;
      RECT 54.69 2.495 54.86 2.665 ;
      RECT 54.585 8.605 54.755 8.775 ;
      RECT 54.515 5.945 54.685 6.115 ;
      RECT 54.45 1.935 54.62 2.105 ;
      RECT 54.445 1.415 54.615 1.585 ;
      RECT 54.445 4.135 54.615 4.305 ;
      RECT 53.985 1.415 54.155 1.585 ;
      RECT 53.985 4.135 54.155 4.305 ;
      RECT 53.69 2.215 53.86 2.385 ;
      RECT 53.525 1.415 53.695 1.585 ;
      RECT 53.525 4.135 53.695 4.305 ;
      RECT 53.45 3.335 53.62 3.505 ;
      RECT 53.21 2.775 53.38 2.945 ;
      RECT 53.065 1.415 53.235 1.585 ;
      RECT 53.065 4.135 53.235 4.305 ;
      RECT 52.73 2.495 52.9 2.665 ;
      RECT 52.605 1.415 52.775 1.585 ;
      RECT 52.605 4.135 52.775 4.305 ;
      RECT 52.49 1.935 52.66 2.105 ;
      RECT 52.49 3.335 52.66 3.505 ;
      RECT 52.145 1.415 52.315 1.585 ;
      RECT 52.145 4.135 52.315 4.305 ;
      RECT 52.01 3.055 52.18 3.225 ;
      RECT 51.685 1.415 51.855 1.585 ;
      RECT 51.685 4.135 51.855 4.305 ;
      RECT 51.49 2.495 51.66 2.665 ;
      RECT 51.25 3.335 51.42 3.505 ;
      RECT 51.225 1.415 51.395 1.585 ;
      RECT 51.225 4.135 51.395 4.305 ;
      RECT 51.01 1.935 51.18 2.105 ;
      RECT 50.77 2.495 50.94 2.665 ;
      RECT 50.77 3.055 50.94 3.225 ;
      RECT 50.765 1.415 50.935 1.585 ;
      RECT 50.765 4.135 50.935 4.305 ;
      RECT 50.305 1.415 50.475 1.585 ;
      RECT 50.305 4.135 50.475 4.305 ;
      RECT 50.05 1.935 50.22 2.105 ;
      RECT 50.05 3.615 50.22 3.785 ;
      RECT 49.845 1.415 50.015 1.585 ;
      RECT 49.845 4.135 50.015 4.305 ;
      RECT 49.57 3.055 49.74 3.225 ;
      RECT 49.385 1.415 49.555 1.585 ;
      RECT 49.385 4.135 49.555 4.305 ;
      RECT 47.96 0.915 48.13 1.085 ;
      RECT 47.96 2.395 48.13 2.565 ;
      RECT 47.96 6.315 48.13 6.485 ;
      RECT 47.96 7.795 48.13 7.965 ;
      RECT 47.61 0.105 47.78 0.275 ;
      RECT 47.61 4.165 47.78 4.335 ;
      RECT 47.61 4.545 47.78 4.715 ;
      RECT 47.61 8.605 47.78 8.775 ;
      RECT 47.59 2.765 47.76 2.935 ;
      RECT 47.59 5.945 47.76 6.115 ;
      RECT 46.97 0.915 47.14 1.085 ;
      RECT 46.97 2.395 47.14 2.565 ;
      RECT 46.97 6.315 47.14 6.485 ;
      RECT 46.97 7.795 47.14 7.965 ;
      RECT 46.62 0.105 46.79 0.275 ;
      RECT 46.62 4.165 46.79 4.335 ;
      RECT 46.62 4.545 46.79 4.715 ;
      RECT 46.62 8.605 46.79 8.775 ;
      RECT 46.6 2.765 46.77 2.935 ;
      RECT 46.6 5.945 46.77 6.115 ;
      RECT 45.915 0.105 46.085 0.275 ;
      RECT 45.915 4.165 46.085 4.335 ;
      RECT 45.915 4.545 46.085 4.715 ;
      RECT 45.915 8.605 46.085 8.775 ;
      RECT 45.605 2.025 45.775 2.195 ;
      RECT 45.605 6.685 45.775 6.855 ;
      RECT 45.235 0.105 45.405 0.275 ;
      RECT 45.235 8.605 45.405 8.775 ;
      RECT 45.175 0.915 45.345 1.085 ;
      RECT 45.175 1.655 45.345 1.825 ;
      RECT 45.175 7.055 45.345 7.225 ;
      RECT 45.175 7.795 45.345 7.965 ;
      RECT 44.8 2.395 44.97 2.565 ;
      RECT 44.8 6.315 44.97 6.485 ;
      RECT 44.555 0.105 44.725 0.275 ;
      RECT 44.555 8.605 44.725 8.775 ;
      RECT 43.875 0.105 44.045 0.275 ;
      RECT 43.875 8.605 44.045 8.775 ;
      RECT 43.805 2.765 43.975 2.935 ;
      RECT 43.805 5.945 43.975 6.115 ;
      RECT 42.26 1.415 42.43 1.585 ;
      RECT 42.26 4.135 42.43 4.305 ;
      RECT 42.005 2.775 42.175 2.945 ;
      RECT 41.8 1.415 41.97 1.585 ;
      RECT 41.8 4.135 41.97 4.305 ;
      RECT 41.525 1.935 41.695 2.105 ;
      RECT 41.34 1.415 41.51 1.585 ;
      RECT 41.34 4.135 41.51 4.305 ;
      RECT 41.285 2.495 41.455 2.665 ;
      RECT 40.88 1.415 41.05 1.585 ;
      RECT 40.88 4.135 41.05 4.305 ;
      RECT 40.805 2.495 40.975 2.665 ;
      RECT 40.565 1.935 40.735 2.105 ;
      RECT 40.565 3.615 40.735 3.785 ;
      RECT 40.42 1.415 40.59 1.585 ;
      RECT 40.42 4.135 40.59 4.305 ;
      RECT 40.3 4.545 40.47 4.715 ;
      RECT 40.3 8.605 40.47 8.775 ;
      RECT 40.045 2.775 40.215 2.945 ;
      RECT 39.99 6.685 40.16 6.855 ;
      RECT 39.96 1.415 40.13 1.585 ;
      RECT 39.96 4.135 40.13 4.305 ;
      RECT 39.805 2.215 39.975 2.385 ;
      RECT 39.62 8.605 39.79 8.775 ;
      RECT 39.565 3.615 39.735 3.785 ;
      RECT 39.56 7.055 39.73 7.225 ;
      RECT 39.56 7.795 39.73 7.965 ;
      RECT 39.5 1.415 39.67 1.585 ;
      RECT 39.5 4.135 39.67 4.305 ;
      RECT 39.325 2.775 39.495 2.945 ;
      RECT 39.185 6.315 39.355 6.485 ;
      RECT 39.04 1.415 39.21 1.585 ;
      RECT 39.04 4.135 39.21 4.305 ;
      RECT 38.94 8.605 39.11 8.775 ;
      RECT 38.845 2.495 39.015 2.665 ;
      RECT 38.58 1.415 38.75 1.585 ;
      RECT 38.58 4.135 38.75 4.305 ;
      RECT 38.365 2.495 38.535 2.665 ;
      RECT 38.26 8.605 38.43 8.775 ;
      RECT 38.19 5.945 38.36 6.115 ;
      RECT 38.125 1.935 38.295 2.105 ;
      RECT 38.12 1.415 38.29 1.585 ;
      RECT 38.12 4.135 38.29 4.305 ;
      RECT 37.66 1.415 37.83 1.585 ;
      RECT 37.66 4.135 37.83 4.305 ;
      RECT 37.365 2.215 37.535 2.385 ;
      RECT 37.2 1.415 37.37 1.585 ;
      RECT 37.2 4.135 37.37 4.305 ;
      RECT 37.125 3.335 37.295 3.505 ;
      RECT 36.885 2.775 37.055 2.945 ;
      RECT 36.74 1.415 36.91 1.585 ;
      RECT 36.74 4.135 36.91 4.305 ;
      RECT 36.405 2.495 36.575 2.665 ;
      RECT 36.28 1.415 36.45 1.585 ;
      RECT 36.28 4.135 36.45 4.305 ;
      RECT 36.165 1.935 36.335 2.105 ;
      RECT 36.165 3.335 36.335 3.505 ;
      RECT 35.82 1.415 35.99 1.585 ;
      RECT 35.82 4.135 35.99 4.305 ;
      RECT 35.685 3.055 35.855 3.225 ;
      RECT 35.36 1.415 35.53 1.585 ;
      RECT 35.36 4.135 35.53 4.305 ;
      RECT 35.165 2.495 35.335 2.665 ;
      RECT 34.925 3.335 35.095 3.505 ;
      RECT 34.9 1.415 35.07 1.585 ;
      RECT 34.9 4.135 35.07 4.305 ;
      RECT 34.685 1.935 34.855 2.105 ;
      RECT 34.445 2.495 34.615 2.665 ;
      RECT 34.445 3.055 34.615 3.225 ;
      RECT 34.44 1.415 34.61 1.585 ;
      RECT 34.44 4.135 34.61 4.305 ;
      RECT 33.98 1.415 34.15 1.585 ;
      RECT 33.98 4.135 34.15 4.305 ;
      RECT 33.725 1.935 33.895 2.105 ;
      RECT 33.725 3.615 33.895 3.785 ;
      RECT 33.52 1.415 33.69 1.585 ;
      RECT 33.52 4.135 33.69 4.305 ;
      RECT 33.245 3.055 33.415 3.225 ;
      RECT 33.06 1.415 33.23 1.585 ;
      RECT 33.06 4.135 33.23 4.305 ;
      RECT 31.635 0.915 31.805 1.085 ;
      RECT 31.635 2.395 31.805 2.565 ;
      RECT 31.635 6.315 31.805 6.485 ;
      RECT 31.635 7.795 31.805 7.965 ;
      RECT 31.285 0.105 31.455 0.275 ;
      RECT 31.285 4.165 31.455 4.335 ;
      RECT 31.285 4.545 31.455 4.715 ;
      RECT 31.285 8.605 31.455 8.775 ;
      RECT 31.265 2.765 31.435 2.935 ;
      RECT 31.265 5.945 31.435 6.115 ;
      RECT 30.645 0.915 30.815 1.085 ;
      RECT 30.645 2.395 30.815 2.565 ;
      RECT 30.645 6.315 30.815 6.485 ;
      RECT 30.645 7.795 30.815 7.965 ;
      RECT 30.295 0.105 30.465 0.275 ;
      RECT 30.295 4.165 30.465 4.335 ;
      RECT 30.295 4.545 30.465 4.715 ;
      RECT 30.295 8.605 30.465 8.775 ;
      RECT 30.275 2.765 30.445 2.935 ;
      RECT 30.275 5.945 30.445 6.115 ;
      RECT 29.59 0.105 29.76 0.275 ;
      RECT 29.59 4.165 29.76 4.335 ;
      RECT 29.59 4.545 29.76 4.715 ;
      RECT 29.59 8.605 29.76 8.775 ;
      RECT 29.28 2.025 29.45 2.195 ;
      RECT 29.28 6.685 29.45 6.855 ;
      RECT 28.91 0.105 29.08 0.275 ;
      RECT 28.91 8.605 29.08 8.775 ;
      RECT 28.85 0.915 29.02 1.085 ;
      RECT 28.85 1.655 29.02 1.825 ;
      RECT 28.85 7.055 29.02 7.225 ;
      RECT 28.85 7.795 29.02 7.965 ;
      RECT 28.475 2.395 28.645 2.565 ;
      RECT 28.475 6.315 28.645 6.485 ;
      RECT 28.23 0.105 28.4 0.275 ;
      RECT 28.23 8.605 28.4 8.775 ;
      RECT 27.55 0.105 27.72 0.275 ;
      RECT 27.55 8.605 27.72 8.775 ;
      RECT 27.48 2.765 27.65 2.935 ;
      RECT 27.48 5.945 27.65 6.115 ;
      RECT 25.935 1.415 26.105 1.585 ;
      RECT 25.935 4.135 26.105 4.305 ;
      RECT 25.68 2.775 25.85 2.945 ;
      RECT 25.475 1.415 25.645 1.585 ;
      RECT 25.475 4.135 25.645 4.305 ;
      RECT 25.2 1.935 25.37 2.105 ;
      RECT 25.015 1.415 25.185 1.585 ;
      RECT 25.015 4.135 25.185 4.305 ;
      RECT 24.96 2.495 25.13 2.665 ;
      RECT 24.555 1.415 24.725 1.585 ;
      RECT 24.555 4.135 24.725 4.305 ;
      RECT 24.48 2.495 24.65 2.665 ;
      RECT 24.24 1.935 24.41 2.105 ;
      RECT 24.24 3.615 24.41 3.785 ;
      RECT 24.095 1.415 24.265 1.585 ;
      RECT 24.095 4.135 24.265 4.305 ;
      RECT 23.975 4.545 24.145 4.715 ;
      RECT 23.975 8.605 24.145 8.775 ;
      RECT 23.72 2.775 23.89 2.945 ;
      RECT 23.665 6.685 23.835 6.855 ;
      RECT 23.635 1.415 23.805 1.585 ;
      RECT 23.635 4.135 23.805 4.305 ;
      RECT 23.48 2.215 23.65 2.385 ;
      RECT 23.295 8.605 23.465 8.775 ;
      RECT 23.24 3.615 23.41 3.785 ;
      RECT 23.235 7.055 23.405 7.225 ;
      RECT 23.235 7.795 23.405 7.965 ;
      RECT 23.175 1.415 23.345 1.585 ;
      RECT 23.175 4.135 23.345 4.305 ;
      RECT 23 2.775 23.17 2.945 ;
      RECT 22.86 6.315 23.03 6.485 ;
      RECT 22.715 1.415 22.885 1.585 ;
      RECT 22.715 4.135 22.885 4.305 ;
      RECT 22.615 8.605 22.785 8.775 ;
      RECT 22.52 2.495 22.69 2.665 ;
      RECT 22.255 1.415 22.425 1.585 ;
      RECT 22.255 4.135 22.425 4.305 ;
      RECT 22.04 2.495 22.21 2.665 ;
      RECT 21.935 8.605 22.105 8.775 ;
      RECT 21.865 5.945 22.035 6.115 ;
      RECT 21.8 1.935 21.97 2.105 ;
      RECT 21.795 1.415 21.965 1.585 ;
      RECT 21.795 4.135 21.965 4.305 ;
      RECT 21.335 1.415 21.505 1.585 ;
      RECT 21.335 4.135 21.505 4.305 ;
      RECT 21.04 2.215 21.21 2.385 ;
      RECT 20.875 1.415 21.045 1.585 ;
      RECT 20.875 4.135 21.045 4.305 ;
      RECT 20.8 3.335 20.97 3.505 ;
      RECT 20.56 2.775 20.73 2.945 ;
      RECT 20.415 1.415 20.585 1.585 ;
      RECT 20.415 4.135 20.585 4.305 ;
      RECT 20.08 2.495 20.25 2.665 ;
      RECT 19.955 1.415 20.125 1.585 ;
      RECT 19.955 4.135 20.125 4.305 ;
      RECT 19.84 1.935 20.01 2.105 ;
      RECT 19.84 3.335 20.01 3.505 ;
      RECT 19.495 1.415 19.665 1.585 ;
      RECT 19.495 4.135 19.665 4.305 ;
      RECT 19.36 3.055 19.53 3.225 ;
      RECT 19.035 1.415 19.205 1.585 ;
      RECT 19.035 4.135 19.205 4.305 ;
      RECT 18.84 2.495 19.01 2.665 ;
      RECT 18.6 3.335 18.77 3.505 ;
      RECT 18.575 1.415 18.745 1.585 ;
      RECT 18.575 4.135 18.745 4.305 ;
      RECT 18.36 1.935 18.53 2.105 ;
      RECT 18.12 2.495 18.29 2.665 ;
      RECT 18.12 3.055 18.29 3.225 ;
      RECT 18.115 1.415 18.285 1.585 ;
      RECT 18.115 4.135 18.285 4.305 ;
      RECT 17.655 1.415 17.825 1.585 ;
      RECT 17.655 4.135 17.825 4.305 ;
      RECT 17.4 1.935 17.57 2.105 ;
      RECT 17.4 3.615 17.57 3.785 ;
      RECT 17.195 1.415 17.365 1.585 ;
      RECT 17.195 4.135 17.365 4.305 ;
      RECT 16.92 3.055 17.09 3.225 ;
      RECT 16.735 1.415 16.905 1.585 ;
      RECT 16.735 4.135 16.905 4.305 ;
      RECT 15.31 0.915 15.48 1.085 ;
      RECT 15.31 2.395 15.48 2.565 ;
      RECT 15.31 6.315 15.48 6.485 ;
      RECT 15.31 7.795 15.48 7.965 ;
      RECT 14.96 0.105 15.13 0.275 ;
      RECT 14.96 4.165 15.13 4.335 ;
      RECT 14.96 4.545 15.13 4.715 ;
      RECT 14.96 8.605 15.13 8.775 ;
      RECT 14.94 2.765 15.11 2.935 ;
      RECT 14.94 5.945 15.11 6.115 ;
      RECT 14.32 0.915 14.49 1.085 ;
      RECT 14.32 2.395 14.49 2.565 ;
      RECT 14.32 6.315 14.49 6.485 ;
      RECT 14.32 7.795 14.49 7.965 ;
      RECT 13.97 0.105 14.14 0.275 ;
      RECT 13.97 4.165 14.14 4.335 ;
      RECT 13.97 4.545 14.14 4.715 ;
      RECT 13.97 8.605 14.14 8.775 ;
      RECT 13.95 2.765 14.12 2.935 ;
      RECT 13.95 5.945 14.12 6.115 ;
      RECT 13.265 0.105 13.435 0.275 ;
      RECT 13.265 4.165 13.435 4.335 ;
      RECT 13.265 4.545 13.435 4.715 ;
      RECT 13.265 8.605 13.435 8.775 ;
      RECT 12.955 2.025 13.125 2.195 ;
      RECT 12.955 6.685 13.125 6.855 ;
      RECT 12.585 0.105 12.755 0.275 ;
      RECT 12.585 8.605 12.755 8.775 ;
      RECT 12.525 0.915 12.695 1.085 ;
      RECT 12.525 1.655 12.695 1.825 ;
      RECT 12.525 7.055 12.695 7.225 ;
      RECT 12.525 7.795 12.695 7.965 ;
      RECT 12.15 2.395 12.32 2.565 ;
      RECT 12.15 6.315 12.32 6.485 ;
      RECT 11.905 0.105 12.075 0.275 ;
      RECT 11.905 8.605 12.075 8.775 ;
      RECT 11.225 0.105 11.395 0.275 ;
      RECT 11.225 8.605 11.395 8.775 ;
      RECT 11.155 2.765 11.325 2.935 ;
      RECT 11.155 5.945 11.325 6.115 ;
      RECT 9.61 1.415 9.78 1.585 ;
      RECT 9.61 4.135 9.78 4.305 ;
      RECT 9.355 2.775 9.525 2.945 ;
      RECT 9.15 1.415 9.32 1.585 ;
      RECT 9.15 4.135 9.32 4.305 ;
      RECT 8.875 1.935 9.045 2.105 ;
      RECT 8.69 1.415 8.86 1.585 ;
      RECT 8.69 4.135 8.86 4.305 ;
      RECT 8.635 2.495 8.805 2.665 ;
      RECT 8.23 1.415 8.4 1.585 ;
      RECT 8.23 4.135 8.4 4.305 ;
      RECT 8.155 2.495 8.325 2.665 ;
      RECT 7.915 1.935 8.085 2.105 ;
      RECT 7.915 3.615 8.085 3.785 ;
      RECT 7.77 1.415 7.94 1.585 ;
      RECT 7.77 4.135 7.94 4.305 ;
      RECT 7.65 4.545 7.82 4.715 ;
      RECT 7.65 8.605 7.82 8.775 ;
      RECT 7.395 2.775 7.565 2.945 ;
      RECT 7.34 6.685 7.51 6.855 ;
      RECT 7.31 1.415 7.48 1.585 ;
      RECT 7.31 4.135 7.48 4.305 ;
      RECT 7.155 2.215 7.325 2.385 ;
      RECT 6.97 8.605 7.14 8.775 ;
      RECT 6.915 3.615 7.085 3.785 ;
      RECT 6.91 7.055 7.08 7.225 ;
      RECT 6.91 7.795 7.08 7.965 ;
      RECT 6.85 1.415 7.02 1.585 ;
      RECT 6.85 4.135 7.02 4.305 ;
      RECT 6.675 2.775 6.845 2.945 ;
      RECT 6.535 6.315 6.705 6.485 ;
      RECT 6.39 1.415 6.56 1.585 ;
      RECT 6.39 4.135 6.56 4.305 ;
      RECT 6.29 8.605 6.46 8.775 ;
      RECT 6.195 2.495 6.365 2.665 ;
      RECT 5.93 1.415 6.1 1.585 ;
      RECT 5.93 4.135 6.1 4.305 ;
      RECT 5.715 2.495 5.885 2.665 ;
      RECT 5.61 8.605 5.78 8.775 ;
      RECT 5.54 5.945 5.71 6.115 ;
      RECT 5.475 1.935 5.645 2.105 ;
      RECT 5.47 1.415 5.64 1.585 ;
      RECT 5.47 4.135 5.64 4.305 ;
      RECT 5.01 1.415 5.18 1.585 ;
      RECT 5.01 4.135 5.18 4.305 ;
      RECT 4.715 2.215 4.885 2.385 ;
      RECT 4.55 1.415 4.72 1.585 ;
      RECT 4.55 4.135 4.72 4.305 ;
      RECT 4.475 3.335 4.645 3.505 ;
      RECT 4.235 2.775 4.405 2.945 ;
      RECT 4.09 1.415 4.26 1.585 ;
      RECT 4.09 4.135 4.26 4.305 ;
      RECT 3.755 2.495 3.925 2.665 ;
      RECT 3.63 1.415 3.8 1.585 ;
      RECT 3.63 4.135 3.8 4.305 ;
      RECT 3.515 1.935 3.685 2.105 ;
      RECT 3.515 3.335 3.685 3.505 ;
      RECT 3.17 1.415 3.34 1.585 ;
      RECT 3.17 4.135 3.34 4.305 ;
      RECT 3.035 3.055 3.205 3.225 ;
      RECT 2.71 1.415 2.88 1.585 ;
      RECT 2.71 4.135 2.88 4.305 ;
      RECT 2.515 2.495 2.685 2.665 ;
      RECT 2.275 3.335 2.445 3.505 ;
      RECT 2.25 1.415 2.42 1.585 ;
      RECT 2.25 4.135 2.42 4.305 ;
      RECT 2.035 1.935 2.205 2.105 ;
      RECT 1.795 2.495 1.965 2.665 ;
      RECT 1.795 3.055 1.965 3.225 ;
      RECT 1.79 1.415 1.96 1.585 ;
      RECT 1.79 4.135 1.96 4.305 ;
      RECT 1.33 1.415 1.5 1.585 ;
      RECT 1.33 4.135 1.5 4.305 ;
      RECT 1.075 1.935 1.245 2.105 ;
      RECT 1.075 3.615 1.245 3.785 ;
      RECT 0.87 1.415 1.04 1.585 ;
      RECT 0.87 4.135 1.04 4.305 ;
      RECT 0.595 3.055 0.765 3.225 ;
      RECT 0.41 1.415 0.58 1.585 ;
      RECT 0.41 4.135 0.58 4.305 ;
      RECT -0.93 4.545 -0.76 4.715 ;
      RECT -0.93 8.605 -0.76 8.775 ;
      RECT -1.24 6.685 -1.07 6.855 ;
      RECT -1.61 8.605 -1.44 8.775 ;
      RECT -1.67 7.055 -1.5 7.225 ;
      RECT -1.67 7.795 -1.5 7.965 ;
      RECT -2.045 6.315 -1.875 6.485 ;
      RECT -2.29 8.605 -2.12 8.775 ;
      RECT -2.97 8.605 -2.8 8.775 ;
      RECT -3.04 5.945 -2.87 6.115 ;
    LAYER li ;
      RECT 73.695 0 73.865 2.085 ;
      RECT 71.735 0 71.905 2.085 ;
      RECT 69.295 0 69.465 2.085 ;
      RECT 68.335 0 68.505 2.085 ;
      RECT 67.815 0 67.985 2.085 ;
      RECT 66.855 0 67.025 2.085 ;
      RECT 65.895 0 66.065 2.085 ;
      RECT 57.37 0 57.54 2.085 ;
      RECT 55.41 0 55.58 2.085 ;
      RECT 52.97 0 53.14 2.085 ;
      RECT 52.01 0 52.18 2.085 ;
      RECT 51.49 0 51.66 2.085 ;
      RECT 50.53 0 50.7 2.085 ;
      RECT 49.57 0 49.74 2.085 ;
      RECT 41.045 0 41.215 2.085 ;
      RECT 39.085 0 39.255 2.085 ;
      RECT 36.645 0 36.815 2.085 ;
      RECT 35.685 0 35.855 2.085 ;
      RECT 35.165 0 35.335 2.085 ;
      RECT 34.205 0 34.375 2.085 ;
      RECT 33.245 0 33.415 2.085 ;
      RECT 24.72 0 24.89 2.085 ;
      RECT 22.76 0 22.93 2.085 ;
      RECT 20.32 0 20.49 2.085 ;
      RECT 19.36 0 19.53 2.085 ;
      RECT 18.84 0 19.01 2.085 ;
      RECT 17.88 0 18.05 2.085 ;
      RECT 16.92 0 17.09 2.085 ;
      RECT 8.395 0 8.565 2.085 ;
      RECT 6.435 0 6.605 2.085 ;
      RECT 3.995 0 4.165 2.085 ;
      RECT 3.035 0 3.205 2.085 ;
      RECT 2.515 0 2.685 2.085 ;
      RECT 1.555 0 1.725 2.085 ;
      RECT 0.595 0 0.765 2.085 ;
      RECT 71.665 0 71.905 1.595 ;
      RECT 70.115 0 70.31 1.595 ;
      RECT 67.99 0 68.185 1.595 ;
      RECT 65.69 0 65.885 1.595 ;
      RECT 55.34 0 55.58 1.595 ;
      RECT 53.79 0 53.985 1.595 ;
      RECT 51.665 0 51.86 1.595 ;
      RECT 49.365 0 49.56 1.595 ;
      RECT 39.015 0 39.255 1.595 ;
      RECT 37.465 0 37.66 1.595 ;
      RECT 35.34 0 35.535 1.595 ;
      RECT 33.04 0 33.235 1.595 ;
      RECT 22.69 0 22.93 1.595 ;
      RECT 21.14 0 21.335 1.595 ;
      RECT 19.015 0 19.21 1.595 ;
      RECT 16.715 0 16.91 1.595 ;
      RECT 6.365 0 6.605 1.595 ;
      RECT 4.815 0 5.01 1.595 ;
      RECT 2.69 0 2.885 1.595 ;
      RECT 0.39 0 0.585 1.595 ;
      RECT 65.565 0 75.38 1.585 ;
      RECT 49.24 0 59.055 1.585 ;
      RECT 32.915 0 42.73 1.585 ;
      RECT 16.59 0 26.405 1.585 ;
      RECT 0.265 0 10.08 1.585 ;
      RECT 80.18 0 80.35 0.935 ;
      RECT 79.19 0 79.36 0.935 ;
      RECT 76.445 0 76.615 0.935 ;
      RECT 63.855 0 64.025 0.935 ;
      RECT 62.865 0 63.035 0.935 ;
      RECT 60.12 0 60.29 0.935 ;
      RECT 47.53 0 47.7 0.935 ;
      RECT 46.54 0 46.71 0.935 ;
      RECT 43.795 0 43.965 0.935 ;
      RECT 31.205 0 31.375 0.935 ;
      RECT 30.215 0 30.385 0.935 ;
      RECT 27.47 0 27.64 0.935 ;
      RECT 14.88 0 15.05 0.935 ;
      RECT 13.89 0 14.06 0.935 ;
      RECT 11.145 0 11.315 0.935 ;
      RECT -3.225 0 81.15 0.305 ;
      RECT -1.24 4.135 -1.07 8.305 ;
      RECT 80.18 3.405 80.35 5.475 ;
      RECT 79.19 3.405 79.36 5.475 ;
      RECT 76.445 3.405 76.615 5.475 ;
      RECT 70.83 4.135 71 5.475 ;
      RECT 63.855 3.405 64.025 5.475 ;
      RECT 62.865 3.405 63.035 5.475 ;
      RECT 60.12 3.405 60.29 5.475 ;
      RECT 54.505 4.135 54.675 5.475 ;
      RECT 47.53 3.405 47.7 5.475 ;
      RECT 46.54 3.405 46.71 5.475 ;
      RECT 43.795 3.405 43.965 5.475 ;
      RECT 38.18 4.135 38.35 5.475 ;
      RECT 31.205 3.405 31.375 5.475 ;
      RECT 30.215 3.405 30.385 5.475 ;
      RECT 27.47 3.405 27.64 5.475 ;
      RECT 21.855 4.135 22.025 5.475 ;
      RECT 14.88 3.405 15.05 5.475 ;
      RECT 13.89 3.405 14.06 5.475 ;
      RECT 11.145 3.405 11.315 5.475 ;
      RECT 5.53 4.135 5.7 5.475 ;
      RECT -3.05 4.135 -2.88 5.475 ;
      RECT -3.225 4.135 81.15 4.745 ;
      RECT 74.655 3.635 74.825 4.745 ;
      RECT 73.695 3.635 73.865 4.745 ;
      RECT 71.255 3.635 71.425 4.745 ;
      RECT 70.255 3.635 70.425 4.745 ;
      RECT 69.295 3.635 69.465 4.745 ;
      RECT 66.855 3.635 67.025 4.745 ;
      RECT 58.33 3.635 58.5 4.745 ;
      RECT 57.37 3.635 57.54 4.745 ;
      RECT 54.93 3.635 55.1 4.745 ;
      RECT 53.93 3.635 54.1 4.745 ;
      RECT 52.97 3.635 53.14 4.745 ;
      RECT 50.53 3.635 50.7 4.745 ;
      RECT 42.005 3.635 42.175 4.745 ;
      RECT 41.045 3.635 41.215 4.745 ;
      RECT 38.605 3.635 38.775 4.745 ;
      RECT 37.605 3.635 37.775 4.745 ;
      RECT 36.645 3.635 36.815 4.745 ;
      RECT 34.205 3.635 34.375 4.745 ;
      RECT 25.68 3.635 25.85 4.745 ;
      RECT 24.72 3.635 24.89 4.745 ;
      RECT 22.28 3.635 22.45 4.745 ;
      RECT 21.28 3.635 21.45 4.745 ;
      RECT 20.32 3.635 20.49 4.745 ;
      RECT 17.88 3.635 18.05 4.745 ;
      RECT 9.355 3.635 9.525 4.745 ;
      RECT 8.395 3.635 8.565 4.745 ;
      RECT 5.955 3.635 6.125 4.745 ;
      RECT 4.955 3.635 5.125 4.745 ;
      RECT 3.995 3.635 4.165 4.745 ;
      RECT 1.555 3.635 1.725 4.745 ;
      RECT -3.225 8.575 81.15 8.88 ;
      RECT 80.18 7.945 80.35 8.88 ;
      RECT 79.19 7.945 79.36 8.88 ;
      RECT 76.445 7.945 76.615 8.88 ;
      RECT 70.83 7.945 71 8.88 ;
      RECT 63.855 7.945 64.025 8.88 ;
      RECT 62.865 7.945 63.035 8.88 ;
      RECT 60.12 7.945 60.29 8.88 ;
      RECT 54.505 7.945 54.675 8.88 ;
      RECT 47.53 7.945 47.7 8.88 ;
      RECT 46.54 7.945 46.71 8.88 ;
      RECT 43.795 7.945 43.965 8.88 ;
      RECT 38.18 7.945 38.35 8.88 ;
      RECT 31.205 7.945 31.375 8.88 ;
      RECT 30.215 7.945 30.385 8.88 ;
      RECT 27.47 7.945 27.64 8.88 ;
      RECT 21.855 7.945 22.025 8.88 ;
      RECT 14.88 7.945 15.05 8.88 ;
      RECT 13.89 7.945 14.06 8.88 ;
      RECT 11.145 7.945 11.315 8.88 ;
      RECT 5.53 7.945 5.7 8.88 ;
      RECT -3.05 7.945 -2.88 8.88 ;
      RECT 80.24 1.74 80.41 2.935 ;
      RECT 80.24 1.74 80.705 1.91 ;
      RECT 80.24 6.97 80.705 7.14 ;
      RECT 80.24 5.945 80.41 7.14 ;
      RECT 79.25 1.74 79.42 2.935 ;
      RECT 79.25 1.74 79.715 1.91 ;
      RECT 79.25 6.97 79.715 7.14 ;
      RECT 79.25 5.945 79.42 7.14 ;
      RECT 77.395 2.635 77.565 3.865 ;
      RECT 77.45 0.855 77.62 2.805 ;
      RECT 77.395 0.575 77.565 1.025 ;
      RECT 77.395 7.855 77.565 8.305 ;
      RECT 77.45 6.075 77.62 8.025 ;
      RECT 77.395 5.015 77.565 6.245 ;
      RECT 76.875 0.575 77.045 3.865 ;
      RECT 76.875 2.075 77.28 2.405 ;
      RECT 76.875 1.235 77.28 1.565 ;
      RECT 76.875 5.015 77.045 8.305 ;
      RECT 76.875 7.315 77.28 7.645 ;
      RECT 76.875 6.475 77.28 6.805 ;
      RECT 74.175 1.835 74.345 2.105 ;
      RECT 74.175 1.835 74.905 2.005 ;
      RECT 74.655 2.575 74.825 2.945 ;
      RECT 74.335 2.575 74.825 2.745 ;
      RECT 74.095 3.225 74.425 3.395 ;
      RECT 73.335 3.055 74.345 3.225 ;
      RECT 73.335 2.575 73.505 3.225 ;
      RECT 73.455 2.495 73.625 2.825 ;
      RECT 72.615 3.225 72.945 3.395 ;
      RECT 70.695 3.225 71.985 3.395 ;
      RECT 71.735 3.14 72.865 3.31 ;
      RECT 72.455 2.215 72.865 2.385 ;
      RECT 72.695 1.755 72.865 2.385 ;
      RECT 72.695 2.575 72.865 2.945 ;
      RECT 72.375 2.575 72.865 2.745 ;
      RECT 71.78 7.855 71.95 8.305 ;
      RECT 71.835 6.075 72.005 8.025 ;
      RECT 71.78 5.015 71.95 6.245 ;
      RECT 71.26 5.015 71.43 8.305 ;
      RECT 71.26 7.315 71.665 7.645 ;
      RECT 71.26 6.475 71.665 6.805 ;
      RECT 69.935 2.575 71.265 2.745 ;
      RECT 71.015 2.495 71.185 2.745 ;
      RECT 70.015 2.175 70.185 2.385 ;
      RECT 70.015 2.175 70.505 2.345 ;
      RECT 68.695 3.335 68.985 3.505 ;
      RECT 68.695 2.575 68.865 3.505 ;
      RECT 68.495 2.575 68.865 2.745 ;
      RECT 67.495 2.575 67.985 2.745 ;
      RECT 67.815 2.495 67.985 2.745 ;
      RECT 67.575 3.335 67.985 3.505 ;
      RECT 67.815 3.145 67.985 3.505 ;
      RECT 66.615 3.055 67.265 3.225 ;
      RECT 66.615 2.495 66.785 3.225 ;
      RECT 66.255 3.615 66.545 3.785 ;
      RECT 66.255 2.575 66.425 3.785 ;
      RECT 66.055 2.575 66.425 2.745 ;
      RECT 63.915 1.74 64.085 2.935 ;
      RECT 63.915 1.74 64.38 1.91 ;
      RECT 63.915 6.97 64.38 7.14 ;
      RECT 63.915 5.945 64.085 7.14 ;
      RECT 62.925 1.74 63.095 2.935 ;
      RECT 62.925 1.74 63.39 1.91 ;
      RECT 62.925 6.97 63.39 7.14 ;
      RECT 62.925 5.945 63.095 7.14 ;
      RECT 61.07 2.635 61.24 3.865 ;
      RECT 61.125 0.855 61.295 2.805 ;
      RECT 61.07 0.575 61.24 1.025 ;
      RECT 61.07 7.855 61.24 8.305 ;
      RECT 61.125 6.075 61.295 8.025 ;
      RECT 61.07 5.015 61.24 6.245 ;
      RECT 60.55 0.575 60.72 3.865 ;
      RECT 60.55 2.075 60.955 2.405 ;
      RECT 60.55 1.235 60.955 1.565 ;
      RECT 60.55 5.015 60.72 8.305 ;
      RECT 60.55 7.315 60.955 7.645 ;
      RECT 60.55 6.475 60.955 6.805 ;
      RECT 57.85 1.835 58.02 2.105 ;
      RECT 57.85 1.835 58.58 2.005 ;
      RECT 58.33 2.575 58.5 2.945 ;
      RECT 58.01 2.575 58.5 2.745 ;
      RECT 57.77 3.225 58.1 3.395 ;
      RECT 57.01 3.055 58.02 3.225 ;
      RECT 57.01 2.575 57.18 3.225 ;
      RECT 57.13 2.495 57.3 2.825 ;
      RECT 56.29 3.225 56.62 3.395 ;
      RECT 54.37 3.225 55.66 3.395 ;
      RECT 55.41 3.14 56.54 3.31 ;
      RECT 56.13 2.215 56.54 2.385 ;
      RECT 56.37 1.755 56.54 2.385 ;
      RECT 56.37 2.575 56.54 2.945 ;
      RECT 56.05 2.575 56.54 2.745 ;
      RECT 55.455 7.855 55.625 8.305 ;
      RECT 55.51 6.075 55.68 8.025 ;
      RECT 55.455 5.015 55.625 6.245 ;
      RECT 54.935 5.015 55.105 8.305 ;
      RECT 54.935 7.315 55.34 7.645 ;
      RECT 54.935 6.475 55.34 6.805 ;
      RECT 53.61 2.575 54.94 2.745 ;
      RECT 54.69 2.495 54.86 2.745 ;
      RECT 53.69 2.175 53.86 2.385 ;
      RECT 53.69 2.175 54.18 2.345 ;
      RECT 52.37 3.335 52.66 3.505 ;
      RECT 52.37 2.575 52.54 3.505 ;
      RECT 52.17 2.575 52.54 2.745 ;
      RECT 51.17 2.575 51.66 2.745 ;
      RECT 51.49 2.495 51.66 2.745 ;
      RECT 51.25 3.335 51.66 3.505 ;
      RECT 51.49 3.145 51.66 3.505 ;
      RECT 50.29 3.055 50.94 3.225 ;
      RECT 50.29 2.495 50.46 3.225 ;
      RECT 49.93 3.615 50.22 3.785 ;
      RECT 49.93 2.575 50.1 3.785 ;
      RECT 49.73 2.575 50.1 2.745 ;
      RECT 47.59 1.74 47.76 2.935 ;
      RECT 47.59 1.74 48.055 1.91 ;
      RECT 47.59 6.97 48.055 7.14 ;
      RECT 47.59 5.945 47.76 7.14 ;
      RECT 46.6 1.74 46.77 2.935 ;
      RECT 46.6 1.74 47.065 1.91 ;
      RECT 46.6 6.97 47.065 7.14 ;
      RECT 46.6 5.945 46.77 7.14 ;
      RECT 44.745 2.635 44.915 3.865 ;
      RECT 44.8 0.855 44.97 2.805 ;
      RECT 44.745 0.575 44.915 1.025 ;
      RECT 44.745 7.855 44.915 8.305 ;
      RECT 44.8 6.075 44.97 8.025 ;
      RECT 44.745 5.015 44.915 6.245 ;
      RECT 44.225 0.575 44.395 3.865 ;
      RECT 44.225 2.075 44.63 2.405 ;
      RECT 44.225 1.235 44.63 1.565 ;
      RECT 44.225 5.015 44.395 8.305 ;
      RECT 44.225 7.315 44.63 7.645 ;
      RECT 44.225 6.475 44.63 6.805 ;
      RECT 41.525 1.835 41.695 2.105 ;
      RECT 41.525 1.835 42.255 2.005 ;
      RECT 42.005 2.575 42.175 2.945 ;
      RECT 41.685 2.575 42.175 2.745 ;
      RECT 41.445 3.225 41.775 3.395 ;
      RECT 40.685 3.055 41.695 3.225 ;
      RECT 40.685 2.575 40.855 3.225 ;
      RECT 40.805 2.495 40.975 2.825 ;
      RECT 39.965 3.225 40.295 3.395 ;
      RECT 38.045 3.225 39.335 3.395 ;
      RECT 39.085 3.14 40.215 3.31 ;
      RECT 39.805 2.215 40.215 2.385 ;
      RECT 40.045 1.755 40.215 2.385 ;
      RECT 40.045 2.575 40.215 2.945 ;
      RECT 39.725 2.575 40.215 2.745 ;
      RECT 39.13 7.855 39.3 8.305 ;
      RECT 39.185 6.075 39.355 8.025 ;
      RECT 39.13 5.015 39.3 6.245 ;
      RECT 38.61 5.015 38.78 8.305 ;
      RECT 38.61 7.315 39.015 7.645 ;
      RECT 38.61 6.475 39.015 6.805 ;
      RECT 37.285 2.575 38.615 2.745 ;
      RECT 38.365 2.495 38.535 2.745 ;
      RECT 37.365 2.175 37.535 2.385 ;
      RECT 37.365 2.175 37.855 2.345 ;
      RECT 36.045 3.335 36.335 3.505 ;
      RECT 36.045 2.575 36.215 3.505 ;
      RECT 35.845 2.575 36.215 2.745 ;
      RECT 34.845 2.575 35.335 2.745 ;
      RECT 35.165 2.495 35.335 2.745 ;
      RECT 34.925 3.335 35.335 3.505 ;
      RECT 35.165 3.145 35.335 3.505 ;
      RECT 33.965 3.055 34.615 3.225 ;
      RECT 33.965 2.495 34.135 3.225 ;
      RECT 33.605 3.615 33.895 3.785 ;
      RECT 33.605 2.575 33.775 3.785 ;
      RECT 33.405 2.575 33.775 2.745 ;
      RECT 31.265 1.74 31.435 2.935 ;
      RECT 31.265 1.74 31.73 1.91 ;
      RECT 31.265 6.97 31.73 7.14 ;
      RECT 31.265 5.945 31.435 7.14 ;
      RECT 30.275 1.74 30.445 2.935 ;
      RECT 30.275 1.74 30.74 1.91 ;
      RECT 30.275 6.97 30.74 7.14 ;
      RECT 30.275 5.945 30.445 7.14 ;
      RECT 28.42 2.635 28.59 3.865 ;
      RECT 28.475 0.855 28.645 2.805 ;
      RECT 28.42 0.575 28.59 1.025 ;
      RECT 28.42 7.855 28.59 8.305 ;
      RECT 28.475 6.075 28.645 8.025 ;
      RECT 28.42 5.015 28.59 6.245 ;
      RECT 27.9 0.575 28.07 3.865 ;
      RECT 27.9 2.075 28.305 2.405 ;
      RECT 27.9 1.235 28.305 1.565 ;
      RECT 27.9 5.015 28.07 8.305 ;
      RECT 27.9 7.315 28.305 7.645 ;
      RECT 27.9 6.475 28.305 6.805 ;
      RECT 25.2 1.835 25.37 2.105 ;
      RECT 25.2 1.835 25.93 2.005 ;
      RECT 25.68 2.575 25.85 2.945 ;
      RECT 25.36 2.575 25.85 2.745 ;
      RECT 25.12 3.225 25.45 3.395 ;
      RECT 24.36 3.055 25.37 3.225 ;
      RECT 24.36 2.575 24.53 3.225 ;
      RECT 24.48 2.495 24.65 2.825 ;
      RECT 23.64 3.225 23.97 3.395 ;
      RECT 21.72 3.225 23.01 3.395 ;
      RECT 22.76 3.14 23.89 3.31 ;
      RECT 23.48 2.215 23.89 2.385 ;
      RECT 23.72 1.755 23.89 2.385 ;
      RECT 23.72 2.575 23.89 2.945 ;
      RECT 23.4 2.575 23.89 2.745 ;
      RECT 22.805 7.855 22.975 8.305 ;
      RECT 22.86 6.075 23.03 8.025 ;
      RECT 22.805 5.015 22.975 6.245 ;
      RECT 22.285 5.015 22.455 8.305 ;
      RECT 22.285 7.315 22.69 7.645 ;
      RECT 22.285 6.475 22.69 6.805 ;
      RECT 20.96 2.575 22.29 2.745 ;
      RECT 22.04 2.495 22.21 2.745 ;
      RECT 21.04 2.175 21.21 2.385 ;
      RECT 21.04 2.175 21.53 2.345 ;
      RECT 19.72 3.335 20.01 3.505 ;
      RECT 19.72 2.575 19.89 3.505 ;
      RECT 19.52 2.575 19.89 2.745 ;
      RECT 18.52 2.575 19.01 2.745 ;
      RECT 18.84 2.495 19.01 2.745 ;
      RECT 18.6 3.335 19.01 3.505 ;
      RECT 18.84 3.145 19.01 3.505 ;
      RECT 17.64 3.055 18.29 3.225 ;
      RECT 17.64 2.495 17.81 3.225 ;
      RECT 17.28 3.615 17.57 3.785 ;
      RECT 17.28 2.575 17.45 3.785 ;
      RECT 17.08 2.575 17.45 2.745 ;
      RECT 14.94 1.74 15.11 2.935 ;
      RECT 14.94 1.74 15.405 1.91 ;
      RECT 14.94 6.97 15.405 7.14 ;
      RECT 14.94 5.945 15.11 7.14 ;
      RECT 13.95 1.74 14.12 2.935 ;
      RECT 13.95 1.74 14.415 1.91 ;
      RECT 13.95 6.97 14.415 7.14 ;
      RECT 13.95 5.945 14.12 7.14 ;
      RECT 12.095 2.635 12.265 3.865 ;
      RECT 12.15 0.855 12.32 2.805 ;
      RECT 12.095 0.575 12.265 1.025 ;
      RECT 12.095 7.855 12.265 8.305 ;
      RECT 12.15 6.075 12.32 8.025 ;
      RECT 12.095 5.015 12.265 6.245 ;
      RECT 11.575 0.575 11.745 3.865 ;
      RECT 11.575 2.075 11.98 2.405 ;
      RECT 11.575 1.235 11.98 1.565 ;
      RECT 11.575 5.015 11.745 8.305 ;
      RECT 11.575 7.315 11.98 7.645 ;
      RECT 11.575 6.475 11.98 6.805 ;
      RECT 8.875 1.835 9.045 2.105 ;
      RECT 8.875 1.835 9.605 2.005 ;
      RECT 9.355 2.575 9.525 2.945 ;
      RECT 9.035 2.575 9.525 2.745 ;
      RECT 8.795 3.225 9.125 3.395 ;
      RECT 8.035 3.055 9.045 3.225 ;
      RECT 8.035 2.575 8.205 3.225 ;
      RECT 8.155 2.495 8.325 2.825 ;
      RECT 7.315 3.225 7.645 3.395 ;
      RECT 5.395 3.225 6.685 3.395 ;
      RECT 6.435 3.14 7.565 3.31 ;
      RECT 7.155 2.215 7.565 2.385 ;
      RECT 7.395 1.755 7.565 2.385 ;
      RECT 7.395 2.575 7.565 2.945 ;
      RECT 7.075 2.575 7.565 2.745 ;
      RECT 6.48 7.855 6.65 8.305 ;
      RECT 6.535 6.075 6.705 8.025 ;
      RECT 6.48 5.015 6.65 6.245 ;
      RECT 5.96 5.015 6.13 8.305 ;
      RECT 5.96 7.315 6.365 7.645 ;
      RECT 5.96 6.475 6.365 6.805 ;
      RECT 4.635 2.575 5.965 2.745 ;
      RECT 5.715 2.495 5.885 2.745 ;
      RECT 4.715 2.175 4.885 2.385 ;
      RECT 4.715 2.175 5.205 2.345 ;
      RECT 3.395 3.335 3.685 3.505 ;
      RECT 3.395 2.575 3.565 3.505 ;
      RECT 3.195 2.575 3.565 2.745 ;
      RECT 2.195 2.575 2.685 2.745 ;
      RECT 2.515 2.495 2.685 2.745 ;
      RECT 2.275 3.335 2.685 3.505 ;
      RECT 2.515 3.145 2.685 3.505 ;
      RECT 1.315 3.055 1.965 3.225 ;
      RECT 1.315 2.495 1.485 3.225 ;
      RECT 0.955 3.615 1.245 3.785 ;
      RECT 0.955 2.575 1.125 3.785 ;
      RECT 0.755 2.575 1.125 2.745 ;
      RECT -2.1 7.855 -1.93 8.305 ;
      RECT -2.045 6.075 -1.875 8.025 ;
      RECT -2.1 5.015 -1.93 6.245 ;
      RECT -2.62 5.015 -2.45 8.305 ;
      RECT -2.62 7.315 -2.215 7.645 ;
      RECT -2.62 6.475 -2.215 6.805 ;
      RECT 80.61 0.575 80.78 1.085 ;
      RECT 80.61 2.395 80.78 3.865 ;
      RECT 80.61 5.015 80.78 6.485 ;
      RECT 80.61 7.795 80.78 8.305 ;
      RECT 79.62 0.575 79.79 1.085 ;
      RECT 79.62 2.395 79.79 3.865 ;
      RECT 79.62 5.015 79.79 6.485 ;
      RECT 79.62 7.795 79.79 8.305 ;
      RECT 78.255 0.575 78.425 3.865 ;
      RECT 78.255 5.015 78.425 8.305 ;
      RECT 77.825 0.575 77.995 1.085 ;
      RECT 77.825 1.655 77.995 3.865 ;
      RECT 77.825 5.015 77.995 7.225 ;
      RECT 77.825 7.795 77.995 8.305 ;
      RECT 76.455 1.66 76.625 2.935 ;
      RECT 76.455 5.945 76.625 7.22 ;
      RECT 73.935 2.495 74.105 2.825 ;
      RECT 73.215 1.755 73.385 2.105 ;
      RECT 73.215 3.485 73.385 3.815 ;
      RECT 72.64 5.015 72.81 8.305 ;
      RECT 72.215 3.485 72.385 3.815 ;
      RECT 72.21 5.015 72.38 7.225 ;
      RECT 72.21 7.795 72.38 8.305 ;
      RECT 71.975 2.495 72.145 2.945 ;
      RECT 71.495 2.495 71.665 2.825 ;
      RECT 70.84 5.945 71.01 7.22 ;
      RECT 70.775 1.755 70.945 2.105 ;
      RECT 69.775 3.145 69.945 3.505 ;
      RECT 69.535 2.495 69.705 2.945 ;
      RECT 69.055 2.495 69.225 2.825 ;
      RECT 68.815 1.755 68.985 2.105 ;
      RECT 68.335 3.055 68.505 3.475 ;
      RECT 67.335 1.755 67.505 2.105 ;
      RECT 67.095 2.495 67.265 2.825 ;
      RECT 66.375 1.755 66.545 2.105 ;
      RECT 65.895 3.055 66.065 3.475 ;
      RECT 64.285 0.575 64.455 1.085 ;
      RECT 64.285 2.395 64.455 3.865 ;
      RECT 64.285 5.015 64.455 6.485 ;
      RECT 64.285 7.795 64.455 8.305 ;
      RECT 63.295 0.575 63.465 1.085 ;
      RECT 63.295 2.395 63.465 3.865 ;
      RECT 63.295 5.015 63.465 6.485 ;
      RECT 63.295 7.795 63.465 8.305 ;
      RECT 61.93 0.575 62.1 3.865 ;
      RECT 61.93 5.015 62.1 8.305 ;
      RECT 61.5 0.575 61.67 1.085 ;
      RECT 61.5 1.655 61.67 3.865 ;
      RECT 61.5 5.015 61.67 7.225 ;
      RECT 61.5 7.795 61.67 8.305 ;
      RECT 60.13 1.66 60.3 2.935 ;
      RECT 60.13 5.945 60.3 7.22 ;
      RECT 57.61 2.495 57.78 2.825 ;
      RECT 56.89 1.755 57.06 2.105 ;
      RECT 56.89 3.485 57.06 3.815 ;
      RECT 56.315 5.015 56.485 8.305 ;
      RECT 55.89 3.485 56.06 3.815 ;
      RECT 55.885 5.015 56.055 7.225 ;
      RECT 55.885 7.795 56.055 8.305 ;
      RECT 55.65 2.495 55.82 2.945 ;
      RECT 55.17 2.495 55.34 2.825 ;
      RECT 54.515 5.945 54.685 7.22 ;
      RECT 54.45 1.755 54.62 2.105 ;
      RECT 53.45 3.145 53.62 3.505 ;
      RECT 53.21 2.495 53.38 2.945 ;
      RECT 52.73 2.495 52.9 2.825 ;
      RECT 52.49 1.755 52.66 2.105 ;
      RECT 52.01 3.055 52.18 3.475 ;
      RECT 51.01 1.755 51.18 2.105 ;
      RECT 50.77 2.495 50.94 2.825 ;
      RECT 50.05 1.755 50.22 2.105 ;
      RECT 49.57 3.055 49.74 3.475 ;
      RECT 47.96 0.575 48.13 1.085 ;
      RECT 47.96 2.395 48.13 3.865 ;
      RECT 47.96 5.015 48.13 6.485 ;
      RECT 47.96 7.795 48.13 8.305 ;
      RECT 46.97 0.575 47.14 1.085 ;
      RECT 46.97 2.395 47.14 3.865 ;
      RECT 46.97 5.015 47.14 6.485 ;
      RECT 46.97 7.795 47.14 8.305 ;
      RECT 45.605 0.575 45.775 3.865 ;
      RECT 45.605 5.015 45.775 8.305 ;
      RECT 45.175 0.575 45.345 1.085 ;
      RECT 45.175 1.655 45.345 3.865 ;
      RECT 45.175 5.015 45.345 7.225 ;
      RECT 45.175 7.795 45.345 8.305 ;
      RECT 43.805 1.66 43.975 2.935 ;
      RECT 43.805 5.945 43.975 7.22 ;
      RECT 41.285 2.495 41.455 2.825 ;
      RECT 40.565 1.755 40.735 2.105 ;
      RECT 40.565 3.485 40.735 3.815 ;
      RECT 39.99 5.015 40.16 8.305 ;
      RECT 39.565 3.485 39.735 3.815 ;
      RECT 39.56 5.015 39.73 7.225 ;
      RECT 39.56 7.795 39.73 8.305 ;
      RECT 39.325 2.495 39.495 2.945 ;
      RECT 38.845 2.495 39.015 2.825 ;
      RECT 38.19 5.945 38.36 7.22 ;
      RECT 38.125 1.755 38.295 2.105 ;
      RECT 37.125 3.145 37.295 3.505 ;
      RECT 36.885 2.495 37.055 2.945 ;
      RECT 36.405 2.495 36.575 2.825 ;
      RECT 36.165 1.755 36.335 2.105 ;
      RECT 35.685 3.055 35.855 3.475 ;
      RECT 34.685 1.755 34.855 2.105 ;
      RECT 34.445 2.495 34.615 2.825 ;
      RECT 33.725 1.755 33.895 2.105 ;
      RECT 33.245 3.055 33.415 3.475 ;
      RECT 31.635 0.575 31.805 1.085 ;
      RECT 31.635 2.395 31.805 3.865 ;
      RECT 31.635 5.015 31.805 6.485 ;
      RECT 31.635 7.795 31.805 8.305 ;
      RECT 30.645 0.575 30.815 1.085 ;
      RECT 30.645 2.395 30.815 3.865 ;
      RECT 30.645 5.015 30.815 6.485 ;
      RECT 30.645 7.795 30.815 8.305 ;
      RECT 29.28 0.575 29.45 3.865 ;
      RECT 29.28 5.015 29.45 8.305 ;
      RECT 28.85 0.575 29.02 1.085 ;
      RECT 28.85 1.655 29.02 3.865 ;
      RECT 28.85 5.015 29.02 7.225 ;
      RECT 28.85 7.795 29.02 8.305 ;
      RECT 27.48 1.66 27.65 2.935 ;
      RECT 27.48 5.945 27.65 7.22 ;
      RECT 24.96 2.495 25.13 2.825 ;
      RECT 24.24 1.755 24.41 2.105 ;
      RECT 24.24 3.485 24.41 3.815 ;
      RECT 23.665 5.015 23.835 8.305 ;
      RECT 23.24 3.485 23.41 3.815 ;
      RECT 23.235 5.015 23.405 7.225 ;
      RECT 23.235 7.795 23.405 8.305 ;
      RECT 23 2.495 23.17 2.945 ;
      RECT 22.52 2.495 22.69 2.825 ;
      RECT 21.865 5.945 22.035 7.22 ;
      RECT 21.8 1.755 21.97 2.105 ;
      RECT 20.8 3.145 20.97 3.505 ;
      RECT 20.56 2.495 20.73 2.945 ;
      RECT 20.08 2.495 20.25 2.825 ;
      RECT 19.84 1.755 20.01 2.105 ;
      RECT 19.36 3.055 19.53 3.475 ;
      RECT 18.36 1.755 18.53 2.105 ;
      RECT 18.12 2.495 18.29 2.825 ;
      RECT 17.4 1.755 17.57 2.105 ;
      RECT 16.92 3.055 17.09 3.475 ;
      RECT 15.31 0.575 15.48 1.085 ;
      RECT 15.31 2.395 15.48 3.865 ;
      RECT 15.31 5.015 15.48 6.485 ;
      RECT 15.31 7.795 15.48 8.305 ;
      RECT 14.32 0.575 14.49 1.085 ;
      RECT 14.32 2.395 14.49 3.865 ;
      RECT 14.32 5.015 14.49 6.485 ;
      RECT 14.32 7.795 14.49 8.305 ;
      RECT 12.955 0.575 13.125 3.865 ;
      RECT 12.955 5.015 13.125 8.305 ;
      RECT 12.525 0.575 12.695 1.085 ;
      RECT 12.525 1.655 12.695 3.865 ;
      RECT 12.525 5.015 12.695 7.225 ;
      RECT 12.525 7.795 12.695 8.305 ;
      RECT 11.155 1.66 11.325 2.935 ;
      RECT 11.155 5.945 11.325 7.22 ;
      RECT 8.635 2.495 8.805 2.825 ;
      RECT 7.915 1.755 8.085 2.105 ;
      RECT 7.915 3.485 8.085 3.815 ;
      RECT 7.34 5.015 7.51 8.305 ;
      RECT 6.915 3.485 7.085 3.815 ;
      RECT 6.91 5.015 7.08 7.225 ;
      RECT 6.91 7.795 7.08 8.305 ;
      RECT 6.675 2.495 6.845 2.945 ;
      RECT 6.195 2.495 6.365 2.825 ;
      RECT 5.54 5.945 5.71 7.22 ;
      RECT 5.475 1.755 5.645 2.105 ;
      RECT 4.475 3.145 4.645 3.505 ;
      RECT 4.235 2.495 4.405 2.945 ;
      RECT 3.755 2.495 3.925 2.825 ;
      RECT 3.515 1.755 3.685 2.105 ;
      RECT 3.035 3.055 3.205 3.475 ;
      RECT 2.035 1.755 2.205 2.105 ;
      RECT 1.795 2.495 1.965 2.825 ;
      RECT 1.075 1.755 1.245 2.105 ;
      RECT 0.595 3.055 0.765 3.475 ;
      RECT -1.67 5.015 -1.5 7.225 ;
      RECT -1.67 7.795 -1.5 8.305 ;
      RECT -3.04 5.945 -2.87 7.22 ;
  END
END sky130_osu_ring_oscillator_mpr2ea_8_b0r1

MACRO sky130_osu_ring_oscillator_mpr2ea_8_b0r2
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 3.27 0 ;
  SIZE 84.42 BY 8.88 ;
  SYMMETRY X Y R90 ;
  SITE CoreSite ;
  OBS
    LAYER met3 ;
      RECT 72.13 7.055 72.5 7.425 ;
      RECT 72.13 7.09 74.115 7.39 ;
      RECT 73.815 2.28 74.115 7.39 ;
      RECT 70.815 2.015 71.145 2.745 ;
      RECT 69.935 2.015 70.265 2.745 ;
      RECT 73.015 2.28 74.305 2.58 ;
      RECT 73.975 1.85 74.305 2.58 ;
      RECT 69.935 2.28 72.075 2.58 ;
      RECT 71.775 1.965 72.075 2.58 ;
      RECT 73.015 1.98 73.32 2.58 ;
      RECT 71.775 1.965 73.135 2.275 ;
      RECT 70.435 3.535 70.765 3.865 ;
      RECT 69.23 3.55 70.765 3.85 ;
      RECT 69.23 2.43 69.53 3.85 ;
      RECT 68.975 2.415 69.305 2.745 ;
      RECT 55.805 7.055 56.175 7.425 ;
      RECT 55.805 7.09 57.79 7.39 ;
      RECT 57.49 2.28 57.79 7.39 ;
      RECT 54.49 2.015 54.82 2.745 ;
      RECT 53.61 2.015 53.94 2.745 ;
      RECT 56.69 2.28 57.98 2.58 ;
      RECT 57.65 1.85 57.98 2.58 ;
      RECT 53.61 2.28 55.75 2.58 ;
      RECT 55.45 1.965 55.75 2.58 ;
      RECT 56.69 1.98 56.995 2.58 ;
      RECT 55.45 1.965 56.81 2.275 ;
      RECT 54.11 3.535 54.44 3.865 ;
      RECT 52.905 3.55 54.44 3.85 ;
      RECT 52.905 2.43 53.205 3.85 ;
      RECT 52.65 2.415 52.98 2.745 ;
      RECT 39.48 7.055 39.85 7.425 ;
      RECT 39.48 7.09 41.465 7.39 ;
      RECT 41.165 2.28 41.465 7.39 ;
      RECT 38.165 2.015 38.495 2.745 ;
      RECT 37.285 2.015 37.615 2.745 ;
      RECT 40.365 2.28 41.655 2.58 ;
      RECT 41.325 1.85 41.655 2.58 ;
      RECT 37.285 2.28 39.425 2.58 ;
      RECT 39.125 1.965 39.425 2.58 ;
      RECT 40.365 1.98 40.67 2.58 ;
      RECT 39.125 1.965 40.485 2.275 ;
      RECT 37.785 3.535 38.115 3.865 ;
      RECT 36.58 3.55 38.115 3.85 ;
      RECT 36.58 2.43 36.88 3.85 ;
      RECT 36.325 2.415 36.655 2.745 ;
      RECT 23.155 7.055 23.525 7.425 ;
      RECT 23.155 7.09 25.14 7.39 ;
      RECT 24.84 2.28 25.14 7.39 ;
      RECT 21.84 2.015 22.17 2.745 ;
      RECT 20.96 2.015 21.29 2.745 ;
      RECT 24.04 2.28 25.33 2.58 ;
      RECT 25 1.85 25.33 2.58 ;
      RECT 20.96 2.28 23.1 2.58 ;
      RECT 22.8 1.965 23.1 2.58 ;
      RECT 24.04 1.98 24.345 2.58 ;
      RECT 22.8 1.965 24.16 2.275 ;
      RECT 21.46 3.535 21.79 3.865 ;
      RECT 20.255 3.55 21.79 3.85 ;
      RECT 20.255 2.43 20.555 3.85 ;
      RECT 20 2.415 20.33 2.745 ;
      RECT 6.83 7.055 7.2 7.425 ;
      RECT 6.83 7.09 8.815 7.39 ;
      RECT 8.515 2.28 8.815 7.39 ;
      RECT 5.515 2.015 5.845 2.745 ;
      RECT 4.635 2.015 4.965 2.745 ;
      RECT 7.715 2.28 9.005 2.58 ;
      RECT 8.675 1.85 9.005 2.58 ;
      RECT 4.635 2.28 6.775 2.58 ;
      RECT 6.475 1.965 6.775 2.58 ;
      RECT 7.715 1.98 8.02 2.58 ;
      RECT 6.475 1.965 7.835 2.275 ;
      RECT 5.135 3.535 5.465 3.865 ;
      RECT 3.93 3.55 5.465 3.85 ;
      RECT 3.93 2.43 4.23 3.85 ;
      RECT 3.675 2.415 4.005 2.745 ;
      RECT 74.455 2.975 74.785 3.705 ;
      RECT 72.375 2.575 72.705 3.305 ;
      RECT 68.255 2.415 68.585 3.145 ;
      RECT 67.255 1.855 67.585 2.585 ;
      RECT 65.815 2.575 66.145 3.305 ;
      RECT 58.13 2.975 58.46 3.705 ;
      RECT 56.05 2.575 56.38 3.305 ;
      RECT 51.93 2.415 52.26 3.145 ;
      RECT 50.93 1.855 51.26 2.585 ;
      RECT 49.49 2.575 49.82 3.305 ;
      RECT 41.805 2.975 42.135 3.705 ;
      RECT 39.725 2.575 40.055 3.305 ;
      RECT 35.605 2.415 35.935 3.145 ;
      RECT 34.605 1.855 34.935 2.585 ;
      RECT 33.165 2.575 33.495 3.305 ;
      RECT 25.48 2.975 25.81 3.705 ;
      RECT 23.4 2.575 23.73 3.305 ;
      RECT 19.28 2.415 19.61 3.145 ;
      RECT 18.28 1.855 18.61 2.585 ;
      RECT 16.84 2.575 17.17 3.305 ;
      RECT 9.155 2.975 9.485 3.705 ;
      RECT 7.075 2.575 7.405 3.305 ;
      RECT 2.955 2.415 3.285 3.145 ;
      RECT 1.955 1.855 2.285 2.585 ;
      RECT 0.515 2.575 0.845 3.305 ;
    LAYER via2 ;
      RECT 74.52 3.04 74.72 3.24 ;
      RECT 74.04 2.315 74.24 2.515 ;
      RECT 72.44 3.04 72.64 3.24 ;
      RECT 72.215 7.14 72.415 7.34 ;
      RECT 70.88 2.48 71.08 2.68 ;
      RECT 70.5 3.6 70.7 3.8 ;
      RECT 70 2.48 70.2 2.68 ;
      RECT 69.04 2.48 69.24 2.68 ;
      RECT 68.32 2.48 68.52 2.68 ;
      RECT 67.32 1.92 67.52 2.12 ;
      RECT 65.88 3.04 66.08 3.24 ;
      RECT 58.195 3.04 58.395 3.24 ;
      RECT 57.715 2.315 57.915 2.515 ;
      RECT 56.115 3.04 56.315 3.24 ;
      RECT 55.89 7.14 56.09 7.34 ;
      RECT 54.555 2.48 54.755 2.68 ;
      RECT 54.175 3.6 54.375 3.8 ;
      RECT 53.675 2.48 53.875 2.68 ;
      RECT 52.715 2.48 52.915 2.68 ;
      RECT 51.995 2.48 52.195 2.68 ;
      RECT 50.995 1.92 51.195 2.12 ;
      RECT 49.555 3.04 49.755 3.24 ;
      RECT 41.87 3.04 42.07 3.24 ;
      RECT 41.39 2.315 41.59 2.515 ;
      RECT 39.79 3.04 39.99 3.24 ;
      RECT 39.565 7.14 39.765 7.34 ;
      RECT 38.23 2.48 38.43 2.68 ;
      RECT 37.85 3.6 38.05 3.8 ;
      RECT 37.35 2.48 37.55 2.68 ;
      RECT 36.39 2.48 36.59 2.68 ;
      RECT 35.67 2.48 35.87 2.68 ;
      RECT 34.67 1.92 34.87 2.12 ;
      RECT 33.23 3.04 33.43 3.24 ;
      RECT 25.545 3.04 25.745 3.24 ;
      RECT 25.065 2.315 25.265 2.515 ;
      RECT 23.465 3.04 23.665 3.24 ;
      RECT 23.24 7.14 23.44 7.34 ;
      RECT 21.905 2.48 22.105 2.68 ;
      RECT 21.525 3.6 21.725 3.8 ;
      RECT 21.025 2.48 21.225 2.68 ;
      RECT 20.065 2.48 20.265 2.68 ;
      RECT 19.345 2.48 19.545 2.68 ;
      RECT 18.345 1.92 18.545 2.12 ;
      RECT 16.905 3.04 17.105 3.24 ;
      RECT 9.22 3.04 9.42 3.24 ;
      RECT 8.74 2.315 8.94 2.515 ;
      RECT 7.14 3.04 7.34 3.24 ;
      RECT 6.915 7.14 7.115 7.34 ;
      RECT 5.58 2.48 5.78 2.68 ;
      RECT 5.2 3.6 5.4 3.8 ;
      RECT 4.7 2.48 4.9 2.68 ;
      RECT 3.74 2.48 3.94 2.68 ;
      RECT 3.02 2.48 3.22 2.68 ;
      RECT 2.02 1.92 2.22 2.12 ;
      RECT 0.58 3.04 0.78 3.24 ;
    LAYER met2 ;
      RECT -2.045 8.4 80.78 8.57 ;
      RECT 80.61 7.275 80.78 8.57 ;
      RECT -2.045 6.255 -1.875 8.57 ;
      RECT 80.58 7.275 80.93 7.625 ;
      RECT -2.105 6.255 -1.815 6.605 ;
      RECT 77.42 6.22 77.74 6.545 ;
      RECT 77.45 5.695 77.62 6.545 ;
      RECT 77.45 5.695 77.625 6.045 ;
      RECT 77.45 5.695 78.425 5.87 ;
      RECT 78.25 1.965 78.425 5.87 ;
      RECT 78.195 1.965 78.545 2.315 ;
      RECT 78.22 6.655 78.545 6.98 ;
      RECT 77.105 6.745 78.545 6.915 ;
      RECT 77.105 2.395 77.265 6.915 ;
      RECT 77.42 2.365 77.74 2.685 ;
      RECT 77.105 2.395 77.74 2.565 ;
      RECT 76.37 5.84 76.71 6.19 ;
      RECT 76.455 2.705 76.625 6.19 ;
      RECT 76.38 2.705 76.72 3.055 ;
      RECT 65.84 2.955 66.12 3.325 ;
      RECT 65.895 1.29 66.065 3.325 ;
      RECT 75.89 1.29 76.06 1.815 ;
      RECT 75.8 1.46 76.14 1.81 ;
      RECT 65.895 1.29 76.06 1.46 ;
      RECT 72.52 2.395 72.8 2.765 ;
      RECT 71.45 2.42 71.71 2.74 ;
      RECT 74 2.23 74.28 2.6 ;
      RECT 74.61 2.14 74.87 2.46 ;
      RECT 71.51 1.58 71.65 2.74 ;
      RECT 72.59 1.58 72.73 2.765 ;
      RECT 73.71 2.23 74.87 2.37 ;
      RECT 73.71 1.58 73.85 2.37 ;
      RECT 71.51 1.58 73.85 1.72 ;
      RECT 74.48 2.955 74.76 3.325 ;
      RECT 74.49 2.7 74.75 3.325 ;
      RECT 71.54 3.72 73.715 3.885 ;
      RECT 73.57 2.6 73.715 3.885 ;
      RECT 70.46 3.515 70.74 3.885 ;
      RECT 70.46 3.63 71.68 3.77 ;
      RECT 73.29 2.6 73.715 2.74 ;
      RECT 73.29 2.42 73.55 2.74 ;
      RECT 66.63 4 70.29 4.14 ;
      RECT 70.15 3.185 70.29 4.14 ;
      RECT 66.63 3.07 66.77 4.14 ;
      RECT 73.17 3.26 73.43 3.58 ;
      RECT 70.15 3.185 72.68 3.325 ;
      RECT 72.4 2.955 72.68 3.325 ;
      RECT 66.63 3.07 67.08 3.325 ;
      RECT 66.8 2.955 67.08 3.325 ;
      RECT 73.17 3.07 73.37 3.58 ;
      RECT 72.4 3.07 73.37 3.21 ;
      RECT 72.97 1.86 73.11 3.21 ;
      RECT 72.91 1.86 73.17 2.18 ;
      RECT 64.23 6.655 64.58 7.005 ;
      RECT 72.785 6.61 73.135 6.96 ;
      RECT 64.23 6.685 73.135 6.885 ;
      RECT 66.81 2.42 67.07 2.74 ;
      RECT 66.81 2.51 67.85 2.65 ;
      RECT 67.71 1.72 67.85 2.65 ;
      RECT 70.47 1.86 70.73 2.18 ;
      RECT 67.71 1.72 70.67 1.86 ;
      RECT 69.85 2.7 70.11 3.02 ;
      RECT 69.85 2.7 70.17 2.93 ;
      RECT 69.96 2.395 70.24 2.765 ;
      RECT 69.55 3.26 69.87 3.58 ;
      RECT 69.55 2.14 69.69 3.58 ;
      RECT 69.49 2.14 69.75 2.46 ;
      RECT 67.05 3.54 67.31 3.86 ;
      RECT 67.05 3.63 68.73 3.77 ;
      RECT 68.59 3.35 68.73 3.77 ;
      RECT 68.59 3.35 69.03 3.58 ;
      RECT 68.77 3.26 69.03 3.58 ;
      RECT 68.09 2.42 68.49 2.93 ;
      RECT 68.28 2.395 68.56 2.765 ;
      RECT 68.03 2.42 68.56 2.74 ;
      RECT 61.095 6.22 61.415 6.545 ;
      RECT 61.125 5.695 61.295 6.545 ;
      RECT 61.125 5.695 61.3 6.045 ;
      RECT 61.125 5.695 62.1 5.87 ;
      RECT 61.925 1.965 62.1 5.87 ;
      RECT 61.87 1.965 62.22 2.315 ;
      RECT 61.895 6.655 62.22 6.98 ;
      RECT 60.78 6.745 62.22 6.915 ;
      RECT 60.78 2.395 60.94 6.915 ;
      RECT 61.095 2.365 61.415 2.685 ;
      RECT 60.78 2.395 61.415 2.565 ;
      RECT 60.045 5.84 60.385 6.19 ;
      RECT 60.13 2.705 60.3 6.19 ;
      RECT 60.055 2.705 60.395 3.055 ;
      RECT 49.515 2.955 49.795 3.325 ;
      RECT 49.57 1.29 49.74 3.325 ;
      RECT 59.565 1.29 59.735 1.815 ;
      RECT 59.475 1.46 59.815 1.81 ;
      RECT 49.57 1.29 59.735 1.46 ;
      RECT 56.195 2.395 56.475 2.765 ;
      RECT 55.125 2.42 55.385 2.74 ;
      RECT 57.675 2.23 57.955 2.6 ;
      RECT 58.285 2.14 58.545 2.46 ;
      RECT 55.185 1.58 55.325 2.74 ;
      RECT 56.265 1.58 56.405 2.765 ;
      RECT 57.385 2.23 58.545 2.37 ;
      RECT 57.385 1.58 57.525 2.37 ;
      RECT 55.185 1.58 57.525 1.72 ;
      RECT 58.155 2.955 58.435 3.325 ;
      RECT 58.165 2.7 58.425 3.325 ;
      RECT 55.215 3.72 57.39 3.885 ;
      RECT 57.245 2.6 57.39 3.885 ;
      RECT 54.135 3.515 54.415 3.885 ;
      RECT 54.135 3.63 55.355 3.77 ;
      RECT 56.965 2.6 57.39 2.74 ;
      RECT 56.965 2.42 57.225 2.74 ;
      RECT 50.305 4 53.965 4.14 ;
      RECT 53.825 3.185 53.965 4.14 ;
      RECT 50.305 3.07 50.445 4.14 ;
      RECT 56.845 3.26 57.105 3.58 ;
      RECT 53.825 3.185 56.355 3.325 ;
      RECT 56.075 2.955 56.355 3.325 ;
      RECT 50.305 3.07 50.755 3.325 ;
      RECT 50.475 2.955 50.755 3.325 ;
      RECT 56.845 3.07 57.045 3.58 ;
      RECT 56.075 3.07 57.045 3.21 ;
      RECT 56.645 1.86 56.785 3.21 ;
      RECT 56.585 1.86 56.845 2.18 ;
      RECT 47.905 6.655 48.255 7.005 ;
      RECT 56.455 6.61 56.805 6.96 ;
      RECT 47.905 6.685 56.805 6.885 ;
      RECT 50.485 2.42 50.745 2.74 ;
      RECT 50.485 2.51 51.525 2.65 ;
      RECT 51.385 1.72 51.525 2.65 ;
      RECT 54.145 1.86 54.405 2.18 ;
      RECT 51.385 1.72 54.345 1.86 ;
      RECT 53.525 2.7 53.785 3.02 ;
      RECT 53.525 2.7 53.845 2.93 ;
      RECT 53.635 2.395 53.915 2.765 ;
      RECT 53.225 3.26 53.545 3.58 ;
      RECT 53.225 2.14 53.365 3.58 ;
      RECT 53.165 2.14 53.425 2.46 ;
      RECT 50.725 3.54 50.985 3.86 ;
      RECT 50.725 3.63 52.405 3.77 ;
      RECT 52.265 3.35 52.405 3.77 ;
      RECT 52.265 3.35 52.705 3.58 ;
      RECT 52.445 3.26 52.705 3.58 ;
      RECT 51.765 2.42 52.165 2.93 ;
      RECT 51.955 2.395 52.235 2.765 ;
      RECT 51.705 2.42 52.235 2.74 ;
      RECT 44.77 6.22 45.09 6.545 ;
      RECT 44.8 5.695 44.97 6.545 ;
      RECT 44.8 5.695 44.975 6.045 ;
      RECT 44.8 5.695 45.775 5.87 ;
      RECT 45.6 1.965 45.775 5.87 ;
      RECT 45.545 1.965 45.895 2.315 ;
      RECT 45.57 6.655 45.895 6.98 ;
      RECT 44.455 6.745 45.895 6.915 ;
      RECT 44.455 2.395 44.615 6.915 ;
      RECT 44.77 2.365 45.09 2.685 ;
      RECT 44.455 2.395 45.09 2.565 ;
      RECT 43.72 5.84 44.06 6.19 ;
      RECT 43.805 2.705 43.975 6.19 ;
      RECT 43.73 2.705 44.07 3.055 ;
      RECT 33.19 2.955 33.47 3.325 ;
      RECT 33.245 1.29 33.415 3.325 ;
      RECT 43.24 1.29 43.41 1.815 ;
      RECT 43.15 1.46 43.49 1.81 ;
      RECT 33.245 1.29 43.41 1.46 ;
      RECT 39.87 2.395 40.15 2.765 ;
      RECT 38.8 2.42 39.06 2.74 ;
      RECT 41.35 2.23 41.63 2.6 ;
      RECT 41.96 2.14 42.22 2.46 ;
      RECT 38.86 1.58 39 2.74 ;
      RECT 39.94 1.58 40.08 2.765 ;
      RECT 41.06 2.23 42.22 2.37 ;
      RECT 41.06 1.58 41.2 2.37 ;
      RECT 38.86 1.58 41.2 1.72 ;
      RECT 41.83 2.955 42.11 3.325 ;
      RECT 41.84 2.7 42.1 3.325 ;
      RECT 38.89 3.72 41.065 3.885 ;
      RECT 40.92 2.6 41.065 3.885 ;
      RECT 37.81 3.515 38.09 3.885 ;
      RECT 37.81 3.63 39.03 3.77 ;
      RECT 40.64 2.6 41.065 2.74 ;
      RECT 40.64 2.42 40.9 2.74 ;
      RECT 33.98 4 37.64 4.14 ;
      RECT 37.5 3.185 37.64 4.14 ;
      RECT 33.98 3.07 34.12 4.14 ;
      RECT 40.52 3.26 40.78 3.58 ;
      RECT 37.5 3.185 40.03 3.325 ;
      RECT 39.75 2.955 40.03 3.325 ;
      RECT 33.98 3.07 34.43 3.325 ;
      RECT 34.15 2.955 34.43 3.325 ;
      RECT 40.52 3.07 40.72 3.58 ;
      RECT 39.75 3.07 40.72 3.21 ;
      RECT 40.32 1.86 40.46 3.21 ;
      RECT 40.26 1.86 40.52 2.18 ;
      RECT 31.625 6.66 31.975 7.01 ;
      RECT 40.13 6.615 40.48 6.965 ;
      RECT 31.625 6.69 40.48 6.89 ;
      RECT 34.16 2.42 34.42 2.74 ;
      RECT 34.16 2.51 35.2 2.65 ;
      RECT 35.06 1.72 35.2 2.65 ;
      RECT 37.82 1.86 38.08 2.18 ;
      RECT 35.06 1.72 38.02 1.86 ;
      RECT 37.2 2.7 37.46 3.02 ;
      RECT 37.2 2.7 37.52 2.93 ;
      RECT 37.31 2.395 37.59 2.765 ;
      RECT 36.9 3.26 37.22 3.58 ;
      RECT 36.9 2.14 37.04 3.58 ;
      RECT 36.84 2.14 37.1 2.46 ;
      RECT 34.4 3.54 34.66 3.86 ;
      RECT 34.4 3.63 36.08 3.77 ;
      RECT 35.94 3.35 36.08 3.77 ;
      RECT 35.94 3.35 36.38 3.58 ;
      RECT 36.12 3.26 36.38 3.58 ;
      RECT 35.44 2.42 35.84 2.93 ;
      RECT 35.63 2.395 35.91 2.765 ;
      RECT 35.38 2.42 35.91 2.74 ;
      RECT 28.445 6.22 28.765 6.545 ;
      RECT 28.475 5.695 28.645 6.545 ;
      RECT 28.475 5.695 28.65 6.045 ;
      RECT 28.475 5.695 29.45 5.87 ;
      RECT 29.275 1.965 29.45 5.87 ;
      RECT 29.22 1.965 29.57 2.315 ;
      RECT 29.245 6.655 29.57 6.98 ;
      RECT 28.13 6.745 29.57 6.915 ;
      RECT 28.13 2.395 28.29 6.915 ;
      RECT 28.445 2.365 28.765 2.685 ;
      RECT 28.13 2.395 28.765 2.565 ;
      RECT 27.395 5.84 27.735 6.19 ;
      RECT 27.48 2.705 27.65 6.19 ;
      RECT 27.405 2.705 27.745 3.055 ;
      RECT 16.865 2.955 17.145 3.325 ;
      RECT 16.92 1.29 17.09 3.325 ;
      RECT 26.915 1.29 27.085 1.815 ;
      RECT 26.825 1.46 27.165 1.81 ;
      RECT 16.92 1.29 27.085 1.46 ;
      RECT 23.545 2.395 23.825 2.765 ;
      RECT 22.475 2.42 22.735 2.74 ;
      RECT 25.025 2.23 25.305 2.6 ;
      RECT 25.635 2.14 25.895 2.46 ;
      RECT 22.535 1.58 22.675 2.74 ;
      RECT 23.615 1.58 23.755 2.765 ;
      RECT 24.735 2.23 25.895 2.37 ;
      RECT 24.735 1.58 24.875 2.37 ;
      RECT 22.535 1.58 24.875 1.72 ;
      RECT 25.505 2.955 25.785 3.325 ;
      RECT 25.515 2.7 25.775 3.325 ;
      RECT 22.565 3.72 24.74 3.885 ;
      RECT 24.595 2.6 24.74 3.885 ;
      RECT 21.485 3.515 21.765 3.885 ;
      RECT 21.485 3.63 22.705 3.77 ;
      RECT 24.315 2.6 24.74 2.74 ;
      RECT 24.315 2.42 24.575 2.74 ;
      RECT 17.655 4 21.315 4.14 ;
      RECT 21.175 3.185 21.315 4.14 ;
      RECT 17.655 3.07 17.795 4.14 ;
      RECT 24.195 3.26 24.455 3.58 ;
      RECT 21.175 3.185 23.705 3.325 ;
      RECT 23.425 2.955 23.705 3.325 ;
      RECT 17.655 3.07 18.105 3.325 ;
      RECT 17.825 2.955 18.105 3.325 ;
      RECT 24.195 3.07 24.395 3.58 ;
      RECT 23.425 3.07 24.395 3.21 ;
      RECT 23.995 1.86 24.135 3.21 ;
      RECT 23.935 1.86 24.195 2.18 ;
      RECT 15.3 6.655 15.65 7.005 ;
      RECT 23.805 6.61 24.155 6.96 ;
      RECT 15.3 6.685 24.155 6.885 ;
      RECT 17.835 2.42 18.095 2.74 ;
      RECT 17.835 2.51 18.875 2.65 ;
      RECT 18.735 1.72 18.875 2.65 ;
      RECT 21.495 1.86 21.755 2.18 ;
      RECT 18.735 1.72 21.695 1.86 ;
      RECT 20.875 2.7 21.135 3.02 ;
      RECT 20.875 2.7 21.195 2.93 ;
      RECT 20.985 2.395 21.265 2.765 ;
      RECT 20.575 3.26 20.895 3.58 ;
      RECT 20.575 2.14 20.715 3.58 ;
      RECT 20.515 2.14 20.775 2.46 ;
      RECT 18.075 3.54 18.335 3.86 ;
      RECT 18.075 3.63 19.755 3.77 ;
      RECT 19.615 3.35 19.755 3.77 ;
      RECT 19.615 3.35 20.055 3.58 ;
      RECT 19.795 3.26 20.055 3.58 ;
      RECT 19.115 2.42 19.515 2.93 ;
      RECT 19.305 2.395 19.585 2.765 ;
      RECT 19.055 2.42 19.585 2.74 ;
      RECT 12.12 6.22 12.44 6.545 ;
      RECT 12.15 5.695 12.32 6.545 ;
      RECT 12.15 5.695 12.325 6.045 ;
      RECT 12.15 5.695 13.125 5.87 ;
      RECT 12.95 1.965 13.125 5.87 ;
      RECT 12.895 1.965 13.245 2.315 ;
      RECT 12.92 6.655 13.245 6.98 ;
      RECT 11.805 6.745 13.245 6.915 ;
      RECT 11.805 2.395 11.965 6.915 ;
      RECT 12.12 2.365 12.44 2.685 ;
      RECT 11.805 2.395 12.44 2.565 ;
      RECT 11.07 5.84 11.41 6.19 ;
      RECT 11.155 2.705 11.325 6.19 ;
      RECT 11.08 2.705 11.42 3.055 ;
      RECT 0.54 2.955 0.82 3.325 ;
      RECT 0.595 1.29 0.765 3.325 ;
      RECT 10.59 1.29 10.76 1.815 ;
      RECT 10.5 1.46 10.84 1.81 ;
      RECT 0.595 1.29 10.76 1.46 ;
      RECT 7.22 2.395 7.5 2.765 ;
      RECT 6.15 2.42 6.41 2.74 ;
      RECT 8.7 2.23 8.98 2.6 ;
      RECT 9.31 2.14 9.57 2.46 ;
      RECT 6.21 1.58 6.35 2.74 ;
      RECT 7.29 1.58 7.43 2.765 ;
      RECT 8.41 2.23 9.57 2.37 ;
      RECT 8.41 1.58 8.55 2.37 ;
      RECT 6.21 1.58 8.55 1.72 ;
      RECT 9.18 2.955 9.46 3.325 ;
      RECT 9.19 2.7 9.45 3.325 ;
      RECT -1.73 6.995 -1.44 7.345 ;
      RECT -1.73 7.05 -0.39 7.22 ;
      RECT -0.56 6.685 -0.39 7.22 ;
      RECT 8.315 6.605 8.665 6.955 ;
      RECT -0.56 6.685 8.665 6.855 ;
      RECT 6.24 3.72 8.415 3.885 ;
      RECT 8.27 2.6 8.415 3.885 ;
      RECT 5.16 3.515 5.44 3.885 ;
      RECT 5.16 3.63 6.38 3.77 ;
      RECT 7.99 2.6 8.415 2.74 ;
      RECT 7.99 2.42 8.25 2.74 ;
      RECT 1.33 4 4.99 4.14 ;
      RECT 4.85 3.185 4.99 4.14 ;
      RECT 1.33 3.07 1.47 4.14 ;
      RECT 7.87 3.26 8.13 3.58 ;
      RECT 4.85 3.185 7.38 3.325 ;
      RECT 7.1 2.955 7.38 3.325 ;
      RECT 1.33 3.07 1.78 3.325 ;
      RECT 1.5 2.955 1.78 3.325 ;
      RECT 7.87 3.07 8.07 3.58 ;
      RECT 7.1 3.07 8.07 3.21 ;
      RECT 7.67 1.86 7.81 3.21 ;
      RECT 7.61 1.86 7.87 2.18 ;
      RECT 1.51 2.42 1.77 2.74 ;
      RECT 1.51 2.51 2.55 2.65 ;
      RECT 2.41 1.72 2.55 2.65 ;
      RECT 5.17 1.86 5.43 2.18 ;
      RECT 2.41 1.72 5.37 1.86 ;
      RECT 4.55 2.7 4.81 3.02 ;
      RECT 4.55 2.7 4.87 2.93 ;
      RECT 4.66 2.395 4.94 2.765 ;
      RECT 4.25 3.26 4.57 3.58 ;
      RECT 4.25 2.14 4.39 3.58 ;
      RECT 4.19 2.14 4.45 2.46 ;
      RECT 1.75 3.54 2.01 3.86 ;
      RECT 1.75 3.63 3.43 3.77 ;
      RECT 3.29 3.35 3.43 3.77 ;
      RECT 3.29 3.35 3.73 3.58 ;
      RECT 3.47 3.26 3.73 3.58 ;
      RECT 2.79 2.42 3.19 2.93 ;
      RECT 2.98 2.395 3.26 2.765 ;
      RECT 2.73 2.42 3.26 2.74 ;
      RECT 72.13 7.055 72.5 7.425 ;
      RECT 70.84 2.395 71.12 2.765 ;
      RECT 69 2.395 69.28 2.765 ;
      RECT 67.28 1.835 67.56 2.205 ;
      RECT 55.805 7.055 56.175 7.425 ;
      RECT 54.515 2.395 54.795 2.765 ;
      RECT 52.675 2.395 52.955 2.765 ;
      RECT 50.955 1.835 51.235 2.205 ;
      RECT 39.48 7.055 39.85 7.425 ;
      RECT 38.19 2.395 38.47 2.765 ;
      RECT 36.35 2.395 36.63 2.765 ;
      RECT 34.63 1.835 34.91 2.205 ;
      RECT 23.155 7.055 23.525 7.425 ;
      RECT 21.865 2.395 22.145 2.765 ;
      RECT 20.025 2.395 20.305 2.765 ;
      RECT 18.305 1.835 18.585 2.205 ;
      RECT 6.83 7.055 7.2 7.425 ;
      RECT 5.54 2.395 5.82 2.765 ;
      RECT 3.7 2.395 3.98 2.765 ;
      RECT 1.98 1.835 2.26 2.205 ;
    LAYER via1 ;
      RECT 80.68 7.375 80.83 7.525 ;
      RECT 78.31 6.74 78.46 6.89 ;
      RECT 78.295 2.065 78.445 2.215 ;
      RECT 77.505 2.45 77.655 2.6 ;
      RECT 77.505 6.325 77.655 6.475 ;
      RECT 76.48 2.805 76.63 2.955 ;
      RECT 76.47 5.94 76.62 6.09 ;
      RECT 75.9 1.56 76.05 1.71 ;
      RECT 74.665 2.225 74.815 2.375 ;
      RECT 74.545 2.785 74.695 2.935 ;
      RECT 73.345 2.505 73.495 2.655 ;
      RECT 73.225 3.345 73.375 3.495 ;
      RECT 72.965 1.945 73.115 2.095 ;
      RECT 72.885 6.71 73.035 6.86 ;
      RECT 72.24 7.165 72.39 7.315 ;
      RECT 71.505 2.505 71.655 2.655 ;
      RECT 70.905 2.505 71.055 2.655 ;
      RECT 70.525 1.945 70.675 2.095 ;
      RECT 69.905 2.785 70.055 2.935 ;
      RECT 69.665 3.345 69.815 3.495 ;
      RECT 69.545 2.225 69.695 2.375 ;
      RECT 69.065 2.505 69.215 2.655 ;
      RECT 68.825 3.345 68.975 3.495 ;
      RECT 68.085 2.505 68.235 2.655 ;
      RECT 67.345 1.945 67.495 2.095 ;
      RECT 67.105 3.625 67.255 3.775 ;
      RECT 66.865 2.505 67.015 2.655 ;
      RECT 66.865 3.065 67.015 3.215 ;
      RECT 65.905 3.065 66.055 3.215 ;
      RECT 64.33 6.755 64.48 6.905 ;
      RECT 61.985 6.74 62.135 6.89 ;
      RECT 61.97 2.065 62.12 2.215 ;
      RECT 61.18 2.45 61.33 2.6 ;
      RECT 61.18 6.325 61.33 6.475 ;
      RECT 60.155 2.805 60.305 2.955 ;
      RECT 60.145 5.94 60.295 6.09 ;
      RECT 59.575 1.56 59.725 1.71 ;
      RECT 58.34 2.225 58.49 2.375 ;
      RECT 58.22 2.785 58.37 2.935 ;
      RECT 57.02 2.505 57.17 2.655 ;
      RECT 56.9 3.345 57.05 3.495 ;
      RECT 56.64 1.945 56.79 2.095 ;
      RECT 56.555 6.71 56.705 6.86 ;
      RECT 55.915 7.165 56.065 7.315 ;
      RECT 55.18 2.505 55.33 2.655 ;
      RECT 54.58 2.505 54.73 2.655 ;
      RECT 54.2 1.945 54.35 2.095 ;
      RECT 53.58 2.785 53.73 2.935 ;
      RECT 53.34 3.345 53.49 3.495 ;
      RECT 53.22 2.225 53.37 2.375 ;
      RECT 52.74 2.505 52.89 2.655 ;
      RECT 52.5 3.345 52.65 3.495 ;
      RECT 51.76 2.505 51.91 2.655 ;
      RECT 51.02 1.945 51.17 2.095 ;
      RECT 50.78 3.625 50.93 3.775 ;
      RECT 50.54 2.505 50.69 2.655 ;
      RECT 50.54 3.065 50.69 3.215 ;
      RECT 49.58 3.065 49.73 3.215 ;
      RECT 48.005 6.755 48.155 6.905 ;
      RECT 45.66 6.74 45.81 6.89 ;
      RECT 45.645 2.065 45.795 2.215 ;
      RECT 44.855 2.45 45.005 2.6 ;
      RECT 44.855 6.325 45.005 6.475 ;
      RECT 43.83 2.805 43.98 2.955 ;
      RECT 43.82 5.94 43.97 6.09 ;
      RECT 43.25 1.56 43.4 1.71 ;
      RECT 42.015 2.225 42.165 2.375 ;
      RECT 41.895 2.785 42.045 2.935 ;
      RECT 40.695 2.505 40.845 2.655 ;
      RECT 40.575 3.345 40.725 3.495 ;
      RECT 40.315 1.945 40.465 2.095 ;
      RECT 40.23 6.715 40.38 6.865 ;
      RECT 39.59 7.165 39.74 7.315 ;
      RECT 38.855 2.505 39.005 2.655 ;
      RECT 38.255 2.505 38.405 2.655 ;
      RECT 37.875 1.945 38.025 2.095 ;
      RECT 37.255 2.785 37.405 2.935 ;
      RECT 37.015 3.345 37.165 3.495 ;
      RECT 36.895 2.225 37.045 2.375 ;
      RECT 36.415 2.505 36.565 2.655 ;
      RECT 36.175 3.345 36.325 3.495 ;
      RECT 35.435 2.505 35.585 2.655 ;
      RECT 34.695 1.945 34.845 2.095 ;
      RECT 34.455 3.625 34.605 3.775 ;
      RECT 34.215 2.505 34.365 2.655 ;
      RECT 34.215 3.065 34.365 3.215 ;
      RECT 33.255 3.065 33.405 3.215 ;
      RECT 31.725 6.76 31.875 6.91 ;
      RECT 29.335 6.74 29.485 6.89 ;
      RECT 29.32 2.065 29.47 2.215 ;
      RECT 28.53 2.45 28.68 2.6 ;
      RECT 28.53 6.325 28.68 6.475 ;
      RECT 27.505 2.805 27.655 2.955 ;
      RECT 27.495 5.94 27.645 6.09 ;
      RECT 26.925 1.56 27.075 1.71 ;
      RECT 25.69 2.225 25.84 2.375 ;
      RECT 25.57 2.785 25.72 2.935 ;
      RECT 24.37 2.505 24.52 2.655 ;
      RECT 24.25 3.345 24.4 3.495 ;
      RECT 23.99 1.945 24.14 2.095 ;
      RECT 23.905 6.71 24.055 6.86 ;
      RECT 23.265 7.165 23.415 7.315 ;
      RECT 22.53 2.505 22.68 2.655 ;
      RECT 21.93 2.505 22.08 2.655 ;
      RECT 21.55 1.945 21.7 2.095 ;
      RECT 20.93 2.785 21.08 2.935 ;
      RECT 20.69 3.345 20.84 3.495 ;
      RECT 20.57 2.225 20.72 2.375 ;
      RECT 20.09 2.505 20.24 2.655 ;
      RECT 19.85 3.345 20 3.495 ;
      RECT 19.11 2.505 19.26 2.655 ;
      RECT 18.37 1.945 18.52 2.095 ;
      RECT 18.13 3.625 18.28 3.775 ;
      RECT 17.89 2.505 18.04 2.655 ;
      RECT 17.89 3.065 18.04 3.215 ;
      RECT 16.93 3.065 17.08 3.215 ;
      RECT 15.4 6.755 15.55 6.905 ;
      RECT 13.01 6.74 13.16 6.89 ;
      RECT 12.995 2.065 13.145 2.215 ;
      RECT 12.205 2.45 12.355 2.6 ;
      RECT 12.205 6.325 12.355 6.475 ;
      RECT 11.18 2.805 11.33 2.955 ;
      RECT 11.17 5.94 11.32 6.09 ;
      RECT 10.6 1.56 10.75 1.71 ;
      RECT 9.365 2.225 9.515 2.375 ;
      RECT 9.245 2.785 9.395 2.935 ;
      RECT 8.415 6.705 8.565 6.855 ;
      RECT 8.045 2.505 8.195 2.655 ;
      RECT 7.925 3.345 8.075 3.495 ;
      RECT 7.665 1.945 7.815 2.095 ;
      RECT 6.94 7.165 7.09 7.315 ;
      RECT 6.205 2.505 6.355 2.655 ;
      RECT 5.605 2.505 5.755 2.655 ;
      RECT 5.225 1.945 5.375 2.095 ;
      RECT 4.605 2.785 4.755 2.935 ;
      RECT 4.365 3.345 4.515 3.495 ;
      RECT 4.245 2.225 4.395 2.375 ;
      RECT 3.765 2.505 3.915 2.655 ;
      RECT 3.525 3.345 3.675 3.495 ;
      RECT 2.785 2.505 2.935 2.655 ;
      RECT 2.045 1.945 2.195 2.095 ;
      RECT 1.805 3.625 1.955 3.775 ;
      RECT 1.565 2.505 1.715 2.655 ;
      RECT 1.565 3.065 1.715 3.215 ;
      RECT 0.605 3.065 0.755 3.215 ;
      RECT -1.66 7.095 -1.51 7.245 ;
      RECT -2.035 6.355 -1.885 6.505 ;
    LAYER met1 ;
      RECT 72.97 2.93 74.57 3.07 ;
      RECT 56.645 2.93 58.245 3.07 ;
      RECT 40.32 2.93 41.92 3.07 ;
      RECT 23.995 2.93 25.595 3.07 ;
      RECT 7.67 2.93 9.27 3.07 ;
      RECT 72.97 2.93 74.735 3.055 ;
      RECT 56.645 2.93 58.41 3.055 ;
      RECT 40.32 2.93 42.085 3.055 ;
      RECT 23.995 2.93 25.76 3.055 ;
      RECT 7.67 2.93 9.435 3.055 ;
      RECT 74.46 2.73 74.78 2.99 ;
      RECT 58.135 2.73 58.455 2.99 ;
      RECT 41.81 2.73 42.13 2.99 ;
      RECT 25.485 2.73 25.805 2.99 ;
      RECT 9.16 2.73 9.48 2.99 ;
      RECT 74.46 2.745 74.885 2.975 ;
      RECT 58.135 2.745 58.56 2.975 ;
      RECT 41.81 2.745 42.235 2.975 ;
      RECT 25.485 2.745 25.91 2.975 ;
      RECT 9.16 2.745 9.585 2.975 ;
      RECT 75.195 0 75.38 2.945 ;
      RECT 58.87 0 59.055 2.945 ;
      RECT 42.545 0 42.73 2.945 ;
      RECT 26.22 0 26.405 2.945 ;
      RECT 9.895 0 10.08 2.945 ;
      RECT 74.43 2.79 75.38 2.945 ;
      RECT 74.46 2.76 75.38 2.945 ;
      RECT 72.635 2.79 73.11 2.975 ;
      RECT 58.105 2.79 59.055 2.945 ;
      RECT 58.135 2.76 59.055 2.945 ;
      RECT 56.31 2.79 56.785 2.975 ;
      RECT 41.78 2.79 42.73 2.945 ;
      RECT 41.81 2.76 42.73 2.945 ;
      RECT 39.985 2.79 40.46 2.975 ;
      RECT 25.455 2.79 26.405 2.945 ;
      RECT 25.485 2.76 26.405 2.945 ;
      RECT 23.66 2.79 24.135 2.975 ;
      RECT 9.13 2.79 10.08 2.945 ;
      RECT 9.16 2.76 10.08 2.945 ;
      RECT 7.335 2.79 7.81 2.975 ;
      RECT 72.635 2.745 72.925 2.975 ;
      RECT 56.31 2.745 56.6 2.975 ;
      RECT 39.985 2.745 40.275 2.975 ;
      RECT 23.66 2.745 23.95 2.975 ;
      RECT 7.335 2.745 7.625 2.975 ;
      RECT 65.565 0 75.38 1.74 ;
      RECT 49.24 0 59.055 1.74 ;
      RECT 32.915 0 42.73 1.74 ;
      RECT 16.59 0 26.405 1.74 ;
      RECT 0.265 0 10.08 1.74 ;
      RECT -3.225 0 81.15 0.305 ;
      RECT -3.225 4.135 81.15 4.745 ;
      RECT 65.565 3.98 75.225 4.745 ;
      RECT 49.24 3.98 58.9 4.745 ;
      RECT 32.915 3.98 42.575 4.745 ;
      RECT 16.59 3.98 26.25 4.745 ;
      RECT 0.265 3.98 9.925 4.745 ;
      RECT -3.23 8.575 81.15 8.88 ;
      RECT 71.4 6.315 71.575 8.88 ;
      RECT 55.075 6.315 55.25 8.88 ;
      RECT 38.75 6.315 38.925 8.88 ;
      RECT 22.425 6.315 22.6 8.88 ;
      RECT 6.1 6.315 6.275 8.88 ;
      RECT 71.775 6.285 72.065 6.515 ;
      RECT 55.45 6.285 55.74 6.515 ;
      RECT 39.125 6.285 39.415 6.515 ;
      RECT 22.8 6.285 23.09 6.515 ;
      RECT 6.475 6.285 6.765 6.515 ;
      RECT 71.4 6.315 72.065 6.485 ;
      RECT 55.075 6.315 55.74 6.485 ;
      RECT 38.75 6.315 39.415 6.485 ;
      RECT 22.425 6.315 23.09 6.485 ;
      RECT 6.1 6.315 6.765 6.485 ;
      RECT 80.55 7.765 80.84 7.995 ;
      RECT 80.61 6.285 80.78 7.995 ;
      RECT 80.58 7.275 80.93 7.625 ;
      RECT 80.55 6.285 80.84 6.515 ;
      RECT 80.55 2.365 80.84 2.595 ;
      RECT 80.61 0.885 80.78 2.595 ;
      RECT 80.55 0.885 80.84 1.115 ;
      RECT 80.14 2.735 80.47 2.965 ;
      RECT 80.14 2.765 80.64 2.935 ;
      RECT 80.14 2.395 80.33 2.965 ;
      RECT 79.56 2.365 79.85 2.595 ;
      RECT 79.56 2.395 80.33 2.565 ;
      RECT 79.62 0.885 79.79 2.595 ;
      RECT 79.56 0.885 79.85 1.115 ;
      RECT 79.56 7.765 79.85 7.995 ;
      RECT 79.62 6.285 79.79 7.995 ;
      RECT 79.56 6.285 79.85 6.515 ;
      RECT 79.56 6.325 80.41 6.485 ;
      RECT 80.24 5.915 80.41 6.485 ;
      RECT 79.56 6.32 79.95 6.485 ;
      RECT 80.18 5.915 80.47 6.145 ;
      RECT 80.18 5.945 80.64 6.115 ;
      RECT 79.19 2.735 79.48 2.965 ;
      RECT 79.19 2.765 79.65 2.935 ;
      RECT 79.25 1.655 79.415 2.965 ;
      RECT 77.765 1.625 78.055 1.855 ;
      RECT 77.765 1.655 79.415 1.825 ;
      RECT 77.825 0.885 77.995 1.855 ;
      RECT 77.765 0.885 78.055 1.115 ;
      RECT 77.765 7.765 78.055 7.995 ;
      RECT 77.825 7.025 77.995 7.995 ;
      RECT 77.825 7.12 79.415 7.29 ;
      RECT 79.245 5.915 79.415 7.29 ;
      RECT 77.765 7.025 78.055 7.255 ;
      RECT 79.19 5.915 79.48 6.145 ;
      RECT 79.19 5.945 79.65 6.115 ;
      RECT 78.195 1.965 78.545 2.315 ;
      RECT 75.89 2.025 78.545 2.195 ;
      RECT 75.89 1.46 76.06 2.195 ;
      RECT 75.8 1.46 76.14 1.81 ;
      RECT 78.22 6.655 78.545 6.98 ;
      RECT 72.785 6.61 73.135 6.96 ;
      RECT 78.195 6.655 78.545 6.885 ;
      RECT 72.58 6.655 73.135 6.885 ;
      RECT 72.41 6.685 78.545 6.855 ;
      RECT 77.42 2.365 77.74 2.685 ;
      RECT 77.39 2.365 77.74 2.595 ;
      RECT 77.22 2.395 77.74 2.565 ;
      RECT 77.42 6.255 77.74 6.545 ;
      RECT 77.39 6.285 77.74 6.515 ;
      RECT 77.22 6.315 77.74 6.485 ;
      RECT 76.38 2.705 76.72 3.055 ;
      RECT 76.38 2.765 76.855 2.935 ;
      RECT 76.37 5.84 76.71 6.19 ;
      RECT 70.78 5.915 71.07 6.145 ;
      RECT 70.78 5.945 76.855 6.115 ;
      RECT 73.875 2.465 74.165 2.695 ;
      RECT 73.875 2.465 74.33 2.65 ;
      RECT 74.19 2.37 74.81 2.51 ;
      RECT 74.58 2.17 74.9 2.43 ;
      RECT 73.26 2.45 73.58 2.71 ;
      RECT 73.26 2.45 73.725 2.695 ;
      RECT 73.585 2.07 73.725 2.695 ;
      RECT 73.585 2.07 73.85 2.21 ;
      RECT 74.115 1.905 74.405 2.135 ;
      RECT 73.71 1.95 74.405 2.09 ;
      RECT 73.155 3.29 73.445 3.815 ;
      RECT 73.14 3.29 73.46 3.55 ;
      RECT 72.88 1.89 73.2 2.15 ;
      RECT 72.88 1.905 73.445 2.135 ;
      RECT 72.155 3.585 72.445 3.815 ;
      RECT 72.35 2.23 72.49 3.77 ;
      RECT 72.395 2.185 72.685 2.415 ;
      RECT 71.99 2.23 72.685 2.37 ;
      RECT 71.99 2.07 72.13 2.37 ;
      RECT 70.53 2.07 72.13 2.21 ;
      RECT 70.44 1.89 70.76 2.15 ;
      RECT 70.44 1.905 71.005 2.15 ;
      RECT 72.15 7.765 72.44 7.995 ;
      RECT 72.21 7.025 72.38 7.995 ;
      RECT 72.13 7.075 72.5 7.425 ;
      RECT 72.13 7.055 72.44 7.425 ;
      RECT 72.15 7.025 72.44 7.425 ;
      RECT 69.55 2.93 72.13 3.07 ;
      RECT 71.915 2.745 72.205 2.975 ;
      RECT 69.475 2.745 70.14 2.975 ;
      RECT 69.82 2.73 70.14 3.07 ;
      RECT 70.82 2.45 71.14 2.71 ;
      RECT 70.82 2.465 71.245 2.695 ;
      RECT 69.46 2.17 69.78 2.43 ;
      RECT 69.955 2.185 70.245 2.415 ;
      RECT 69.46 2.23 70.245 2.37 ;
      RECT 69.58 3.29 69.9 3.55 ;
      RECT 68.74 3.29 69.06 3.55 ;
      RECT 69.58 3.305 70.005 3.535 ;
      RECT 68.74 3.35 70.005 3.49 ;
      RECT 68.275 3.025 68.565 3.255 ;
      RECT 68.35 1.95 68.49 3.255 ;
      RECT 68 2.45 68.49 2.71 ;
      RECT 67.755 2.465 68.49 2.695 ;
      RECT 68.755 1.905 69.045 2.135 ;
      RECT 68.35 1.95 69.045 2.09 ;
      RECT 67.515 3.305 67.805 3.535 ;
      RECT 67.515 3.305 67.97 3.49 ;
      RECT 67.83 2.93 67.97 3.49 ;
      RECT 67.47 2.93 67.97 3.07 ;
      RECT 67.47 1.95 67.61 3.07 ;
      RECT 67.26 1.89 67.58 2.15 ;
      RECT 67.02 3.57 67.34 3.83 ;
      RECT 66.315 3.585 66.605 3.815 ;
      RECT 66.315 3.63 67.34 3.77 ;
      RECT 66.39 3.58 66.65 3.77 ;
      RECT 66.78 2.45 67.1 2.71 ;
      RECT 66.78 2.465 67.325 2.695 ;
      RECT 66.78 3.01 67.1 3.27 ;
      RECT 66.78 3.025 67.325 3.255 ;
      RECT 65.82 3.01 66.14 3.27 ;
      RECT 65.91 1.95 66.05 3.27 ;
      RECT 66.315 1.905 66.605 2.135 ;
      RECT 65.91 1.95 66.605 2.09 ;
      RECT 64.225 7.765 64.515 7.995 ;
      RECT 64.285 6.285 64.455 7.995 ;
      RECT 64.23 6.655 64.58 7.005 ;
      RECT 64.225 6.285 64.515 6.515 ;
      RECT 64.225 2.365 64.515 2.595 ;
      RECT 64.285 0.885 64.455 2.595 ;
      RECT 64.225 0.885 64.515 1.115 ;
      RECT 63.815 2.735 64.145 2.965 ;
      RECT 63.815 2.765 64.315 2.935 ;
      RECT 63.815 2.395 64.005 2.965 ;
      RECT 63.235 2.365 63.525 2.595 ;
      RECT 63.235 2.395 64.005 2.565 ;
      RECT 63.295 0.885 63.465 2.595 ;
      RECT 63.235 0.885 63.525 1.115 ;
      RECT 63.235 7.765 63.525 7.995 ;
      RECT 63.295 6.285 63.465 7.995 ;
      RECT 63.235 6.285 63.525 6.515 ;
      RECT 63.235 6.325 64.085 6.485 ;
      RECT 63.915 5.915 64.085 6.485 ;
      RECT 63.235 6.32 63.625 6.485 ;
      RECT 63.855 5.915 64.145 6.145 ;
      RECT 63.855 5.945 64.315 6.115 ;
      RECT 62.865 2.735 63.155 2.965 ;
      RECT 62.865 2.765 63.325 2.935 ;
      RECT 62.925 1.655 63.09 2.965 ;
      RECT 61.44 1.625 61.73 1.855 ;
      RECT 61.44 1.655 63.09 1.825 ;
      RECT 61.5 0.885 61.67 1.855 ;
      RECT 61.44 0.885 61.73 1.115 ;
      RECT 61.44 7.765 61.73 7.995 ;
      RECT 61.5 7.025 61.67 7.995 ;
      RECT 61.5 7.12 63.09 7.29 ;
      RECT 62.92 5.915 63.09 7.29 ;
      RECT 61.44 7.025 61.73 7.255 ;
      RECT 62.865 5.915 63.155 6.145 ;
      RECT 62.865 5.945 63.325 6.115 ;
      RECT 61.87 1.965 62.22 2.315 ;
      RECT 59.565 2.025 62.22 2.195 ;
      RECT 59.565 1.46 59.735 2.195 ;
      RECT 59.475 1.46 59.815 1.81 ;
      RECT 61.895 6.655 62.22 6.98 ;
      RECT 56.455 6.61 56.805 6.96 ;
      RECT 61.87 6.655 62.22 6.885 ;
      RECT 56.255 6.655 56.805 6.885 ;
      RECT 56.085 6.685 62.22 6.855 ;
      RECT 61.095 2.365 61.415 2.685 ;
      RECT 61.065 2.365 61.415 2.595 ;
      RECT 60.895 2.395 61.415 2.565 ;
      RECT 61.095 6.255 61.415 6.545 ;
      RECT 61.065 6.285 61.415 6.515 ;
      RECT 60.895 6.315 61.415 6.485 ;
      RECT 60.055 2.705 60.395 3.055 ;
      RECT 60.055 2.765 60.53 2.935 ;
      RECT 60.045 5.84 60.385 6.19 ;
      RECT 54.455 5.915 54.745 6.145 ;
      RECT 54.455 5.945 60.53 6.115 ;
      RECT 57.55 2.465 57.84 2.695 ;
      RECT 57.55 2.465 58.005 2.65 ;
      RECT 57.865 2.37 58.485 2.51 ;
      RECT 58.255 2.17 58.575 2.43 ;
      RECT 56.935 2.45 57.255 2.71 ;
      RECT 56.935 2.45 57.4 2.695 ;
      RECT 57.26 2.07 57.4 2.695 ;
      RECT 57.26 2.07 57.525 2.21 ;
      RECT 57.79 1.905 58.08 2.135 ;
      RECT 57.385 1.95 58.08 2.09 ;
      RECT 56.83 3.29 57.12 3.815 ;
      RECT 56.815 3.29 57.135 3.55 ;
      RECT 56.555 1.89 56.875 2.15 ;
      RECT 56.555 1.905 57.12 2.135 ;
      RECT 55.83 3.585 56.12 3.815 ;
      RECT 56.025 2.23 56.165 3.77 ;
      RECT 56.07 2.185 56.36 2.415 ;
      RECT 55.665 2.23 56.36 2.37 ;
      RECT 55.665 2.07 55.805 2.37 ;
      RECT 54.205 2.07 55.805 2.21 ;
      RECT 54.115 1.89 54.435 2.15 ;
      RECT 54.115 1.905 54.68 2.15 ;
      RECT 55.825 7.765 56.115 7.995 ;
      RECT 55.885 7.025 56.055 7.995 ;
      RECT 55.805 7.075 56.175 7.425 ;
      RECT 55.805 7.055 56.115 7.425 ;
      RECT 55.825 7.025 56.115 7.425 ;
      RECT 53.225 2.93 55.805 3.07 ;
      RECT 55.59 2.745 55.88 2.975 ;
      RECT 53.15 2.745 53.815 2.975 ;
      RECT 53.495 2.73 53.815 3.07 ;
      RECT 54.495 2.45 54.815 2.71 ;
      RECT 54.495 2.465 54.92 2.695 ;
      RECT 53.135 2.17 53.455 2.43 ;
      RECT 53.63 2.185 53.92 2.415 ;
      RECT 53.135 2.23 53.92 2.37 ;
      RECT 53.255 3.29 53.575 3.55 ;
      RECT 52.415 3.29 52.735 3.55 ;
      RECT 53.255 3.305 53.68 3.535 ;
      RECT 52.415 3.35 53.68 3.49 ;
      RECT 51.95 3.025 52.24 3.255 ;
      RECT 52.025 1.95 52.165 3.255 ;
      RECT 51.675 2.45 52.165 2.71 ;
      RECT 51.43 2.465 52.165 2.695 ;
      RECT 52.43 1.905 52.72 2.135 ;
      RECT 52.025 1.95 52.72 2.09 ;
      RECT 51.19 3.305 51.48 3.535 ;
      RECT 51.19 3.305 51.645 3.49 ;
      RECT 51.505 2.93 51.645 3.49 ;
      RECT 51.145 2.93 51.645 3.07 ;
      RECT 51.145 1.95 51.285 3.07 ;
      RECT 50.935 1.89 51.255 2.15 ;
      RECT 50.695 3.57 51.015 3.83 ;
      RECT 49.99 3.585 50.28 3.815 ;
      RECT 49.99 3.63 51.015 3.77 ;
      RECT 50.065 3.58 50.325 3.77 ;
      RECT 50.455 2.45 50.775 2.71 ;
      RECT 50.455 2.465 51 2.695 ;
      RECT 50.455 3.01 50.775 3.27 ;
      RECT 50.455 3.025 51 3.255 ;
      RECT 49.495 3.01 49.815 3.27 ;
      RECT 49.585 1.95 49.725 3.27 ;
      RECT 49.99 1.905 50.28 2.135 ;
      RECT 49.585 1.95 50.28 2.09 ;
      RECT 47.9 7.765 48.19 7.995 ;
      RECT 47.96 6.285 48.13 7.995 ;
      RECT 47.905 6.655 48.255 7.005 ;
      RECT 47.9 6.285 48.19 6.515 ;
      RECT 47.9 2.365 48.19 2.595 ;
      RECT 47.96 0.885 48.13 2.595 ;
      RECT 47.9 0.885 48.19 1.115 ;
      RECT 47.49 2.735 47.82 2.965 ;
      RECT 47.49 2.765 47.99 2.935 ;
      RECT 47.49 2.395 47.68 2.965 ;
      RECT 46.91 2.365 47.2 2.595 ;
      RECT 46.91 2.395 47.68 2.565 ;
      RECT 46.97 0.885 47.14 2.595 ;
      RECT 46.91 0.885 47.2 1.115 ;
      RECT 46.91 7.765 47.2 7.995 ;
      RECT 46.97 6.285 47.14 7.995 ;
      RECT 46.91 6.285 47.2 6.515 ;
      RECT 46.91 6.325 47.76 6.485 ;
      RECT 47.59 5.915 47.76 6.485 ;
      RECT 46.91 6.32 47.3 6.485 ;
      RECT 47.53 5.915 47.82 6.145 ;
      RECT 47.53 5.945 47.99 6.115 ;
      RECT 46.54 2.735 46.83 2.965 ;
      RECT 46.54 2.765 47 2.935 ;
      RECT 46.6 1.655 46.765 2.965 ;
      RECT 45.115 1.625 45.405 1.855 ;
      RECT 45.115 1.655 46.765 1.825 ;
      RECT 45.175 0.885 45.345 1.855 ;
      RECT 45.115 0.885 45.405 1.115 ;
      RECT 45.115 7.765 45.405 7.995 ;
      RECT 45.175 7.025 45.345 7.995 ;
      RECT 45.175 7.12 46.765 7.29 ;
      RECT 46.595 5.915 46.765 7.29 ;
      RECT 45.115 7.025 45.405 7.255 ;
      RECT 46.54 5.915 46.83 6.145 ;
      RECT 46.54 5.945 47 6.115 ;
      RECT 45.545 1.965 45.895 2.315 ;
      RECT 43.24 2.025 45.895 2.195 ;
      RECT 43.24 1.46 43.41 2.195 ;
      RECT 43.15 1.46 43.49 1.81 ;
      RECT 45.57 6.655 45.895 6.98 ;
      RECT 40.13 6.615 40.48 6.965 ;
      RECT 45.545 6.655 45.895 6.885 ;
      RECT 39.93 6.655 40.48 6.885 ;
      RECT 39.76 6.685 45.895 6.855 ;
      RECT 44.77 2.365 45.09 2.685 ;
      RECT 44.74 2.365 45.09 2.595 ;
      RECT 44.57 2.395 45.09 2.565 ;
      RECT 44.77 6.255 45.09 6.545 ;
      RECT 44.74 6.285 45.09 6.515 ;
      RECT 44.57 6.315 45.09 6.485 ;
      RECT 43.73 2.705 44.07 3.055 ;
      RECT 43.73 2.765 44.205 2.935 ;
      RECT 43.72 5.84 44.06 6.19 ;
      RECT 38.13 5.915 38.42 6.145 ;
      RECT 38.13 5.945 44.205 6.115 ;
      RECT 41.225 2.465 41.515 2.695 ;
      RECT 41.225 2.465 41.68 2.65 ;
      RECT 41.54 2.37 42.16 2.51 ;
      RECT 41.93 2.17 42.25 2.43 ;
      RECT 40.61 2.45 40.93 2.71 ;
      RECT 40.61 2.45 41.075 2.695 ;
      RECT 40.935 2.07 41.075 2.695 ;
      RECT 40.935 2.07 41.2 2.21 ;
      RECT 41.465 1.905 41.755 2.135 ;
      RECT 41.06 1.95 41.755 2.09 ;
      RECT 40.505 3.29 40.795 3.815 ;
      RECT 40.49 3.29 40.81 3.55 ;
      RECT 40.23 1.89 40.55 2.15 ;
      RECT 40.23 1.905 40.795 2.135 ;
      RECT 39.505 3.585 39.795 3.815 ;
      RECT 39.7 2.23 39.84 3.77 ;
      RECT 39.745 2.185 40.035 2.415 ;
      RECT 39.34 2.23 40.035 2.37 ;
      RECT 39.34 2.07 39.48 2.37 ;
      RECT 37.88 2.07 39.48 2.21 ;
      RECT 37.79 1.89 38.11 2.15 ;
      RECT 37.79 1.905 38.355 2.15 ;
      RECT 39.5 7.765 39.79 7.995 ;
      RECT 39.56 7.025 39.73 7.995 ;
      RECT 39.48 7.075 39.85 7.425 ;
      RECT 39.48 7.055 39.79 7.425 ;
      RECT 39.5 7.025 39.79 7.425 ;
      RECT 36.9 2.93 39.48 3.07 ;
      RECT 39.265 2.745 39.555 2.975 ;
      RECT 36.825 2.745 37.49 2.975 ;
      RECT 37.17 2.73 37.49 3.07 ;
      RECT 38.17 2.45 38.49 2.71 ;
      RECT 38.17 2.465 38.595 2.695 ;
      RECT 36.81 2.17 37.13 2.43 ;
      RECT 37.305 2.185 37.595 2.415 ;
      RECT 36.81 2.23 37.595 2.37 ;
      RECT 36.93 3.29 37.25 3.55 ;
      RECT 36.09 3.29 36.41 3.55 ;
      RECT 36.93 3.305 37.355 3.535 ;
      RECT 36.09 3.35 37.355 3.49 ;
      RECT 35.625 3.025 35.915 3.255 ;
      RECT 35.7 1.95 35.84 3.255 ;
      RECT 35.35 2.45 35.84 2.71 ;
      RECT 35.105 2.465 35.84 2.695 ;
      RECT 36.105 1.905 36.395 2.135 ;
      RECT 35.7 1.95 36.395 2.09 ;
      RECT 34.865 3.305 35.155 3.535 ;
      RECT 34.865 3.305 35.32 3.49 ;
      RECT 35.18 2.93 35.32 3.49 ;
      RECT 34.82 2.93 35.32 3.07 ;
      RECT 34.82 1.95 34.96 3.07 ;
      RECT 34.61 1.89 34.93 2.15 ;
      RECT 34.37 3.57 34.69 3.83 ;
      RECT 33.665 3.585 33.955 3.815 ;
      RECT 33.665 3.63 34.69 3.77 ;
      RECT 33.74 3.58 34 3.77 ;
      RECT 34.13 2.45 34.45 2.71 ;
      RECT 34.13 2.465 34.675 2.695 ;
      RECT 34.13 3.01 34.45 3.27 ;
      RECT 34.13 3.025 34.675 3.255 ;
      RECT 33.17 3.01 33.49 3.27 ;
      RECT 33.26 1.95 33.4 3.27 ;
      RECT 33.665 1.905 33.955 2.135 ;
      RECT 33.26 1.95 33.955 2.09 ;
      RECT 31.575 7.765 31.865 7.995 ;
      RECT 31.635 6.285 31.805 7.995 ;
      RECT 31.62 6.66 31.975 7.015 ;
      RECT 31.575 6.285 31.865 6.515 ;
      RECT 31.575 2.365 31.865 2.595 ;
      RECT 31.635 0.885 31.805 2.595 ;
      RECT 31.575 0.885 31.865 1.115 ;
      RECT 31.165 2.735 31.495 2.965 ;
      RECT 31.165 2.765 31.665 2.935 ;
      RECT 31.165 2.395 31.355 2.965 ;
      RECT 30.585 2.365 30.875 2.595 ;
      RECT 30.585 2.395 31.355 2.565 ;
      RECT 30.645 0.885 30.815 2.595 ;
      RECT 30.585 0.885 30.875 1.115 ;
      RECT 30.585 7.765 30.875 7.995 ;
      RECT 30.645 6.285 30.815 7.995 ;
      RECT 30.585 6.285 30.875 6.515 ;
      RECT 30.585 6.325 31.435 6.485 ;
      RECT 31.265 5.915 31.435 6.485 ;
      RECT 30.585 6.32 30.975 6.485 ;
      RECT 31.205 5.915 31.495 6.145 ;
      RECT 31.205 5.945 31.665 6.115 ;
      RECT 30.215 2.735 30.505 2.965 ;
      RECT 30.215 2.765 30.675 2.935 ;
      RECT 30.275 1.655 30.44 2.965 ;
      RECT 28.79 1.625 29.08 1.855 ;
      RECT 28.79 1.655 30.44 1.825 ;
      RECT 28.85 0.885 29.02 1.855 ;
      RECT 28.79 0.885 29.08 1.115 ;
      RECT 28.79 7.765 29.08 7.995 ;
      RECT 28.85 7.025 29.02 7.995 ;
      RECT 28.85 7.12 30.44 7.29 ;
      RECT 30.27 5.915 30.44 7.29 ;
      RECT 28.79 7.025 29.08 7.255 ;
      RECT 30.215 5.915 30.505 6.145 ;
      RECT 30.215 5.945 30.675 6.115 ;
      RECT 29.22 1.965 29.57 2.315 ;
      RECT 26.915 2.025 29.57 2.195 ;
      RECT 26.915 1.46 27.085 2.195 ;
      RECT 26.825 1.46 27.165 1.81 ;
      RECT 29.245 6.655 29.57 6.98 ;
      RECT 23.805 6.61 24.155 6.96 ;
      RECT 29.22 6.655 29.57 6.885 ;
      RECT 23.605 6.655 24.155 6.885 ;
      RECT 23.435 6.685 29.57 6.855 ;
      RECT 28.445 2.365 28.765 2.685 ;
      RECT 28.415 2.365 28.765 2.595 ;
      RECT 28.245 2.395 28.765 2.565 ;
      RECT 28.445 6.255 28.765 6.545 ;
      RECT 28.415 6.285 28.765 6.515 ;
      RECT 28.245 6.315 28.765 6.485 ;
      RECT 27.405 2.705 27.745 3.055 ;
      RECT 27.405 2.765 27.88 2.935 ;
      RECT 27.395 5.84 27.735 6.19 ;
      RECT 21.805 5.915 22.095 6.145 ;
      RECT 21.805 5.945 27.88 6.115 ;
      RECT 24.9 2.465 25.19 2.695 ;
      RECT 24.9 2.465 25.355 2.65 ;
      RECT 25.215 2.37 25.835 2.51 ;
      RECT 25.605 2.17 25.925 2.43 ;
      RECT 24.285 2.45 24.605 2.71 ;
      RECT 24.285 2.45 24.75 2.695 ;
      RECT 24.61 2.07 24.75 2.695 ;
      RECT 24.61 2.07 24.875 2.21 ;
      RECT 25.14 1.905 25.43 2.135 ;
      RECT 24.735 1.95 25.43 2.09 ;
      RECT 24.18 3.29 24.47 3.815 ;
      RECT 24.165 3.29 24.485 3.55 ;
      RECT 23.905 1.89 24.225 2.15 ;
      RECT 23.905 1.905 24.47 2.135 ;
      RECT 23.18 3.585 23.47 3.815 ;
      RECT 23.375 2.23 23.515 3.77 ;
      RECT 23.42 2.185 23.71 2.415 ;
      RECT 23.015 2.23 23.71 2.37 ;
      RECT 23.015 2.07 23.155 2.37 ;
      RECT 21.555 2.07 23.155 2.21 ;
      RECT 21.465 1.89 21.785 2.15 ;
      RECT 21.465 1.905 22.03 2.15 ;
      RECT 23.175 7.765 23.465 7.995 ;
      RECT 23.235 7.025 23.405 7.995 ;
      RECT 23.155 7.075 23.525 7.425 ;
      RECT 23.155 7.055 23.465 7.425 ;
      RECT 23.175 7.025 23.465 7.425 ;
      RECT 20.575 2.93 23.155 3.07 ;
      RECT 22.94 2.745 23.23 2.975 ;
      RECT 20.5 2.745 21.165 2.975 ;
      RECT 20.845 2.73 21.165 3.07 ;
      RECT 21.845 2.45 22.165 2.71 ;
      RECT 21.845 2.465 22.27 2.695 ;
      RECT 20.485 2.17 20.805 2.43 ;
      RECT 20.98 2.185 21.27 2.415 ;
      RECT 20.485 2.23 21.27 2.37 ;
      RECT 20.605 3.29 20.925 3.55 ;
      RECT 19.765 3.29 20.085 3.55 ;
      RECT 20.605 3.305 21.03 3.535 ;
      RECT 19.765 3.35 21.03 3.49 ;
      RECT 19.3 3.025 19.59 3.255 ;
      RECT 19.375 1.95 19.515 3.255 ;
      RECT 19.025 2.45 19.515 2.71 ;
      RECT 18.78 2.465 19.515 2.695 ;
      RECT 19.78 1.905 20.07 2.135 ;
      RECT 19.375 1.95 20.07 2.09 ;
      RECT 18.54 3.305 18.83 3.535 ;
      RECT 18.54 3.305 18.995 3.49 ;
      RECT 18.855 2.93 18.995 3.49 ;
      RECT 18.495 2.93 18.995 3.07 ;
      RECT 18.495 1.95 18.635 3.07 ;
      RECT 18.285 1.89 18.605 2.15 ;
      RECT 18.045 3.57 18.365 3.83 ;
      RECT 17.34 3.585 17.63 3.815 ;
      RECT 17.34 3.63 18.365 3.77 ;
      RECT 17.415 3.58 17.675 3.77 ;
      RECT 17.805 2.45 18.125 2.71 ;
      RECT 17.805 2.465 18.35 2.695 ;
      RECT 17.805 3.01 18.125 3.27 ;
      RECT 17.805 3.025 18.35 3.255 ;
      RECT 16.845 3.01 17.165 3.27 ;
      RECT 16.935 1.95 17.075 3.27 ;
      RECT 17.34 1.905 17.63 2.135 ;
      RECT 16.935 1.95 17.63 2.09 ;
      RECT 15.25 7.765 15.54 7.995 ;
      RECT 15.31 6.285 15.48 7.995 ;
      RECT 15.3 6.655 15.65 7.005 ;
      RECT 15.25 6.285 15.54 6.515 ;
      RECT 15.25 2.365 15.54 2.595 ;
      RECT 15.31 0.885 15.48 2.595 ;
      RECT 15.25 0.885 15.54 1.115 ;
      RECT 14.84 2.735 15.17 2.965 ;
      RECT 14.84 2.765 15.34 2.935 ;
      RECT 14.84 2.395 15.03 2.965 ;
      RECT 14.26 2.365 14.55 2.595 ;
      RECT 14.26 2.395 15.03 2.565 ;
      RECT 14.32 0.885 14.49 2.595 ;
      RECT 14.26 0.885 14.55 1.115 ;
      RECT 14.26 7.765 14.55 7.995 ;
      RECT 14.32 6.285 14.49 7.995 ;
      RECT 14.26 6.285 14.55 6.515 ;
      RECT 14.26 6.325 15.11 6.485 ;
      RECT 14.94 5.915 15.11 6.485 ;
      RECT 14.26 6.32 14.65 6.485 ;
      RECT 14.88 5.915 15.17 6.145 ;
      RECT 14.88 5.945 15.34 6.115 ;
      RECT 13.89 2.735 14.18 2.965 ;
      RECT 13.89 2.765 14.35 2.935 ;
      RECT 13.95 1.655 14.115 2.965 ;
      RECT 12.465 1.625 12.755 1.855 ;
      RECT 12.465 1.655 14.115 1.825 ;
      RECT 12.525 0.885 12.695 1.855 ;
      RECT 12.465 0.885 12.755 1.115 ;
      RECT 12.465 7.765 12.755 7.995 ;
      RECT 12.525 7.025 12.695 7.995 ;
      RECT 12.525 7.12 14.115 7.29 ;
      RECT 13.945 5.915 14.115 7.29 ;
      RECT 12.465 7.025 12.755 7.255 ;
      RECT 13.89 5.915 14.18 6.145 ;
      RECT 13.89 5.945 14.35 6.115 ;
      RECT 12.895 1.965 13.245 2.315 ;
      RECT 10.59 2.025 13.245 2.195 ;
      RECT 10.59 1.46 10.76 2.195 ;
      RECT 10.5 1.46 10.84 1.81 ;
      RECT 12.92 6.655 13.245 6.98 ;
      RECT 8.315 6.605 8.665 6.955 ;
      RECT 12.895 6.655 13.245 6.885 ;
      RECT 7.28 6.655 7.57 6.885 ;
      RECT 7.11 6.685 13.245 6.855 ;
      RECT 12.12 2.365 12.44 2.685 ;
      RECT 12.09 2.365 12.44 2.595 ;
      RECT 11.92 2.395 12.44 2.565 ;
      RECT 12.12 6.255 12.44 6.545 ;
      RECT 12.09 6.285 12.44 6.515 ;
      RECT 11.92 6.315 12.44 6.485 ;
      RECT 11.08 2.705 11.42 3.055 ;
      RECT 11.08 2.765 11.555 2.935 ;
      RECT 11.07 5.84 11.41 6.19 ;
      RECT 5.48 5.915 5.77 6.145 ;
      RECT 5.48 5.945 11.555 6.115 ;
      RECT 8.575 2.465 8.865 2.695 ;
      RECT 8.575 2.465 9.03 2.65 ;
      RECT 8.89 2.37 9.51 2.51 ;
      RECT 9.28 2.17 9.6 2.43 ;
      RECT 7.96 2.45 8.28 2.71 ;
      RECT 7.96 2.45 8.425 2.695 ;
      RECT 8.285 2.07 8.425 2.695 ;
      RECT 8.285 2.07 8.55 2.21 ;
      RECT 8.815 1.905 9.105 2.135 ;
      RECT 8.41 1.95 9.105 2.09 ;
      RECT 7.855 3.29 8.145 3.815 ;
      RECT 7.84 3.29 8.16 3.55 ;
      RECT 7.58 1.89 7.9 2.15 ;
      RECT 7.58 1.905 8.145 2.135 ;
      RECT 6.855 3.585 7.145 3.815 ;
      RECT 7.05 2.23 7.19 3.77 ;
      RECT 7.095 2.185 7.385 2.415 ;
      RECT 6.69 2.23 7.385 2.37 ;
      RECT 6.69 2.07 6.83 2.37 ;
      RECT 5.23 2.07 6.83 2.21 ;
      RECT 5.14 1.89 5.46 2.15 ;
      RECT 5.14 1.905 5.705 2.15 ;
      RECT 6.85 7.765 7.14 7.995 ;
      RECT 6.91 7.025 7.08 7.995 ;
      RECT 6.83 7.075 7.2 7.425 ;
      RECT 6.83 7.055 7.14 7.425 ;
      RECT 6.85 7.025 7.14 7.425 ;
      RECT 4.25 2.93 6.83 3.07 ;
      RECT 6.615 2.745 6.905 2.975 ;
      RECT 4.175 2.745 4.84 2.975 ;
      RECT 4.52 2.73 4.84 3.07 ;
      RECT 5.52 2.45 5.84 2.71 ;
      RECT 5.52 2.465 5.945 2.695 ;
      RECT 4.16 2.17 4.48 2.43 ;
      RECT 4.655 2.185 4.945 2.415 ;
      RECT 4.16 2.23 4.945 2.37 ;
      RECT 4.28 3.29 4.6 3.55 ;
      RECT 3.44 3.29 3.76 3.55 ;
      RECT 4.28 3.305 4.705 3.535 ;
      RECT 3.44 3.35 4.705 3.49 ;
      RECT 2.975 3.025 3.265 3.255 ;
      RECT 3.05 1.95 3.19 3.255 ;
      RECT 2.7 2.45 3.19 2.71 ;
      RECT 2.455 2.465 3.19 2.695 ;
      RECT 3.455 1.905 3.745 2.135 ;
      RECT 3.05 1.95 3.745 2.09 ;
      RECT 2.215 3.305 2.505 3.535 ;
      RECT 2.215 3.305 2.67 3.49 ;
      RECT 2.53 2.93 2.67 3.49 ;
      RECT 2.17 2.93 2.67 3.07 ;
      RECT 2.17 1.95 2.31 3.07 ;
      RECT 1.96 1.89 2.28 2.15 ;
      RECT 1.72 3.57 2.04 3.83 ;
      RECT 1.015 3.585 1.305 3.815 ;
      RECT 1.015 3.63 2.04 3.77 ;
      RECT 1.09 3.58 1.35 3.77 ;
      RECT 1.48 2.45 1.8 2.71 ;
      RECT 1.48 2.465 2.025 2.695 ;
      RECT 1.48 3.01 1.8 3.27 ;
      RECT 1.48 3.025 2.025 3.255 ;
      RECT 0.52 3.01 0.84 3.27 ;
      RECT 0.61 1.95 0.75 3.27 ;
      RECT 1.015 1.905 1.305 2.135 ;
      RECT 0.61 1.95 1.305 2.09 ;
      RECT -1.3 6.655 -1.01 6.885 ;
      RECT -1.47 6.685 -1.01 6.855 ;
      RECT -1.73 7.765 -1.44 7.995 ;
      RECT -1.67 7.025 -1.5 7.995 ;
      RECT -1.76 7.025 -1.41 7.315 ;
      RECT -2.135 6.285 -1.785 6.575 ;
      RECT -2.275 6.315 -1.785 6.485 ;
      RECT -3.1 5.915 -2.81 6.145 ;
      RECT -3.1 5.945 -2.64 6.115 ;
      RECT 71.42 2.45 71.74 2.71 ;
      RECT 68.98 2.45 69.3 2.71 ;
      RECT 55.095 2.45 55.415 2.71 ;
      RECT 52.655 2.45 52.975 2.71 ;
      RECT 38.77 2.45 39.09 2.71 ;
      RECT 36.33 2.45 36.65 2.71 ;
      RECT 22.445 2.45 22.765 2.71 ;
      RECT 20.005 2.45 20.325 2.71 ;
      RECT 6.12 2.45 6.44 2.71 ;
      RECT 3.68 2.45 4 2.71 ;
    LAYER mcon ;
      RECT 80.61 0.915 80.78 1.085 ;
      RECT 80.61 2.395 80.78 2.565 ;
      RECT 80.61 6.315 80.78 6.485 ;
      RECT 80.61 7.795 80.78 7.965 ;
      RECT 80.26 0.105 80.43 0.275 ;
      RECT 80.26 4.165 80.43 4.335 ;
      RECT 80.26 4.545 80.43 4.715 ;
      RECT 80.26 8.605 80.43 8.775 ;
      RECT 80.24 2.765 80.41 2.935 ;
      RECT 80.24 5.945 80.41 6.115 ;
      RECT 79.62 0.915 79.79 1.085 ;
      RECT 79.62 2.395 79.79 2.565 ;
      RECT 79.62 6.315 79.79 6.485 ;
      RECT 79.62 7.795 79.79 7.965 ;
      RECT 79.27 0.105 79.44 0.275 ;
      RECT 79.27 4.165 79.44 4.335 ;
      RECT 79.27 4.545 79.44 4.715 ;
      RECT 79.27 8.605 79.44 8.775 ;
      RECT 79.25 2.765 79.42 2.935 ;
      RECT 79.25 5.945 79.42 6.115 ;
      RECT 78.565 0.105 78.735 0.275 ;
      RECT 78.565 4.165 78.735 4.335 ;
      RECT 78.565 4.545 78.735 4.715 ;
      RECT 78.565 8.605 78.735 8.775 ;
      RECT 78.255 2.025 78.425 2.195 ;
      RECT 78.255 6.685 78.425 6.855 ;
      RECT 77.885 0.105 78.055 0.275 ;
      RECT 77.885 8.605 78.055 8.775 ;
      RECT 77.825 0.915 77.995 1.085 ;
      RECT 77.825 1.655 77.995 1.825 ;
      RECT 77.825 7.055 77.995 7.225 ;
      RECT 77.825 7.795 77.995 7.965 ;
      RECT 77.45 2.395 77.62 2.565 ;
      RECT 77.45 6.315 77.62 6.485 ;
      RECT 77.205 0.105 77.375 0.275 ;
      RECT 77.205 8.605 77.375 8.775 ;
      RECT 76.525 0.105 76.695 0.275 ;
      RECT 76.525 8.605 76.695 8.775 ;
      RECT 76.455 2.765 76.625 2.935 ;
      RECT 76.455 5.945 76.625 6.115 ;
      RECT 74.91 1.415 75.08 1.585 ;
      RECT 74.91 4.135 75.08 4.305 ;
      RECT 74.655 2.775 74.825 2.945 ;
      RECT 74.45 1.415 74.62 1.585 ;
      RECT 74.45 4.135 74.62 4.305 ;
      RECT 74.175 1.935 74.345 2.105 ;
      RECT 73.99 1.415 74.16 1.585 ;
      RECT 73.99 4.135 74.16 4.305 ;
      RECT 73.935 2.495 74.105 2.665 ;
      RECT 73.53 1.415 73.7 1.585 ;
      RECT 73.53 4.135 73.7 4.305 ;
      RECT 73.455 2.495 73.625 2.665 ;
      RECT 73.215 1.935 73.385 2.105 ;
      RECT 73.215 3.615 73.385 3.785 ;
      RECT 73.07 1.415 73.24 1.585 ;
      RECT 73.07 4.135 73.24 4.305 ;
      RECT 72.95 4.545 73.12 4.715 ;
      RECT 72.95 8.605 73.12 8.775 ;
      RECT 72.695 2.775 72.865 2.945 ;
      RECT 72.64 6.685 72.81 6.855 ;
      RECT 72.61 1.415 72.78 1.585 ;
      RECT 72.61 4.135 72.78 4.305 ;
      RECT 72.455 2.215 72.625 2.385 ;
      RECT 72.27 8.605 72.44 8.775 ;
      RECT 72.215 3.615 72.385 3.785 ;
      RECT 72.21 7.055 72.38 7.225 ;
      RECT 72.21 7.795 72.38 7.965 ;
      RECT 72.15 1.415 72.32 1.585 ;
      RECT 72.15 4.135 72.32 4.305 ;
      RECT 71.975 2.775 72.145 2.945 ;
      RECT 71.835 6.315 72.005 6.485 ;
      RECT 71.69 1.415 71.86 1.585 ;
      RECT 71.69 4.135 71.86 4.305 ;
      RECT 71.59 8.605 71.76 8.775 ;
      RECT 71.495 2.495 71.665 2.665 ;
      RECT 71.23 1.415 71.4 1.585 ;
      RECT 71.23 4.135 71.4 4.305 ;
      RECT 71.015 2.495 71.185 2.665 ;
      RECT 70.91 8.605 71.08 8.775 ;
      RECT 70.84 5.945 71.01 6.115 ;
      RECT 70.775 1.935 70.945 2.105 ;
      RECT 70.77 1.415 70.94 1.585 ;
      RECT 70.77 4.135 70.94 4.305 ;
      RECT 70.31 1.415 70.48 1.585 ;
      RECT 70.31 4.135 70.48 4.305 ;
      RECT 70.015 2.215 70.185 2.385 ;
      RECT 69.85 1.415 70.02 1.585 ;
      RECT 69.85 4.135 70.02 4.305 ;
      RECT 69.775 3.335 69.945 3.505 ;
      RECT 69.535 2.775 69.705 2.945 ;
      RECT 69.39 1.415 69.56 1.585 ;
      RECT 69.39 4.135 69.56 4.305 ;
      RECT 69.055 2.495 69.225 2.665 ;
      RECT 68.93 1.415 69.1 1.585 ;
      RECT 68.93 4.135 69.1 4.305 ;
      RECT 68.815 1.935 68.985 2.105 ;
      RECT 68.815 3.335 68.985 3.505 ;
      RECT 68.47 1.415 68.64 1.585 ;
      RECT 68.47 4.135 68.64 4.305 ;
      RECT 68.335 3.055 68.505 3.225 ;
      RECT 68.01 1.415 68.18 1.585 ;
      RECT 68.01 4.135 68.18 4.305 ;
      RECT 67.815 2.495 67.985 2.665 ;
      RECT 67.575 3.335 67.745 3.505 ;
      RECT 67.55 1.415 67.72 1.585 ;
      RECT 67.55 4.135 67.72 4.305 ;
      RECT 67.335 1.935 67.505 2.105 ;
      RECT 67.095 2.495 67.265 2.665 ;
      RECT 67.095 3.055 67.265 3.225 ;
      RECT 67.09 1.415 67.26 1.585 ;
      RECT 67.09 4.135 67.26 4.305 ;
      RECT 66.63 1.415 66.8 1.585 ;
      RECT 66.63 4.135 66.8 4.305 ;
      RECT 66.375 1.935 66.545 2.105 ;
      RECT 66.375 3.615 66.545 3.785 ;
      RECT 66.17 1.415 66.34 1.585 ;
      RECT 66.17 4.135 66.34 4.305 ;
      RECT 65.895 3.055 66.065 3.225 ;
      RECT 65.71 1.415 65.88 1.585 ;
      RECT 65.71 4.135 65.88 4.305 ;
      RECT 64.285 0.915 64.455 1.085 ;
      RECT 64.285 2.395 64.455 2.565 ;
      RECT 64.285 6.315 64.455 6.485 ;
      RECT 64.285 7.795 64.455 7.965 ;
      RECT 63.935 0.105 64.105 0.275 ;
      RECT 63.935 4.165 64.105 4.335 ;
      RECT 63.935 4.545 64.105 4.715 ;
      RECT 63.935 8.605 64.105 8.775 ;
      RECT 63.915 2.765 64.085 2.935 ;
      RECT 63.915 5.945 64.085 6.115 ;
      RECT 63.295 0.915 63.465 1.085 ;
      RECT 63.295 2.395 63.465 2.565 ;
      RECT 63.295 6.315 63.465 6.485 ;
      RECT 63.295 7.795 63.465 7.965 ;
      RECT 62.945 0.105 63.115 0.275 ;
      RECT 62.945 4.165 63.115 4.335 ;
      RECT 62.945 4.545 63.115 4.715 ;
      RECT 62.945 8.605 63.115 8.775 ;
      RECT 62.925 2.765 63.095 2.935 ;
      RECT 62.925 5.945 63.095 6.115 ;
      RECT 62.24 0.105 62.41 0.275 ;
      RECT 62.24 4.165 62.41 4.335 ;
      RECT 62.24 4.545 62.41 4.715 ;
      RECT 62.24 8.605 62.41 8.775 ;
      RECT 61.93 2.025 62.1 2.195 ;
      RECT 61.93 6.685 62.1 6.855 ;
      RECT 61.56 0.105 61.73 0.275 ;
      RECT 61.56 8.605 61.73 8.775 ;
      RECT 61.5 0.915 61.67 1.085 ;
      RECT 61.5 1.655 61.67 1.825 ;
      RECT 61.5 7.055 61.67 7.225 ;
      RECT 61.5 7.795 61.67 7.965 ;
      RECT 61.125 2.395 61.295 2.565 ;
      RECT 61.125 6.315 61.295 6.485 ;
      RECT 60.88 0.105 61.05 0.275 ;
      RECT 60.88 8.605 61.05 8.775 ;
      RECT 60.2 0.105 60.37 0.275 ;
      RECT 60.2 8.605 60.37 8.775 ;
      RECT 60.13 2.765 60.3 2.935 ;
      RECT 60.13 5.945 60.3 6.115 ;
      RECT 58.585 1.415 58.755 1.585 ;
      RECT 58.585 4.135 58.755 4.305 ;
      RECT 58.33 2.775 58.5 2.945 ;
      RECT 58.125 1.415 58.295 1.585 ;
      RECT 58.125 4.135 58.295 4.305 ;
      RECT 57.85 1.935 58.02 2.105 ;
      RECT 57.665 1.415 57.835 1.585 ;
      RECT 57.665 4.135 57.835 4.305 ;
      RECT 57.61 2.495 57.78 2.665 ;
      RECT 57.205 1.415 57.375 1.585 ;
      RECT 57.205 4.135 57.375 4.305 ;
      RECT 57.13 2.495 57.3 2.665 ;
      RECT 56.89 1.935 57.06 2.105 ;
      RECT 56.89 3.615 57.06 3.785 ;
      RECT 56.745 1.415 56.915 1.585 ;
      RECT 56.745 4.135 56.915 4.305 ;
      RECT 56.625 4.545 56.795 4.715 ;
      RECT 56.625 8.605 56.795 8.775 ;
      RECT 56.37 2.775 56.54 2.945 ;
      RECT 56.315 6.685 56.485 6.855 ;
      RECT 56.285 1.415 56.455 1.585 ;
      RECT 56.285 4.135 56.455 4.305 ;
      RECT 56.13 2.215 56.3 2.385 ;
      RECT 55.945 8.605 56.115 8.775 ;
      RECT 55.89 3.615 56.06 3.785 ;
      RECT 55.885 7.055 56.055 7.225 ;
      RECT 55.885 7.795 56.055 7.965 ;
      RECT 55.825 1.415 55.995 1.585 ;
      RECT 55.825 4.135 55.995 4.305 ;
      RECT 55.65 2.775 55.82 2.945 ;
      RECT 55.51 6.315 55.68 6.485 ;
      RECT 55.365 1.415 55.535 1.585 ;
      RECT 55.365 4.135 55.535 4.305 ;
      RECT 55.265 8.605 55.435 8.775 ;
      RECT 55.17 2.495 55.34 2.665 ;
      RECT 54.905 1.415 55.075 1.585 ;
      RECT 54.905 4.135 55.075 4.305 ;
      RECT 54.69 2.495 54.86 2.665 ;
      RECT 54.585 8.605 54.755 8.775 ;
      RECT 54.515 5.945 54.685 6.115 ;
      RECT 54.45 1.935 54.62 2.105 ;
      RECT 54.445 1.415 54.615 1.585 ;
      RECT 54.445 4.135 54.615 4.305 ;
      RECT 53.985 1.415 54.155 1.585 ;
      RECT 53.985 4.135 54.155 4.305 ;
      RECT 53.69 2.215 53.86 2.385 ;
      RECT 53.525 1.415 53.695 1.585 ;
      RECT 53.525 4.135 53.695 4.305 ;
      RECT 53.45 3.335 53.62 3.505 ;
      RECT 53.21 2.775 53.38 2.945 ;
      RECT 53.065 1.415 53.235 1.585 ;
      RECT 53.065 4.135 53.235 4.305 ;
      RECT 52.73 2.495 52.9 2.665 ;
      RECT 52.605 1.415 52.775 1.585 ;
      RECT 52.605 4.135 52.775 4.305 ;
      RECT 52.49 1.935 52.66 2.105 ;
      RECT 52.49 3.335 52.66 3.505 ;
      RECT 52.145 1.415 52.315 1.585 ;
      RECT 52.145 4.135 52.315 4.305 ;
      RECT 52.01 3.055 52.18 3.225 ;
      RECT 51.685 1.415 51.855 1.585 ;
      RECT 51.685 4.135 51.855 4.305 ;
      RECT 51.49 2.495 51.66 2.665 ;
      RECT 51.25 3.335 51.42 3.505 ;
      RECT 51.225 1.415 51.395 1.585 ;
      RECT 51.225 4.135 51.395 4.305 ;
      RECT 51.01 1.935 51.18 2.105 ;
      RECT 50.77 2.495 50.94 2.665 ;
      RECT 50.77 3.055 50.94 3.225 ;
      RECT 50.765 1.415 50.935 1.585 ;
      RECT 50.765 4.135 50.935 4.305 ;
      RECT 50.305 1.415 50.475 1.585 ;
      RECT 50.305 4.135 50.475 4.305 ;
      RECT 50.05 1.935 50.22 2.105 ;
      RECT 50.05 3.615 50.22 3.785 ;
      RECT 49.845 1.415 50.015 1.585 ;
      RECT 49.845 4.135 50.015 4.305 ;
      RECT 49.57 3.055 49.74 3.225 ;
      RECT 49.385 1.415 49.555 1.585 ;
      RECT 49.385 4.135 49.555 4.305 ;
      RECT 47.96 0.915 48.13 1.085 ;
      RECT 47.96 2.395 48.13 2.565 ;
      RECT 47.96 6.315 48.13 6.485 ;
      RECT 47.96 7.795 48.13 7.965 ;
      RECT 47.61 0.105 47.78 0.275 ;
      RECT 47.61 4.165 47.78 4.335 ;
      RECT 47.61 4.545 47.78 4.715 ;
      RECT 47.61 8.605 47.78 8.775 ;
      RECT 47.59 2.765 47.76 2.935 ;
      RECT 47.59 5.945 47.76 6.115 ;
      RECT 46.97 0.915 47.14 1.085 ;
      RECT 46.97 2.395 47.14 2.565 ;
      RECT 46.97 6.315 47.14 6.485 ;
      RECT 46.97 7.795 47.14 7.965 ;
      RECT 46.62 0.105 46.79 0.275 ;
      RECT 46.62 4.165 46.79 4.335 ;
      RECT 46.62 4.545 46.79 4.715 ;
      RECT 46.62 8.605 46.79 8.775 ;
      RECT 46.6 2.765 46.77 2.935 ;
      RECT 46.6 5.945 46.77 6.115 ;
      RECT 45.915 0.105 46.085 0.275 ;
      RECT 45.915 4.165 46.085 4.335 ;
      RECT 45.915 4.545 46.085 4.715 ;
      RECT 45.915 8.605 46.085 8.775 ;
      RECT 45.605 2.025 45.775 2.195 ;
      RECT 45.605 6.685 45.775 6.855 ;
      RECT 45.235 0.105 45.405 0.275 ;
      RECT 45.235 8.605 45.405 8.775 ;
      RECT 45.175 0.915 45.345 1.085 ;
      RECT 45.175 1.655 45.345 1.825 ;
      RECT 45.175 7.055 45.345 7.225 ;
      RECT 45.175 7.795 45.345 7.965 ;
      RECT 44.8 2.395 44.97 2.565 ;
      RECT 44.8 6.315 44.97 6.485 ;
      RECT 44.555 0.105 44.725 0.275 ;
      RECT 44.555 8.605 44.725 8.775 ;
      RECT 43.875 0.105 44.045 0.275 ;
      RECT 43.875 8.605 44.045 8.775 ;
      RECT 43.805 2.765 43.975 2.935 ;
      RECT 43.805 5.945 43.975 6.115 ;
      RECT 42.26 1.415 42.43 1.585 ;
      RECT 42.26 4.135 42.43 4.305 ;
      RECT 42.005 2.775 42.175 2.945 ;
      RECT 41.8 1.415 41.97 1.585 ;
      RECT 41.8 4.135 41.97 4.305 ;
      RECT 41.525 1.935 41.695 2.105 ;
      RECT 41.34 1.415 41.51 1.585 ;
      RECT 41.34 4.135 41.51 4.305 ;
      RECT 41.285 2.495 41.455 2.665 ;
      RECT 40.88 1.415 41.05 1.585 ;
      RECT 40.88 4.135 41.05 4.305 ;
      RECT 40.805 2.495 40.975 2.665 ;
      RECT 40.565 1.935 40.735 2.105 ;
      RECT 40.565 3.615 40.735 3.785 ;
      RECT 40.42 1.415 40.59 1.585 ;
      RECT 40.42 4.135 40.59 4.305 ;
      RECT 40.3 4.545 40.47 4.715 ;
      RECT 40.3 8.605 40.47 8.775 ;
      RECT 40.045 2.775 40.215 2.945 ;
      RECT 39.99 6.685 40.16 6.855 ;
      RECT 39.96 1.415 40.13 1.585 ;
      RECT 39.96 4.135 40.13 4.305 ;
      RECT 39.805 2.215 39.975 2.385 ;
      RECT 39.62 8.605 39.79 8.775 ;
      RECT 39.565 3.615 39.735 3.785 ;
      RECT 39.56 7.055 39.73 7.225 ;
      RECT 39.56 7.795 39.73 7.965 ;
      RECT 39.5 1.415 39.67 1.585 ;
      RECT 39.5 4.135 39.67 4.305 ;
      RECT 39.325 2.775 39.495 2.945 ;
      RECT 39.185 6.315 39.355 6.485 ;
      RECT 39.04 1.415 39.21 1.585 ;
      RECT 39.04 4.135 39.21 4.305 ;
      RECT 38.94 8.605 39.11 8.775 ;
      RECT 38.845 2.495 39.015 2.665 ;
      RECT 38.58 1.415 38.75 1.585 ;
      RECT 38.58 4.135 38.75 4.305 ;
      RECT 38.365 2.495 38.535 2.665 ;
      RECT 38.26 8.605 38.43 8.775 ;
      RECT 38.19 5.945 38.36 6.115 ;
      RECT 38.125 1.935 38.295 2.105 ;
      RECT 38.12 1.415 38.29 1.585 ;
      RECT 38.12 4.135 38.29 4.305 ;
      RECT 37.66 1.415 37.83 1.585 ;
      RECT 37.66 4.135 37.83 4.305 ;
      RECT 37.365 2.215 37.535 2.385 ;
      RECT 37.2 1.415 37.37 1.585 ;
      RECT 37.2 4.135 37.37 4.305 ;
      RECT 37.125 3.335 37.295 3.505 ;
      RECT 36.885 2.775 37.055 2.945 ;
      RECT 36.74 1.415 36.91 1.585 ;
      RECT 36.74 4.135 36.91 4.305 ;
      RECT 36.405 2.495 36.575 2.665 ;
      RECT 36.28 1.415 36.45 1.585 ;
      RECT 36.28 4.135 36.45 4.305 ;
      RECT 36.165 1.935 36.335 2.105 ;
      RECT 36.165 3.335 36.335 3.505 ;
      RECT 35.82 1.415 35.99 1.585 ;
      RECT 35.82 4.135 35.99 4.305 ;
      RECT 35.685 3.055 35.855 3.225 ;
      RECT 35.36 1.415 35.53 1.585 ;
      RECT 35.36 4.135 35.53 4.305 ;
      RECT 35.165 2.495 35.335 2.665 ;
      RECT 34.925 3.335 35.095 3.505 ;
      RECT 34.9 1.415 35.07 1.585 ;
      RECT 34.9 4.135 35.07 4.305 ;
      RECT 34.685 1.935 34.855 2.105 ;
      RECT 34.445 2.495 34.615 2.665 ;
      RECT 34.445 3.055 34.615 3.225 ;
      RECT 34.44 1.415 34.61 1.585 ;
      RECT 34.44 4.135 34.61 4.305 ;
      RECT 33.98 1.415 34.15 1.585 ;
      RECT 33.98 4.135 34.15 4.305 ;
      RECT 33.725 1.935 33.895 2.105 ;
      RECT 33.725 3.615 33.895 3.785 ;
      RECT 33.52 1.415 33.69 1.585 ;
      RECT 33.52 4.135 33.69 4.305 ;
      RECT 33.245 3.055 33.415 3.225 ;
      RECT 33.06 1.415 33.23 1.585 ;
      RECT 33.06 4.135 33.23 4.305 ;
      RECT 31.635 0.915 31.805 1.085 ;
      RECT 31.635 2.395 31.805 2.565 ;
      RECT 31.635 6.315 31.805 6.485 ;
      RECT 31.635 7.795 31.805 7.965 ;
      RECT 31.285 0.105 31.455 0.275 ;
      RECT 31.285 4.165 31.455 4.335 ;
      RECT 31.285 4.545 31.455 4.715 ;
      RECT 31.285 8.605 31.455 8.775 ;
      RECT 31.265 2.765 31.435 2.935 ;
      RECT 31.265 5.945 31.435 6.115 ;
      RECT 30.645 0.915 30.815 1.085 ;
      RECT 30.645 2.395 30.815 2.565 ;
      RECT 30.645 6.315 30.815 6.485 ;
      RECT 30.645 7.795 30.815 7.965 ;
      RECT 30.295 0.105 30.465 0.275 ;
      RECT 30.295 4.165 30.465 4.335 ;
      RECT 30.295 4.545 30.465 4.715 ;
      RECT 30.295 8.605 30.465 8.775 ;
      RECT 30.275 2.765 30.445 2.935 ;
      RECT 30.275 5.945 30.445 6.115 ;
      RECT 29.59 0.105 29.76 0.275 ;
      RECT 29.59 4.165 29.76 4.335 ;
      RECT 29.59 4.545 29.76 4.715 ;
      RECT 29.59 8.605 29.76 8.775 ;
      RECT 29.28 2.025 29.45 2.195 ;
      RECT 29.28 6.685 29.45 6.855 ;
      RECT 28.91 0.105 29.08 0.275 ;
      RECT 28.91 8.605 29.08 8.775 ;
      RECT 28.85 0.915 29.02 1.085 ;
      RECT 28.85 1.655 29.02 1.825 ;
      RECT 28.85 7.055 29.02 7.225 ;
      RECT 28.85 7.795 29.02 7.965 ;
      RECT 28.475 2.395 28.645 2.565 ;
      RECT 28.475 6.315 28.645 6.485 ;
      RECT 28.23 0.105 28.4 0.275 ;
      RECT 28.23 8.605 28.4 8.775 ;
      RECT 27.55 0.105 27.72 0.275 ;
      RECT 27.55 8.605 27.72 8.775 ;
      RECT 27.48 2.765 27.65 2.935 ;
      RECT 27.48 5.945 27.65 6.115 ;
      RECT 25.935 1.415 26.105 1.585 ;
      RECT 25.935 4.135 26.105 4.305 ;
      RECT 25.68 2.775 25.85 2.945 ;
      RECT 25.475 1.415 25.645 1.585 ;
      RECT 25.475 4.135 25.645 4.305 ;
      RECT 25.2 1.935 25.37 2.105 ;
      RECT 25.015 1.415 25.185 1.585 ;
      RECT 25.015 4.135 25.185 4.305 ;
      RECT 24.96 2.495 25.13 2.665 ;
      RECT 24.555 1.415 24.725 1.585 ;
      RECT 24.555 4.135 24.725 4.305 ;
      RECT 24.48 2.495 24.65 2.665 ;
      RECT 24.24 1.935 24.41 2.105 ;
      RECT 24.24 3.615 24.41 3.785 ;
      RECT 24.095 1.415 24.265 1.585 ;
      RECT 24.095 4.135 24.265 4.305 ;
      RECT 23.975 4.545 24.145 4.715 ;
      RECT 23.975 8.605 24.145 8.775 ;
      RECT 23.72 2.775 23.89 2.945 ;
      RECT 23.665 6.685 23.835 6.855 ;
      RECT 23.635 1.415 23.805 1.585 ;
      RECT 23.635 4.135 23.805 4.305 ;
      RECT 23.48 2.215 23.65 2.385 ;
      RECT 23.295 8.605 23.465 8.775 ;
      RECT 23.24 3.615 23.41 3.785 ;
      RECT 23.235 7.055 23.405 7.225 ;
      RECT 23.235 7.795 23.405 7.965 ;
      RECT 23.175 1.415 23.345 1.585 ;
      RECT 23.175 4.135 23.345 4.305 ;
      RECT 23 2.775 23.17 2.945 ;
      RECT 22.86 6.315 23.03 6.485 ;
      RECT 22.715 1.415 22.885 1.585 ;
      RECT 22.715 4.135 22.885 4.305 ;
      RECT 22.615 8.605 22.785 8.775 ;
      RECT 22.52 2.495 22.69 2.665 ;
      RECT 22.255 1.415 22.425 1.585 ;
      RECT 22.255 4.135 22.425 4.305 ;
      RECT 22.04 2.495 22.21 2.665 ;
      RECT 21.935 8.605 22.105 8.775 ;
      RECT 21.865 5.945 22.035 6.115 ;
      RECT 21.8 1.935 21.97 2.105 ;
      RECT 21.795 1.415 21.965 1.585 ;
      RECT 21.795 4.135 21.965 4.305 ;
      RECT 21.335 1.415 21.505 1.585 ;
      RECT 21.335 4.135 21.505 4.305 ;
      RECT 21.04 2.215 21.21 2.385 ;
      RECT 20.875 1.415 21.045 1.585 ;
      RECT 20.875 4.135 21.045 4.305 ;
      RECT 20.8 3.335 20.97 3.505 ;
      RECT 20.56 2.775 20.73 2.945 ;
      RECT 20.415 1.415 20.585 1.585 ;
      RECT 20.415 4.135 20.585 4.305 ;
      RECT 20.08 2.495 20.25 2.665 ;
      RECT 19.955 1.415 20.125 1.585 ;
      RECT 19.955 4.135 20.125 4.305 ;
      RECT 19.84 1.935 20.01 2.105 ;
      RECT 19.84 3.335 20.01 3.505 ;
      RECT 19.495 1.415 19.665 1.585 ;
      RECT 19.495 4.135 19.665 4.305 ;
      RECT 19.36 3.055 19.53 3.225 ;
      RECT 19.035 1.415 19.205 1.585 ;
      RECT 19.035 4.135 19.205 4.305 ;
      RECT 18.84 2.495 19.01 2.665 ;
      RECT 18.6 3.335 18.77 3.505 ;
      RECT 18.575 1.415 18.745 1.585 ;
      RECT 18.575 4.135 18.745 4.305 ;
      RECT 18.36 1.935 18.53 2.105 ;
      RECT 18.12 2.495 18.29 2.665 ;
      RECT 18.12 3.055 18.29 3.225 ;
      RECT 18.115 1.415 18.285 1.585 ;
      RECT 18.115 4.135 18.285 4.305 ;
      RECT 17.655 1.415 17.825 1.585 ;
      RECT 17.655 4.135 17.825 4.305 ;
      RECT 17.4 1.935 17.57 2.105 ;
      RECT 17.4 3.615 17.57 3.785 ;
      RECT 17.195 1.415 17.365 1.585 ;
      RECT 17.195 4.135 17.365 4.305 ;
      RECT 16.92 3.055 17.09 3.225 ;
      RECT 16.735 1.415 16.905 1.585 ;
      RECT 16.735 4.135 16.905 4.305 ;
      RECT 15.31 0.915 15.48 1.085 ;
      RECT 15.31 2.395 15.48 2.565 ;
      RECT 15.31 6.315 15.48 6.485 ;
      RECT 15.31 7.795 15.48 7.965 ;
      RECT 14.96 0.105 15.13 0.275 ;
      RECT 14.96 4.165 15.13 4.335 ;
      RECT 14.96 4.545 15.13 4.715 ;
      RECT 14.96 8.605 15.13 8.775 ;
      RECT 14.94 2.765 15.11 2.935 ;
      RECT 14.94 5.945 15.11 6.115 ;
      RECT 14.32 0.915 14.49 1.085 ;
      RECT 14.32 2.395 14.49 2.565 ;
      RECT 14.32 6.315 14.49 6.485 ;
      RECT 14.32 7.795 14.49 7.965 ;
      RECT 13.97 0.105 14.14 0.275 ;
      RECT 13.97 4.165 14.14 4.335 ;
      RECT 13.97 4.545 14.14 4.715 ;
      RECT 13.97 8.605 14.14 8.775 ;
      RECT 13.95 2.765 14.12 2.935 ;
      RECT 13.95 5.945 14.12 6.115 ;
      RECT 13.265 0.105 13.435 0.275 ;
      RECT 13.265 4.165 13.435 4.335 ;
      RECT 13.265 4.545 13.435 4.715 ;
      RECT 13.265 8.605 13.435 8.775 ;
      RECT 12.955 2.025 13.125 2.195 ;
      RECT 12.955 6.685 13.125 6.855 ;
      RECT 12.585 0.105 12.755 0.275 ;
      RECT 12.585 8.605 12.755 8.775 ;
      RECT 12.525 0.915 12.695 1.085 ;
      RECT 12.525 1.655 12.695 1.825 ;
      RECT 12.525 7.055 12.695 7.225 ;
      RECT 12.525 7.795 12.695 7.965 ;
      RECT 12.15 2.395 12.32 2.565 ;
      RECT 12.15 6.315 12.32 6.485 ;
      RECT 11.905 0.105 12.075 0.275 ;
      RECT 11.905 8.605 12.075 8.775 ;
      RECT 11.225 0.105 11.395 0.275 ;
      RECT 11.225 8.605 11.395 8.775 ;
      RECT 11.155 2.765 11.325 2.935 ;
      RECT 11.155 5.945 11.325 6.115 ;
      RECT 9.61 1.415 9.78 1.585 ;
      RECT 9.61 4.135 9.78 4.305 ;
      RECT 9.355 2.775 9.525 2.945 ;
      RECT 9.15 1.415 9.32 1.585 ;
      RECT 9.15 4.135 9.32 4.305 ;
      RECT 8.875 1.935 9.045 2.105 ;
      RECT 8.69 1.415 8.86 1.585 ;
      RECT 8.69 4.135 8.86 4.305 ;
      RECT 8.635 2.495 8.805 2.665 ;
      RECT 8.23 1.415 8.4 1.585 ;
      RECT 8.23 4.135 8.4 4.305 ;
      RECT 8.155 2.495 8.325 2.665 ;
      RECT 7.915 1.935 8.085 2.105 ;
      RECT 7.915 3.615 8.085 3.785 ;
      RECT 7.77 1.415 7.94 1.585 ;
      RECT 7.77 4.135 7.94 4.305 ;
      RECT 7.65 4.545 7.82 4.715 ;
      RECT 7.65 8.605 7.82 8.775 ;
      RECT 7.395 2.775 7.565 2.945 ;
      RECT 7.34 6.685 7.51 6.855 ;
      RECT 7.31 1.415 7.48 1.585 ;
      RECT 7.31 4.135 7.48 4.305 ;
      RECT 7.155 2.215 7.325 2.385 ;
      RECT 6.97 8.605 7.14 8.775 ;
      RECT 6.915 3.615 7.085 3.785 ;
      RECT 6.91 7.055 7.08 7.225 ;
      RECT 6.91 7.795 7.08 7.965 ;
      RECT 6.85 1.415 7.02 1.585 ;
      RECT 6.85 4.135 7.02 4.305 ;
      RECT 6.675 2.775 6.845 2.945 ;
      RECT 6.535 6.315 6.705 6.485 ;
      RECT 6.39 1.415 6.56 1.585 ;
      RECT 6.39 4.135 6.56 4.305 ;
      RECT 6.29 8.605 6.46 8.775 ;
      RECT 6.195 2.495 6.365 2.665 ;
      RECT 5.93 1.415 6.1 1.585 ;
      RECT 5.93 4.135 6.1 4.305 ;
      RECT 5.715 2.495 5.885 2.665 ;
      RECT 5.61 8.605 5.78 8.775 ;
      RECT 5.54 5.945 5.71 6.115 ;
      RECT 5.475 1.935 5.645 2.105 ;
      RECT 5.47 1.415 5.64 1.585 ;
      RECT 5.47 4.135 5.64 4.305 ;
      RECT 5.01 1.415 5.18 1.585 ;
      RECT 5.01 4.135 5.18 4.305 ;
      RECT 4.715 2.215 4.885 2.385 ;
      RECT 4.55 1.415 4.72 1.585 ;
      RECT 4.55 4.135 4.72 4.305 ;
      RECT 4.475 3.335 4.645 3.505 ;
      RECT 4.235 2.775 4.405 2.945 ;
      RECT 4.09 1.415 4.26 1.585 ;
      RECT 4.09 4.135 4.26 4.305 ;
      RECT 3.755 2.495 3.925 2.665 ;
      RECT 3.63 1.415 3.8 1.585 ;
      RECT 3.63 4.135 3.8 4.305 ;
      RECT 3.515 1.935 3.685 2.105 ;
      RECT 3.515 3.335 3.685 3.505 ;
      RECT 3.17 1.415 3.34 1.585 ;
      RECT 3.17 4.135 3.34 4.305 ;
      RECT 3.035 3.055 3.205 3.225 ;
      RECT 2.71 1.415 2.88 1.585 ;
      RECT 2.71 4.135 2.88 4.305 ;
      RECT 2.515 2.495 2.685 2.665 ;
      RECT 2.275 3.335 2.445 3.505 ;
      RECT 2.25 1.415 2.42 1.585 ;
      RECT 2.25 4.135 2.42 4.305 ;
      RECT 2.035 1.935 2.205 2.105 ;
      RECT 1.795 2.495 1.965 2.665 ;
      RECT 1.795 3.055 1.965 3.225 ;
      RECT 1.79 1.415 1.96 1.585 ;
      RECT 1.79 4.135 1.96 4.305 ;
      RECT 1.33 1.415 1.5 1.585 ;
      RECT 1.33 4.135 1.5 4.305 ;
      RECT 1.075 1.935 1.245 2.105 ;
      RECT 1.075 3.615 1.245 3.785 ;
      RECT 0.87 1.415 1.04 1.585 ;
      RECT 0.87 4.135 1.04 4.305 ;
      RECT 0.595 3.055 0.765 3.225 ;
      RECT 0.41 1.415 0.58 1.585 ;
      RECT 0.41 4.135 0.58 4.305 ;
      RECT -0.93 4.545 -0.76 4.715 ;
      RECT -0.93 8.605 -0.76 8.775 ;
      RECT -1.24 6.685 -1.07 6.855 ;
      RECT -1.61 8.605 -1.44 8.775 ;
      RECT -1.67 7.055 -1.5 7.225 ;
      RECT -1.67 7.795 -1.5 7.965 ;
      RECT -2.045 6.315 -1.875 6.485 ;
      RECT -2.29 8.605 -2.12 8.775 ;
      RECT -2.97 8.605 -2.8 8.775 ;
      RECT -3.04 5.945 -2.87 6.115 ;
    LAYER li ;
      RECT 73.695 0 73.865 2.085 ;
      RECT 71.735 0 71.905 2.085 ;
      RECT 69.295 0 69.465 2.085 ;
      RECT 68.335 0 68.505 2.085 ;
      RECT 67.815 0 67.985 2.085 ;
      RECT 66.855 0 67.025 2.085 ;
      RECT 65.895 0 66.065 2.085 ;
      RECT 57.37 0 57.54 2.085 ;
      RECT 55.41 0 55.58 2.085 ;
      RECT 52.97 0 53.14 2.085 ;
      RECT 52.01 0 52.18 2.085 ;
      RECT 51.49 0 51.66 2.085 ;
      RECT 50.53 0 50.7 2.085 ;
      RECT 49.57 0 49.74 2.085 ;
      RECT 41.045 0 41.215 2.085 ;
      RECT 39.085 0 39.255 2.085 ;
      RECT 36.645 0 36.815 2.085 ;
      RECT 35.685 0 35.855 2.085 ;
      RECT 35.165 0 35.335 2.085 ;
      RECT 34.205 0 34.375 2.085 ;
      RECT 33.245 0 33.415 2.085 ;
      RECT 24.72 0 24.89 2.085 ;
      RECT 22.76 0 22.93 2.085 ;
      RECT 20.32 0 20.49 2.085 ;
      RECT 19.36 0 19.53 2.085 ;
      RECT 18.84 0 19.01 2.085 ;
      RECT 17.88 0 18.05 2.085 ;
      RECT 16.92 0 17.09 2.085 ;
      RECT 8.395 0 8.565 2.085 ;
      RECT 6.435 0 6.605 2.085 ;
      RECT 3.995 0 4.165 2.085 ;
      RECT 3.035 0 3.205 2.085 ;
      RECT 2.515 0 2.685 2.085 ;
      RECT 1.555 0 1.725 2.085 ;
      RECT 0.595 0 0.765 2.085 ;
      RECT 71.665 0 71.905 1.595 ;
      RECT 70.115 0 70.31 1.595 ;
      RECT 67.99 0 68.185 1.595 ;
      RECT 65.69 0 65.885 1.595 ;
      RECT 55.34 0 55.58 1.595 ;
      RECT 53.79 0 53.985 1.595 ;
      RECT 51.665 0 51.86 1.595 ;
      RECT 49.365 0 49.56 1.595 ;
      RECT 39.015 0 39.255 1.595 ;
      RECT 37.465 0 37.66 1.595 ;
      RECT 35.34 0 35.535 1.595 ;
      RECT 33.04 0 33.235 1.595 ;
      RECT 22.69 0 22.93 1.595 ;
      RECT 21.14 0 21.335 1.595 ;
      RECT 19.015 0 19.21 1.595 ;
      RECT 16.715 0 16.91 1.595 ;
      RECT 6.365 0 6.605 1.595 ;
      RECT 4.815 0 5.01 1.595 ;
      RECT 2.69 0 2.885 1.595 ;
      RECT 0.39 0 0.585 1.595 ;
      RECT 65.565 0 75.38 1.585 ;
      RECT 49.24 0 59.055 1.585 ;
      RECT 32.915 0 42.73 1.585 ;
      RECT 16.59 0 26.405 1.585 ;
      RECT 0.265 0 10.08 1.585 ;
      RECT 80.18 0 80.35 0.935 ;
      RECT 79.19 0 79.36 0.935 ;
      RECT 76.445 0 76.615 0.935 ;
      RECT 63.855 0 64.025 0.935 ;
      RECT 62.865 0 63.035 0.935 ;
      RECT 60.12 0 60.29 0.935 ;
      RECT 47.53 0 47.7 0.935 ;
      RECT 46.54 0 46.71 0.935 ;
      RECT 43.795 0 43.965 0.935 ;
      RECT 31.205 0 31.375 0.935 ;
      RECT 30.215 0 30.385 0.935 ;
      RECT 27.47 0 27.64 0.935 ;
      RECT 14.88 0 15.05 0.935 ;
      RECT 13.89 0 14.06 0.935 ;
      RECT 11.145 0 11.315 0.935 ;
      RECT -3.225 0 81.15 0.305 ;
      RECT -1.24 4.135 -1.07 8.305 ;
      RECT 80.18 3.405 80.35 5.475 ;
      RECT 79.19 3.405 79.36 5.475 ;
      RECT 76.445 3.405 76.615 5.475 ;
      RECT 70.83 4.135 71 5.475 ;
      RECT 63.855 3.405 64.025 5.475 ;
      RECT 62.865 3.405 63.035 5.475 ;
      RECT 60.12 3.405 60.29 5.475 ;
      RECT 54.505 4.135 54.675 5.475 ;
      RECT 47.53 3.405 47.7 5.475 ;
      RECT 46.54 3.405 46.71 5.475 ;
      RECT 43.795 3.405 43.965 5.475 ;
      RECT 38.18 4.135 38.35 5.475 ;
      RECT 31.205 3.405 31.375 5.475 ;
      RECT 30.215 3.405 30.385 5.475 ;
      RECT 27.47 3.405 27.64 5.475 ;
      RECT 21.855 4.135 22.025 5.475 ;
      RECT 14.88 3.405 15.05 5.475 ;
      RECT 13.89 3.405 14.06 5.475 ;
      RECT 11.145 3.405 11.315 5.475 ;
      RECT 5.53 4.135 5.7 5.475 ;
      RECT -3.05 4.135 -2.88 5.475 ;
      RECT -3.225 4.135 81.15 4.745 ;
      RECT 74.655 3.635 74.825 4.745 ;
      RECT 73.695 3.635 73.865 4.745 ;
      RECT 71.255 3.635 71.425 4.745 ;
      RECT 70.255 3.635 70.425 4.745 ;
      RECT 69.295 3.635 69.465 4.745 ;
      RECT 66.855 3.635 67.025 4.745 ;
      RECT 58.33 3.635 58.5 4.745 ;
      RECT 57.37 3.635 57.54 4.745 ;
      RECT 54.93 3.635 55.1 4.745 ;
      RECT 53.93 3.635 54.1 4.745 ;
      RECT 52.97 3.635 53.14 4.745 ;
      RECT 50.53 3.635 50.7 4.745 ;
      RECT 42.005 3.635 42.175 4.745 ;
      RECT 41.045 3.635 41.215 4.745 ;
      RECT 38.605 3.635 38.775 4.745 ;
      RECT 37.605 3.635 37.775 4.745 ;
      RECT 36.645 3.635 36.815 4.745 ;
      RECT 34.205 3.635 34.375 4.745 ;
      RECT 25.68 3.635 25.85 4.745 ;
      RECT 24.72 3.635 24.89 4.745 ;
      RECT 22.28 3.635 22.45 4.745 ;
      RECT 21.28 3.635 21.45 4.745 ;
      RECT 20.32 3.635 20.49 4.745 ;
      RECT 17.88 3.635 18.05 4.745 ;
      RECT 9.355 3.635 9.525 4.745 ;
      RECT 8.395 3.635 8.565 4.745 ;
      RECT 5.955 3.635 6.125 4.745 ;
      RECT 4.955 3.635 5.125 4.745 ;
      RECT 3.995 3.635 4.165 4.745 ;
      RECT 1.555 3.635 1.725 4.745 ;
      RECT -3.23 8.575 81.15 8.88 ;
      RECT 80.18 7.945 80.35 8.88 ;
      RECT 79.19 7.945 79.36 8.88 ;
      RECT 76.445 7.945 76.615 8.88 ;
      RECT 70.83 7.945 71 8.88 ;
      RECT 63.855 7.945 64.025 8.88 ;
      RECT 62.865 7.945 63.035 8.88 ;
      RECT 60.12 7.945 60.29 8.88 ;
      RECT 54.505 7.945 54.675 8.88 ;
      RECT 47.53 7.945 47.7 8.88 ;
      RECT 46.54 7.945 46.71 8.88 ;
      RECT 43.795 7.945 43.965 8.88 ;
      RECT 38.18 7.945 38.35 8.88 ;
      RECT 31.205 7.945 31.375 8.88 ;
      RECT 30.215 7.945 30.385 8.88 ;
      RECT 27.47 7.945 27.64 8.88 ;
      RECT 21.855 7.945 22.025 8.88 ;
      RECT 14.88 7.945 15.05 8.88 ;
      RECT 13.89 7.945 14.06 8.88 ;
      RECT 11.145 7.945 11.315 8.88 ;
      RECT 5.53 7.945 5.7 8.88 ;
      RECT -3.05 7.945 -2.88 8.88 ;
      RECT 80.24 1.74 80.41 2.935 ;
      RECT 80.24 1.74 80.705 1.91 ;
      RECT 80.24 6.97 80.705 7.14 ;
      RECT 80.24 5.945 80.41 7.14 ;
      RECT 79.25 1.74 79.42 2.935 ;
      RECT 79.25 1.74 79.715 1.91 ;
      RECT 79.25 6.97 79.715 7.14 ;
      RECT 79.25 5.945 79.42 7.14 ;
      RECT 77.395 2.635 77.565 3.865 ;
      RECT 77.45 0.855 77.62 2.805 ;
      RECT 77.395 0.575 77.565 1.025 ;
      RECT 77.395 7.855 77.565 8.305 ;
      RECT 77.45 6.075 77.62 8.025 ;
      RECT 77.395 5.015 77.565 6.245 ;
      RECT 76.875 0.575 77.045 3.865 ;
      RECT 76.875 2.075 77.28 2.405 ;
      RECT 76.875 1.235 77.28 1.565 ;
      RECT 76.875 5.015 77.045 8.305 ;
      RECT 76.875 7.315 77.28 7.645 ;
      RECT 76.875 6.475 77.28 6.805 ;
      RECT 74.175 1.835 74.345 2.105 ;
      RECT 74.175 1.835 74.905 2.005 ;
      RECT 74.655 2.575 74.825 2.945 ;
      RECT 74.335 2.575 74.825 2.745 ;
      RECT 74.095 3.225 74.425 3.395 ;
      RECT 73.335 3.055 74.345 3.225 ;
      RECT 73.335 2.575 73.505 3.225 ;
      RECT 73.455 2.495 73.625 2.825 ;
      RECT 72.615 3.225 72.945 3.395 ;
      RECT 70.695 3.225 71.985 3.395 ;
      RECT 71.735 3.14 72.865 3.31 ;
      RECT 72.455 2.215 72.865 2.385 ;
      RECT 72.695 1.755 72.865 2.385 ;
      RECT 72.695 2.575 72.865 2.945 ;
      RECT 72.375 2.575 72.865 2.745 ;
      RECT 71.78 7.855 71.95 8.305 ;
      RECT 71.835 6.075 72.005 8.025 ;
      RECT 71.78 5.015 71.95 6.245 ;
      RECT 71.26 5.015 71.43 8.305 ;
      RECT 71.26 7.315 71.665 7.645 ;
      RECT 71.26 6.475 71.665 6.805 ;
      RECT 69.935 2.575 71.265 2.745 ;
      RECT 71.015 2.495 71.185 2.745 ;
      RECT 70.015 2.175 70.185 2.385 ;
      RECT 70.015 2.175 70.505 2.345 ;
      RECT 68.695 3.335 68.985 3.505 ;
      RECT 68.695 2.575 68.865 3.505 ;
      RECT 68.495 2.575 68.865 2.745 ;
      RECT 67.495 2.575 67.985 2.745 ;
      RECT 67.815 2.495 67.985 2.745 ;
      RECT 67.575 3.335 67.985 3.505 ;
      RECT 67.815 3.145 67.985 3.505 ;
      RECT 66.615 3.055 67.265 3.225 ;
      RECT 66.615 2.495 66.785 3.225 ;
      RECT 66.255 3.615 66.545 3.785 ;
      RECT 66.255 2.575 66.425 3.785 ;
      RECT 66.055 2.575 66.425 2.745 ;
      RECT 63.915 1.74 64.085 2.935 ;
      RECT 63.915 1.74 64.38 1.91 ;
      RECT 63.915 6.97 64.38 7.14 ;
      RECT 63.915 5.945 64.085 7.14 ;
      RECT 62.925 1.74 63.095 2.935 ;
      RECT 62.925 1.74 63.39 1.91 ;
      RECT 62.925 6.97 63.39 7.14 ;
      RECT 62.925 5.945 63.095 7.14 ;
      RECT 61.07 2.635 61.24 3.865 ;
      RECT 61.125 0.855 61.295 2.805 ;
      RECT 61.07 0.575 61.24 1.025 ;
      RECT 61.07 7.855 61.24 8.305 ;
      RECT 61.125 6.075 61.295 8.025 ;
      RECT 61.07 5.015 61.24 6.245 ;
      RECT 60.55 0.575 60.72 3.865 ;
      RECT 60.55 2.075 60.955 2.405 ;
      RECT 60.55 1.235 60.955 1.565 ;
      RECT 60.55 5.015 60.72 8.305 ;
      RECT 60.55 7.315 60.955 7.645 ;
      RECT 60.55 6.475 60.955 6.805 ;
      RECT 57.85 1.835 58.02 2.105 ;
      RECT 57.85 1.835 58.58 2.005 ;
      RECT 58.33 2.575 58.5 2.945 ;
      RECT 58.01 2.575 58.5 2.745 ;
      RECT 57.77 3.225 58.1 3.395 ;
      RECT 57.01 3.055 58.02 3.225 ;
      RECT 57.01 2.575 57.18 3.225 ;
      RECT 57.13 2.495 57.3 2.825 ;
      RECT 56.29 3.225 56.62 3.395 ;
      RECT 54.37 3.225 55.66 3.395 ;
      RECT 55.41 3.14 56.54 3.31 ;
      RECT 56.13 2.215 56.54 2.385 ;
      RECT 56.37 1.755 56.54 2.385 ;
      RECT 56.37 2.575 56.54 2.945 ;
      RECT 56.05 2.575 56.54 2.745 ;
      RECT 55.455 7.855 55.625 8.305 ;
      RECT 55.51 6.075 55.68 8.025 ;
      RECT 55.455 5.015 55.625 6.245 ;
      RECT 54.935 5.015 55.105 8.305 ;
      RECT 54.935 7.315 55.34 7.645 ;
      RECT 54.935 6.475 55.34 6.805 ;
      RECT 53.61 2.575 54.94 2.745 ;
      RECT 54.69 2.495 54.86 2.745 ;
      RECT 53.69 2.175 53.86 2.385 ;
      RECT 53.69 2.175 54.18 2.345 ;
      RECT 52.37 3.335 52.66 3.505 ;
      RECT 52.37 2.575 52.54 3.505 ;
      RECT 52.17 2.575 52.54 2.745 ;
      RECT 51.17 2.575 51.66 2.745 ;
      RECT 51.49 2.495 51.66 2.745 ;
      RECT 51.25 3.335 51.66 3.505 ;
      RECT 51.49 3.145 51.66 3.505 ;
      RECT 50.29 3.055 50.94 3.225 ;
      RECT 50.29 2.495 50.46 3.225 ;
      RECT 49.93 3.615 50.22 3.785 ;
      RECT 49.93 2.575 50.1 3.785 ;
      RECT 49.73 2.575 50.1 2.745 ;
      RECT 47.59 1.74 47.76 2.935 ;
      RECT 47.59 1.74 48.055 1.91 ;
      RECT 47.59 6.97 48.055 7.14 ;
      RECT 47.59 5.945 47.76 7.14 ;
      RECT 46.6 1.74 46.77 2.935 ;
      RECT 46.6 1.74 47.065 1.91 ;
      RECT 46.6 6.97 47.065 7.14 ;
      RECT 46.6 5.945 46.77 7.14 ;
      RECT 44.745 2.635 44.915 3.865 ;
      RECT 44.8 0.855 44.97 2.805 ;
      RECT 44.745 0.575 44.915 1.025 ;
      RECT 44.745 7.855 44.915 8.305 ;
      RECT 44.8 6.075 44.97 8.025 ;
      RECT 44.745 5.015 44.915 6.245 ;
      RECT 44.225 0.575 44.395 3.865 ;
      RECT 44.225 2.075 44.63 2.405 ;
      RECT 44.225 1.235 44.63 1.565 ;
      RECT 44.225 5.015 44.395 8.305 ;
      RECT 44.225 7.315 44.63 7.645 ;
      RECT 44.225 6.475 44.63 6.805 ;
      RECT 41.525 1.835 41.695 2.105 ;
      RECT 41.525 1.835 42.255 2.005 ;
      RECT 42.005 2.575 42.175 2.945 ;
      RECT 41.685 2.575 42.175 2.745 ;
      RECT 41.445 3.225 41.775 3.395 ;
      RECT 40.685 3.055 41.695 3.225 ;
      RECT 40.685 2.575 40.855 3.225 ;
      RECT 40.805 2.495 40.975 2.825 ;
      RECT 39.965 3.225 40.295 3.395 ;
      RECT 38.045 3.225 39.335 3.395 ;
      RECT 39.085 3.14 40.215 3.31 ;
      RECT 39.805 2.215 40.215 2.385 ;
      RECT 40.045 1.755 40.215 2.385 ;
      RECT 40.045 2.575 40.215 2.945 ;
      RECT 39.725 2.575 40.215 2.745 ;
      RECT 39.13 7.855 39.3 8.305 ;
      RECT 39.185 6.075 39.355 8.025 ;
      RECT 39.13 5.015 39.3 6.245 ;
      RECT 38.61 5.015 38.78 8.305 ;
      RECT 38.61 7.315 39.015 7.645 ;
      RECT 38.61 6.475 39.015 6.805 ;
      RECT 37.285 2.575 38.615 2.745 ;
      RECT 38.365 2.495 38.535 2.745 ;
      RECT 37.365 2.175 37.535 2.385 ;
      RECT 37.365 2.175 37.855 2.345 ;
      RECT 36.045 3.335 36.335 3.505 ;
      RECT 36.045 2.575 36.215 3.505 ;
      RECT 35.845 2.575 36.215 2.745 ;
      RECT 34.845 2.575 35.335 2.745 ;
      RECT 35.165 2.495 35.335 2.745 ;
      RECT 34.925 3.335 35.335 3.505 ;
      RECT 35.165 3.145 35.335 3.505 ;
      RECT 33.965 3.055 34.615 3.225 ;
      RECT 33.965 2.495 34.135 3.225 ;
      RECT 33.605 3.615 33.895 3.785 ;
      RECT 33.605 2.575 33.775 3.785 ;
      RECT 33.405 2.575 33.775 2.745 ;
      RECT 31.265 1.74 31.435 2.935 ;
      RECT 31.265 1.74 31.73 1.91 ;
      RECT 31.265 6.97 31.73 7.14 ;
      RECT 31.265 5.945 31.435 7.14 ;
      RECT 30.275 1.74 30.445 2.935 ;
      RECT 30.275 1.74 30.74 1.91 ;
      RECT 30.275 6.97 30.74 7.14 ;
      RECT 30.275 5.945 30.445 7.14 ;
      RECT 28.42 2.635 28.59 3.865 ;
      RECT 28.475 0.855 28.645 2.805 ;
      RECT 28.42 0.575 28.59 1.025 ;
      RECT 28.42 7.855 28.59 8.305 ;
      RECT 28.475 6.075 28.645 8.025 ;
      RECT 28.42 5.015 28.59 6.245 ;
      RECT 27.9 0.575 28.07 3.865 ;
      RECT 27.9 2.075 28.305 2.405 ;
      RECT 27.9 1.235 28.305 1.565 ;
      RECT 27.9 5.015 28.07 8.305 ;
      RECT 27.9 7.315 28.305 7.645 ;
      RECT 27.9 6.475 28.305 6.805 ;
      RECT 25.2 1.835 25.37 2.105 ;
      RECT 25.2 1.835 25.93 2.005 ;
      RECT 25.68 2.575 25.85 2.945 ;
      RECT 25.36 2.575 25.85 2.745 ;
      RECT 25.12 3.225 25.45 3.395 ;
      RECT 24.36 3.055 25.37 3.225 ;
      RECT 24.36 2.575 24.53 3.225 ;
      RECT 24.48 2.495 24.65 2.825 ;
      RECT 23.64 3.225 23.97 3.395 ;
      RECT 21.72 3.225 23.01 3.395 ;
      RECT 22.76 3.14 23.89 3.31 ;
      RECT 23.48 2.215 23.89 2.385 ;
      RECT 23.72 1.755 23.89 2.385 ;
      RECT 23.72 2.575 23.89 2.945 ;
      RECT 23.4 2.575 23.89 2.745 ;
      RECT 22.805 7.855 22.975 8.305 ;
      RECT 22.86 6.075 23.03 8.025 ;
      RECT 22.805 5.015 22.975 6.245 ;
      RECT 22.285 5.015 22.455 8.305 ;
      RECT 22.285 7.315 22.69 7.645 ;
      RECT 22.285 6.475 22.69 6.805 ;
      RECT 20.96 2.575 22.29 2.745 ;
      RECT 22.04 2.495 22.21 2.745 ;
      RECT 21.04 2.175 21.21 2.385 ;
      RECT 21.04 2.175 21.53 2.345 ;
      RECT 19.72 3.335 20.01 3.505 ;
      RECT 19.72 2.575 19.89 3.505 ;
      RECT 19.52 2.575 19.89 2.745 ;
      RECT 18.52 2.575 19.01 2.745 ;
      RECT 18.84 2.495 19.01 2.745 ;
      RECT 18.6 3.335 19.01 3.505 ;
      RECT 18.84 3.145 19.01 3.505 ;
      RECT 17.64 3.055 18.29 3.225 ;
      RECT 17.64 2.495 17.81 3.225 ;
      RECT 17.28 3.615 17.57 3.785 ;
      RECT 17.28 2.575 17.45 3.785 ;
      RECT 17.08 2.575 17.45 2.745 ;
      RECT 14.94 1.74 15.11 2.935 ;
      RECT 14.94 1.74 15.405 1.91 ;
      RECT 14.94 6.97 15.405 7.14 ;
      RECT 14.94 5.945 15.11 7.14 ;
      RECT 13.95 1.74 14.12 2.935 ;
      RECT 13.95 1.74 14.415 1.91 ;
      RECT 13.95 6.97 14.415 7.14 ;
      RECT 13.95 5.945 14.12 7.14 ;
      RECT 12.095 2.635 12.265 3.865 ;
      RECT 12.15 0.855 12.32 2.805 ;
      RECT 12.095 0.575 12.265 1.025 ;
      RECT 12.095 7.855 12.265 8.305 ;
      RECT 12.15 6.075 12.32 8.025 ;
      RECT 12.095 5.015 12.265 6.245 ;
      RECT 11.575 0.575 11.745 3.865 ;
      RECT 11.575 2.075 11.98 2.405 ;
      RECT 11.575 1.235 11.98 1.565 ;
      RECT 11.575 5.015 11.745 8.305 ;
      RECT 11.575 7.315 11.98 7.645 ;
      RECT 11.575 6.475 11.98 6.805 ;
      RECT 8.875 1.835 9.045 2.105 ;
      RECT 8.875 1.835 9.605 2.005 ;
      RECT 9.355 2.575 9.525 2.945 ;
      RECT 9.035 2.575 9.525 2.745 ;
      RECT 8.795 3.225 9.125 3.395 ;
      RECT 8.035 3.055 9.045 3.225 ;
      RECT 8.035 2.575 8.205 3.225 ;
      RECT 8.155 2.495 8.325 2.825 ;
      RECT 7.315 3.225 7.645 3.395 ;
      RECT 5.395 3.225 6.685 3.395 ;
      RECT 6.435 3.14 7.565 3.31 ;
      RECT 7.155 2.215 7.565 2.385 ;
      RECT 7.395 1.755 7.565 2.385 ;
      RECT 7.395 2.575 7.565 2.945 ;
      RECT 7.075 2.575 7.565 2.745 ;
      RECT 6.48 7.855 6.65 8.305 ;
      RECT 6.535 6.075 6.705 8.025 ;
      RECT 6.48 5.015 6.65 6.245 ;
      RECT 5.96 5.015 6.13 8.305 ;
      RECT 5.96 7.315 6.365 7.645 ;
      RECT 5.96 6.475 6.365 6.805 ;
      RECT 4.635 2.575 5.965 2.745 ;
      RECT 5.715 2.495 5.885 2.745 ;
      RECT 4.715 2.175 4.885 2.385 ;
      RECT 4.715 2.175 5.205 2.345 ;
      RECT 3.395 3.335 3.685 3.505 ;
      RECT 3.395 2.575 3.565 3.505 ;
      RECT 3.195 2.575 3.565 2.745 ;
      RECT 2.195 2.575 2.685 2.745 ;
      RECT 2.515 2.495 2.685 2.745 ;
      RECT 2.275 3.335 2.685 3.505 ;
      RECT 2.515 3.145 2.685 3.505 ;
      RECT 1.315 3.055 1.965 3.225 ;
      RECT 1.315 2.495 1.485 3.225 ;
      RECT 0.955 3.615 1.245 3.785 ;
      RECT 0.955 2.575 1.125 3.785 ;
      RECT 0.755 2.575 1.125 2.745 ;
      RECT -2.1 7.855 -1.93 8.305 ;
      RECT -2.045 6.075 -1.875 8.025 ;
      RECT -2.1 5.015 -1.93 6.245 ;
      RECT -2.62 5.015 -2.45 8.305 ;
      RECT -2.62 7.315 -2.215 7.645 ;
      RECT -2.62 6.475 -2.215 6.805 ;
      RECT 80.61 0.575 80.78 1.085 ;
      RECT 80.61 2.395 80.78 3.865 ;
      RECT 80.61 5.015 80.78 6.485 ;
      RECT 80.61 7.795 80.78 8.305 ;
      RECT 79.62 0.575 79.79 1.085 ;
      RECT 79.62 2.395 79.79 3.865 ;
      RECT 79.62 5.015 79.79 6.485 ;
      RECT 79.62 7.795 79.79 8.305 ;
      RECT 78.255 0.575 78.425 3.865 ;
      RECT 78.255 5.015 78.425 8.305 ;
      RECT 77.825 0.575 77.995 1.085 ;
      RECT 77.825 1.655 77.995 3.865 ;
      RECT 77.825 5.015 77.995 7.225 ;
      RECT 77.825 7.795 77.995 8.305 ;
      RECT 76.455 1.66 76.625 2.935 ;
      RECT 76.455 5.945 76.625 7.22 ;
      RECT 73.935 2.495 74.105 2.825 ;
      RECT 73.215 1.755 73.385 2.105 ;
      RECT 73.215 3.485 73.385 3.815 ;
      RECT 72.64 5.015 72.81 8.305 ;
      RECT 72.215 3.485 72.385 3.815 ;
      RECT 72.21 5.015 72.38 7.225 ;
      RECT 72.21 7.795 72.38 8.305 ;
      RECT 71.975 2.495 72.145 2.945 ;
      RECT 71.495 2.495 71.665 2.825 ;
      RECT 70.84 5.945 71.01 7.22 ;
      RECT 70.775 1.755 70.945 2.105 ;
      RECT 69.775 3.145 69.945 3.505 ;
      RECT 69.535 2.495 69.705 2.945 ;
      RECT 69.055 2.495 69.225 2.825 ;
      RECT 68.815 1.755 68.985 2.105 ;
      RECT 68.335 3.055 68.505 3.475 ;
      RECT 67.335 1.755 67.505 2.105 ;
      RECT 67.095 2.495 67.265 2.825 ;
      RECT 66.375 1.755 66.545 2.105 ;
      RECT 65.895 3.055 66.065 3.475 ;
      RECT 64.285 0.575 64.455 1.085 ;
      RECT 64.285 2.395 64.455 3.865 ;
      RECT 64.285 5.015 64.455 6.485 ;
      RECT 64.285 7.795 64.455 8.305 ;
      RECT 63.295 0.575 63.465 1.085 ;
      RECT 63.295 2.395 63.465 3.865 ;
      RECT 63.295 5.015 63.465 6.485 ;
      RECT 63.295 7.795 63.465 8.305 ;
      RECT 61.93 0.575 62.1 3.865 ;
      RECT 61.93 5.015 62.1 8.305 ;
      RECT 61.5 0.575 61.67 1.085 ;
      RECT 61.5 1.655 61.67 3.865 ;
      RECT 61.5 5.015 61.67 7.225 ;
      RECT 61.5 7.795 61.67 8.305 ;
      RECT 60.13 1.66 60.3 2.935 ;
      RECT 60.13 5.945 60.3 7.22 ;
      RECT 57.61 2.495 57.78 2.825 ;
      RECT 56.89 1.755 57.06 2.105 ;
      RECT 56.89 3.485 57.06 3.815 ;
      RECT 56.315 5.015 56.485 8.305 ;
      RECT 55.89 3.485 56.06 3.815 ;
      RECT 55.885 5.015 56.055 7.225 ;
      RECT 55.885 7.795 56.055 8.305 ;
      RECT 55.65 2.495 55.82 2.945 ;
      RECT 55.17 2.495 55.34 2.825 ;
      RECT 54.515 5.945 54.685 7.22 ;
      RECT 54.45 1.755 54.62 2.105 ;
      RECT 53.45 3.145 53.62 3.505 ;
      RECT 53.21 2.495 53.38 2.945 ;
      RECT 52.73 2.495 52.9 2.825 ;
      RECT 52.49 1.755 52.66 2.105 ;
      RECT 52.01 3.055 52.18 3.475 ;
      RECT 51.01 1.755 51.18 2.105 ;
      RECT 50.77 2.495 50.94 2.825 ;
      RECT 50.05 1.755 50.22 2.105 ;
      RECT 49.57 3.055 49.74 3.475 ;
      RECT 47.96 0.575 48.13 1.085 ;
      RECT 47.96 2.395 48.13 3.865 ;
      RECT 47.96 5.015 48.13 6.485 ;
      RECT 47.96 7.795 48.13 8.305 ;
      RECT 46.97 0.575 47.14 1.085 ;
      RECT 46.97 2.395 47.14 3.865 ;
      RECT 46.97 5.015 47.14 6.485 ;
      RECT 46.97 7.795 47.14 8.305 ;
      RECT 45.605 0.575 45.775 3.865 ;
      RECT 45.605 5.015 45.775 8.305 ;
      RECT 45.175 0.575 45.345 1.085 ;
      RECT 45.175 1.655 45.345 3.865 ;
      RECT 45.175 5.015 45.345 7.225 ;
      RECT 45.175 7.795 45.345 8.305 ;
      RECT 43.805 1.66 43.975 2.935 ;
      RECT 43.805 5.945 43.975 7.22 ;
      RECT 41.285 2.495 41.455 2.825 ;
      RECT 40.565 1.755 40.735 2.105 ;
      RECT 40.565 3.485 40.735 3.815 ;
      RECT 39.99 5.015 40.16 8.305 ;
      RECT 39.565 3.485 39.735 3.815 ;
      RECT 39.56 5.015 39.73 7.225 ;
      RECT 39.56 7.795 39.73 8.305 ;
      RECT 39.325 2.495 39.495 2.945 ;
      RECT 38.845 2.495 39.015 2.825 ;
      RECT 38.19 5.945 38.36 7.22 ;
      RECT 38.125 1.755 38.295 2.105 ;
      RECT 37.125 3.145 37.295 3.505 ;
      RECT 36.885 2.495 37.055 2.945 ;
      RECT 36.405 2.495 36.575 2.825 ;
      RECT 36.165 1.755 36.335 2.105 ;
      RECT 35.685 3.055 35.855 3.475 ;
      RECT 34.685 1.755 34.855 2.105 ;
      RECT 34.445 2.495 34.615 2.825 ;
      RECT 33.725 1.755 33.895 2.105 ;
      RECT 33.245 3.055 33.415 3.475 ;
      RECT 31.635 0.575 31.805 1.085 ;
      RECT 31.635 2.395 31.805 3.865 ;
      RECT 31.635 5.015 31.805 6.485 ;
      RECT 31.635 7.795 31.805 8.305 ;
      RECT 30.645 0.575 30.815 1.085 ;
      RECT 30.645 2.395 30.815 3.865 ;
      RECT 30.645 5.015 30.815 6.485 ;
      RECT 30.645 7.795 30.815 8.305 ;
      RECT 29.28 0.575 29.45 3.865 ;
      RECT 29.28 5.015 29.45 8.305 ;
      RECT 28.85 0.575 29.02 1.085 ;
      RECT 28.85 1.655 29.02 3.865 ;
      RECT 28.85 5.015 29.02 7.225 ;
      RECT 28.85 7.795 29.02 8.305 ;
      RECT 27.48 1.66 27.65 2.935 ;
      RECT 27.48 5.945 27.65 7.22 ;
      RECT 24.96 2.495 25.13 2.825 ;
      RECT 24.24 1.755 24.41 2.105 ;
      RECT 24.24 3.485 24.41 3.815 ;
      RECT 23.665 5.015 23.835 8.305 ;
      RECT 23.24 3.485 23.41 3.815 ;
      RECT 23.235 5.015 23.405 7.225 ;
      RECT 23.235 7.795 23.405 8.305 ;
      RECT 23 2.495 23.17 2.945 ;
      RECT 22.52 2.495 22.69 2.825 ;
      RECT 21.865 5.945 22.035 7.22 ;
      RECT 21.8 1.755 21.97 2.105 ;
      RECT 20.8 3.145 20.97 3.505 ;
      RECT 20.56 2.495 20.73 2.945 ;
      RECT 20.08 2.495 20.25 2.825 ;
      RECT 19.84 1.755 20.01 2.105 ;
      RECT 19.36 3.055 19.53 3.475 ;
      RECT 18.36 1.755 18.53 2.105 ;
      RECT 18.12 2.495 18.29 2.825 ;
      RECT 17.4 1.755 17.57 2.105 ;
      RECT 16.92 3.055 17.09 3.475 ;
      RECT 15.31 0.575 15.48 1.085 ;
      RECT 15.31 2.395 15.48 3.865 ;
      RECT 15.31 5.015 15.48 6.485 ;
      RECT 15.31 7.795 15.48 8.305 ;
      RECT 14.32 0.575 14.49 1.085 ;
      RECT 14.32 2.395 14.49 3.865 ;
      RECT 14.32 5.015 14.49 6.485 ;
      RECT 14.32 7.795 14.49 8.305 ;
      RECT 12.955 0.575 13.125 3.865 ;
      RECT 12.955 5.015 13.125 8.305 ;
      RECT 12.525 0.575 12.695 1.085 ;
      RECT 12.525 1.655 12.695 3.865 ;
      RECT 12.525 5.015 12.695 7.225 ;
      RECT 12.525 7.795 12.695 8.305 ;
      RECT 11.155 1.66 11.325 2.935 ;
      RECT 11.155 5.945 11.325 7.22 ;
      RECT 8.635 2.495 8.805 2.825 ;
      RECT 7.915 1.755 8.085 2.105 ;
      RECT 7.915 3.485 8.085 3.815 ;
      RECT 7.34 5.015 7.51 8.305 ;
      RECT 6.915 3.485 7.085 3.815 ;
      RECT 6.91 5.015 7.08 7.225 ;
      RECT 6.91 7.795 7.08 8.305 ;
      RECT 6.675 2.495 6.845 2.945 ;
      RECT 6.195 2.495 6.365 2.825 ;
      RECT 5.54 5.945 5.71 7.22 ;
      RECT 5.475 1.755 5.645 2.105 ;
      RECT 4.475 3.145 4.645 3.505 ;
      RECT 4.235 2.495 4.405 2.945 ;
      RECT 3.755 2.495 3.925 2.825 ;
      RECT 3.515 1.755 3.685 2.105 ;
      RECT 3.035 3.055 3.205 3.475 ;
      RECT 2.035 1.755 2.205 2.105 ;
      RECT 1.795 2.495 1.965 2.825 ;
      RECT 1.075 1.755 1.245 2.105 ;
      RECT 0.595 3.055 0.765 3.475 ;
      RECT -1.67 5.015 -1.5 7.225 ;
      RECT -1.67 7.795 -1.5 8.305 ;
      RECT -3.04 5.945 -2.87 7.22 ;
  END
END sky130_osu_ring_oscillator_mpr2ea_8_b0r2

MACRO sky130_osu_ring_oscillator_mpr2et_8_b0r1
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 5.505 0 ;
  SIZE 95.595 BY 8.88 ;
  SYMMETRY X Y R90 ;
  SITE CoreSite ;
  OBS
    LAYER met3 ;
      RECT 81.58 3.535 82.135 3.865 ;
      RECT 81.58 1.87 81.88 3.865 ;
      RECT 77.645 2.975 78.2 3.305 ;
      RECT 77.9 1.87 78.2 3.305 ;
      RECT 77.9 1.87 81.88 2.17 ;
      RECT 81.05 7.055 81.425 7.425 ;
      RECT 81.05 7.095 82.055 7.395 ;
      RECT 81.755 4.405 82.055 7.395 ;
      RECT 71.925 4.405 82.055 4.705 ;
      RECT 76.43 2.415 76.73 4.705 ;
      RECT 74.995 2.975 75.295 4.705 ;
      RECT 71.925 2.42 72.225 4.705 ;
      RECT 74.965 2.975 75.695 3.305 ;
      RECT 76.405 2.415 77.135 2.745 ;
      RECT 72.855 2.415 73.585 2.745 ;
      RECT 71.925 2.42 73.585 2.72 ;
      RECT 63.02 3.535 63.575 3.865 ;
      RECT 63.02 1.87 63.32 3.865 ;
      RECT 59.085 2.975 59.64 3.305 ;
      RECT 59.34 1.87 59.64 3.305 ;
      RECT 59.34 1.87 63.32 2.17 ;
      RECT 62.49 7.055 62.865 7.425 ;
      RECT 62.49 7.095 63.495 7.395 ;
      RECT 63.195 4.405 63.495 7.395 ;
      RECT 53.365 4.405 63.495 4.705 ;
      RECT 57.87 2.415 58.17 4.705 ;
      RECT 56.435 2.975 56.735 4.705 ;
      RECT 53.365 2.42 53.665 4.705 ;
      RECT 56.405 2.975 57.135 3.305 ;
      RECT 57.845 2.415 58.575 2.745 ;
      RECT 54.295 2.415 55.025 2.745 ;
      RECT 53.365 2.42 55.025 2.72 ;
      RECT 44.46 3.535 45.015 3.865 ;
      RECT 44.46 1.87 44.76 3.865 ;
      RECT 40.525 2.975 41.08 3.305 ;
      RECT 40.78 1.87 41.08 3.305 ;
      RECT 40.78 1.87 44.76 2.17 ;
      RECT 43.93 7.055 44.305 7.425 ;
      RECT 43.93 7.095 44.935 7.395 ;
      RECT 44.635 4.405 44.935 7.395 ;
      RECT 34.805 4.405 44.935 4.705 ;
      RECT 39.31 2.415 39.61 4.705 ;
      RECT 37.875 2.975 38.175 4.705 ;
      RECT 34.805 2.42 35.105 4.705 ;
      RECT 37.845 2.975 38.575 3.305 ;
      RECT 39.285 2.415 40.015 2.745 ;
      RECT 35.735 2.415 36.465 2.745 ;
      RECT 34.805 2.42 36.465 2.72 ;
      RECT 25.9 3.535 26.455 3.865 ;
      RECT 25.9 1.87 26.2 3.865 ;
      RECT 21.965 2.975 22.52 3.305 ;
      RECT 22.22 1.87 22.52 3.305 ;
      RECT 22.22 1.87 26.2 2.17 ;
      RECT 25.37 7.055 25.745 7.425 ;
      RECT 25.37 7.095 26.375 7.395 ;
      RECT 26.075 4.405 26.375 7.395 ;
      RECT 16.245 4.405 26.375 4.705 ;
      RECT 20.75 2.415 21.05 4.705 ;
      RECT 19.315 2.975 19.615 4.705 ;
      RECT 16.245 2.42 16.545 4.705 ;
      RECT 19.285 2.975 20.015 3.305 ;
      RECT 20.725 2.415 21.455 2.745 ;
      RECT 17.175 2.415 17.905 2.745 ;
      RECT 16.245 2.42 17.905 2.72 ;
      RECT 7.34 3.535 7.895 3.865 ;
      RECT 7.34 1.87 7.64 3.865 ;
      RECT 3.405 2.975 3.96 3.305 ;
      RECT 3.66 1.87 3.96 3.305 ;
      RECT 3.66 1.87 7.64 2.17 ;
      RECT 6.81 7.055 7.185 7.425 ;
      RECT 6.81 7.095 7.815 7.395 ;
      RECT 7.515 4.405 7.815 7.395 ;
      RECT -5.46 4.145 -0.245 4.75 ;
      RECT -5.46 4.405 7.815 4.705 ;
      RECT 2.19 2.415 2.49 4.705 ;
      RECT 0.755 2.975 1.055 4.705 ;
      RECT -2.315 2.42 -2.015 4.75 ;
      RECT 0.725 2.975 1.455 3.305 ;
      RECT 2.165 2.415 2.895 2.745 ;
      RECT -1.385 2.415 -0.655 2.745 ;
      RECT -2.315 2.42 -0.655 2.72 ;
      RECT 82.765 1.855 83.495 2.185 ;
      RECT 80.545 3.535 81.275 3.865 ;
      RECT 78.845 3.535 79.575 3.865 ;
      RECT 73.89 2.415 74.62 2.745 ;
      RECT 72.525 3.535 73.255 3.865 ;
      RECT 64.205 1.855 64.935 2.185 ;
      RECT 61.985 3.535 62.715 3.865 ;
      RECT 60.285 3.535 61.015 3.865 ;
      RECT 55.33 2.415 56.06 2.745 ;
      RECT 53.965 3.535 54.695 3.865 ;
      RECT 45.645 1.855 46.375 2.185 ;
      RECT 43.425 3.535 44.155 3.865 ;
      RECT 41.725 3.535 42.455 3.865 ;
      RECT 36.77 2.415 37.5 2.745 ;
      RECT 35.405 3.535 36.135 3.865 ;
      RECT 27.085 1.855 27.815 2.185 ;
      RECT 24.865 3.535 25.595 3.865 ;
      RECT 23.165 3.535 23.895 3.865 ;
      RECT 18.21 2.415 18.94 2.745 ;
      RECT 16.845 3.535 17.575 3.865 ;
      RECT 8.525 1.855 9.255 2.185 ;
      RECT 6.305 3.535 7.035 3.865 ;
      RECT 4.605 3.535 5.335 3.865 ;
      RECT -0.35 2.415 0.38 2.745 ;
      RECT -1.715 3.535 -0.985 3.865 ;
    LAYER via2 ;
      RECT 82.83 1.92 83.03 2.12 ;
      RECT 81.87 3.6 82.07 3.8 ;
      RECT 81.135 7.14 81.335 7.34 ;
      RECT 80.87 3.6 81.07 3.8 ;
      RECT 78.91 3.6 79.11 3.8 ;
      RECT 77.71 3.04 77.91 3.24 ;
      RECT 76.47 2.48 76.67 2.68 ;
      RECT 75.03 3.04 75.23 3.24 ;
      RECT 74.29 2.48 74.49 2.68 ;
      RECT 73.07 2.48 73.27 2.68 ;
      RECT 72.59 3.6 72.79 3.8 ;
      RECT 64.27 1.92 64.47 2.12 ;
      RECT 63.31 3.6 63.51 3.8 ;
      RECT 62.575 7.14 62.775 7.34 ;
      RECT 62.31 3.6 62.51 3.8 ;
      RECT 60.35 3.6 60.55 3.8 ;
      RECT 59.15 3.04 59.35 3.24 ;
      RECT 57.91 2.48 58.11 2.68 ;
      RECT 56.47 3.04 56.67 3.24 ;
      RECT 55.73 2.48 55.93 2.68 ;
      RECT 54.51 2.48 54.71 2.68 ;
      RECT 54.03 3.6 54.23 3.8 ;
      RECT 45.71 1.92 45.91 2.12 ;
      RECT 44.75 3.6 44.95 3.8 ;
      RECT 44.015 7.14 44.215 7.34 ;
      RECT 43.75 3.6 43.95 3.8 ;
      RECT 41.79 3.6 41.99 3.8 ;
      RECT 40.59 3.04 40.79 3.24 ;
      RECT 39.35 2.48 39.55 2.68 ;
      RECT 37.91 3.04 38.11 3.24 ;
      RECT 37.17 2.48 37.37 2.68 ;
      RECT 35.95 2.48 36.15 2.68 ;
      RECT 35.47 3.6 35.67 3.8 ;
      RECT 27.15 1.92 27.35 2.12 ;
      RECT 26.19 3.6 26.39 3.8 ;
      RECT 25.455 7.14 25.655 7.34 ;
      RECT 25.19 3.6 25.39 3.8 ;
      RECT 23.23 3.6 23.43 3.8 ;
      RECT 22.03 3.04 22.23 3.24 ;
      RECT 20.79 2.48 20.99 2.68 ;
      RECT 19.35 3.04 19.55 3.24 ;
      RECT 18.61 2.48 18.81 2.68 ;
      RECT 17.39 2.48 17.59 2.68 ;
      RECT 16.91 3.6 17.11 3.8 ;
      RECT 8.59 1.92 8.79 2.12 ;
      RECT 7.63 3.6 7.83 3.8 ;
      RECT 6.895 7.14 7.095 7.34 ;
      RECT 6.63 3.6 6.83 3.8 ;
      RECT 4.67 3.6 4.87 3.8 ;
      RECT 3.47 3.04 3.67 3.24 ;
      RECT 2.23 2.48 2.43 2.68 ;
      RECT 0.79 3.04 0.99 3.24 ;
      RECT 0.05 2.48 0.25 2.68 ;
      RECT -1.17 2.48 -0.97 2.68 ;
      RECT -1.65 3.6 -1.45 3.8 ;
    LAYER met2 ;
      RECT -4.275 8.4 89.72 8.57 ;
      RECT 89.55 7.275 89.72 8.57 ;
      RECT -4.275 6.255 -4.105 8.57 ;
      RECT 89.52 7.275 89.87 7.625 ;
      RECT -4.34 6.255 -4.05 6.605 ;
      RECT 86.36 6.22 86.68 6.545 ;
      RECT 86.39 5.695 86.56 6.545 ;
      RECT 86.39 5.695 86.565 6.045 ;
      RECT 86.39 5.695 87.365 5.87 ;
      RECT 87.19 1.965 87.365 5.87 ;
      RECT 87.135 1.965 87.485 2.315 ;
      RECT 87.16 6.655 87.485 6.98 ;
      RECT 86.045 6.745 87.485 6.915 ;
      RECT 86.045 2.395 86.205 6.915 ;
      RECT 86.36 2.365 86.68 2.685 ;
      RECT 86.045 2.395 86.68 2.565 ;
      RECT 85.31 5.845 85.65 6.195 ;
      RECT 85.395 2.705 85.565 6.195 ;
      RECT 85.32 2.705 85.66 3.055 ;
      RECT 80.88 4.135 85.015 4.325 ;
      RECT 84.845 3.145 85.015 4.325 ;
      RECT 84.825 3.15 85.015 4.325 ;
      RECT 80.88 3.515 81.07 4.325 ;
      RECT 80.83 3.515 81.11 3.885 ;
      RECT 84.755 3.15 85.095 3.5 ;
      RECT 70.935 6.655 71.285 7.005 ;
      RECT 81.72 6.61 82.07 6.96 ;
      RECT 70.935 6.685 82.07 6.885 ;
      RECT 81.36 2.98 81.62 3.3 ;
      RECT 81.42 1.86 81.56 3.3 ;
      RECT 81.36 1.86 81.62 2.18 ;
      RECT 80.36 3.54 80.62 3.86 ;
      RECT 80.36 2.955 80.56 3.86 ;
      RECT 80.3 1.86 80.44 3.49 ;
      RECT 80.3 2.955 80.8 3.325 ;
      RECT 80.24 1.86 80.5 2.18 ;
      RECT 79.88 3.54 80.14 3.86 ;
      RECT 79.94 1.95 80.08 3.86 ;
      RECT 79.64 1.95 80.08 2.18 ;
      RECT 79.64 1.86 79.9 2.18 ;
      RECT 79.4 2.42 79.66 2.74 ;
      RECT 78.82 2.51 79.66 2.65 ;
      RECT 78.82 1.57 78.96 2.65 ;
      RECT 75.48 1.86 75.74 2.18 ;
      RECT 75.48 1.95 76.52 2.09 ;
      RECT 76.38 1.57 76.52 2.09 ;
      RECT 76.38 1.57 78.96 1.71 ;
      RECT 78.87 3.515 79.15 3.885 ;
      RECT 78.94 3.07 79.08 3.885 ;
      RECT 78.75 2.955 79.03 3.325 ;
      RECT 78.46 3.07 79.08 3.21 ;
      RECT 78.46 1.86 78.6 3.21 ;
      RECT 78.4 1.86 78.66 2.18 ;
      RECT 77.67 2.955 77.95 3.325 ;
      RECT 77.74 1.86 77.88 3.325 ;
      RECT 77.68 1.86 77.94 2.18 ;
      RECT 77.32 3.54 77.58 3.86 ;
      RECT 77.38 1.95 77.52 3.86 ;
      RECT 76.96 1.86 77.22 2.18 ;
      RECT 76.96 1.95 77.52 2.09 ;
      RECT 74.99 2.955 75.27 3.325 ;
      RECT 76.96 2.98 77.22 3.3 ;
      RECT 74.64 2.98 75.27 3.3 ;
      RECT 74.64 3.07 77.22 3.21 ;
      RECT 76.43 2.395 76.71 2.765 ;
      RECT 76.43 2.42 76.96 2.74 ;
      RECT 74 2.98 74.26 3.3 ;
      RECT 73.94 2.51 74.08 3.21 ;
      RECT 74.25 2.395 74.53 2.765 ;
      RECT 75.72 2.42 75.98 2.74 ;
      RECT 73.94 2.51 75.98 2.65 ;
      RECT 74.345 1 74.515 2.765 ;
      RECT 74.32 1 74.66 1.34 ;
      RECT 73.52 2.98 73.78 3.3 ;
      RECT 73.58 1.86 73.72 3.3 ;
      RECT 73.52 1.86 73.78 2.18 ;
      RECT 72.55 3.515 72.83 3.885 ;
      RECT 72.56 3.26 72.82 3.885 ;
      RECT 67.8 6.22 68.12 6.545 ;
      RECT 67.83 5.695 68 6.545 ;
      RECT 67.83 5.695 68.005 6.045 ;
      RECT 67.83 5.695 68.805 5.87 ;
      RECT 68.63 1.965 68.805 5.87 ;
      RECT 68.575 1.965 68.925 2.315 ;
      RECT 68.6 6.655 68.925 6.98 ;
      RECT 67.485 6.745 68.925 6.915 ;
      RECT 67.485 2.395 67.645 6.915 ;
      RECT 67.8 2.365 68.12 2.685 ;
      RECT 67.485 2.395 68.12 2.565 ;
      RECT 66.75 5.845 67.09 6.195 ;
      RECT 66.835 2.705 67.005 6.195 ;
      RECT 66.76 2.705 67.1 3.055 ;
      RECT 62.32 4.135 66.455 4.325 ;
      RECT 66.285 3.145 66.455 4.325 ;
      RECT 66.265 3.15 66.455 4.325 ;
      RECT 62.32 3.515 62.51 4.325 ;
      RECT 62.27 3.515 62.55 3.885 ;
      RECT 66.195 3.15 66.535 3.5 ;
      RECT 52.375 6.655 52.725 7.005 ;
      RECT 63.16 6.61 63.51 6.96 ;
      RECT 52.375 6.685 63.51 6.885 ;
      RECT 62.8 2.98 63.06 3.3 ;
      RECT 62.86 1.86 63 3.3 ;
      RECT 62.8 1.86 63.06 2.18 ;
      RECT 61.8 3.54 62.06 3.86 ;
      RECT 61.8 2.955 62 3.86 ;
      RECT 61.74 1.86 61.88 3.49 ;
      RECT 61.74 2.955 62.24 3.325 ;
      RECT 61.68 1.86 61.94 2.18 ;
      RECT 61.32 3.54 61.58 3.86 ;
      RECT 61.38 1.95 61.52 3.86 ;
      RECT 61.08 1.95 61.52 2.18 ;
      RECT 61.08 1.86 61.34 2.18 ;
      RECT 60.84 2.42 61.1 2.74 ;
      RECT 60.26 2.51 61.1 2.65 ;
      RECT 60.26 1.57 60.4 2.65 ;
      RECT 56.92 1.86 57.18 2.18 ;
      RECT 56.92 1.95 57.96 2.09 ;
      RECT 57.82 1.57 57.96 2.09 ;
      RECT 57.82 1.57 60.4 1.71 ;
      RECT 60.31 3.515 60.59 3.885 ;
      RECT 60.38 3.07 60.52 3.885 ;
      RECT 60.19 2.955 60.47 3.325 ;
      RECT 59.9 3.07 60.52 3.21 ;
      RECT 59.9 1.86 60.04 3.21 ;
      RECT 59.84 1.86 60.1 2.18 ;
      RECT 59.11 2.955 59.39 3.325 ;
      RECT 59.18 1.86 59.32 3.325 ;
      RECT 59.12 1.86 59.38 2.18 ;
      RECT 58.76 3.54 59.02 3.86 ;
      RECT 58.82 1.95 58.96 3.86 ;
      RECT 58.4 1.86 58.66 2.18 ;
      RECT 58.4 1.95 58.96 2.09 ;
      RECT 56.43 2.955 56.71 3.325 ;
      RECT 58.4 2.98 58.66 3.3 ;
      RECT 56.08 2.98 56.71 3.3 ;
      RECT 56.08 3.07 58.66 3.21 ;
      RECT 57.87 2.395 58.15 2.765 ;
      RECT 57.87 2.42 58.4 2.74 ;
      RECT 55.44 2.98 55.7 3.3 ;
      RECT 55.38 2.51 55.52 3.21 ;
      RECT 55.69 2.395 55.97 2.765 ;
      RECT 57.16 2.42 57.42 2.74 ;
      RECT 55.38 2.51 57.42 2.65 ;
      RECT 55.785 1 55.955 2.765 ;
      RECT 55.76 1 56.1 1.34 ;
      RECT 54.96 2.98 55.22 3.3 ;
      RECT 55.02 1.86 55.16 3.3 ;
      RECT 54.96 1.86 55.22 2.18 ;
      RECT 53.99 3.515 54.27 3.885 ;
      RECT 54 3.26 54.26 3.885 ;
      RECT 49.24 6.22 49.56 6.545 ;
      RECT 49.27 5.695 49.44 6.545 ;
      RECT 49.27 5.695 49.445 6.045 ;
      RECT 49.27 5.695 50.245 5.87 ;
      RECT 50.07 1.965 50.245 5.87 ;
      RECT 50.015 1.965 50.365 2.315 ;
      RECT 50.04 6.655 50.365 6.98 ;
      RECT 48.925 6.745 50.365 6.915 ;
      RECT 48.925 2.395 49.085 6.915 ;
      RECT 49.24 2.365 49.56 2.685 ;
      RECT 48.925 2.395 49.56 2.565 ;
      RECT 48.19 5.845 48.53 6.195 ;
      RECT 48.275 2.705 48.445 6.195 ;
      RECT 48.2 2.705 48.54 3.055 ;
      RECT 43.76 4.135 47.895 4.325 ;
      RECT 47.725 3.145 47.895 4.325 ;
      RECT 47.705 3.15 47.895 4.325 ;
      RECT 43.76 3.515 43.95 4.325 ;
      RECT 43.71 3.515 43.99 3.885 ;
      RECT 47.635 3.15 47.975 3.5 ;
      RECT 33.86 6.66 34.21 7.01 ;
      RECT 44.6 6.615 44.95 6.965 ;
      RECT 33.86 6.69 44.95 6.89 ;
      RECT 44.24 2.98 44.5 3.3 ;
      RECT 44.3 1.86 44.44 3.3 ;
      RECT 44.24 1.86 44.5 2.18 ;
      RECT 43.24 3.54 43.5 3.86 ;
      RECT 43.24 2.955 43.44 3.86 ;
      RECT 43.18 1.86 43.32 3.49 ;
      RECT 43.18 2.955 43.68 3.325 ;
      RECT 43.12 1.86 43.38 2.18 ;
      RECT 42.76 3.54 43.02 3.86 ;
      RECT 42.82 1.95 42.96 3.86 ;
      RECT 42.52 1.95 42.96 2.18 ;
      RECT 42.52 1.86 42.78 2.18 ;
      RECT 42.28 2.42 42.54 2.74 ;
      RECT 41.7 2.51 42.54 2.65 ;
      RECT 41.7 1.57 41.84 2.65 ;
      RECT 38.36 1.86 38.62 2.18 ;
      RECT 38.36 1.95 39.4 2.09 ;
      RECT 39.26 1.57 39.4 2.09 ;
      RECT 39.26 1.57 41.84 1.71 ;
      RECT 41.75 3.515 42.03 3.885 ;
      RECT 41.82 3.07 41.96 3.885 ;
      RECT 41.63 2.955 41.91 3.325 ;
      RECT 41.34 3.07 41.96 3.21 ;
      RECT 41.34 1.86 41.48 3.21 ;
      RECT 41.28 1.86 41.54 2.18 ;
      RECT 40.55 2.955 40.83 3.325 ;
      RECT 40.62 1.86 40.76 3.325 ;
      RECT 40.56 1.86 40.82 2.18 ;
      RECT 40.2 3.54 40.46 3.86 ;
      RECT 40.26 1.95 40.4 3.86 ;
      RECT 39.84 1.86 40.1 2.18 ;
      RECT 39.84 1.95 40.4 2.09 ;
      RECT 37.87 2.955 38.15 3.325 ;
      RECT 39.84 2.98 40.1 3.3 ;
      RECT 37.52 2.98 38.15 3.3 ;
      RECT 37.52 3.07 40.1 3.21 ;
      RECT 39.31 2.395 39.59 2.765 ;
      RECT 39.31 2.42 39.84 2.74 ;
      RECT 36.88 2.98 37.14 3.3 ;
      RECT 36.82 2.51 36.96 3.21 ;
      RECT 37.13 2.395 37.41 2.765 ;
      RECT 38.6 2.42 38.86 2.74 ;
      RECT 36.82 2.51 38.86 2.65 ;
      RECT 37.225 1 37.395 2.765 ;
      RECT 37.2 1 37.54 1.34 ;
      RECT 36.4 2.98 36.66 3.3 ;
      RECT 36.46 1.86 36.6 3.3 ;
      RECT 36.4 1.86 36.66 2.18 ;
      RECT 35.43 3.515 35.71 3.885 ;
      RECT 35.44 3.26 35.7 3.885 ;
      RECT 30.68 6.22 31 6.545 ;
      RECT 30.71 5.695 30.88 6.545 ;
      RECT 30.71 5.695 30.885 6.045 ;
      RECT 30.71 5.695 31.685 5.87 ;
      RECT 31.51 1.965 31.685 5.87 ;
      RECT 31.455 1.965 31.805 2.315 ;
      RECT 31.48 6.655 31.805 6.98 ;
      RECT 30.365 6.745 31.805 6.915 ;
      RECT 30.365 2.395 30.525 6.915 ;
      RECT 30.68 2.365 31 2.685 ;
      RECT 30.365 2.395 31 2.565 ;
      RECT 29.63 5.845 29.97 6.195 ;
      RECT 29.715 2.705 29.885 6.195 ;
      RECT 29.64 2.705 29.98 3.055 ;
      RECT 25.2 4.135 29.335 4.325 ;
      RECT 29.165 3.145 29.335 4.325 ;
      RECT 29.145 3.15 29.335 4.325 ;
      RECT 25.2 3.515 25.39 4.325 ;
      RECT 25.15 3.515 25.43 3.885 ;
      RECT 29.075 3.15 29.415 3.5 ;
      RECT 15.3 6.655 15.65 7.005 ;
      RECT 26.045 6.61 26.395 6.96 ;
      RECT 15.3 6.685 26.395 6.885 ;
      RECT 25.68 2.98 25.94 3.3 ;
      RECT 25.74 1.86 25.88 3.3 ;
      RECT 25.68 1.86 25.94 2.18 ;
      RECT 24.68 3.54 24.94 3.86 ;
      RECT 24.68 2.955 24.88 3.86 ;
      RECT 24.62 1.86 24.76 3.49 ;
      RECT 24.62 2.955 25.12 3.325 ;
      RECT 24.56 1.86 24.82 2.18 ;
      RECT 24.2 3.54 24.46 3.86 ;
      RECT 24.26 1.95 24.4 3.86 ;
      RECT 23.96 1.95 24.4 2.18 ;
      RECT 23.96 1.86 24.22 2.18 ;
      RECT 23.72 2.42 23.98 2.74 ;
      RECT 23.14 2.51 23.98 2.65 ;
      RECT 23.14 1.57 23.28 2.65 ;
      RECT 19.8 1.86 20.06 2.18 ;
      RECT 19.8 1.95 20.84 2.09 ;
      RECT 20.7 1.57 20.84 2.09 ;
      RECT 20.7 1.57 23.28 1.71 ;
      RECT 23.19 3.515 23.47 3.885 ;
      RECT 23.26 3.07 23.4 3.885 ;
      RECT 23.07 2.955 23.35 3.325 ;
      RECT 22.78 3.07 23.4 3.21 ;
      RECT 22.78 1.86 22.92 3.21 ;
      RECT 22.72 1.86 22.98 2.18 ;
      RECT 21.99 2.955 22.27 3.325 ;
      RECT 22.06 1.86 22.2 3.325 ;
      RECT 22 1.86 22.26 2.18 ;
      RECT 21.64 3.54 21.9 3.86 ;
      RECT 21.7 1.95 21.84 3.86 ;
      RECT 21.28 1.86 21.54 2.18 ;
      RECT 21.28 1.95 21.84 2.09 ;
      RECT 19.31 2.955 19.59 3.325 ;
      RECT 21.28 2.98 21.54 3.3 ;
      RECT 18.96 2.98 19.59 3.3 ;
      RECT 18.96 3.07 21.54 3.21 ;
      RECT 20.75 2.395 21.03 2.765 ;
      RECT 20.75 2.42 21.28 2.74 ;
      RECT 18.32 2.98 18.58 3.3 ;
      RECT 18.26 2.51 18.4 3.21 ;
      RECT 18.57 2.395 18.85 2.765 ;
      RECT 20.04 2.42 20.3 2.74 ;
      RECT 18.26 2.51 20.3 2.65 ;
      RECT 18.665 1 18.835 2.765 ;
      RECT 18.64 1 18.98 1.34 ;
      RECT 17.84 2.98 18.1 3.3 ;
      RECT 17.9 1.86 18.04 3.3 ;
      RECT 17.84 1.86 18.1 2.18 ;
      RECT 16.87 3.515 17.15 3.885 ;
      RECT 16.88 3.26 17.14 3.885 ;
      RECT 12.12 6.22 12.44 6.545 ;
      RECT 12.15 5.695 12.32 6.545 ;
      RECT 12.15 5.695 12.325 6.045 ;
      RECT 12.15 5.695 13.125 5.87 ;
      RECT 12.95 1.965 13.125 5.87 ;
      RECT 12.895 1.965 13.245 2.315 ;
      RECT 12.92 6.655 13.245 6.98 ;
      RECT 11.805 6.745 13.245 6.915 ;
      RECT 11.805 2.395 11.965 6.915 ;
      RECT 12.12 2.365 12.44 2.685 ;
      RECT 11.805 2.395 12.44 2.565 ;
      RECT 11.07 5.845 11.41 6.195 ;
      RECT 11.155 2.705 11.325 6.195 ;
      RECT 11.08 2.705 11.42 3.055 ;
      RECT 6.64 4.135 10.775 4.325 ;
      RECT 10.605 3.145 10.775 4.325 ;
      RECT 10.585 3.15 10.775 4.325 ;
      RECT 6.64 3.515 6.83 4.325 ;
      RECT 6.59 3.515 6.87 3.885 ;
      RECT 10.515 3.15 10.855 3.5 ;
      RECT -3.965 6.995 -3.675 7.345 ;
      RECT -3.965 7.05 -2.65 7.22 ;
      RECT -2.82 6.685 -2.65 7.22 ;
      RECT 7.485 6.605 7.835 6.955 ;
      RECT -2.82 6.685 7.835 6.855 ;
      RECT 7.12 2.98 7.38 3.3 ;
      RECT 7.18 1.86 7.32 3.3 ;
      RECT 7.12 1.86 7.38 2.18 ;
      RECT 6.12 3.54 6.38 3.86 ;
      RECT 6.12 2.955 6.32 3.86 ;
      RECT 6.06 1.86 6.2 3.49 ;
      RECT 6.06 2.955 6.56 3.325 ;
      RECT 6 1.86 6.26 2.18 ;
      RECT 5.64 3.54 5.9 3.86 ;
      RECT 5.7 1.95 5.84 3.86 ;
      RECT 5.4 1.95 5.84 2.18 ;
      RECT 5.4 1.86 5.66 2.18 ;
      RECT 5.16 2.42 5.42 2.74 ;
      RECT 4.58 2.51 5.42 2.65 ;
      RECT 4.58 1.57 4.72 2.65 ;
      RECT 1.24 1.86 1.5 2.18 ;
      RECT 1.24 1.95 2.28 2.09 ;
      RECT 2.14 1.57 2.28 2.09 ;
      RECT 2.14 1.57 4.72 1.71 ;
      RECT 4.63 3.515 4.91 3.885 ;
      RECT 4.7 3.07 4.84 3.885 ;
      RECT 4.51 2.955 4.79 3.325 ;
      RECT 4.22 3.07 4.84 3.21 ;
      RECT 4.22 1.86 4.36 3.21 ;
      RECT 4.16 1.86 4.42 2.18 ;
      RECT 3.43 2.955 3.71 3.325 ;
      RECT 3.5 1.86 3.64 3.325 ;
      RECT 3.44 1.86 3.7 2.18 ;
      RECT 3.08 3.54 3.34 3.86 ;
      RECT 3.14 1.95 3.28 3.86 ;
      RECT 2.72 1.86 2.98 2.18 ;
      RECT 2.72 1.95 3.28 2.09 ;
      RECT 0.75 2.955 1.03 3.325 ;
      RECT 2.72 2.98 2.98 3.3 ;
      RECT 0.4 2.98 1.03 3.3 ;
      RECT 0.4 3.07 2.98 3.21 ;
      RECT 2.19 2.395 2.47 2.765 ;
      RECT 2.19 2.42 2.72 2.74 ;
      RECT -0.24 2.98 0.02 3.3 ;
      RECT -0.3 2.51 -0.16 3.21 ;
      RECT 0.01 2.395 0.29 2.765 ;
      RECT 1.48 2.42 1.74 2.74 ;
      RECT -0.3 2.51 1.74 2.65 ;
      RECT 0.105 1 0.275 2.765 ;
      RECT 0.08 1 0.42 1.34 ;
      RECT -0.72 2.98 -0.46 3.3 ;
      RECT -0.66 1.86 -0.52 3.3 ;
      RECT -0.72 1.86 -0.46 2.18 ;
      RECT -1.69 3.515 -1.41 3.885 ;
      RECT -1.68 3.26 -1.42 3.885 ;
      RECT 82.79 1.835 83.07 2.205 ;
      RECT 81.83 3.515 82.11 3.885 ;
      RECT 81.05 7.055 81.425 7.425 ;
      RECT 73.03 2.395 73.31 2.765 ;
      RECT 64.23 1.835 64.51 2.205 ;
      RECT 63.27 3.515 63.55 3.885 ;
      RECT 62.49 7.055 62.865 7.425 ;
      RECT 54.47 2.395 54.75 2.765 ;
      RECT 45.67 1.835 45.95 2.205 ;
      RECT 44.71 3.515 44.99 3.885 ;
      RECT 43.93 7.055 44.305 7.425 ;
      RECT 35.91 2.395 36.19 2.765 ;
      RECT 27.11 1.835 27.39 2.205 ;
      RECT 26.15 3.515 26.43 3.885 ;
      RECT 25.37 7.055 25.745 7.425 ;
      RECT 17.35 2.395 17.63 2.765 ;
      RECT 8.55 1.835 8.83 2.205 ;
      RECT 7.59 3.515 7.87 3.885 ;
      RECT 6.81 7.055 7.185 7.425 ;
      RECT -1.21 2.395 -0.93 2.765 ;
    LAYER via1 ;
      RECT 89.62 7.375 89.77 7.525 ;
      RECT 87.25 6.74 87.4 6.89 ;
      RECT 87.235 2.065 87.385 2.215 ;
      RECT 86.445 2.45 86.595 2.6 ;
      RECT 86.445 6.325 86.595 6.475 ;
      RECT 85.42 2.805 85.57 2.955 ;
      RECT 85.41 5.945 85.56 6.095 ;
      RECT 84.855 3.25 85.005 3.4 ;
      RECT 82.855 1.945 83.005 2.095 ;
      RECT 81.895 3.625 82.045 3.775 ;
      RECT 81.82 6.71 81.97 6.86 ;
      RECT 81.415 1.945 81.565 2.095 ;
      RECT 81.415 3.065 81.565 3.215 ;
      RECT 81.16 7.165 81.31 7.315 ;
      RECT 80.895 3.625 81.045 3.775 ;
      RECT 80.415 3.625 80.565 3.775 ;
      RECT 80.295 1.945 80.445 2.095 ;
      RECT 79.935 3.625 80.085 3.775 ;
      RECT 79.695 1.945 79.845 2.095 ;
      RECT 79.455 2.505 79.605 2.655 ;
      RECT 78.935 3.625 79.085 3.775 ;
      RECT 78.455 1.945 78.605 2.095 ;
      RECT 77.735 1.945 77.885 2.095 ;
      RECT 77.735 3.065 77.885 3.215 ;
      RECT 77.375 3.625 77.525 3.775 ;
      RECT 77.015 1.945 77.165 2.095 ;
      RECT 77.015 3.065 77.165 3.215 ;
      RECT 76.755 2.505 76.905 2.655 ;
      RECT 75.775 2.505 75.925 2.655 ;
      RECT 75.535 1.945 75.685 2.095 ;
      RECT 74.695 3.065 74.845 3.215 ;
      RECT 74.415 1.095 74.565 1.245 ;
      RECT 74.055 3.065 74.205 3.215 ;
      RECT 73.575 1.945 73.725 2.095 ;
      RECT 73.575 3.065 73.725 3.215 ;
      RECT 73.095 2.505 73.245 2.655 ;
      RECT 72.615 3.345 72.765 3.495 ;
      RECT 71.035 6.755 71.185 6.905 ;
      RECT 68.69 6.74 68.84 6.89 ;
      RECT 68.675 2.065 68.825 2.215 ;
      RECT 67.885 2.45 68.035 2.6 ;
      RECT 67.885 6.325 68.035 6.475 ;
      RECT 66.86 2.805 67.01 2.955 ;
      RECT 66.85 5.945 67 6.095 ;
      RECT 66.295 3.25 66.445 3.4 ;
      RECT 64.295 1.945 64.445 2.095 ;
      RECT 63.335 3.625 63.485 3.775 ;
      RECT 63.26 6.71 63.41 6.86 ;
      RECT 62.855 1.945 63.005 2.095 ;
      RECT 62.855 3.065 63.005 3.215 ;
      RECT 62.6 7.165 62.75 7.315 ;
      RECT 62.335 3.625 62.485 3.775 ;
      RECT 61.855 3.625 62.005 3.775 ;
      RECT 61.735 1.945 61.885 2.095 ;
      RECT 61.375 3.625 61.525 3.775 ;
      RECT 61.135 1.945 61.285 2.095 ;
      RECT 60.895 2.505 61.045 2.655 ;
      RECT 60.375 3.625 60.525 3.775 ;
      RECT 59.895 1.945 60.045 2.095 ;
      RECT 59.175 1.945 59.325 2.095 ;
      RECT 59.175 3.065 59.325 3.215 ;
      RECT 58.815 3.625 58.965 3.775 ;
      RECT 58.455 1.945 58.605 2.095 ;
      RECT 58.455 3.065 58.605 3.215 ;
      RECT 58.195 2.505 58.345 2.655 ;
      RECT 57.215 2.505 57.365 2.655 ;
      RECT 56.975 1.945 57.125 2.095 ;
      RECT 56.135 3.065 56.285 3.215 ;
      RECT 55.855 1.095 56.005 1.245 ;
      RECT 55.495 3.065 55.645 3.215 ;
      RECT 55.015 1.945 55.165 2.095 ;
      RECT 55.015 3.065 55.165 3.215 ;
      RECT 54.535 2.505 54.685 2.655 ;
      RECT 54.055 3.345 54.205 3.495 ;
      RECT 52.475 6.755 52.625 6.905 ;
      RECT 50.13 6.74 50.28 6.89 ;
      RECT 50.115 2.065 50.265 2.215 ;
      RECT 49.325 2.45 49.475 2.6 ;
      RECT 49.325 6.325 49.475 6.475 ;
      RECT 48.3 2.805 48.45 2.955 ;
      RECT 48.29 5.945 48.44 6.095 ;
      RECT 47.735 3.25 47.885 3.4 ;
      RECT 45.735 1.945 45.885 2.095 ;
      RECT 44.775 3.625 44.925 3.775 ;
      RECT 44.7 6.715 44.85 6.865 ;
      RECT 44.295 1.945 44.445 2.095 ;
      RECT 44.295 3.065 44.445 3.215 ;
      RECT 44.04 7.165 44.19 7.315 ;
      RECT 43.775 3.625 43.925 3.775 ;
      RECT 43.295 3.625 43.445 3.775 ;
      RECT 43.175 1.945 43.325 2.095 ;
      RECT 42.815 3.625 42.965 3.775 ;
      RECT 42.575 1.945 42.725 2.095 ;
      RECT 42.335 2.505 42.485 2.655 ;
      RECT 41.815 3.625 41.965 3.775 ;
      RECT 41.335 1.945 41.485 2.095 ;
      RECT 40.615 1.945 40.765 2.095 ;
      RECT 40.615 3.065 40.765 3.215 ;
      RECT 40.255 3.625 40.405 3.775 ;
      RECT 39.895 1.945 40.045 2.095 ;
      RECT 39.895 3.065 40.045 3.215 ;
      RECT 39.635 2.505 39.785 2.655 ;
      RECT 38.655 2.505 38.805 2.655 ;
      RECT 38.415 1.945 38.565 2.095 ;
      RECT 37.575 3.065 37.725 3.215 ;
      RECT 37.295 1.095 37.445 1.245 ;
      RECT 36.935 3.065 37.085 3.215 ;
      RECT 36.455 1.945 36.605 2.095 ;
      RECT 36.455 3.065 36.605 3.215 ;
      RECT 35.975 2.505 36.125 2.655 ;
      RECT 35.495 3.345 35.645 3.495 ;
      RECT 33.96 6.76 34.11 6.91 ;
      RECT 31.57 6.74 31.72 6.89 ;
      RECT 31.555 2.065 31.705 2.215 ;
      RECT 30.765 2.45 30.915 2.6 ;
      RECT 30.765 6.325 30.915 6.475 ;
      RECT 29.74 2.805 29.89 2.955 ;
      RECT 29.73 5.945 29.88 6.095 ;
      RECT 29.175 3.25 29.325 3.4 ;
      RECT 27.175 1.945 27.325 2.095 ;
      RECT 26.215 3.625 26.365 3.775 ;
      RECT 26.145 6.71 26.295 6.86 ;
      RECT 25.735 1.945 25.885 2.095 ;
      RECT 25.735 3.065 25.885 3.215 ;
      RECT 25.48 7.165 25.63 7.315 ;
      RECT 25.215 3.625 25.365 3.775 ;
      RECT 24.735 3.625 24.885 3.775 ;
      RECT 24.615 1.945 24.765 2.095 ;
      RECT 24.255 3.625 24.405 3.775 ;
      RECT 24.015 1.945 24.165 2.095 ;
      RECT 23.775 2.505 23.925 2.655 ;
      RECT 23.255 3.625 23.405 3.775 ;
      RECT 22.775 1.945 22.925 2.095 ;
      RECT 22.055 1.945 22.205 2.095 ;
      RECT 22.055 3.065 22.205 3.215 ;
      RECT 21.695 3.625 21.845 3.775 ;
      RECT 21.335 1.945 21.485 2.095 ;
      RECT 21.335 3.065 21.485 3.215 ;
      RECT 21.075 2.505 21.225 2.655 ;
      RECT 20.095 2.505 20.245 2.655 ;
      RECT 19.855 1.945 20.005 2.095 ;
      RECT 19.015 3.065 19.165 3.215 ;
      RECT 18.735 1.095 18.885 1.245 ;
      RECT 18.375 3.065 18.525 3.215 ;
      RECT 17.895 1.945 18.045 2.095 ;
      RECT 17.895 3.065 18.045 3.215 ;
      RECT 17.415 2.505 17.565 2.655 ;
      RECT 16.935 3.345 17.085 3.495 ;
      RECT 15.4 6.755 15.55 6.905 ;
      RECT 13.01 6.74 13.16 6.89 ;
      RECT 12.995 2.065 13.145 2.215 ;
      RECT 12.205 2.45 12.355 2.6 ;
      RECT 12.205 6.325 12.355 6.475 ;
      RECT 11.18 2.805 11.33 2.955 ;
      RECT 11.17 5.945 11.32 6.095 ;
      RECT 10.615 3.25 10.765 3.4 ;
      RECT 8.615 1.945 8.765 2.095 ;
      RECT 7.655 3.625 7.805 3.775 ;
      RECT 7.585 6.705 7.735 6.855 ;
      RECT 7.175 1.945 7.325 2.095 ;
      RECT 7.175 3.065 7.325 3.215 ;
      RECT 6.92 7.165 7.07 7.315 ;
      RECT 6.655 3.625 6.805 3.775 ;
      RECT 6.175 3.625 6.325 3.775 ;
      RECT 6.055 1.945 6.205 2.095 ;
      RECT 5.695 3.625 5.845 3.775 ;
      RECT 5.455 1.945 5.605 2.095 ;
      RECT 5.215 2.505 5.365 2.655 ;
      RECT 4.695 3.625 4.845 3.775 ;
      RECT 4.215 1.945 4.365 2.095 ;
      RECT 3.495 1.945 3.645 2.095 ;
      RECT 3.495 3.065 3.645 3.215 ;
      RECT 3.135 3.625 3.285 3.775 ;
      RECT 2.775 1.945 2.925 2.095 ;
      RECT 2.775 3.065 2.925 3.215 ;
      RECT 2.515 2.505 2.665 2.655 ;
      RECT 1.535 2.505 1.685 2.655 ;
      RECT 1.295 1.945 1.445 2.095 ;
      RECT 0.455 3.065 0.605 3.215 ;
      RECT 0.175 1.095 0.325 1.245 ;
      RECT -0.185 3.065 -0.035 3.215 ;
      RECT -0.665 1.945 -0.515 2.095 ;
      RECT -0.665 3.065 -0.515 3.215 ;
      RECT -1.145 2.505 -0.995 2.655 ;
      RECT -1.625 3.345 -1.475 3.495 ;
      RECT -3.895 7.095 -3.745 7.245 ;
      RECT -4.27 6.355 -4.12 6.505 ;
    LAYER met1 ;
      RECT 72.275 0 84.235 1.74 ;
      RECT 53.715 0 65.675 1.74 ;
      RECT 35.155 0 47.115 1.74 ;
      RECT 16.595 0 28.555 1.74 ;
      RECT -1.965 0 9.995 1.74 ;
      RECT 72.275 0 84.32 1.585 ;
      RECT 53.715 0 65.76 1.585 ;
      RECT 35.155 0 47.2 1.585 ;
      RECT 16.595 0 28.64 1.585 ;
      RECT -1.965 0 10.08 1.585 ;
      RECT -5.465 0 90.09 0.305 ;
      RECT 71.53 4.145 73.995 4.75 ;
      RECT 52.97 4.145 55.435 4.75 ;
      RECT 34.41 4.145 36.875 4.75 ;
      RECT 15.85 4.145 18.315 4.75 ;
      RECT -5.46 4.145 -0.245 4.75 ;
      RECT 72.275 4.135 90.09 4.745 ;
      RECT 53.715 4.135 71.53 4.745 ;
      RECT 35.155 4.135 52.97 4.745 ;
      RECT 16.595 4.135 34.41 4.745 ;
      RECT -1.965 4.135 15.85 4.745 ;
      RECT 72.275 3.98 84.235 4.745 ;
      RECT 53.715 3.98 65.675 4.745 ;
      RECT 35.155 3.98 47.115 4.745 ;
      RECT 16.595 3.98 28.555 4.745 ;
      RECT -1.965 3.98 9.995 4.745 ;
      RECT -5.465 8.575 90.09 8.88 ;
      RECT 80.28 6.315 80.45 8.88 ;
      RECT 61.72 6.315 61.89 8.88 ;
      RECT 43.16 6.315 43.33 8.88 ;
      RECT 24.6 6.315 24.77 8.88 ;
      RECT 6.04 6.315 6.21 8.88 ;
      RECT 80.715 6.285 81.005 6.515 ;
      RECT 62.155 6.285 62.445 6.515 ;
      RECT 43.595 6.285 43.885 6.515 ;
      RECT 25.035 6.285 25.325 6.515 ;
      RECT 6.475 6.285 6.765 6.515 ;
      RECT 80.28 6.315 81.005 6.485 ;
      RECT 61.72 6.315 62.445 6.485 ;
      RECT 43.16 6.315 43.885 6.485 ;
      RECT 24.6 6.315 25.325 6.485 ;
      RECT 6.04 6.315 6.765 6.485 ;
      RECT 89.49 7.765 89.78 7.995 ;
      RECT 89.55 6.285 89.72 7.995 ;
      RECT 89.52 7.275 89.87 7.625 ;
      RECT 89.49 6.285 89.78 6.515 ;
      RECT 89.49 2.365 89.78 2.595 ;
      RECT 89.55 0.885 89.72 2.595 ;
      RECT 89.49 0.885 89.78 1.115 ;
      RECT 89.08 2.735 89.41 2.965 ;
      RECT 89.08 2.765 89.58 2.935 ;
      RECT 89.08 2.395 89.27 2.965 ;
      RECT 88.5 2.365 88.79 2.595 ;
      RECT 88.5 2.395 89.27 2.565 ;
      RECT 88.56 0.885 88.73 2.595 ;
      RECT 88.5 0.885 88.79 1.115 ;
      RECT 88.5 7.765 88.79 7.995 ;
      RECT 88.56 6.285 88.73 7.995 ;
      RECT 88.5 6.285 88.79 6.515 ;
      RECT 88.5 6.325 89.35 6.485 ;
      RECT 89.18 5.915 89.35 6.485 ;
      RECT 88.5 6.32 88.89 6.485 ;
      RECT 89.12 5.915 89.41 6.145 ;
      RECT 89.12 5.945 89.58 6.115 ;
      RECT 88.13 2.735 88.42 2.965 ;
      RECT 88.13 2.765 88.59 2.935 ;
      RECT 88.19 1.655 88.355 2.965 ;
      RECT 86.705 1.625 86.995 1.855 ;
      RECT 86.705 1.655 88.355 1.825 ;
      RECT 86.765 0.885 86.935 1.855 ;
      RECT 86.705 0.885 86.995 1.115 ;
      RECT 86.705 7.765 86.995 7.995 ;
      RECT 86.765 7.025 86.935 7.995 ;
      RECT 86.765 7.12 88.355 7.29 ;
      RECT 88.185 5.915 88.355 7.29 ;
      RECT 86.705 7.025 86.995 7.255 ;
      RECT 88.13 5.915 88.42 6.145 ;
      RECT 88.13 5.945 88.59 6.115 ;
      RECT 84.755 3.15 85.095 3.5 ;
      RECT 84.845 2.025 85.015 3.5 ;
      RECT 87.135 1.965 87.485 2.315 ;
      RECT 84.845 2.025 87.485 2.195 ;
      RECT 87.16 6.655 87.485 6.98 ;
      RECT 81.72 6.61 82.07 6.96 ;
      RECT 87.135 6.655 87.485 6.885 ;
      RECT 81.52 6.655 82.07 6.885 ;
      RECT 81.35 6.685 87.485 6.855 ;
      RECT 86.36 2.365 86.68 2.685 ;
      RECT 86.33 2.365 86.68 2.595 ;
      RECT 86.16 2.395 86.68 2.565 ;
      RECT 86.36 6.255 86.68 6.545 ;
      RECT 86.33 6.285 86.68 6.515 ;
      RECT 86.16 6.315 86.68 6.485 ;
      RECT 85.32 2.705 85.66 3.055 ;
      RECT 85.32 2.765 85.795 2.935 ;
      RECT 85.31 5.845 85.65 6.195 ;
      RECT 79.72 5.915 80.01 6.145 ;
      RECT 79.72 5.945 85.795 6.115 ;
      RECT 81.81 3.57 82.13 3.83 ;
      RECT 83.1 2.745 83.24 3.605 ;
      RECT 81.9 3.465 83.24 3.605 ;
      RECT 81.9 3.025 82.04 3.83 ;
      RECT 81.825 3.025 82.115 3.255 ;
      RECT 83.025 2.745 83.315 2.975 ;
      RECT 82.545 3.025 82.835 3.255 ;
      RECT 82.74 1.95 82.88 3.21 ;
      RECT 82.77 1.89 83.09 2.15 ;
      RECT 79.37 2.45 79.69 2.71 ;
      RECT 82.065 2.465 82.355 2.695 ;
      RECT 79.46 2.37 82.28 2.51 ;
      RECT 81.33 1.89 81.65 2.15 ;
      RECT 81.825 1.905 82.115 2.135 ;
      RECT 81.33 1.95 82.115 2.09 ;
      RECT 81.33 3.01 81.65 3.27 ;
      RECT 81.33 2.79 81.56 3.27 ;
      RECT 80.825 2.745 81.115 2.975 ;
      RECT 80.825 2.79 81.56 2.93 ;
      RECT 81.09 7.765 81.38 7.995 ;
      RECT 81.15 7.025 81.32 7.995 ;
      RECT 81.05 7.055 81.43 7.425 ;
      RECT 81.09 7.025 81.38 7.425 ;
      RECT 79.85 3.57 80.17 3.83 ;
      RECT 79.385 3.585 79.675 3.815 ;
      RECT 79.385 3.63 80.17 3.77 ;
      RECT 78.145 2.465 78.435 2.695 ;
      RECT 78.145 2.51 79.08 2.65 ;
      RECT 78.94 1.95 79.08 2.65 ;
      RECT 79.61 1.89 79.93 2.15 ;
      RECT 79.385 1.905 79.93 2.135 ;
      RECT 78.94 1.95 79.93 2.09 ;
      RECT 77.29 3.57 77.61 3.83 ;
      RECT 77.29 3.63 78.36 3.77 ;
      RECT 78.22 3.07 78.36 3.77 ;
      RECT 79.385 3.025 79.675 3.255 ;
      RECT 78.22 3.07 79.675 3.21 ;
      RECT 77.65 1.89 77.97 2.15 ;
      RECT 77.425 1.905 77.97 2.135 ;
      RECT 76.67 2.45 76.99 2.71 ;
      RECT 77.665 2.465 77.955 2.695 ;
      RECT 76.425 2.465 76.99 2.695 ;
      RECT 76.425 2.51 77.955 2.65 ;
      RECT 75.945 3.025 76.235 3.255 ;
      RECT 76.14 1.95 76.28 3.21 ;
      RECT 76.93 1.89 77.25 2.15 ;
      RECT 75.945 1.905 76.235 2.135 ;
      RECT 75.945 1.95 77.25 2.09 ;
      RECT 75.54 3.465 76.64 3.605 ;
      RECT 76.425 3.305 76.715 3.535 ;
      RECT 75.465 3.305 75.755 3.535 ;
      RECT 75.705 2.37 75.995 2.74 ;
      RECT 74.94 2.37 75.995 2.51 ;
      RECT 75.45 1.89 75.77 2.15 ;
      RECT 73.49 1.89 73.81 2.15 ;
      RECT 73.49 1.95 75.77 2.09 ;
      RECT 74.61 3.01 74.93 3.27 ;
      RECT 74.61 3.01 75.44 3.15 ;
      RECT 75.225 2.745 75.44 3.15 ;
      RECT 75.225 2.745 75.515 2.975 ;
      RECT 73.01 2.45 73.33 2.71 ;
      RECT 74.42 2.465 74.71 2.695 ;
      RECT 73.01 2.465 73.555 2.695 ;
      RECT 73.01 2.55 73.96 2.69 ;
      RECT 73.82 2.37 73.96 2.69 ;
      RECT 74.32 2.465 74.71 2.65 ;
      RECT 73.82 2.37 74.46 2.51 ;
      RECT 72.53 3.26 72.85 3.675 ;
      RECT 72.61 1.905 72.765 3.675 ;
      RECT 72.545 1.905 72.835 2.135 ;
      RECT 70.93 7.765 71.22 7.995 ;
      RECT 70.99 6.285 71.16 7.995 ;
      RECT 70.935 6.655 71.285 7.005 ;
      RECT 70.93 6.285 71.22 6.515 ;
      RECT 70.93 2.365 71.22 2.595 ;
      RECT 70.99 0.885 71.16 2.595 ;
      RECT 70.93 0.885 71.22 1.115 ;
      RECT 70.52 2.735 70.85 2.965 ;
      RECT 70.52 2.765 71.02 2.935 ;
      RECT 70.52 2.395 70.71 2.965 ;
      RECT 69.94 2.365 70.23 2.595 ;
      RECT 69.94 2.395 70.71 2.565 ;
      RECT 70 0.885 70.17 2.595 ;
      RECT 69.94 0.885 70.23 1.115 ;
      RECT 69.94 7.765 70.23 7.995 ;
      RECT 70 6.285 70.17 7.995 ;
      RECT 69.94 6.285 70.23 6.515 ;
      RECT 69.94 6.325 70.79 6.485 ;
      RECT 70.62 5.915 70.79 6.485 ;
      RECT 69.94 6.32 70.33 6.485 ;
      RECT 70.56 5.915 70.85 6.145 ;
      RECT 70.56 5.945 71.02 6.115 ;
      RECT 69.57 2.735 69.86 2.965 ;
      RECT 69.57 2.765 70.03 2.935 ;
      RECT 69.63 1.655 69.795 2.965 ;
      RECT 68.145 1.625 68.435 1.855 ;
      RECT 68.145 1.655 69.795 1.825 ;
      RECT 68.205 0.885 68.375 1.855 ;
      RECT 68.145 0.885 68.435 1.115 ;
      RECT 68.145 7.765 68.435 7.995 ;
      RECT 68.205 7.025 68.375 7.995 ;
      RECT 68.205 7.12 69.795 7.29 ;
      RECT 69.625 5.915 69.795 7.29 ;
      RECT 68.145 7.025 68.435 7.255 ;
      RECT 69.57 5.915 69.86 6.145 ;
      RECT 69.57 5.945 70.03 6.115 ;
      RECT 66.195 3.15 66.535 3.5 ;
      RECT 66.285 2.025 66.455 3.5 ;
      RECT 68.575 1.965 68.925 2.315 ;
      RECT 66.285 2.025 68.925 2.195 ;
      RECT 68.6 6.655 68.925 6.98 ;
      RECT 63.16 6.61 63.51 6.96 ;
      RECT 68.575 6.655 68.925 6.885 ;
      RECT 62.96 6.655 63.51 6.885 ;
      RECT 62.79 6.685 68.925 6.855 ;
      RECT 67.8 2.365 68.12 2.685 ;
      RECT 67.77 2.365 68.12 2.595 ;
      RECT 67.6 2.395 68.12 2.565 ;
      RECT 67.8 6.255 68.12 6.545 ;
      RECT 67.77 6.285 68.12 6.515 ;
      RECT 67.6 6.315 68.12 6.485 ;
      RECT 66.76 2.705 67.1 3.055 ;
      RECT 66.76 2.765 67.235 2.935 ;
      RECT 66.75 5.845 67.09 6.195 ;
      RECT 61.16 5.915 61.45 6.145 ;
      RECT 61.16 5.945 67.235 6.115 ;
      RECT 63.25 3.57 63.57 3.83 ;
      RECT 64.54 2.745 64.68 3.605 ;
      RECT 63.34 3.465 64.68 3.605 ;
      RECT 63.34 3.025 63.48 3.83 ;
      RECT 63.265 3.025 63.555 3.255 ;
      RECT 64.465 2.745 64.755 2.975 ;
      RECT 63.985 3.025 64.275 3.255 ;
      RECT 64.18 1.95 64.32 3.21 ;
      RECT 64.21 1.89 64.53 2.15 ;
      RECT 60.81 2.45 61.13 2.71 ;
      RECT 63.505 2.465 63.795 2.695 ;
      RECT 60.9 2.37 63.72 2.51 ;
      RECT 62.77 1.89 63.09 2.15 ;
      RECT 63.265 1.905 63.555 2.135 ;
      RECT 62.77 1.95 63.555 2.09 ;
      RECT 62.77 3.01 63.09 3.27 ;
      RECT 62.77 2.79 63 3.27 ;
      RECT 62.265 2.745 62.555 2.975 ;
      RECT 62.265 2.79 63 2.93 ;
      RECT 62.53 7.765 62.82 7.995 ;
      RECT 62.59 7.025 62.76 7.995 ;
      RECT 62.49 7.055 62.87 7.425 ;
      RECT 62.53 7.025 62.82 7.425 ;
      RECT 61.29 3.57 61.61 3.83 ;
      RECT 60.825 3.585 61.115 3.815 ;
      RECT 60.825 3.63 61.61 3.77 ;
      RECT 59.585 2.465 59.875 2.695 ;
      RECT 59.585 2.51 60.52 2.65 ;
      RECT 60.38 1.95 60.52 2.65 ;
      RECT 61.05 1.89 61.37 2.15 ;
      RECT 60.825 1.905 61.37 2.135 ;
      RECT 60.38 1.95 61.37 2.09 ;
      RECT 58.73 3.57 59.05 3.83 ;
      RECT 58.73 3.63 59.8 3.77 ;
      RECT 59.66 3.07 59.8 3.77 ;
      RECT 60.825 3.025 61.115 3.255 ;
      RECT 59.66 3.07 61.115 3.21 ;
      RECT 59.09 1.89 59.41 2.15 ;
      RECT 58.865 1.905 59.41 2.135 ;
      RECT 58.11 2.45 58.43 2.71 ;
      RECT 59.105 2.465 59.395 2.695 ;
      RECT 57.865 2.465 58.43 2.695 ;
      RECT 57.865 2.51 59.395 2.65 ;
      RECT 57.385 3.025 57.675 3.255 ;
      RECT 57.58 1.95 57.72 3.21 ;
      RECT 58.37 1.89 58.69 2.15 ;
      RECT 57.385 1.905 57.675 2.135 ;
      RECT 57.385 1.95 58.69 2.09 ;
      RECT 56.98 3.465 58.08 3.605 ;
      RECT 57.865 3.305 58.155 3.535 ;
      RECT 56.905 3.305 57.195 3.535 ;
      RECT 57.145 2.37 57.435 2.74 ;
      RECT 56.38 2.37 57.435 2.51 ;
      RECT 56.89 1.89 57.21 2.15 ;
      RECT 54.93 1.89 55.25 2.15 ;
      RECT 54.93 1.95 57.21 2.09 ;
      RECT 56.05 3.01 56.37 3.27 ;
      RECT 56.05 3.01 56.88 3.15 ;
      RECT 56.665 2.745 56.88 3.15 ;
      RECT 56.665 2.745 56.955 2.975 ;
      RECT 54.45 2.45 54.77 2.71 ;
      RECT 55.86 2.465 56.15 2.695 ;
      RECT 54.45 2.465 54.995 2.695 ;
      RECT 54.45 2.55 55.4 2.69 ;
      RECT 55.26 2.37 55.4 2.69 ;
      RECT 55.76 2.465 56.15 2.65 ;
      RECT 55.26 2.37 55.9 2.51 ;
      RECT 53.97 3.26 54.29 3.675 ;
      RECT 54.05 1.905 54.205 3.675 ;
      RECT 53.985 1.905 54.275 2.135 ;
      RECT 52.37 7.765 52.66 7.995 ;
      RECT 52.43 6.285 52.6 7.995 ;
      RECT 52.375 6.655 52.725 7.005 ;
      RECT 52.37 6.285 52.66 6.515 ;
      RECT 52.37 2.365 52.66 2.595 ;
      RECT 52.43 0.885 52.6 2.595 ;
      RECT 52.37 0.885 52.66 1.115 ;
      RECT 51.96 2.735 52.29 2.965 ;
      RECT 51.96 2.765 52.46 2.935 ;
      RECT 51.96 2.395 52.15 2.965 ;
      RECT 51.38 2.365 51.67 2.595 ;
      RECT 51.38 2.395 52.15 2.565 ;
      RECT 51.44 0.885 51.61 2.595 ;
      RECT 51.38 0.885 51.67 1.115 ;
      RECT 51.38 7.765 51.67 7.995 ;
      RECT 51.44 6.285 51.61 7.995 ;
      RECT 51.38 6.285 51.67 6.515 ;
      RECT 51.38 6.325 52.23 6.485 ;
      RECT 52.06 5.915 52.23 6.485 ;
      RECT 51.38 6.32 51.77 6.485 ;
      RECT 52 5.915 52.29 6.145 ;
      RECT 52 5.945 52.46 6.115 ;
      RECT 51.01 2.735 51.3 2.965 ;
      RECT 51.01 2.765 51.47 2.935 ;
      RECT 51.07 1.655 51.235 2.965 ;
      RECT 49.585 1.625 49.875 1.855 ;
      RECT 49.585 1.655 51.235 1.825 ;
      RECT 49.645 0.885 49.815 1.855 ;
      RECT 49.585 0.885 49.875 1.115 ;
      RECT 49.585 7.765 49.875 7.995 ;
      RECT 49.645 7.025 49.815 7.995 ;
      RECT 49.645 7.12 51.235 7.29 ;
      RECT 51.065 5.915 51.235 7.29 ;
      RECT 49.585 7.025 49.875 7.255 ;
      RECT 51.01 5.915 51.3 6.145 ;
      RECT 51.01 5.945 51.47 6.115 ;
      RECT 47.635 3.15 47.975 3.5 ;
      RECT 47.725 2.025 47.895 3.5 ;
      RECT 50.015 1.965 50.365 2.315 ;
      RECT 47.725 2.025 50.365 2.195 ;
      RECT 50.04 6.655 50.365 6.98 ;
      RECT 44.6 6.615 44.95 6.965 ;
      RECT 50.015 6.655 50.365 6.885 ;
      RECT 44.4 6.655 44.95 6.885 ;
      RECT 44.23 6.685 50.365 6.855 ;
      RECT 49.24 2.365 49.56 2.685 ;
      RECT 49.21 2.365 49.56 2.595 ;
      RECT 49.04 2.395 49.56 2.565 ;
      RECT 49.24 6.255 49.56 6.545 ;
      RECT 49.21 6.285 49.56 6.515 ;
      RECT 49.04 6.315 49.56 6.485 ;
      RECT 48.2 2.705 48.54 3.055 ;
      RECT 48.2 2.765 48.675 2.935 ;
      RECT 48.19 5.845 48.53 6.195 ;
      RECT 42.6 5.915 42.89 6.145 ;
      RECT 42.6 5.945 48.675 6.115 ;
      RECT 44.69 3.57 45.01 3.83 ;
      RECT 45.98 2.745 46.12 3.605 ;
      RECT 44.78 3.465 46.12 3.605 ;
      RECT 44.78 3.025 44.92 3.83 ;
      RECT 44.705 3.025 44.995 3.255 ;
      RECT 45.905 2.745 46.195 2.975 ;
      RECT 45.425 3.025 45.715 3.255 ;
      RECT 45.62 1.95 45.76 3.21 ;
      RECT 45.65 1.89 45.97 2.15 ;
      RECT 42.25 2.45 42.57 2.71 ;
      RECT 44.945 2.465 45.235 2.695 ;
      RECT 42.34 2.37 45.16 2.51 ;
      RECT 44.21 1.89 44.53 2.15 ;
      RECT 44.705 1.905 44.995 2.135 ;
      RECT 44.21 1.95 44.995 2.09 ;
      RECT 44.21 3.01 44.53 3.27 ;
      RECT 44.21 2.79 44.44 3.27 ;
      RECT 43.705 2.745 43.995 2.975 ;
      RECT 43.705 2.79 44.44 2.93 ;
      RECT 43.97 7.765 44.26 7.995 ;
      RECT 44.03 7.025 44.2 7.995 ;
      RECT 43.93 7.055 44.31 7.425 ;
      RECT 43.97 7.025 44.26 7.425 ;
      RECT 42.73 3.57 43.05 3.83 ;
      RECT 42.265 3.585 42.555 3.815 ;
      RECT 42.265 3.63 43.05 3.77 ;
      RECT 41.025 2.465 41.315 2.695 ;
      RECT 41.025 2.51 41.96 2.65 ;
      RECT 41.82 1.95 41.96 2.65 ;
      RECT 42.49 1.89 42.81 2.15 ;
      RECT 42.265 1.905 42.81 2.135 ;
      RECT 41.82 1.95 42.81 2.09 ;
      RECT 40.17 3.57 40.49 3.83 ;
      RECT 40.17 3.63 41.24 3.77 ;
      RECT 41.1 3.07 41.24 3.77 ;
      RECT 42.265 3.025 42.555 3.255 ;
      RECT 41.1 3.07 42.555 3.21 ;
      RECT 40.53 1.89 40.85 2.15 ;
      RECT 40.305 1.905 40.85 2.135 ;
      RECT 39.55 2.45 39.87 2.71 ;
      RECT 40.545 2.465 40.835 2.695 ;
      RECT 39.305 2.465 39.87 2.695 ;
      RECT 39.305 2.51 40.835 2.65 ;
      RECT 38.825 3.025 39.115 3.255 ;
      RECT 39.02 1.95 39.16 3.21 ;
      RECT 39.81 1.89 40.13 2.15 ;
      RECT 38.825 1.905 39.115 2.135 ;
      RECT 38.825 1.95 40.13 2.09 ;
      RECT 38.42 3.465 39.52 3.605 ;
      RECT 39.305 3.305 39.595 3.535 ;
      RECT 38.345 3.305 38.635 3.535 ;
      RECT 38.585 2.37 38.875 2.74 ;
      RECT 37.82 2.37 38.875 2.51 ;
      RECT 38.33 1.89 38.65 2.15 ;
      RECT 36.37 1.89 36.69 2.15 ;
      RECT 36.37 1.95 38.65 2.09 ;
      RECT 37.49 3.01 37.81 3.27 ;
      RECT 37.49 3.01 38.32 3.15 ;
      RECT 38.105 2.745 38.32 3.15 ;
      RECT 38.105 2.745 38.395 2.975 ;
      RECT 35.89 2.45 36.21 2.71 ;
      RECT 37.3 2.465 37.59 2.695 ;
      RECT 35.89 2.465 36.435 2.695 ;
      RECT 35.89 2.55 36.84 2.69 ;
      RECT 36.7 2.37 36.84 2.69 ;
      RECT 37.2 2.465 37.59 2.65 ;
      RECT 36.7 2.37 37.34 2.51 ;
      RECT 35.41 3.26 35.73 3.675 ;
      RECT 35.49 1.905 35.645 3.675 ;
      RECT 35.425 1.905 35.715 2.135 ;
      RECT 33.81 7.765 34.1 7.995 ;
      RECT 33.87 6.285 34.04 7.995 ;
      RECT 33.855 6.66 34.21 7.015 ;
      RECT 33.81 6.285 34.1 6.515 ;
      RECT 33.81 2.365 34.1 2.595 ;
      RECT 33.87 0.885 34.04 2.595 ;
      RECT 33.81 0.885 34.1 1.115 ;
      RECT 33.4 2.735 33.73 2.965 ;
      RECT 33.4 2.765 33.9 2.935 ;
      RECT 33.4 2.395 33.59 2.965 ;
      RECT 32.82 2.365 33.11 2.595 ;
      RECT 32.82 2.395 33.59 2.565 ;
      RECT 32.88 0.885 33.05 2.595 ;
      RECT 32.82 0.885 33.11 1.115 ;
      RECT 32.82 7.765 33.11 7.995 ;
      RECT 32.88 6.285 33.05 7.995 ;
      RECT 32.82 6.285 33.11 6.515 ;
      RECT 32.82 6.325 33.67 6.485 ;
      RECT 33.5 5.915 33.67 6.485 ;
      RECT 32.82 6.32 33.21 6.485 ;
      RECT 33.44 5.915 33.73 6.145 ;
      RECT 33.44 5.945 33.9 6.115 ;
      RECT 32.45 2.735 32.74 2.965 ;
      RECT 32.45 2.765 32.91 2.935 ;
      RECT 32.51 1.655 32.675 2.965 ;
      RECT 31.025 1.625 31.315 1.855 ;
      RECT 31.025 1.655 32.675 1.825 ;
      RECT 31.085 0.885 31.255 1.855 ;
      RECT 31.025 0.885 31.315 1.115 ;
      RECT 31.025 7.765 31.315 7.995 ;
      RECT 31.085 7.025 31.255 7.995 ;
      RECT 31.085 7.12 32.675 7.29 ;
      RECT 32.505 5.915 32.675 7.29 ;
      RECT 31.025 7.025 31.315 7.255 ;
      RECT 32.45 5.915 32.74 6.145 ;
      RECT 32.45 5.945 32.91 6.115 ;
      RECT 29.075 3.15 29.415 3.5 ;
      RECT 29.165 2.025 29.335 3.5 ;
      RECT 31.455 1.965 31.805 2.315 ;
      RECT 29.165 2.025 31.805 2.195 ;
      RECT 31.48 6.655 31.805 6.98 ;
      RECT 26.045 6.61 26.395 6.96 ;
      RECT 31.455 6.655 31.805 6.885 ;
      RECT 25.84 6.655 26.395 6.885 ;
      RECT 25.67 6.685 31.805 6.855 ;
      RECT 30.68 2.365 31 2.685 ;
      RECT 30.65 2.365 31 2.595 ;
      RECT 30.48 2.395 31 2.565 ;
      RECT 30.68 6.255 31 6.545 ;
      RECT 30.65 6.285 31 6.515 ;
      RECT 30.48 6.315 31 6.485 ;
      RECT 29.64 2.705 29.98 3.055 ;
      RECT 29.64 2.765 30.115 2.935 ;
      RECT 29.63 5.845 29.97 6.195 ;
      RECT 24.04 5.915 24.33 6.145 ;
      RECT 24.04 5.945 30.115 6.115 ;
      RECT 26.13 3.57 26.45 3.83 ;
      RECT 27.42 2.745 27.56 3.605 ;
      RECT 26.22 3.465 27.56 3.605 ;
      RECT 26.22 3.025 26.36 3.83 ;
      RECT 26.145 3.025 26.435 3.255 ;
      RECT 27.345 2.745 27.635 2.975 ;
      RECT 26.865 3.025 27.155 3.255 ;
      RECT 27.06 1.95 27.2 3.21 ;
      RECT 27.09 1.89 27.41 2.15 ;
      RECT 23.69 2.45 24.01 2.71 ;
      RECT 26.385 2.465 26.675 2.695 ;
      RECT 23.78 2.37 26.6 2.51 ;
      RECT 25.65 1.89 25.97 2.15 ;
      RECT 26.145 1.905 26.435 2.135 ;
      RECT 25.65 1.95 26.435 2.09 ;
      RECT 25.65 3.01 25.97 3.27 ;
      RECT 25.65 2.79 25.88 3.27 ;
      RECT 25.145 2.745 25.435 2.975 ;
      RECT 25.145 2.79 25.88 2.93 ;
      RECT 25.41 7.765 25.7 7.995 ;
      RECT 25.47 7.025 25.64 7.995 ;
      RECT 25.37 7.055 25.75 7.425 ;
      RECT 25.41 7.025 25.7 7.425 ;
      RECT 24.17 3.57 24.49 3.83 ;
      RECT 23.705 3.585 23.995 3.815 ;
      RECT 23.705 3.63 24.49 3.77 ;
      RECT 22.465 2.465 22.755 2.695 ;
      RECT 22.465 2.51 23.4 2.65 ;
      RECT 23.26 1.95 23.4 2.65 ;
      RECT 23.93 1.89 24.25 2.15 ;
      RECT 23.705 1.905 24.25 2.135 ;
      RECT 23.26 1.95 24.25 2.09 ;
      RECT 21.61 3.57 21.93 3.83 ;
      RECT 21.61 3.63 22.68 3.77 ;
      RECT 22.54 3.07 22.68 3.77 ;
      RECT 23.705 3.025 23.995 3.255 ;
      RECT 22.54 3.07 23.995 3.21 ;
      RECT 21.97 1.89 22.29 2.15 ;
      RECT 21.745 1.905 22.29 2.135 ;
      RECT 20.99 2.45 21.31 2.71 ;
      RECT 21.985 2.465 22.275 2.695 ;
      RECT 20.745 2.465 21.31 2.695 ;
      RECT 20.745 2.51 22.275 2.65 ;
      RECT 20.265 3.025 20.555 3.255 ;
      RECT 20.46 1.95 20.6 3.21 ;
      RECT 21.25 1.89 21.57 2.15 ;
      RECT 20.265 1.905 20.555 2.135 ;
      RECT 20.265 1.95 21.57 2.09 ;
      RECT 19.86 3.465 20.96 3.605 ;
      RECT 20.745 3.305 21.035 3.535 ;
      RECT 19.785 3.305 20.075 3.535 ;
      RECT 20.025 2.37 20.315 2.74 ;
      RECT 19.26 2.37 20.315 2.51 ;
      RECT 19.77 1.89 20.09 2.15 ;
      RECT 17.81 1.89 18.13 2.15 ;
      RECT 17.81 1.95 20.09 2.09 ;
      RECT 18.93 3.01 19.25 3.27 ;
      RECT 18.93 3.01 19.76 3.15 ;
      RECT 19.545 2.745 19.76 3.15 ;
      RECT 19.545 2.745 19.835 2.975 ;
      RECT 17.33 2.45 17.65 2.71 ;
      RECT 18.74 2.465 19.03 2.695 ;
      RECT 17.33 2.465 17.875 2.695 ;
      RECT 17.33 2.55 18.28 2.69 ;
      RECT 18.14 2.37 18.28 2.69 ;
      RECT 18.64 2.465 19.03 2.65 ;
      RECT 18.14 2.37 18.78 2.51 ;
      RECT 16.85 3.26 17.17 3.675 ;
      RECT 16.93 1.905 17.085 3.675 ;
      RECT 16.865 1.905 17.155 2.135 ;
      RECT 15.25 7.765 15.54 7.995 ;
      RECT 15.31 6.285 15.48 7.995 ;
      RECT 15.3 6.655 15.65 7.005 ;
      RECT 15.25 6.285 15.54 6.515 ;
      RECT 15.25 2.365 15.54 2.595 ;
      RECT 15.31 0.885 15.48 2.595 ;
      RECT 15.25 0.885 15.54 1.115 ;
      RECT 14.84 2.735 15.17 2.965 ;
      RECT 14.84 2.765 15.34 2.935 ;
      RECT 14.84 2.395 15.03 2.965 ;
      RECT 14.26 2.365 14.55 2.595 ;
      RECT 14.26 2.395 15.03 2.565 ;
      RECT 14.32 0.885 14.49 2.595 ;
      RECT 14.26 0.885 14.55 1.115 ;
      RECT 14.26 7.765 14.55 7.995 ;
      RECT 14.32 6.285 14.49 7.995 ;
      RECT 14.26 6.285 14.55 6.515 ;
      RECT 14.26 6.325 15.11 6.485 ;
      RECT 14.94 5.915 15.11 6.485 ;
      RECT 14.26 6.32 14.65 6.485 ;
      RECT 14.88 5.915 15.17 6.145 ;
      RECT 14.88 5.945 15.34 6.115 ;
      RECT 13.89 2.735 14.18 2.965 ;
      RECT 13.89 2.765 14.35 2.935 ;
      RECT 13.95 1.655 14.115 2.965 ;
      RECT 12.465 1.625 12.755 1.855 ;
      RECT 12.465 1.655 14.115 1.825 ;
      RECT 12.525 0.885 12.695 1.855 ;
      RECT 12.465 0.885 12.755 1.115 ;
      RECT 12.465 7.765 12.755 7.995 ;
      RECT 12.525 7.025 12.695 7.995 ;
      RECT 12.525 7.12 14.115 7.29 ;
      RECT 13.945 5.915 14.115 7.29 ;
      RECT 12.465 7.025 12.755 7.255 ;
      RECT 13.89 5.915 14.18 6.145 ;
      RECT 13.89 5.945 14.35 6.115 ;
      RECT 10.515 3.15 10.855 3.5 ;
      RECT 10.605 2.025 10.775 3.5 ;
      RECT 12.895 1.965 13.245 2.315 ;
      RECT 10.605 2.025 13.245 2.195 ;
      RECT 12.92 6.655 13.245 6.98 ;
      RECT 7.485 6.605 7.835 6.955 ;
      RECT 12.895 6.655 13.245 6.885 ;
      RECT 7.28 6.655 7.835 6.885 ;
      RECT 7.11 6.685 13.245 6.855 ;
      RECT 12.12 2.365 12.44 2.685 ;
      RECT 12.09 2.365 12.44 2.595 ;
      RECT 11.92 2.395 12.44 2.565 ;
      RECT 12.12 6.255 12.44 6.545 ;
      RECT 12.09 6.285 12.44 6.515 ;
      RECT 11.92 6.315 12.44 6.485 ;
      RECT 11.08 2.705 11.42 3.055 ;
      RECT 11.08 2.765 11.555 2.935 ;
      RECT 11.07 5.845 11.41 6.195 ;
      RECT 5.48 5.915 5.77 6.145 ;
      RECT 5.48 5.945 11.555 6.115 ;
      RECT 7.57 3.57 7.89 3.83 ;
      RECT 8.86 2.745 9 3.605 ;
      RECT 7.66 3.465 9 3.605 ;
      RECT 7.66 3.025 7.8 3.83 ;
      RECT 7.585 3.025 7.875 3.255 ;
      RECT 8.785 2.745 9.075 2.975 ;
      RECT 8.305 3.025 8.595 3.255 ;
      RECT 8.5 1.95 8.64 3.21 ;
      RECT 8.53 1.89 8.85 2.15 ;
      RECT 5.13 2.45 5.45 2.71 ;
      RECT 7.825 2.465 8.115 2.695 ;
      RECT 5.22 2.37 8.04 2.51 ;
      RECT 7.09 1.89 7.41 2.15 ;
      RECT 7.585 1.905 7.875 2.135 ;
      RECT 7.09 1.95 7.875 2.09 ;
      RECT 7.09 3.01 7.41 3.27 ;
      RECT 7.09 2.79 7.32 3.27 ;
      RECT 6.585 2.745 6.875 2.975 ;
      RECT 6.585 2.79 7.32 2.93 ;
      RECT 6.85 7.765 7.14 7.995 ;
      RECT 6.91 7.025 7.08 7.995 ;
      RECT 6.81 7.055 7.19 7.425 ;
      RECT 6.85 7.025 7.14 7.425 ;
      RECT 5.61 3.57 5.93 3.83 ;
      RECT 5.145 3.585 5.435 3.815 ;
      RECT 5.145 3.63 5.93 3.77 ;
      RECT 3.905 2.465 4.195 2.695 ;
      RECT 3.905 2.51 4.84 2.65 ;
      RECT 4.7 1.95 4.84 2.65 ;
      RECT 5.37 1.89 5.69 2.15 ;
      RECT 5.145 1.905 5.69 2.135 ;
      RECT 4.7 1.95 5.69 2.09 ;
      RECT 3.05 3.57 3.37 3.83 ;
      RECT 3.05 3.63 4.12 3.77 ;
      RECT 3.98 3.07 4.12 3.77 ;
      RECT 5.145 3.025 5.435 3.255 ;
      RECT 3.98 3.07 5.435 3.21 ;
      RECT 3.41 1.89 3.73 2.15 ;
      RECT 3.185 1.905 3.73 2.135 ;
      RECT 2.43 2.45 2.75 2.71 ;
      RECT 3.425 2.465 3.715 2.695 ;
      RECT 2.185 2.465 2.75 2.695 ;
      RECT 2.185 2.51 3.715 2.65 ;
      RECT 1.705 3.025 1.995 3.255 ;
      RECT 1.9 1.95 2.04 3.21 ;
      RECT 2.69 1.89 3.01 2.15 ;
      RECT 1.705 1.905 1.995 2.135 ;
      RECT 1.705 1.95 3.01 2.09 ;
      RECT 1.3 3.465 2.4 3.605 ;
      RECT 2.185 3.305 2.475 3.535 ;
      RECT 1.225 3.305 1.515 3.535 ;
      RECT 1.465 2.37 1.755 2.74 ;
      RECT 0.7 2.37 1.755 2.51 ;
      RECT 1.21 1.89 1.53 2.15 ;
      RECT -0.75 1.89 -0.43 2.15 ;
      RECT -0.75 1.95 1.53 2.09 ;
      RECT 0.37 3.01 0.69 3.27 ;
      RECT 0.37 3.01 1.2 3.15 ;
      RECT 0.985 2.745 1.2 3.15 ;
      RECT 0.985 2.745 1.275 2.975 ;
      RECT -1.23 2.45 -0.91 2.71 ;
      RECT 0.18 2.465 0.47 2.695 ;
      RECT -1.23 2.465 -0.685 2.695 ;
      RECT -1.23 2.55 -0.28 2.69 ;
      RECT -0.42 2.37 -0.28 2.69 ;
      RECT 0.08 2.465 0.47 2.65 ;
      RECT -0.42 2.37 0.22 2.51 ;
      RECT -1.71 3.26 -1.39 3.675 ;
      RECT -1.63 1.905 -1.475 3.675 ;
      RECT -1.695 1.905 -1.405 2.135 ;
      RECT -3.535 6.655 -3.245 6.885 ;
      RECT -3.705 6.685 -3.245 6.855 ;
      RECT -3.965 7.765 -3.675 7.995 ;
      RECT -3.905 7.025 -3.735 7.995 ;
      RECT -3.995 7.025 -3.645 7.315 ;
      RECT -4.37 6.285 -4.02 6.575 ;
      RECT -4.51 6.315 -4.02 6.485 ;
      RECT -5.335 5.915 -5.045 6.145 ;
      RECT -5.335 5.945 -4.875 6.115 ;
      RECT 80.81 3.57 81.13 3.83 ;
      RECT 80.21 1.89 80.89 2.15 ;
      RECT 80.33 3.57 80.65 3.83 ;
      RECT 78.85 3.57 79.17 3.83 ;
      RECT 78.37 1.89 78.69 2.15 ;
      RECT 77.65 3.01 77.97 3.27 ;
      RECT 76.93 3.01 77.25 3.27 ;
      RECT 73.97 3.01 74.29 3.27 ;
      RECT 73.49 3.01 73.81 3.27 ;
      RECT 62.25 3.57 62.57 3.83 ;
      RECT 61.65 1.89 62.33 2.15 ;
      RECT 61.77 3.57 62.09 3.83 ;
      RECT 60.29 3.57 60.61 3.83 ;
      RECT 59.81 1.89 60.13 2.15 ;
      RECT 59.09 3.01 59.41 3.27 ;
      RECT 58.37 3.01 58.69 3.27 ;
      RECT 55.41 3.01 55.73 3.27 ;
      RECT 54.93 3.01 55.25 3.27 ;
      RECT 43.69 3.57 44.01 3.83 ;
      RECT 43.09 1.89 43.77 2.15 ;
      RECT 43.21 3.57 43.53 3.83 ;
      RECT 41.73 3.57 42.05 3.83 ;
      RECT 41.25 1.89 41.57 2.15 ;
      RECT 40.53 3.01 40.85 3.27 ;
      RECT 39.81 3.01 40.13 3.27 ;
      RECT 36.85 3.01 37.17 3.27 ;
      RECT 36.37 3.01 36.69 3.27 ;
      RECT 25.13 3.57 25.45 3.83 ;
      RECT 24.53 1.89 25.21 2.15 ;
      RECT 24.65 3.57 24.97 3.83 ;
      RECT 23.17 3.57 23.49 3.83 ;
      RECT 22.69 1.89 23.01 2.15 ;
      RECT 21.97 3.01 22.29 3.27 ;
      RECT 21.25 3.01 21.57 3.27 ;
      RECT 18.29 3.01 18.61 3.27 ;
      RECT 17.81 3.01 18.13 3.27 ;
      RECT 6.57 3.57 6.89 3.83 ;
      RECT 5.97 1.89 6.65 2.15 ;
      RECT 6.09 3.57 6.41 3.83 ;
      RECT 4.61 3.57 4.93 3.83 ;
      RECT 4.13 1.89 4.45 2.15 ;
      RECT 3.41 3.01 3.73 3.27 ;
      RECT 2.69 3.01 3.01 3.27 ;
      RECT -0.27 3.01 0.05 3.27 ;
      RECT -0.75 3.01 -0.43 3.27 ;
    LAYER mcon ;
      RECT 89.55 0.915 89.72 1.085 ;
      RECT 89.55 2.395 89.72 2.565 ;
      RECT 89.55 6.315 89.72 6.485 ;
      RECT 89.55 7.795 89.72 7.965 ;
      RECT 89.2 0.105 89.37 0.275 ;
      RECT 89.2 4.165 89.37 4.335 ;
      RECT 89.2 4.545 89.37 4.715 ;
      RECT 89.2 8.605 89.37 8.775 ;
      RECT 89.18 2.765 89.35 2.935 ;
      RECT 89.18 5.945 89.35 6.115 ;
      RECT 88.56 0.915 88.73 1.085 ;
      RECT 88.56 2.395 88.73 2.565 ;
      RECT 88.56 6.315 88.73 6.485 ;
      RECT 88.56 7.795 88.73 7.965 ;
      RECT 88.21 0.105 88.38 0.275 ;
      RECT 88.21 4.165 88.38 4.335 ;
      RECT 88.21 4.545 88.38 4.715 ;
      RECT 88.21 8.605 88.38 8.775 ;
      RECT 88.19 2.765 88.36 2.935 ;
      RECT 88.19 5.945 88.36 6.115 ;
      RECT 87.505 0.105 87.675 0.275 ;
      RECT 87.505 4.165 87.675 4.335 ;
      RECT 87.505 4.545 87.675 4.715 ;
      RECT 87.505 8.605 87.675 8.775 ;
      RECT 87.195 2.025 87.365 2.195 ;
      RECT 87.195 6.685 87.365 6.855 ;
      RECT 86.825 0.105 86.995 0.275 ;
      RECT 86.825 8.605 86.995 8.775 ;
      RECT 86.765 0.915 86.935 1.085 ;
      RECT 86.765 1.655 86.935 1.825 ;
      RECT 86.765 7.055 86.935 7.225 ;
      RECT 86.765 7.795 86.935 7.965 ;
      RECT 86.39 2.395 86.56 2.565 ;
      RECT 86.39 6.315 86.56 6.485 ;
      RECT 86.145 0.105 86.315 0.275 ;
      RECT 86.145 8.605 86.315 8.775 ;
      RECT 85.465 0.105 85.635 0.275 ;
      RECT 85.465 8.605 85.635 8.775 ;
      RECT 85.395 2.765 85.565 2.935 ;
      RECT 85.395 5.945 85.565 6.115 ;
      RECT 83.92 1.415 84.09 1.585 ;
      RECT 83.92 4.135 84.09 4.305 ;
      RECT 83.46 1.415 83.63 1.585 ;
      RECT 83.46 4.135 83.63 4.305 ;
      RECT 83.085 2.775 83.255 2.945 ;
      RECT 83 1.415 83.17 1.585 ;
      RECT 83 4.135 83.17 4.305 ;
      RECT 82.845 1.935 83.015 2.105 ;
      RECT 82.605 3.055 82.775 3.225 ;
      RECT 82.54 1.415 82.71 1.585 ;
      RECT 82.54 4.135 82.71 4.305 ;
      RECT 82.125 2.495 82.295 2.665 ;
      RECT 82.08 1.415 82.25 1.585 ;
      RECT 82.08 4.135 82.25 4.305 ;
      RECT 81.89 4.545 82.06 4.715 ;
      RECT 81.89 8.605 82.06 8.775 ;
      RECT 81.885 1.935 82.055 2.105 ;
      RECT 81.885 3.055 82.055 3.225 ;
      RECT 81.885 3.615 82.055 3.785 ;
      RECT 81.62 1.415 81.79 1.585 ;
      RECT 81.62 4.135 81.79 4.305 ;
      RECT 81.58 6.685 81.75 6.855 ;
      RECT 81.405 3.055 81.575 3.225 ;
      RECT 81.21 8.605 81.38 8.775 ;
      RECT 81.16 1.415 81.33 1.585 ;
      RECT 81.16 4.135 81.33 4.305 ;
      RECT 81.15 7.055 81.32 7.225 ;
      RECT 81.15 7.795 81.32 7.965 ;
      RECT 80.885 2.775 81.055 2.945 ;
      RECT 80.885 3.615 81.055 3.785 ;
      RECT 80.775 6.315 80.945 6.485 ;
      RECT 80.7 1.415 80.87 1.585 ;
      RECT 80.7 4.135 80.87 4.305 ;
      RECT 80.53 8.605 80.7 8.775 ;
      RECT 80.405 1.935 80.575 2.105 ;
      RECT 80.405 3.615 80.575 3.785 ;
      RECT 80.24 1.415 80.41 1.585 ;
      RECT 80.24 4.135 80.41 4.305 ;
      RECT 79.85 8.605 80.02 8.775 ;
      RECT 79.78 1.415 79.95 1.585 ;
      RECT 79.78 4.135 79.95 4.305 ;
      RECT 79.78 5.945 79.95 6.115 ;
      RECT 79.445 1.935 79.615 2.105 ;
      RECT 79.445 2.495 79.615 2.665 ;
      RECT 79.445 3.055 79.615 3.225 ;
      RECT 79.445 3.615 79.615 3.785 ;
      RECT 79.32 1.415 79.49 1.585 ;
      RECT 79.32 4.135 79.49 4.305 ;
      RECT 78.925 3.615 79.095 3.785 ;
      RECT 78.86 1.415 79.03 1.585 ;
      RECT 78.86 4.135 79.03 4.305 ;
      RECT 78.445 1.935 78.615 2.105 ;
      RECT 78.4 1.415 78.57 1.585 ;
      RECT 78.4 4.135 78.57 4.305 ;
      RECT 78.205 2.495 78.375 2.665 ;
      RECT 77.94 1.415 78.11 1.585 ;
      RECT 77.94 4.135 78.11 4.305 ;
      RECT 77.725 2.495 77.895 2.665 ;
      RECT 77.725 3.055 77.895 3.225 ;
      RECT 77.485 1.935 77.655 2.105 ;
      RECT 77.48 1.415 77.65 1.585 ;
      RECT 77.48 4.135 77.65 4.305 ;
      RECT 77.02 1.415 77.19 1.585 ;
      RECT 77.02 4.135 77.19 4.305 ;
      RECT 77.005 3.055 77.175 3.225 ;
      RECT 76.56 1.415 76.73 1.585 ;
      RECT 76.56 4.135 76.73 4.305 ;
      RECT 76.485 2.495 76.655 2.665 ;
      RECT 76.485 3.335 76.655 3.505 ;
      RECT 76.1 1.415 76.27 1.585 ;
      RECT 76.1 4.135 76.27 4.305 ;
      RECT 76.005 1.935 76.175 2.105 ;
      RECT 76.005 3.055 76.175 3.225 ;
      RECT 75.765 2.495 75.935 2.665 ;
      RECT 75.64 1.415 75.81 1.585 ;
      RECT 75.64 4.135 75.81 4.305 ;
      RECT 75.525 3.335 75.695 3.505 ;
      RECT 75.285 2.775 75.455 2.945 ;
      RECT 75.18 1.415 75.35 1.585 ;
      RECT 75.18 4.135 75.35 4.305 ;
      RECT 74.72 1.415 74.89 1.585 ;
      RECT 74.72 4.135 74.89 4.305 ;
      RECT 74.48 2.495 74.65 2.665 ;
      RECT 74.26 1.415 74.43 1.585 ;
      RECT 74.26 4.135 74.43 4.305 ;
      RECT 74.045 3.055 74.215 3.225 ;
      RECT 73.8 1.415 73.97 1.585 ;
      RECT 73.8 4.135 73.97 4.305 ;
      RECT 73.565 1.935 73.735 2.105 ;
      RECT 73.565 3.055 73.735 3.225 ;
      RECT 73.34 1.415 73.51 1.585 ;
      RECT 73.34 4.135 73.51 4.305 ;
      RECT 73.325 2.495 73.495 2.665 ;
      RECT 72.88 1.415 73.05 1.585 ;
      RECT 72.88 4.135 73.05 4.305 ;
      RECT 72.605 1.935 72.775 2.105 ;
      RECT 72.605 3.475 72.775 3.645 ;
      RECT 72.42 1.415 72.59 1.585 ;
      RECT 72.42 4.135 72.59 4.305 ;
      RECT 70.99 0.915 71.16 1.085 ;
      RECT 70.99 2.395 71.16 2.565 ;
      RECT 70.99 6.315 71.16 6.485 ;
      RECT 70.99 7.795 71.16 7.965 ;
      RECT 70.64 0.105 70.81 0.275 ;
      RECT 70.64 4.165 70.81 4.335 ;
      RECT 70.64 4.545 70.81 4.715 ;
      RECT 70.64 8.605 70.81 8.775 ;
      RECT 70.62 2.765 70.79 2.935 ;
      RECT 70.62 5.945 70.79 6.115 ;
      RECT 70 0.915 70.17 1.085 ;
      RECT 70 2.395 70.17 2.565 ;
      RECT 70 6.315 70.17 6.485 ;
      RECT 70 7.795 70.17 7.965 ;
      RECT 69.65 0.105 69.82 0.275 ;
      RECT 69.65 4.165 69.82 4.335 ;
      RECT 69.65 4.545 69.82 4.715 ;
      RECT 69.65 8.605 69.82 8.775 ;
      RECT 69.63 2.765 69.8 2.935 ;
      RECT 69.63 5.945 69.8 6.115 ;
      RECT 68.945 0.105 69.115 0.275 ;
      RECT 68.945 4.165 69.115 4.335 ;
      RECT 68.945 4.545 69.115 4.715 ;
      RECT 68.945 8.605 69.115 8.775 ;
      RECT 68.635 2.025 68.805 2.195 ;
      RECT 68.635 6.685 68.805 6.855 ;
      RECT 68.265 0.105 68.435 0.275 ;
      RECT 68.265 8.605 68.435 8.775 ;
      RECT 68.205 0.915 68.375 1.085 ;
      RECT 68.205 1.655 68.375 1.825 ;
      RECT 68.205 7.055 68.375 7.225 ;
      RECT 68.205 7.795 68.375 7.965 ;
      RECT 67.83 2.395 68 2.565 ;
      RECT 67.83 6.315 68 6.485 ;
      RECT 67.585 0.105 67.755 0.275 ;
      RECT 67.585 8.605 67.755 8.775 ;
      RECT 66.905 0.105 67.075 0.275 ;
      RECT 66.905 8.605 67.075 8.775 ;
      RECT 66.835 2.765 67.005 2.935 ;
      RECT 66.835 5.945 67.005 6.115 ;
      RECT 65.36 1.415 65.53 1.585 ;
      RECT 65.36 4.135 65.53 4.305 ;
      RECT 64.9 1.415 65.07 1.585 ;
      RECT 64.9 4.135 65.07 4.305 ;
      RECT 64.525 2.775 64.695 2.945 ;
      RECT 64.44 1.415 64.61 1.585 ;
      RECT 64.44 4.135 64.61 4.305 ;
      RECT 64.285 1.935 64.455 2.105 ;
      RECT 64.045 3.055 64.215 3.225 ;
      RECT 63.98 1.415 64.15 1.585 ;
      RECT 63.98 4.135 64.15 4.305 ;
      RECT 63.565 2.495 63.735 2.665 ;
      RECT 63.52 1.415 63.69 1.585 ;
      RECT 63.52 4.135 63.69 4.305 ;
      RECT 63.33 4.545 63.5 4.715 ;
      RECT 63.33 8.605 63.5 8.775 ;
      RECT 63.325 1.935 63.495 2.105 ;
      RECT 63.325 3.055 63.495 3.225 ;
      RECT 63.325 3.615 63.495 3.785 ;
      RECT 63.06 1.415 63.23 1.585 ;
      RECT 63.06 4.135 63.23 4.305 ;
      RECT 63.02 6.685 63.19 6.855 ;
      RECT 62.845 3.055 63.015 3.225 ;
      RECT 62.65 8.605 62.82 8.775 ;
      RECT 62.6 1.415 62.77 1.585 ;
      RECT 62.6 4.135 62.77 4.305 ;
      RECT 62.59 7.055 62.76 7.225 ;
      RECT 62.59 7.795 62.76 7.965 ;
      RECT 62.325 2.775 62.495 2.945 ;
      RECT 62.325 3.615 62.495 3.785 ;
      RECT 62.215 6.315 62.385 6.485 ;
      RECT 62.14 1.415 62.31 1.585 ;
      RECT 62.14 4.135 62.31 4.305 ;
      RECT 61.97 8.605 62.14 8.775 ;
      RECT 61.845 1.935 62.015 2.105 ;
      RECT 61.845 3.615 62.015 3.785 ;
      RECT 61.68 1.415 61.85 1.585 ;
      RECT 61.68 4.135 61.85 4.305 ;
      RECT 61.29 8.605 61.46 8.775 ;
      RECT 61.22 1.415 61.39 1.585 ;
      RECT 61.22 4.135 61.39 4.305 ;
      RECT 61.22 5.945 61.39 6.115 ;
      RECT 60.885 1.935 61.055 2.105 ;
      RECT 60.885 2.495 61.055 2.665 ;
      RECT 60.885 3.055 61.055 3.225 ;
      RECT 60.885 3.615 61.055 3.785 ;
      RECT 60.76 1.415 60.93 1.585 ;
      RECT 60.76 4.135 60.93 4.305 ;
      RECT 60.365 3.615 60.535 3.785 ;
      RECT 60.3 1.415 60.47 1.585 ;
      RECT 60.3 4.135 60.47 4.305 ;
      RECT 59.885 1.935 60.055 2.105 ;
      RECT 59.84 1.415 60.01 1.585 ;
      RECT 59.84 4.135 60.01 4.305 ;
      RECT 59.645 2.495 59.815 2.665 ;
      RECT 59.38 1.415 59.55 1.585 ;
      RECT 59.38 4.135 59.55 4.305 ;
      RECT 59.165 2.495 59.335 2.665 ;
      RECT 59.165 3.055 59.335 3.225 ;
      RECT 58.925 1.935 59.095 2.105 ;
      RECT 58.92 1.415 59.09 1.585 ;
      RECT 58.92 4.135 59.09 4.305 ;
      RECT 58.46 1.415 58.63 1.585 ;
      RECT 58.46 4.135 58.63 4.305 ;
      RECT 58.445 3.055 58.615 3.225 ;
      RECT 58 1.415 58.17 1.585 ;
      RECT 58 4.135 58.17 4.305 ;
      RECT 57.925 2.495 58.095 2.665 ;
      RECT 57.925 3.335 58.095 3.505 ;
      RECT 57.54 1.415 57.71 1.585 ;
      RECT 57.54 4.135 57.71 4.305 ;
      RECT 57.445 1.935 57.615 2.105 ;
      RECT 57.445 3.055 57.615 3.225 ;
      RECT 57.205 2.495 57.375 2.665 ;
      RECT 57.08 1.415 57.25 1.585 ;
      RECT 57.08 4.135 57.25 4.305 ;
      RECT 56.965 3.335 57.135 3.505 ;
      RECT 56.725 2.775 56.895 2.945 ;
      RECT 56.62 1.415 56.79 1.585 ;
      RECT 56.62 4.135 56.79 4.305 ;
      RECT 56.16 1.415 56.33 1.585 ;
      RECT 56.16 4.135 56.33 4.305 ;
      RECT 55.92 2.495 56.09 2.665 ;
      RECT 55.7 1.415 55.87 1.585 ;
      RECT 55.7 4.135 55.87 4.305 ;
      RECT 55.485 3.055 55.655 3.225 ;
      RECT 55.24 1.415 55.41 1.585 ;
      RECT 55.24 4.135 55.41 4.305 ;
      RECT 55.005 1.935 55.175 2.105 ;
      RECT 55.005 3.055 55.175 3.225 ;
      RECT 54.78 1.415 54.95 1.585 ;
      RECT 54.78 4.135 54.95 4.305 ;
      RECT 54.765 2.495 54.935 2.665 ;
      RECT 54.32 1.415 54.49 1.585 ;
      RECT 54.32 4.135 54.49 4.305 ;
      RECT 54.045 1.935 54.215 2.105 ;
      RECT 54.045 3.475 54.215 3.645 ;
      RECT 53.86 1.415 54.03 1.585 ;
      RECT 53.86 4.135 54.03 4.305 ;
      RECT 52.43 0.915 52.6 1.085 ;
      RECT 52.43 2.395 52.6 2.565 ;
      RECT 52.43 6.315 52.6 6.485 ;
      RECT 52.43 7.795 52.6 7.965 ;
      RECT 52.08 0.105 52.25 0.275 ;
      RECT 52.08 4.165 52.25 4.335 ;
      RECT 52.08 4.545 52.25 4.715 ;
      RECT 52.08 8.605 52.25 8.775 ;
      RECT 52.06 2.765 52.23 2.935 ;
      RECT 52.06 5.945 52.23 6.115 ;
      RECT 51.44 0.915 51.61 1.085 ;
      RECT 51.44 2.395 51.61 2.565 ;
      RECT 51.44 6.315 51.61 6.485 ;
      RECT 51.44 7.795 51.61 7.965 ;
      RECT 51.09 0.105 51.26 0.275 ;
      RECT 51.09 4.165 51.26 4.335 ;
      RECT 51.09 4.545 51.26 4.715 ;
      RECT 51.09 8.605 51.26 8.775 ;
      RECT 51.07 2.765 51.24 2.935 ;
      RECT 51.07 5.945 51.24 6.115 ;
      RECT 50.385 0.105 50.555 0.275 ;
      RECT 50.385 4.165 50.555 4.335 ;
      RECT 50.385 4.545 50.555 4.715 ;
      RECT 50.385 8.605 50.555 8.775 ;
      RECT 50.075 2.025 50.245 2.195 ;
      RECT 50.075 6.685 50.245 6.855 ;
      RECT 49.705 0.105 49.875 0.275 ;
      RECT 49.705 8.605 49.875 8.775 ;
      RECT 49.645 0.915 49.815 1.085 ;
      RECT 49.645 1.655 49.815 1.825 ;
      RECT 49.645 7.055 49.815 7.225 ;
      RECT 49.645 7.795 49.815 7.965 ;
      RECT 49.27 2.395 49.44 2.565 ;
      RECT 49.27 6.315 49.44 6.485 ;
      RECT 49.025 0.105 49.195 0.275 ;
      RECT 49.025 8.605 49.195 8.775 ;
      RECT 48.345 0.105 48.515 0.275 ;
      RECT 48.345 8.605 48.515 8.775 ;
      RECT 48.275 2.765 48.445 2.935 ;
      RECT 48.275 5.945 48.445 6.115 ;
      RECT 46.8 1.415 46.97 1.585 ;
      RECT 46.8 4.135 46.97 4.305 ;
      RECT 46.34 1.415 46.51 1.585 ;
      RECT 46.34 4.135 46.51 4.305 ;
      RECT 45.965 2.775 46.135 2.945 ;
      RECT 45.88 1.415 46.05 1.585 ;
      RECT 45.88 4.135 46.05 4.305 ;
      RECT 45.725 1.935 45.895 2.105 ;
      RECT 45.485 3.055 45.655 3.225 ;
      RECT 45.42 1.415 45.59 1.585 ;
      RECT 45.42 4.135 45.59 4.305 ;
      RECT 45.005 2.495 45.175 2.665 ;
      RECT 44.96 1.415 45.13 1.585 ;
      RECT 44.96 4.135 45.13 4.305 ;
      RECT 44.77 4.545 44.94 4.715 ;
      RECT 44.77 8.605 44.94 8.775 ;
      RECT 44.765 1.935 44.935 2.105 ;
      RECT 44.765 3.055 44.935 3.225 ;
      RECT 44.765 3.615 44.935 3.785 ;
      RECT 44.5 1.415 44.67 1.585 ;
      RECT 44.5 4.135 44.67 4.305 ;
      RECT 44.46 6.685 44.63 6.855 ;
      RECT 44.285 3.055 44.455 3.225 ;
      RECT 44.09 8.605 44.26 8.775 ;
      RECT 44.04 1.415 44.21 1.585 ;
      RECT 44.04 4.135 44.21 4.305 ;
      RECT 44.03 7.055 44.2 7.225 ;
      RECT 44.03 7.795 44.2 7.965 ;
      RECT 43.765 2.775 43.935 2.945 ;
      RECT 43.765 3.615 43.935 3.785 ;
      RECT 43.655 6.315 43.825 6.485 ;
      RECT 43.58 1.415 43.75 1.585 ;
      RECT 43.58 4.135 43.75 4.305 ;
      RECT 43.41 8.605 43.58 8.775 ;
      RECT 43.285 1.935 43.455 2.105 ;
      RECT 43.285 3.615 43.455 3.785 ;
      RECT 43.12 1.415 43.29 1.585 ;
      RECT 43.12 4.135 43.29 4.305 ;
      RECT 42.73 8.605 42.9 8.775 ;
      RECT 42.66 1.415 42.83 1.585 ;
      RECT 42.66 4.135 42.83 4.305 ;
      RECT 42.66 5.945 42.83 6.115 ;
      RECT 42.325 1.935 42.495 2.105 ;
      RECT 42.325 2.495 42.495 2.665 ;
      RECT 42.325 3.055 42.495 3.225 ;
      RECT 42.325 3.615 42.495 3.785 ;
      RECT 42.2 1.415 42.37 1.585 ;
      RECT 42.2 4.135 42.37 4.305 ;
      RECT 41.805 3.615 41.975 3.785 ;
      RECT 41.74 1.415 41.91 1.585 ;
      RECT 41.74 4.135 41.91 4.305 ;
      RECT 41.325 1.935 41.495 2.105 ;
      RECT 41.28 1.415 41.45 1.585 ;
      RECT 41.28 4.135 41.45 4.305 ;
      RECT 41.085 2.495 41.255 2.665 ;
      RECT 40.82 1.415 40.99 1.585 ;
      RECT 40.82 4.135 40.99 4.305 ;
      RECT 40.605 2.495 40.775 2.665 ;
      RECT 40.605 3.055 40.775 3.225 ;
      RECT 40.365 1.935 40.535 2.105 ;
      RECT 40.36 1.415 40.53 1.585 ;
      RECT 40.36 4.135 40.53 4.305 ;
      RECT 39.9 1.415 40.07 1.585 ;
      RECT 39.9 4.135 40.07 4.305 ;
      RECT 39.885 3.055 40.055 3.225 ;
      RECT 39.44 1.415 39.61 1.585 ;
      RECT 39.44 4.135 39.61 4.305 ;
      RECT 39.365 2.495 39.535 2.665 ;
      RECT 39.365 3.335 39.535 3.505 ;
      RECT 38.98 1.415 39.15 1.585 ;
      RECT 38.98 4.135 39.15 4.305 ;
      RECT 38.885 1.935 39.055 2.105 ;
      RECT 38.885 3.055 39.055 3.225 ;
      RECT 38.645 2.495 38.815 2.665 ;
      RECT 38.52 1.415 38.69 1.585 ;
      RECT 38.52 4.135 38.69 4.305 ;
      RECT 38.405 3.335 38.575 3.505 ;
      RECT 38.165 2.775 38.335 2.945 ;
      RECT 38.06 1.415 38.23 1.585 ;
      RECT 38.06 4.135 38.23 4.305 ;
      RECT 37.6 1.415 37.77 1.585 ;
      RECT 37.6 4.135 37.77 4.305 ;
      RECT 37.36 2.495 37.53 2.665 ;
      RECT 37.14 1.415 37.31 1.585 ;
      RECT 37.14 4.135 37.31 4.305 ;
      RECT 36.925 3.055 37.095 3.225 ;
      RECT 36.68 1.415 36.85 1.585 ;
      RECT 36.68 4.135 36.85 4.305 ;
      RECT 36.445 1.935 36.615 2.105 ;
      RECT 36.445 3.055 36.615 3.225 ;
      RECT 36.22 1.415 36.39 1.585 ;
      RECT 36.22 4.135 36.39 4.305 ;
      RECT 36.205 2.495 36.375 2.665 ;
      RECT 35.76 1.415 35.93 1.585 ;
      RECT 35.76 4.135 35.93 4.305 ;
      RECT 35.485 1.935 35.655 2.105 ;
      RECT 35.485 3.475 35.655 3.645 ;
      RECT 35.3 1.415 35.47 1.585 ;
      RECT 35.3 4.135 35.47 4.305 ;
      RECT 33.87 0.915 34.04 1.085 ;
      RECT 33.87 2.395 34.04 2.565 ;
      RECT 33.87 6.315 34.04 6.485 ;
      RECT 33.87 7.795 34.04 7.965 ;
      RECT 33.52 0.105 33.69 0.275 ;
      RECT 33.52 4.165 33.69 4.335 ;
      RECT 33.52 4.545 33.69 4.715 ;
      RECT 33.52 8.605 33.69 8.775 ;
      RECT 33.5 2.765 33.67 2.935 ;
      RECT 33.5 5.945 33.67 6.115 ;
      RECT 32.88 0.915 33.05 1.085 ;
      RECT 32.88 2.395 33.05 2.565 ;
      RECT 32.88 6.315 33.05 6.485 ;
      RECT 32.88 7.795 33.05 7.965 ;
      RECT 32.53 0.105 32.7 0.275 ;
      RECT 32.53 4.165 32.7 4.335 ;
      RECT 32.53 4.545 32.7 4.715 ;
      RECT 32.53 8.605 32.7 8.775 ;
      RECT 32.51 2.765 32.68 2.935 ;
      RECT 32.51 5.945 32.68 6.115 ;
      RECT 31.825 0.105 31.995 0.275 ;
      RECT 31.825 4.165 31.995 4.335 ;
      RECT 31.825 4.545 31.995 4.715 ;
      RECT 31.825 8.605 31.995 8.775 ;
      RECT 31.515 2.025 31.685 2.195 ;
      RECT 31.515 6.685 31.685 6.855 ;
      RECT 31.145 0.105 31.315 0.275 ;
      RECT 31.145 8.605 31.315 8.775 ;
      RECT 31.085 0.915 31.255 1.085 ;
      RECT 31.085 1.655 31.255 1.825 ;
      RECT 31.085 7.055 31.255 7.225 ;
      RECT 31.085 7.795 31.255 7.965 ;
      RECT 30.71 2.395 30.88 2.565 ;
      RECT 30.71 6.315 30.88 6.485 ;
      RECT 30.465 0.105 30.635 0.275 ;
      RECT 30.465 8.605 30.635 8.775 ;
      RECT 29.785 0.105 29.955 0.275 ;
      RECT 29.785 8.605 29.955 8.775 ;
      RECT 29.715 2.765 29.885 2.935 ;
      RECT 29.715 5.945 29.885 6.115 ;
      RECT 28.24 1.415 28.41 1.585 ;
      RECT 28.24 4.135 28.41 4.305 ;
      RECT 27.78 1.415 27.95 1.585 ;
      RECT 27.78 4.135 27.95 4.305 ;
      RECT 27.405 2.775 27.575 2.945 ;
      RECT 27.32 1.415 27.49 1.585 ;
      RECT 27.32 4.135 27.49 4.305 ;
      RECT 27.165 1.935 27.335 2.105 ;
      RECT 26.925 3.055 27.095 3.225 ;
      RECT 26.86 1.415 27.03 1.585 ;
      RECT 26.86 4.135 27.03 4.305 ;
      RECT 26.445 2.495 26.615 2.665 ;
      RECT 26.4 1.415 26.57 1.585 ;
      RECT 26.4 4.135 26.57 4.305 ;
      RECT 26.21 4.545 26.38 4.715 ;
      RECT 26.21 8.605 26.38 8.775 ;
      RECT 26.205 1.935 26.375 2.105 ;
      RECT 26.205 3.055 26.375 3.225 ;
      RECT 26.205 3.615 26.375 3.785 ;
      RECT 25.94 1.415 26.11 1.585 ;
      RECT 25.94 4.135 26.11 4.305 ;
      RECT 25.9 6.685 26.07 6.855 ;
      RECT 25.725 3.055 25.895 3.225 ;
      RECT 25.53 8.605 25.7 8.775 ;
      RECT 25.48 1.415 25.65 1.585 ;
      RECT 25.48 4.135 25.65 4.305 ;
      RECT 25.47 7.055 25.64 7.225 ;
      RECT 25.47 7.795 25.64 7.965 ;
      RECT 25.205 2.775 25.375 2.945 ;
      RECT 25.205 3.615 25.375 3.785 ;
      RECT 25.095 6.315 25.265 6.485 ;
      RECT 25.02 1.415 25.19 1.585 ;
      RECT 25.02 4.135 25.19 4.305 ;
      RECT 24.85 8.605 25.02 8.775 ;
      RECT 24.725 1.935 24.895 2.105 ;
      RECT 24.725 3.615 24.895 3.785 ;
      RECT 24.56 1.415 24.73 1.585 ;
      RECT 24.56 4.135 24.73 4.305 ;
      RECT 24.17 8.605 24.34 8.775 ;
      RECT 24.1 1.415 24.27 1.585 ;
      RECT 24.1 4.135 24.27 4.305 ;
      RECT 24.1 5.945 24.27 6.115 ;
      RECT 23.765 1.935 23.935 2.105 ;
      RECT 23.765 2.495 23.935 2.665 ;
      RECT 23.765 3.055 23.935 3.225 ;
      RECT 23.765 3.615 23.935 3.785 ;
      RECT 23.64 1.415 23.81 1.585 ;
      RECT 23.64 4.135 23.81 4.305 ;
      RECT 23.245 3.615 23.415 3.785 ;
      RECT 23.18 1.415 23.35 1.585 ;
      RECT 23.18 4.135 23.35 4.305 ;
      RECT 22.765 1.935 22.935 2.105 ;
      RECT 22.72 1.415 22.89 1.585 ;
      RECT 22.72 4.135 22.89 4.305 ;
      RECT 22.525 2.495 22.695 2.665 ;
      RECT 22.26 1.415 22.43 1.585 ;
      RECT 22.26 4.135 22.43 4.305 ;
      RECT 22.045 2.495 22.215 2.665 ;
      RECT 22.045 3.055 22.215 3.225 ;
      RECT 21.805 1.935 21.975 2.105 ;
      RECT 21.8 1.415 21.97 1.585 ;
      RECT 21.8 4.135 21.97 4.305 ;
      RECT 21.34 1.415 21.51 1.585 ;
      RECT 21.34 4.135 21.51 4.305 ;
      RECT 21.325 3.055 21.495 3.225 ;
      RECT 20.88 1.415 21.05 1.585 ;
      RECT 20.88 4.135 21.05 4.305 ;
      RECT 20.805 2.495 20.975 2.665 ;
      RECT 20.805 3.335 20.975 3.505 ;
      RECT 20.42 1.415 20.59 1.585 ;
      RECT 20.42 4.135 20.59 4.305 ;
      RECT 20.325 1.935 20.495 2.105 ;
      RECT 20.325 3.055 20.495 3.225 ;
      RECT 20.085 2.495 20.255 2.665 ;
      RECT 19.96 1.415 20.13 1.585 ;
      RECT 19.96 4.135 20.13 4.305 ;
      RECT 19.845 3.335 20.015 3.505 ;
      RECT 19.605 2.775 19.775 2.945 ;
      RECT 19.5 1.415 19.67 1.585 ;
      RECT 19.5 4.135 19.67 4.305 ;
      RECT 19.04 1.415 19.21 1.585 ;
      RECT 19.04 4.135 19.21 4.305 ;
      RECT 18.8 2.495 18.97 2.665 ;
      RECT 18.58 1.415 18.75 1.585 ;
      RECT 18.58 4.135 18.75 4.305 ;
      RECT 18.365 3.055 18.535 3.225 ;
      RECT 18.12 1.415 18.29 1.585 ;
      RECT 18.12 4.135 18.29 4.305 ;
      RECT 17.885 1.935 18.055 2.105 ;
      RECT 17.885 3.055 18.055 3.225 ;
      RECT 17.66 1.415 17.83 1.585 ;
      RECT 17.66 4.135 17.83 4.305 ;
      RECT 17.645 2.495 17.815 2.665 ;
      RECT 17.2 1.415 17.37 1.585 ;
      RECT 17.2 4.135 17.37 4.305 ;
      RECT 16.925 1.935 17.095 2.105 ;
      RECT 16.925 3.475 17.095 3.645 ;
      RECT 16.74 1.415 16.91 1.585 ;
      RECT 16.74 4.135 16.91 4.305 ;
      RECT 15.31 0.915 15.48 1.085 ;
      RECT 15.31 2.395 15.48 2.565 ;
      RECT 15.31 6.315 15.48 6.485 ;
      RECT 15.31 7.795 15.48 7.965 ;
      RECT 14.96 0.105 15.13 0.275 ;
      RECT 14.96 4.165 15.13 4.335 ;
      RECT 14.96 4.545 15.13 4.715 ;
      RECT 14.96 8.605 15.13 8.775 ;
      RECT 14.94 2.765 15.11 2.935 ;
      RECT 14.94 5.945 15.11 6.115 ;
      RECT 14.32 0.915 14.49 1.085 ;
      RECT 14.32 2.395 14.49 2.565 ;
      RECT 14.32 6.315 14.49 6.485 ;
      RECT 14.32 7.795 14.49 7.965 ;
      RECT 13.97 0.105 14.14 0.275 ;
      RECT 13.97 4.165 14.14 4.335 ;
      RECT 13.97 4.545 14.14 4.715 ;
      RECT 13.97 8.605 14.14 8.775 ;
      RECT 13.95 2.765 14.12 2.935 ;
      RECT 13.95 5.945 14.12 6.115 ;
      RECT 13.265 0.105 13.435 0.275 ;
      RECT 13.265 4.165 13.435 4.335 ;
      RECT 13.265 4.545 13.435 4.715 ;
      RECT 13.265 8.605 13.435 8.775 ;
      RECT 12.955 2.025 13.125 2.195 ;
      RECT 12.955 6.685 13.125 6.855 ;
      RECT 12.585 0.105 12.755 0.275 ;
      RECT 12.585 8.605 12.755 8.775 ;
      RECT 12.525 0.915 12.695 1.085 ;
      RECT 12.525 1.655 12.695 1.825 ;
      RECT 12.525 7.055 12.695 7.225 ;
      RECT 12.525 7.795 12.695 7.965 ;
      RECT 12.15 2.395 12.32 2.565 ;
      RECT 12.15 6.315 12.32 6.485 ;
      RECT 11.905 0.105 12.075 0.275 ;
      RECT 11.905 8.605 12.075 8.775 ;
      RECT 11.225 0.105 11.395 0.275 ;
      RECT 11.225 8.605 11.395 8.775 ;
      RECT 11.155 2.765 11.325 2.935 ;
      RECT 11.155 5.945 11.325 6.115 ;
      RECT 9.68 1.415 9.85 1.585 ;
      RECT 9.68 4.135 9.85 4.305 ;
      RECT 9.22 1.415 9.39 1.585 ;
      RECT 9.22 4.135 9.39 4.305 ;
      RECT 8.845 2.775 9.015 2.945 ;
      RECT 8.76 1.415 8.93 1.585 ;
      RECT 8.76 4.135 8.93 4.305 ;
      RECT 8.605 1.935 8.775 2.105 ;
      RECT 8.365 3.055 8.535 3.225 ;
      RECT 8.3 1.415 8.47 1.585 ;
      RECT 8.3 4.135 8.47 4.305 ;
      RECT 7.885 2.495 8.055 2.665 ;
      RECT 7.84 1.415 8.01 1.585 ;
      RECT 7.84 4.135 8.01 4.305 ;
      RECT 7.65 4.545 7.82 4.715 ;
      RECT 7.65 8.605 7.82 8.775 ;
      RECT 7.645 1.935 7.815 2.105 ;
      RECT 7.645 3.055 7.815 3.225 ;
      RECT 7.645 3.615 7.815 3.785 ;
      RECT 7.38 1.415 7.55 1.585 ;
      RECT 7.38 4.135 7.55 4.305 ;
      RECT 7.34 6.685 7.51 6.855 ;
      RECT 7.165 3.055 7.335 3.225 ;
      RECT 6.97 8.605 7.14 8.775 ;
      RECT 6.92 1.415 7.09 1.585 ;
      RECT 6.92 4.135 7.09 4.305 ;
      RECT 6.91 7.055 7.08 7.225 ;
      RECT 6.91 7.795 7.08 7.965 ;
      RECT 6.645 2.775 6.815 2.945 ;
      RECT 6.645 3.615 6.815 3.785 ;
      RECT 6.535 6.315 6.705 6.485 ;
      RECT 6.46 1.415 6.63 1.585 ;
      RECT 6.46 4.135 6.63 4.305 ;
      RECT 6.29 8.605 6.46 8.775 ;
      RECT 6.165 1.935 6.335 2.105 ;
      RECT 6.165 3.615 6.335 3.785 ;
      RECT 6 1.415 6.17 1.585 ;
      RECT 6 4.135 6.17 4.305 ;
      RECT 5.61 8.605 5.78 8.775 ;
      RECT 5.54 1.415 5.71 1.585 ;
      RECT 5.54 4.135 5.71 4.305 ;
      RECT 5.54 5.945 5.71 6.115 ;
      RECT 5.205 1.935 5.375 2.105 ;
      RECT 5.205 2.495 5.375 2.665 ;
      RECT 5.205 3.055 5.375 3.225 ;
      RECT 5.205 3.615 5.375 3.785 ;
      RECT 5.08 1.415 5.25 1.585 ;
      RECT 5.08 4.135 5.25 4.305 ;
      RECT 4.685 3.615 4.855 3.785 ;
      RECT 4.62 1.415 4.79 1.585 ;
      RECT 4.62 4.135 4.79 4.305 ;
      RECT 4.205 1.935 4.375 2.105 ;
      RECT 4.16 1.415 4.33 1.585 ;
      RECT 4.16 4.135 4.33 4.305 ;
      RECT 3.965 2.495 4.135 2.665 ;
      RECT 3.7 1.415 3.87 1.585 ;
      RECT 3.7 4.135 3.87 4.305 ;
      RECT 3.485 2.495 3.655 2.665 ;
      RECT 3.485 3.055 3.655 3.225 ;
      RECT 3.245 1.935 3.415 2.105 ;
      RECT 3.24 1.415 3.41 1.585 ;
      RECT 3.24 4.135 3.41 4.305 ;
      RECT 2.78 1.415 2.95 1.585 ;
      RECT 2.78 4.135 2.95 4.305 ;
      RECT 2.765 3.055 2.935 3.225 ;
      RECT 2.32 1.415 2.49 1.585 ;
      RECT 2.32 4.135 2.49 4.305 ;
      RECT 2.245 2.495 2.415 2.665 ;
      RECT 2.245 3.335 2.415 3.505 ;
      RECT 1.86 1.415 2.03 1.585 ;
      RECT 1.86 4.135 2.03 4.305 ;
      RECT 1.765 1.935 1.935 2.105 ;
      RECT 1.765 3.055 1.935 3.225 ;
      RECT 1.525 2.495 1.695 2.665 ;
      RECT 1.4 1.415 1.57 1.585 ;
      RECT 1.4 4.135 1.57 4.305 ;
      RECT 1.285 3.335 1.455 3.505 ;
      RECT 1.045 2.775 1.215 2.945 ;
      RECT 0.94 1.415 1.11 1.585 ;
      RECT 0.94 4.135 1.11 4.305 ;
      RECT 0.48 1.415 0.65 1.585 ;
      RECT 0.48 4.135 0.65 4.305 ;
      RECT 0.24 2.495 0.41 2.665 ;
      RECT 0.02 1.415 0.19 1.585 ;
      RECT 0.02 4.135 0.19 4.305 ;
      RECT -0.195 3.055 -0.025 3.225 ;
      RECT -0.44 1.415 -0.27 1.585 ;
      RECT -0.44 4.135 -0.27 4.305 ;
      RECT -0.675 1.935 -0.505 2.105 ;
      RECT -0.675 3.055 -0.505 3.225 ;
      RECT -0.9 1.415 -0.73 1.585 ;
      RECT -0.9 4.135 -0.73 4.305 ;
      RECT -0.915 2.495 -0.745 2.665 ;
      RECT -1.36 1.415 -1.19 1.585 ;
      RECT -1.36 4.135 -1.19 4.305 ;
      RECT -1.635 1.935 -1.465 2.105 ;
      RECT -1.635 3.475 -1.465 3.645 ;
      RECT -1.82 1.415 -1.65 1.585 ;
      RECT -1.82 4.135 -1.65 4.305 ;
      RECT -3.165 4.545 -2.995 4.715 ;
      RECT -3.165 8.605 -2.995 8.775 ;
      RECT -3.475 6.685 -3.305 6.855 ;
      RECT -3.845 8.605 -3.675 8.775 ;
      RECT -3.905 7.055 -3.735 7.225 ;
      RECT -3.905 7.795 -3.735 7.965 ;
      RECT -4.28 6.315 -4.11 6.485 ;
      RECT -4.525 8.605 -4.355 8.775 ;
      RECT -5.205 8.605 -5.035 8.775 ;
      RECT -5.275 5.945 -5.105 6.115 ;
    LAYER li ;
      RECT 83.325 0 83.495 2.085 ;
      RECT 82.365 0 82.535 2.085 ;
      RECT 81.405 0 81.575 2.085 ;
      RECT 80.885 0 81.055 2.085 ;
      RECT 79.925 0 80.095 2.085 ;
      RECT 78.925 0 79.095 2.085 ;
      RECT 77.965 0 78.135 2.085 ;
      RECT 76.485 0 76.655 2.085 ;
      RECT 74.565 0 74.735 2.085 ;
      RECT 73.085 0 73.255 2.085 ;
      RECT 64.765 0 64.935 2.085 ;
      RECT 63.805 0 63.975 2.085 ;
      RECT 62.845 0 63.015 2.085 ;
      RECT 62.325 0 62.495 2.085 ;
      RECT 61.365 0 61.535 2.085 ;
      RECT 60.365 0 60.535 2.085 ;
      RECT 59.405 0 59.575 2.085 ;
      RECT 57.925 0 58.095 2.085 ;
      RECT 56.005 0 56.175 2.085 ;
      RECT 54.525 0 54.695 2.085 ;
      RECT 46.205 0 46.375 2.085 ;
      RECT 45.245 0 45.415 2.085 ;
      RECT 44.285 0 44.455 2.085 ;
      RECT 43.765 0 43.935 2.085 ;
      RECT 42.805 0 42.975 2.085 ;
      RECT 41.805 0 41.975 2.085 ;
      RECT 40.845 0 41.015 2.085 ;
      RECT 39.365 0 39.535 2.085 ;
      RECT 37.445 0 37.615 2.085 ;
      RECT 35.965 0 36.135 2.085 ;
      RECT 27.645 0 27.815 2.085 ;
      RECT 26.685 0 26.855 2.085 ;
      RECT 25.725 0 25.895 2.085 ;
      RECT 25.205 0 25.375 2.085 ;
      RECT 24.245 0 24.415 2.085 ;
      RECT 23.245 0 23.415 2.085 ;
      RECT 22.285 0 22.455 2.085 ;
      RECT 20.805 0 20.975 2.085 ;
      RECT 18.885 0 19.055 2.085 ;
      RECT 17.405 0 17.575 2.085 ;
      RECT 9.085 0 9.255 2.085 ;
      RECT 8.125 0 8.295 2.085 ;
      RECT 7.165 0 7.335 2.085 ;
      RECT 6.645 0 6.815 2.085 ;
      RECT 5.685 0 5.855 2.085 ;
      RECT 4.685 0 4.855 2.085 ;
      RECT 3.725 0 3.895 2.085 ;
      RECT 2.245 0 2.415 2.085 ;
      RECT 0.325 0 0.495 2.085 ;
      RECT -1.155 0 -0.985 2.085 ;
      RECT 80.605 0 80.8 1.595 ;
      RECT 76.93 0 77.125 1.595 ;
      RECT 74.565 0 74.825 1.595 ;
      RECT 62.045 0 62.24 1.595 ;
      RECT 58.37 0 58.565 1.595 ;
      RECT 56.005 0 56.265 1.595 ;
      RECT 43.485 0 43.68 1.595 ;
      RECT 39.81 0 40.005 1.595 ;
      RECT 37.445 0 37.705 1.595 ;
      RECT 24.925 0 25.12 1.595 ;
      RECT 21.25 0 21.445 1.595 ;
      RECT 18.885 0 19.145 1.595 ;
      RECT 6.365 0 6.56 1.595 ;
      RECT 2.69 0 2.885 1.595 ;
      RECT 0.325 0 0.585 1.595 ;
      RECT 72.275 0 84.32 1.585 ;
      RECT 53.715 0 65.76 1.585 ;
      RECT 35.155 0 47.2 1.585 ;
      RECT 16.595 0 28.64 1.585 ;
      RECT -1.965 0 10.08 1.585 ;
      RECT 89.12 0 89.29 0.935 ;
      RECT 88.13 0 88.3 0.935 ;
      RECT 85.385 0 85.555 0.935 ;
      RECT 70.56 0 70.73 0.935 ;
      RECT 69.57 0 69.74 0.935 ;
      RECT 66.825 0 66.995 0.935 ;
      RECT 52 0 52.17 0.935 ;
      RECT 51.01 0 51.18 0.935 ;
      RECT 48.265 0 48.435 0.935 ;
      RECT 33.44 0 33.61 0.935 ;
      RECT 32.45 0 32.62 0.935 ;
      RECT 29.705 0 29.875 0.935 ;
      RECT 14.88 0 15.05 0.935 ;
      RECT 13.89 0 14.06 0.935 ;
      RECT 11.145 0 11.315 0.935 ;
      RECT -5.465 0 90.09 0.305 ;
      RECT -3.475 4.145 -3.305 8.305 ;
      RECT 89.12 3.405 89.29 5.475 ;
      RECT 88.13 3.405 88.3 5.475 ;
      RECT 85.385 3.405 85.555 5.475 ;
      RECT 79.77 4.135 79.94 5.475 ;
      RECT 70.56 3.405 70.73 5.475 ;
      RECT 69.57 3.405 69.74 5.475 ;
      RECT 66.825 3.405 66.995 5.475 ;
      RECT 61.21 4.135 61.38 5.475 ;
      RECT 52 3.405 52.17 5.475 ;
      RECT 51.01 3.405 51.18 5.475 ;
      RECT 48.265 3.405 48.435 5.475 ;
      RECT 42.65 4.135 42.82 5.475 ;
      RECT 33.44 3.405 33.61 5.475 ;
      RECT 32.45 3.405 32.62 5.475 ;
      RECT 29.705 3.405 29.875 5.475 ;
      RECT 24.09 4.135 24.26 5.475 ;
      RECT 14.88 3.405 15.05 5.475 ;
      RECT 13.89 3.405 14.06 5.475 ;
      RECT 11.145 3.405 11.315 5.475 ;
      RECT 5.53 4.135 5.7 5.475 ;
      RECT -5.285 4.145 -5.115 5.475 ;
      RECT 71.53 4.145 73.995 4.75 ;
      RECT 52.97 4.145 55.435 4.75 ;
      RECT 34.41 4.145 36.875 4.75 ;
      RECT 15.85 4.145 18.315 4.75 ;
      RECT -5.46 4.145 -0.245 4.75 ;
      RECT 72.275 4.135 90.09 4.745 ;
      RECT 53.715 4.135 71.53 4.745 ;
      RECT 35.155 4.135 52.97 4.745 ;
      RECT 16.595 4.135 34.41 4.745 ;
      RECT -1.965 4.135 15.85 4.745 ;
      RECT 82.365 3.635 82.535 4.745 ;
      RECT 79.925 3.635 80.095 4.745 ;
      RECT 77.965 3.635 78.135 4.745 ;
      RECT 77.005 3.635 77.175 4.745 ;
      RECT 75.045 3.635 75.215 4.745 ;
      RECT 74.045 3.635 74.215 4.745 ;
      RECT 73.085 3.635 73.255 4.75 ;
      RECT 63.805 3.635 63.975 4.745 ;
      RECT 61.365 3.635 61.535 4.745 ;
      RECT 59.405 3.635 59.575 4.745 ;
      RECT 58.445 3.635 58.615 4.745 ;
      RECT 56.485 3.635 56.655 4.745 ;
      RECT 55.485 3.635 55.655 4.745 ;
      RECT 54.525 3.635 54.695 4.75 ;
      RECT 45.245 3.635 45.415 4.745 ;
      RECT 42.805 3.635 42.975 4.745 ;
      RECT 40.845 3.635 41.015 4.745 ;
      RECT 39.885 3.635 40.055 4.745 ;
      RECT 37.925 3.635 38.095 4.745 ;
      RECT 36.925 3.635 37.095 4.745 ;
      RECT 35.965 3.635 36.135 4.75 ;
      RECT 26.685 3.635 26.855 4.745 ;
      RECT 24.245 3.635 24.415 4.745 ;
      RECT 22.285 3.635 22.455 4.745 ;
      RECT 21.325 3.635 21.495 4.745 ;
      RECT 19.365 3.635 19.535 4.745 ;
      RECT 18.365 3.635 18.535 4.745 ;
      RECT 17.405 3.635 17.575 4.75 ;
      RECT 8.125 3.635 8.295 4.745 ;
      RECT 5.685 3.635 5.855 4.745 ;
      RECT 3.725 3.635 3.895 4.745 ;
      RECT 2.765 3.635 2.935 4.745 ;
      RECT 0.805 3.635 0.975 4.745 ;
      RECT -0.195 3.635 -0.025 4.745 ;
      RECT -1.155 3.635 -0.985 4.75 ;
      RECT -5.465 8.575 90.09 8.88 ;
      RECT 89.12 7.945 89.29 8.88 ;
      RECT 88.13 7.945 88.3 8.88 ;
      RECT 85.385 7.945 85.555 8.88 ;
      RECT 79.77 7.945 79.94 8.88 ;
      RECT 70.56 7.945 70.73 8.88 ;
      RECT 69.57 7.945 69.74 8.88 ;
      RECT 66.825 7.945 66.995 8.88 ;
      RECT 61.21 7.945 61.38 8.88 ;
      RECT 52 7.945 52.17 8.88 ;
      RECT 51.01 7.945 51.18 8.88 ;
      RECT 48.265 7.945 48.435 8.88 ;
      RECT 42.65 7.945 42.82 8.88 ;
      RECT 33.44 7.945 33.61 8.88 ;
      RECT 32.45 7.945 32.62 8.88 ;
      RECT 29.705 7.945 29.875 8.88 ;
      RECT 24.09 7.945 24.26 8.88 ;
      RECT 14.88 7.945 15.05 8.88 ;
      RECT 13.89 7.945 14.06 8.88 ;
      RECT 11.145 7.945 11.315 8.88 ;
      RECT 5.53 7.945 5.7 8.88 ;
      RECT -5.285 7.945 -5.115 8.88 ;
      RECT 89.18 1.74 89.35 2.935 ;
      RECT 89.18 1.74 89.645 1.91 ;
      RECT 89.18 6.97 89.645 7.14 ;
      RECT 89.18 5.945 89.35 7.14 ;
      RECT 88.19 1.74 88.36 2.935 ;
      RECT 88.19 1.74 88.655 1.91 ;
      RECT 88.19 6.97 88.655 7.14 ;
      RECT 88.19 5.945 88.36 7.14 ;
      RECT 86.335 2.635 86.505 3.865 ;
      RECT 86.39 0.855 86.56 2.805 ;
      RECT 86.335 0.575 86.505 1.025 ;
      RECT 86.335 7.855 86.505 8.305 ;
      RECT 86.39 6.075 86.56 8.025 ;
      RECT 86.335 5.015 86.505 6.245 ;
      RECT 85.815 0.575 85.985 3.865 ;
      RECT 85.815 2.075 86.22 2.405 ;
      RECT 85.815 1.235 86.22 1.565 ;
      RECT 85.815 5.015 85.985 8.305 ;
      RECT 85.815 7.315 86.22 7.645 ;
      RECT 85.815 6.475 86.22 6.805 ;
      RECT 82.605 3.225 83.575 3.395 ;
      RECT 82.605 3.055 82.775 3.395 ;
      RECT 82.125 2.495 82.295 2.825 ;
      RECT 82.125 2.575 82.855 2.745 ;
      RECT 81.765 3.615 82.055 3.785 ;
      RECT 81.765 2.575 81.935 3.785 ;
      RECT 81.765 3.055 82.055 3.225 ;
      RECT 81.565 2.575 81.935 2.745 ;
      RECT 80.885 2.675 81.055 2.945 ;
      RECT 80.645 2.675 81.055 2.845 ;
      RECT 80.565 2.575 80.895 2.745 ;
      RECT 80.405 3.615 81.055 3.785 ;
      RECT 80.885 3.145 81.055 3.785 ;
      RECT 80.765 3.225 81.055 3.785 ;
      RECT 80.72 7.855 80.89 8.305 ;
      RECT 80.775 6.075 80.945 8.025 ;
      RECT 80.72 5.015 80.89 6.245 ;
      RECT 80.2 5.015 80.37 8.305 ;
      RECT 80.2 7.315 80.605 7.645 ;
      RECT 80.2 6.475 80.605 6.805 ;
      RECT 79.445 2.915 79.615 3.225 ;
      RECT 79.445 2.915 80.335 3.085 ;
      RECT 80.165 2.495 80.335 3.085 ;
      RECT 79.445 2.575 79.935 2.745 ;
      RECT 79.445 2.495 79.615 2.745 ;
      RECT 77.405 3.225 77.895 3.395 ;
      RECT 78.565 2.575 78.735 3.225 ;
      RECT 77.725 3.055 78.735 3.225 ;
      RECT 78.685 2.495 78.855 2.825 ;
      RECT 77.485 1.835 77.655 2.105 ;
      RECT 76.925 1.835 77.655 2.005 ;
      RECT 77.005 2.575 77.175 3.225 ;
      RECT 77.005 2.575 77.495 2.745 ;
      RECT 76.165 2.575 76.655 2.745 ;
      RECT 76.485 2.495 76.655 2.745 ;
      RECT 76.005 1.835 76.175 2.105 ;
      RECT 75.445 1.835 76.175 2.005 ;
      RECT 75.525 3.225 75.695 3.505 ;
      RECT 74.485 3.225 75.775 3.395 ;
      RECT 74.48 2.575 75.055 2.745 ;
      RECT 74.48 2.495 74.65 2.745 ;
      RECT 73.565 1.835 73.735 2.105 ;
      RECT 73.565 1.835 74.295 2.005 ;
      RECT 73.925 3.055 74.215 3.225 ;
      RECT 73.925 2.575 74.095 3.225 ;
      RECT 73.725 2.575 74.095 2.745 ;
      RECT 73.565 3.055 73.735 3.475 ;
      RECT 72.945 3.14 73.735 3.31 ;
      RECT 72.945 2.915 73.115 3.31 ;
      RECT 72.845 2.495 73.015 3.085 ;
      RECT 72.605 2.575 73.015 2.845 ;
      RECT 70.62 1.74 70.79 2.935 ;
      RECT 70.62 1.74 71.085 1.91 ;
      RECT 70.62 6.97 71.085 7.14 ;
      RECT 70.62 5.945 70.79 7.14 ;
      RECT 69.63 1.74 69.8 2.935 ;
      RECT 69.63 1.74 70.095 1.91 ;
      RECT 69.63 6.97 70.095 7.14 ;
      RECT 69.63 5.945 69.8 7.14 ;
      RECT 67.775 2.635 67.945 3.865 ;
      RECT 67.83 0.855 68 2.805 ;
      RECT 67.775 0.575 67.945 1.025 ;
      RECT 67.775 7.855 67.945 8.305 ;
      RECT 67.83 6.075 68 8.025 ;
      RECT 67.775 5.015 67.945 6.245 ;
      RECT 67.255 0.575 67.425 3.865 ;
      RECT 67.255 2.075 67.66 2.405 ;
      RECT 67.255 1.235 67.66 1.565 ;
      RECT 67.255 5.015 67.425 8.305 ;
      RECT 67.255 7.315 67.66 7.645 ;
      RECT 67.255 6.475 67.66 6.805 ;
      RECT 64.045 3.225 65.015 3.395 ;
      RECT 64.045 3.055 64.215 3.395 ;
      RECT 63.565 2.495 63.735 2.825 ;
      RECT 63.565 2.575 64.295 2.745 ;
      RECT 63.205 3.615 63.495 3.785 ;
      RECT 63.205 2.575 63.375 3.785 ;
      RECT 63.205 3.055 63.495 3.225 ;
      RECT 63.005 2.575 63.375 2.745 ;
      RECT 62.325 2.675 62.495 2.945 ;
      RECT 62.085 2.675 62.495 2.845 ;
      RECT 62.005 2.575 62.335 2.745 ;
      RECT 61.845 3.615 62.495 3.785 ;
      RECT 62.325 3.145 62.495 3.785 ;
      RECT 62.205 3.225 62.495 3.785 ;
      RECT 62.16 7.855 62.33 8.305 ;
      RECT 62.215 6.075 62.385 8.025 ;
      RECT 62.16 5.015 62.33 6.245 ;
      RECT 61.64 5.015 61.81 8.305 ;
      RECT 61.64 7.315 62.045 7.645 ;
      RECT 61.64 6.475 62.045 6.805 ;
      RECT 60.885 2.915 61.055 3.225 ;
      RECT 60.885 2.915 61.775 3.085 ;
      RECT 61.605 2.495 61.775 3.085 ;
      RECT 60.885 2.575 61.375 2.745 ;
      RECT 60.885 2.495 61.055 2.745 ;
      RECT 58.845 3.225 59.335 3.395 ;
      RECT 60.005 2.575 60.175 3.225 ;
      RECT 59.165 3.055 60.175 3.225 ;
      RECT 60.125 2.495 60.295 2.825 ;
      RECT 58.925 1.835 59.095 2.105 ;
      RECT 58.365 1.835 59.095 2.005 ;
      RECT 58.445 2.575 58.615 3.225 ;
      RECT 58.445 2.575 58.935 2.745 ;
      RECT 57.605 2.575 58.095 2.745 ;
      RECT 57.925 2.495 58.095 2.745 ;
      RECT 57.445 1.835 57.615 2.105 ;
      RECT 56.885 1.835 57.615 2.005 ;
      RECT 56.965 3.225 57.135 3.505 ;
      RECT 55.925 3.225 57.215 3.395 ;
      RECT 55.92 2.575 56.495 2.745 ;
      RECT 55.92 2.495 56.09 2.745 ;
      RECT 55.005 1.835 55.175 2.105 ;
      RECT 55.005 1.835 55.735 2.005 ;
      RECT 55.365 3.055 55.655 3.225 ;
      RECT 55.365 2.575 55.535 3.225 ;
      RECT 55.165 2.575 55.535 2.745 ;
      RECT 55.005 3.055 55.175 3.475 ;
      RECT 54.385 3.14 55.175 3.31 ;
      RECT 54.385 2.915 54.555 3.31 ;
      RECT 54.285 2.495 54.455 3.085 ;
      RECT 54.045 2.575 54.455 2.845 ;
      RECT 52.06 1.74 52.23 2.935 ;
      RECT 52.06 1.74 52.525 1.91 ;
      RECT 52.06 6.97 52.525 7.14 ;
      RECT 52.06 5.945 52.23 7.14 ;
      RECT 51.07 1.74 51.24 2.935 ;
      RECT 51.07 1.74 51.535 1.91 ;
      RECT 51.07 6.97 51.535 7.14 ;
      RECT 51.07 5.945 51.24 7.14 ;
      RECT 49.215 2.635 49.385 3.865 ;
      RECT 49.27 0.855 49.44 2.805 ;
      RECT 49.215 0.575 49.385 1.025 ;
      RECT 49.215 7.855 49.385 8.305 ;
      RECT 49.27 6.075 49.44 8.025 ;
      RECT 49.215 5.015 49.385 6.245 ;
      RECT 48.695 0.575 48.865 3.865 ;
      RECT 48.695 2.075 49.1 2.405 ;
      RECT 48.695 1.235 49.1 1.565 ;
      RECT 48.695 5.015 48.865 8.305 ;
      RECT 48.695 7.315 49.1 7.645 ;
      RECT 48.695 6.475 49.1 6.805 ;
      RECT 45.485 3.225 46.455 3.395 ;
      RECT 45.485 3.055 45.655 3.395 ;
      RECT 45.005 2.495 45.175 2.825 ;
      RECT 45.005 2.575 45.735 2.745 ;
      RECT 44.645 3.615 44.935 3.785 ;
      RECT 44.645 2.575 44.815 3.785 ;
      RECT 44.645 3.055 44.935 3.225 ;
      RECT 44.445 2.575 44.815 2.745 ;
      RECT 43.765 2.675 43.935 2.945 ;
      RECT 43.525 2.675 43.935 2.845 ;
      RECT 43.445 2.575 43.775 2.745 ;
      RECT 43.285 3.615 43.935 3.785 ;
      RECT 43.765 3.145 43.935 3.785 ;
      RECT 43.645 3.225 43.935 3.785 ;
      RECT 43.6 7.855 43.77 8.305 ;
      RECT 43.655 6.075 43.825 8.025 ;
      RECT 43.6 5.015 43.77 6.245 ;
      RECT 43.08 5.015 43.25 8.305 ;
      RECT 43.08 7.315 43.485 7.645 ;
      RECT 43.08 6.475 43.485 6.805 ;
      RECT 42.325 2.915 42.495 3.225 ;
      RECT 42.325 2.915 43.215 3.085 ;
      RECT 43.045 2.495 43.215 3.085 ;
      RECT 42.325 2.575 42.815 2.745 ;
      RECT 42.325 2.495 42.495 2.745 ;
      RECT 40.285 3.225 40.775 3.395 ;
      RECT 41.445 2.575 41.615 3.225 ;
      RECT 40.605 3.055 41.615 3.225 ;
      RECT 41.565 2.495 41.735 2.825 ;
      RECT 40.365 1.835 40.535 2.105 ;
      RECT 39.805 1.835 40.535 2.005 ;
      RECT 39.885 2.575 40.055 3.225 ;
      RECT 39.885 2.575 40.375 2.745 ;
      RECT 39.045 2.575 39.535 2.745 ;
      RECT 39.365 2.495 39.535 2.745 ;
      RECT 38.885 1.835 39.055 2.105 ;
      RECT 38.325 1.835 39.055 2.005 ;
      RECT 38.405 3.225 38.575 3.505 ;
      RECT 37.365 3.225 38.655 3.395 ;
      RECT 37.36 2.575 37.935 2.745 ;
      RECT 37.36 2.495 37.53 2.745 ;
      RECT 36.445 1.835 36.615 2.105 ;
      RECT 36.445 1.835 37.175 2.005 ;
      RECT 36.805 3.055 37.095 3.225 ;
      RECT 36.805 2.575 36.975 3.225 ;
      RECT 36.605 2.575 36.975 2.745 ;
      RECT 36.445 3.055 36.615 3.475 ;
      RECT 35.825 3.14 36.615 3.31 ;
      RECT 35.825 2.915 35.995 3.31 ;
      RECT 35.725 2.495 35.895 3.085 ;
      RECT 35.485 2.575 35.895 2.845 ;
      RECT 33.5 1.74 33.67 2.935 ;
      RECT 33.5 1.74 33.965 1.91 ;
      RECT 33.5 6.97 33.965 7.14 ;
      RECT 33.5 5.945 33.67 7.14 ;
      RECT 32.51 1.74 32.68 2.935 ;
      RECT 32.51 1.74 32.975 1.91 ;
      RECT 32.51 6.97 32.975 7.14 ;
      RECT 32.51 5.945 32.68 7.14 ;
      RECT 30.655 2.635 30.825 3.865 ;
      RECT 30.71 0.855 30.88 2.805 ;
      RECT 30.655 0.575 30.825 1.025 ;
      RECT 30.655 7.855 30.825 8.305 ;
      RECT 30.71 6.075 30.88 8.025 ;
      RECT 30.655 5.015 30.825 6.245 ;
      RECT 30.135 0.575 30.305 3.865 ;
      RECT 30.135 2.075 30.54 2.405 ;
      RECT 30.135 1.235 30.54 1.565 ;
      RECT 30.135 5.015 30.305 8.305 ;
      RECT 30.135 7.315 30.54 7.645 ;
      RECT 30.135 6.475 30.54 6.805 ;
      RECT 26.925 3.225 27.895 3.395 ;
      RECT 26.925 3.055 27.095 3.395 ;
      RECT 26.445 2.495 26.615 2.825 ;
      RECT 26.445 2.575 27.175 2.745 ;
      RECT 26.085 3.615 26.375 3.785 ;
      RECT 26.085 2.575 26.255 3.785 ;
      RECT 26.085 3.055 26.375 3.225 ;
      RECT 25.885 2.575 26.255 2.745 ;
      RECT 25.205 2.675 25.375 2.945 ;
      RECT 24.965 2.675 25.375 2.845 ;
      RECT 24.885 2.575 25.215 2.745 ;
      RECT 24.725 3.615 25.375 3.785 ;
      RECT 25.205 3.145 25.375 3.785 ;
      RECT 25.085 3.225 25.375 3.785 ;
      RECT 25.04 7.855 25.21 8.305 ;
      RECT 25.095 6.075 25.265 8.025 ;
      RECT 25.04 5.015 25.21 6.245 ;
      RECT 24.52 5.015 24.69 8.305 ;
      RECT 24.52 7.315 24.925 7.645 ;
      RECT 24.52 6.475 24.925 6.805 ;
      RECT 23.765 2.915 23.935 3.225 ;
      RECT 23.765 2.915 24.655 3.085 ;
      RECT 24.485 2.495 24.655 3.085 ;
      RECT 23.765 2.575 24.255 2.745 ;
      RECT 23.765 2.495 23.935 2.745 ;
      RECT 21.725 3.225 22.215 3.395 ;
      RECT 22.885 2.575 23.055 3.225 ;
      RECT 22.045 3.055 23.055 3.225 ;
      RECT 23.005 2.495 23.175 2.825 ;
      RECT 21.805 1.835 21.975 2.105 ;
      RECT 21.245 1.835 21.975 2.005 ;
      RECT 21.325 2.575 21.495 3.225 ;
      RECT 21.325 2.575 21.815 2.745 ;
      RECT 20.485 2.575 20.975 2.745 ;
      RECT 20.805 2.495 20.975 2.745 ;
      RECT 20.325 1.835 20.495 2.105 ;
      RECT 19.765 1.835 20.495 2.005 ;
      RECT 19.845 3.225 20.015 3.505 ;
      RECT 18.805 3.225 20.095 3.395 ;
      RECT 18.8 2.575 19.375 2.745 ;
      RECT 18.8 2.495 18.97 2.745 ;
      RECT 17.885 1.835 18.055 2.105 ;
      RECT 17.885 1.835 18.615 2.005 ;
      RECT 18.245 3.055 18.535 3.225 ;
      RECT 18.245 2.575 18.415 3.225 ;
      RECT 18.045 2.575 18.415 2.745 ;
      RECT 17.885 3.055 18.055 3.475 ;
      RECT 17.265 3.14 18.055 3.31 ;
      RECT 17.265 2.915 17.435 3.31 ;
      RECT 17.165 2.495 17.335 3.085 ;
      RECT 16.925 2.575 17.335 2.845 ;
      RECT 14.94 1.74 15.11 2.935 ;
      RECT 14.94 1.74 15.405 1.91 ;
      RECT 14.94 6.97 15.405 7.14 ;
      RECT 14.94 5.945 15.11 7.14 ;
      RECT 13.95 1.74 14.12 2.935 ;
      RECT 13.95 1.74 14.415 1.91 ;
      RECT 13.95 6.97 14.415 7.14 ;
      RECT 13.95 5.945 14.12 7.14 ;
      RECT 12.095 2.635 12.265 3.865 ;
      RECT 12.15 0.855 12.32 2.805 ;
      RECT 12.095 0.575 12.265 1.025 ;
      RECT 12.095 7.855 12.265 8.305 ;
      RECT 12.15 6.075 12.32 8.025 ;
      RECT 12.095 5.015 12.265 6.245 ;
      RECT 11.575 0.575 11.745 3.865 ;
      RECT 11.575 2.075 11.98 2.405 ;
      RECT 11.575 1.235 11.98 1.565 ;
      RECT 11.575 5.015 11.745 8.305 ;
      RECT 11.575 7.315 11.98 7.645 ;
      RECT 11.575 6.475 11.98 6.805 ;
      RECT 8.365 3.225 9.335 3.395 ;
      RECT 8.365 3.055 8.535 3.395 ;
      RECT 7.885 2.495 8.055 2.825 ;
      RECT 7.885 2.575 8.615 2.745 ;
      RECT 7.525 3.615 7.815 3.785 ;
      RECT 7.525 2.575 7.695 3.785 ;
      RECT 7.525 3.055 7.815 3.225 ;
      RECT 7.325 2.575 7.695 2.745 ;
      RECT 6.645 2.675 6.815 2.945 ;
      RECT 6.405 2.675 6.815 2.845 ;
      RECT 6.325 2.575 6.655 2.745 ;
      RECT 6.165 3.615 6.815 3.785 ;
      RECT 6.645 3.145 6.815 3.785 ;
      RECT 6.525 3.225 6.815 3.785 ;
      RECT 6.48 7.855 6.65 8.305 ;
      RECT 6.535 6.075 6.705 8.025 ;
      RECT 6.48 5.015 6.65 6.245 ;
      RECT 5.96 5.015 6.13 8.305 ;
      RECT 5.96 7.315 6.365 7.645 ;
      RECT 5.96 6.475 6.365 6.805 ;
      RECT 5.205 2.915 5.375 3.225 ;
      RECT 5.205 2.915 6.095 3.085 ;
      RECT 5.925 2.495 6.095 3.085 ;
      RECT 5.205 2.575 5.695 2.745 ;
      RECT 5.205 2.495 5.375 2.745 ;
      RECT 3.165 3.225 3.655 3.395 ;
      RECT 4.325 2.575 4.495 3.225 ;
      RECT 3.485 3.055 4.495 3.225 ;
      RECT 4.445 2.495 4.615 2.825 ;
      RECT 3.245 1.835 3.415 2.105 ;
      RECT 2.685 1.835 3.415 2.005 ;
      RECT 2.765 2.575 2.935 3.225 ;
      RECT 2.765 2.575 3.255 2.745 ;
      RECT 1.925 2.575 2.415 2.745 ;
      RECT 2.245 2.495 2.415 2.745 ;
      RECT 1.765 1.835 1.935 2.105 ;
      RECT 1.205 1.835 1.935 2.005 ;
      RECT 1.285 3.225 1.455 3.505 ;
      RECT 0.245 3.225 1.535 3.395 ;
      RECT 0.24 2.575 0.815 2.745 ;
      RECT 0.24 2.495 0.41 2.745 ;
      RECT -0.675 1.835 -0.505 2.105 ;
      RECT -0.675 1.835 0.055 2.005 ;
      RECT -0.315 3.055 -0.025 3.225 ;
      RECT -0.315 2.575 -0.145 3.225 ;
      RECT -0.515 2.575 -0.145 2.745 ;
      RECT -0.675 3.055 -0.505 3.475 ;
      RECT -1.295 3.14 -0.505 3.31 ;
      RECT -1.295 2.915 -1.125 3.31 ;
      RECT -1.395 2.495 -1.225 3.085 ;
      RECT -1.635 2.575 -1.225 2.845 ;
      RECT -4.335 7.855 -4.165 8.305 ;
      RECT -4.28 6.075 -4.11 8.025 ;
      RECT -4.335 5.015 -4.165 6.245 ;
      RECT -4.855 5.015 -4.685 8.305 ;
      RECT -4.855 7.315 -4.45 7.645 ;
      RECT -4.855 6.475 -4.45 6.805 ;
      RECT 89.55 0.575 89.72 1.085 ;
      RECT 89.55 2.395 89.72 3.865 ;
      RECT 89.55 5.015 89.72 6.485 ;
      RECT 89.55 7.795 89.72 8.305 ;
      RECT 88.56 0.575 88.73 1.085 ;
      RECT 88.56 2.395 88.73 3.865 ;
      RECT 88.56 5.015 88.73 6.485 ;
      RECT 88.56 7.795 88.73 8.305 ;
      RECT 87.195 0.575 87.365 3.865 ;
      RECT 87.195 5.015 87.365 8.305 ;
      RECT 86.765 0.575 86.935 1.085 ;
      RECT 86.765 1.655 86.935 3.865 ;
      RECT 86.765 5.015 86.935 7.225 ;
      RECT 86.765 7.795 86.935 8.305 ;
      RECT 85.395 1.66 85.565 2.935 ;
      RECT 85.395 5.945 85.565 7.22 ;
      RECT 83.085 2.495 83.255 2.945 ;
      RECT 82.845 1.755 83.015 2.105 ;
      RECT 81.885 1.755 82.055 2.105 ;
      RECT 81.58 5.015 81.75 8.305 ;
      RECT 81.405 3.055 81.575 3.475 ;
      RECT 81.15 5.015 81.32 7.225 ;
      RECT 81.15 7.795 81.32 8.305 ;
      RECT 80.405 1.755 80.575 2.105 ;
      RECT 79.78 5.945 79.95 7.22 ;
      RECT 79.445 1.755 79.615 2.105 ;
      RECT 79.445 3.485 79.615 3.815 ;
      RECT 78.925 3.145 79.095 3.785 ;
      RECT 78.445 1.755 78.615 2.105 ;
      RECT 78.205 2.495 78.375 2.825 ;
      RECT 77.725 2.495 77.895 2.825 ;
      RECT 76.485 3.145 76.655 3.505 ;
      RECT 76.005 3.055 76.175 3.475 ;
      RECT 75.765 2.495 75.935 2.825 ;
      RECT 75.285 2.495 75.455 2.945 ;
      RECT 73.325 2.495 73.495 2.825 ;
      RECT 72.605 1.755 72.775 2.105 ;
      RECT 72.605 3.285 72.775 3.645 ;
      RECT 70.99 0.575 71.16 1.085 ;
      RECT 70.99 2.395 71.16 3.865 ;
      RECT 70.99 5.015 71.16 6.485 ;
      RECT 70.99 7.795 71.16 8.305 ;
      RECT 70 0.575 70.17 1.085 ;
      RECT 70 2.395 70.17 3.865 ;
      RECT 70 5.015 70.17 6.485 ;
      RECT 70 7.795 70.17 8.305 ;
      RECT 68.635 0.575 68.805 3.865 ;
      RECT 68.635 5.015 68.805 8.305 ;
      RECT 68.205 0.575 68.375 1.085 ;
      RECT 68.205 1.655 68.375 3.865 ;
      RECT 68.205 5.015 68.375 7.225 ;
      RECT 68.205 7.795 68.375 8.305 ;
      RECT 66.835 1.66 67.005 2.935 ;
      RECT 66.835 5.945 67.005 7.22 ;
      RECT 64.525 2.495 64.695 2.945 ;
      RECT 64.285 1.755 64.455 2.105 ;
      RECT 63.325 1.755 63.495 2.105 ;
      RECT 63.02 5.015 63.19 8.305 ;
      RECT 62.845 3.055 63.015 3.475 ;
      RECT 62.59 5.015 62.76 7.225 ;
      RECT 62.59 7.795 62.76 8.305 ;
      RECT 61.845 1.755 62.015 2.105 ;
      RECT 61.22 5.945 61.39 7.22 ;
      RECT 60.885 1.755 61.055 2.105 ;
      RECT 60.885 3.485 61.055 3.815 ;
      RECT 60.365 3.145 60.535 3.785 ;
      RECT 59.885 1.755 60.055 2.105 ;
      RECT 59.645 2.495 59.815 2.825 ;
      RECT 59.165 2.495 59.335 2.825 ;
      RECT 57.925 3.145 58.095 3.505 ;
      RECT 57.445 3.055 57.615 3.475 ;
      RECT 57.205 2.495 57.375 2.825 ;
      RECT 56.725 2.495 56.895 2.945 ;
      RECT 54.765 2.495 54.935 2.825 ;
      RECT 54.045 1.755 54.215 2.105 ;
      RECT 54.045 3.285 54.215 3.645 ;
      RECT 52.43 0.575 52.6 1.085 ;
      RECT 52.43 2.395 52.6 3.865 ;
      RECT 52.43 5.015 52.6 6.485 ;
      RECT 52.43 7.795 52.6 8.305 ;
      RECT 51.44 0.575 51.61 1.085 ;
      RECT 51.44 2.395 51.61 3.865 ;
      RECT 51.44 5.015 51.61 6.485 ;
      RECT 51.44 7.795 51.61 8.305 ;
      RECT 50.075 0.575 50.245 3.865 ;
      RECT 50.075 5.015 50.245 8.305 ;
      RECT 49.645 0.575 49.815 1.085 ;
      RECT 49.645 1.655 49.815 3.865 ;
      RECT 49.645 5.015 49.815 7.225 ;
      RECT 49.645 7.795 49.815 8.305 ;
      RECT 48.275 1.66 48.445 2.935 ;
      RECT 48.275 5.945 48.445 7.22 ;
      RECT 45.965 2.495 46.135 2.945 ;
      RECT 45.725 1.755 45.895 2.105 ;
      RECT 44.765 1.755 44.935 2.105 ;
      RECT 44.46 5.015 44.63 8.305 ;
      RECT 44.285 3.055 44.455 3.475 ;
      RECT 44.03 5.015 44.2 7.225 ;
      RECT 44.03 7.795 44.2 8.305 ;
      RECT 43.285 1.755 43.455 2.105 ;
      RECT 42.66 5.945 42.83 7.22 ;
      RECT 42.325 1.755 42.495 2.105 ;
      RECT 42.325 3.485 42.495 3.815 ;
      RECT 41.805 3.145 41.975 3.785 ;
      RECT 41.325 1.755 41.495 2.105 ;
      RECT 41.085 2.495 41.255 2.825 ;
      RECT 40.605 2.495 40.775 2.825 ;
      RECT 39.365 3.145 39.535 3.505 ;
      RECT 38.885 3.055 39.055 3.475 ;
      RECT 38.645 2.495 38.815 2.825 ;
      RECT 38.165 2.495 38.335 2.945 ;
      RECT 36.205 2.495 36.375 2.825 ;
      RECT 35.485 1.755 35.655 2.105 ;
      RECT 35.485 3.285 35.655 3.645 ;
      RECT 33.87 0.575 34.04 1.085 ;
      RECT 33.87 2.395 34.04 3.865 ;
      RECT 33.87 5.015 34.04 6.485 ;
      RECT 33.87 7.795 34.04 8.305 ;
      RECT 32.88 0.575 33.05 1.085 ;
      RECT 32.88 2.395 33.05 3.865 ;
      RECT 32.88 5.015 33.05 6.485 ;
      RECT 32.88 7.795 33.05 8.305 ;
      RECT 31.515 0.575 31.685 3.865 ;
      RECT 31.515 5.015 31.685 8.305 ;
      RECT 31.085 0.575 31.255 1.085 ;
      RECT 31.085 1.655 31.255 3.865 ;
      RECT 31.085 5.015 31.255 7.225 ;
      RECT 31.085 7.795 31.255 8.305 ;
      RECT 29.715 1.66 29.885 2.935 ;
      RECT 29.715 5.945 29.885 7.22 ;
      RECT 27.405 2.495 27.575 2.945 ;
      RECT 27.165 1.755 27.335 2.105 ;
      RECT 26.205 1.755 26.375 2.105 ;
      RECT 25.9 5.015 26.07 8.305 ;
      RECT 25.725 3.055 25.895 3.475 ;
      RECT 25.47 5.015 25.64 7.225 ;
      RECT 25.47 7.795 25.64 8.305 ;
      RECT 24.725 1.755 24.895 2.105 ;
      RECT 24.1 5.945 24.27 7.22 ;
      RECT 23.765 1.755 23.935 2.105 ;
      RECT 23.765 3.485 23.935 3.815 ;
      RECT 23.245 3.145 23.415 3.785 ;
      RECT 22.765 1.755 22.935 2.105 ;
      RECT 22.525 2.495 22.695 2.825 ;
      RECT 22.045 2.495 22.215 2.825 ;
      RECT 20.805 3.145 20.975 3.505 ;
      RECT 20.325 3.055 20.495 3.475 ;
      RECT 20.085 2.495 20.255 2.825 ;
      RECT 19.605 2.495 19.775 2.945 ;
      RECT 17.645 2.495 17.815 2.825 ;
      RECT 16.925 1.755 17.095 2.105 ;
      RECT 16.925 3.285 17.095 3.645 ;
      RECT 15.31 0.575 15.48 1.085 ;
      RECT 15.31 2.395 15.48 3.865 ;
      RECT 15.31 5.015 15.48 6.485 ;
      RECT 15.31 7.795 15.48 8.305 ;
      RECT 14.32 0.575 14.49 1.085 ;
      RECT 14.32 2.395 14.49 3.865 ;
      RECT 14.32 5.015 14.49 6.485 ;
      RECT 14.32 7.795 14.49 8.305 ;
      RECT 12.955 0.575 13.125 3.865 ;
      RECT 12.955 5.015 13.125 8.305 ;
      RECT 12.525 0.575 12.695 1.085 ;
      RECT 12.525 1.655 12.695 3.865 ;
      RECT 12.525 5.015 12.695 7.225 ;
      RECT 12.525 7.795 12.695 8.305 ;
      RECT 11.155 1.66 11.325 2.935 ;
      RECT 11.155 5.945 11.325 7.22 ;
      RECT 8.845 2.495 9.015 2.945 ;
      RECT 8.605 1.755 8.775 2.105 ;
      RECT 7.645 1.755 7.815 2.105 ;
      RECT 7.34 5.015 7.51 8.305 ;
      RECT 7.165 3.055 7.335 3.475 ;
      RECT 6.91 5.015 7.08 7.225 ;
      RECT 6.91 7.795 7.08 8.305 ;
      RECT 6.165 1.755 6.335 2.105 ;
      RECT 5.54 5.945 5.71 7.22 ;
      RECT 5.205 1.755 5.375 2.105 ;
      RECT 5.205 3.485 5.375 3.815 ;
      RECT 4.685 3.145 4.855 3.785 ;
      RECT 4.205 1.755 4.375 2.105 ;
      RECT 3.965 2.495 4.135 2.825 ;
      RECT 3.485 2.495 3.655 2.825 ;
      RECT 2.245 3.145 2.415 3.505 ;
      RECT 1.765 3.055 1.935 3.475 ;
      RECT 1.525 2.495 1.695 2.825 ;
      RECT 1.045 2.495 1.215 2.945 ;
      RECT -0.915 2.495 -0.745 2.825 ;
      RECT -1.635 1.755 -1.465 2.105 ;
      RECT -1.635 3.285 -1.465 3.645 ;
      RECT -3.905 5.015 -3.735 7.225 ;
      RECT -3.905 7.795 -3.735 8.305 ;
      RECT -5.275 5.945 -5.105 7.22 ;
  END
END sky130_osu_ring_oscillator_mpr2et_8_b0r1

MACRO sky130_osu_ring_oscillator_mpr2et_8_b0r2
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 5.505 0 ;
  SIZE 95.595 BY 8.88 ;
  SYMMETRY X Y R90 ;
  SITE CoreSite ;
  OBS
    LAYER met3 ;
      RECT 81.58 3.535 82.135 3.865 ;
      RECT 81.58 1.87 81.88 3.865 ;
      RECT 77.645 2.975 78.2 3.305 ;
      RECT 77.9 1.87 78.2 3.305 ;
      RECT 77.9 1.87 81.88 2.17 ;
      RECT 81.05 7.055 81.425 7.425 ;
      RECT 81.05 7.095 82.055 7.395 ;
      RECT 81.755 4.405 82.055 7.395 ;
      RECT 71.925 4.405 82.055 4.705 ;
      RECT 76.43 2.415 76.73 4.705 ;
      RECT 74.995 2.975 75.295 4.705 ;
      RECT 71.925 2.42 72.225 4.705 ;
      RECT 74.965 2.975 75.695 3.305 ;
      RECT 76.405 2.415 77.135 2.745 ;
      RECT 72.855 2.415 73.585 2.745 ;
      RECT 71.925 2.42 73.585 2.72 ;
      RECT 63.02 3.535 63.575 3.865 ;
      RECT 63.02 1.87 63.32 3.865 ;
      RECT 59.085 2.975 59.64 3.305 ;
      RECT 59.34 1.87 59.64 3.305 ;
      RECT 59.34 1.87 63.32 2.17 ;
      RECT 62.49 7.055 62.865 7.425 ;
      RECT 62.49 7.095 63.495 7.395 ;
      RECT 63.195 4.405 63.495 7.395 ;
      RECT 53.365 4.405 63.495 4.705 ;
      RECT 57.87 2.415 58.17 4.705 ;
      RECT 56.435 2.975 56.735 4.705 ;
      RECT 53.365 2.42 53.665 4.705 ;
      RECT 56.405 2.975 57.135 3.305 ;
      RECT 57.845 2.415 58.575 2.745 ;
      RECT 54.295 2.415 55.025 2.745 ;
      RECT 53.365 2.42 55.025 2.72 ;
      RECT 44.46 3.535 45.015 3.865 ;
      RECT 44.46 1.87 44.76 3.865 ;
      RECT 40.525 2.975 41.08 3.305 ;
      RECT 40.78 1.87 41.08 3.305 ;
      RECT 40.78 1.87 44.76 2.17 ;
      RECT 43.93 7.055 44.305 7.425 ;
      RECT 43.93 7.095 44.935 7.395 ;
      RECT 44.635 4.405 44.935 7.395 ;
      RECT 34.805 4.405 44.935 4.705 ;
      RECT 39.31 2.415 39.61 4.705 ;
      RECT 37.875 2.975 38.175 4.705 ;
      RECT 34.805 2.42 35.105 4.705 ;
      RECT 37.845 2.975 38.575 3.305 ;
      RECT 39.285 2.415 40.015 2.745 ;
      RECT 35.735 2.415 36.465 2.745 ;
      RECT 34.805 2.42 36.465 2.72 ;
      RECT 25.9 3.535 26.455 3.865 ;
      RECT 25.9 1.87 26.2 3.865 ;
      RECT 21.965 2.975 22.52 3.305 ;
      RECT 22.22 1.87 22.52 3.305 ;
      RECT 22.22 1.87 26.2 2.17 ;
      RECT 25.37 7.055 25.745 7.425 ;
      RECT 25.37 7.095 26.375 7.395 ;
      RECT 26.075 4.405 26.375 7.395 ;
      RECT 16.245 4.405 26.375 4.705 ;
      RECT 20.75 2.415 21.05 4.705 ;
      RECT 19.315 2.975 19.615 4.705 ;
      RECT 16.245 2.42 16.545 4.705 ;
      RECT 19.285 2.975 20.015 3.305 ;
      RECT 20.725 2.415 21.455 2.745 ;
      RECT 17.175 2.415 17.905 2.745 ;
      RECT 16.245 2.42 17.905 2.72 ;
      RECT 7.34 3.535 7.895 3.865 ;
      RECT 7.34 1.87 7.64 3.865 ;
      RECT 3.405 2.975 3.96 3.305 ;
      RECT 3.66 1.87 3.96 3.305 ;
      RECT 3.66 1.87 7.64 2.17 ;
      RECT 6.81 7.055 7.185 7.425 ;
      RECT 6.81 7.095 7.815 7.395 ;
      RECT 7.515 4.405 7.815 7.395 ;
      RECT -2.315 4.405 7.815 4.705 ;
      RECT 2.19 2.415 2.49 4.705 ;
      RECT 0.755 2.975 1.055 4.705 ;
      RECT -2.315 2.42 -2.015 4.705 ;
      RECT 0.725 2.975 1.455 3.305 ;
      RECT 2.165 2.415 2.895 2.745 ;
      RECT -1.385 2.415 -0.655 2.745 ;
      RECT -2.315 2.42 -0.655 2.72 ;
      RECT 82.765 1.855 83.495 2.185 ;
      RECT 80.545 3.535 81.275 3.865 ;
      RECT 78.845 3.535 79.575 3.865 ;
      RECT 73.89 2.415 74.62 2.745 ;
      RECT 72.525 3.535 73.255 3.865 ;
      RECT 64.205 1.855 64.935 2.185 ;
      RECT 61.985 3.535 62.715 3.865 ;
      RECT 60.285 3.535 61.015 3.865 ;
      RECT 55.33 2.415 56.06 2.745 ;
      RECT 53.965 3.535 54.695 3.865 ;
      RECT 45.645 1.855 46.375 2.185 ;
      RECT 43.425 3.535 44.155 3.865 ;
      RECT 41.725 3.535 42.455 3.865 ;
      RECT 36.77 2.415 37.5 2.745 ;
      RECT 35.405 3.535 36.135 3.865 ;
      RECT 27.085 1.855 27.815 2.185 ;
      RECT 24.865 3.535 25.595 3.865 ;
      RECT 23.165 3.535 23.895 3.865 ;
      RECT 18.21 2.415 18.94 2.745 ;
      RECT 16.845 3.535 17.575 3.865 ;
      RECT 8.525 1.855 9.255 2.185 ;
      RECT 6.305 3.535 7.035 3.865 ;
      RECT 4.605 3.535 5.335 3.865 ;
      RECT -0.35 2.415 0.38 2.745 ;
      RECT -1.715 3.535 -0.985 3.865 ;
    LAYER via2 ;
      RECT 82.83 1.92 83.03 2.12 ;
      RECT 81.87 3.6 82.07 3.8 ;
      RECT 81.135 7.14 81.335 7.34 ;
      RECT 80.87 3.6 81.07 3.8 ;
      RECT 78.91 3.6 79.11 3.8 ;
      RECT 77.71 3.04 77.91 3.24 ;
      RECT 76.47 2.48 76.67 2.68 ;
      RECT 75.03 3.04 75.23 3.24 ;
      RECT 74.29 2.48 74.49 2.68 ;
      RECT 73.07 2.48 73.27 2.68 ;
      RECT 72.59 3.6 72.79 3.8 ;
      RECT 64.27 1.92 64.47 2.12 ;
      RECT 63.31 3.6 63.51 3.8 ;
      RECT 62.575 7.14 62.775 7.34 ;
      RECT 62.31 3.6 62.51 3.8 ;
      RECT 60.35 3.6 60.55 3.8 ;
      RECT 59.15 3.04 59.35 3.24 ;
      RECT 57.91 2.48 58.11 2.68 ;
      RECT 56.47 3.04 56.67 3.24 ;
      RECT 55.73 2.48 55.93 2.68 ;
      RECT 54.51 2.48 54.71 2.68 ;
      RECT 54.03 3.6 54.23 3.8 ;
      RECT 45.71 1.92 45.91 2.12 ;
      RECT 44.75 3.6 44.95 3.8 ;
      RECT 44.015 7.14 44.215 7.34 ;
      RECT 43.75 3.6 43.95 3.8 ;
      RECT 41.79 3.6 41.99 3.8 ;
      RECT 40.59 3.04 40.79 3.24 ;
      RECT 39.35 2.48 39.55 2.68 ;
      RECT 37.91 3.04 38.11 3.24 ;
      RECT 37.17 2.48 37.37 2.68 ;
      RECT 35.95 2.48 36.15 2.68 ;
      RECT 35.47 3.6 35.67 3.8 ;
      RECT 27.15 1.92 27.35 2.12 ;
      RECT 26.19 3.6 26.39 3.8 ;
      RECT 25.455 7.14 25.655 7.34 ;
      RECT 25.19 3.6 25.39 3.8 ;
      RECT 23.23 3.6 23.43 3.8 ;
      RECT 22.03 3.04 22.23 3.24 ;
      RECT 20.79 2.48 20.99 2.68 ;
      RECT 19.35 3.04 19.55 3.24 ;
      RECT 18.61 2.48 18.81 2.68 ;
      RECT 17.39 2.48 17.59 2.68 ;
      RECT 16.91 3.6 17.11 3.8 ;
      RECT 8.59 1.92 8.79 2.12 ;
      RECT 7.63 3.6 7.83 3.8 ;
      RECT 6.895 7.14 7.095 7.34 ;
      RECT 6.63 3.6 6.83 3.8 ;
      RECT 4.67 3.6 4.87 3.8 ;
      RECT 3.47 3.04 3.67 3.24 ;
      RECT 2.23 2.48 2.43 2.68 ;
      RECT 0.79 3.04 0.99 3.24 ;
      RECT 0.05 2.48 0.25 2.68 ;
      RECT -1.17 2.48 -0.97 2.68 ;
      RECT -1.65 3.6 -1.45 3.8 ;
    LAYER met2 ;
      RECT -4.28 8.4 89.72 8.57 ;
      RECT 89.55 7.275 89.72 8.57 ;
      RECT -4.28 6.255 -4.11 8.57 ;
      RECT 89.52 7.275 89.87 7.625 ;
      RECT -4.34 6.255 -4.05 6.605 ;
      RECT 86.36 6.22 86.68 6.545 ;
      RECT 86.39 5.695 86.56 6.545 ;
      RECT 86.39 5.695 86.565 6.045 ;
      RECT 86.39 5.695 87.365 5.87 ;
      RECT 87.19 1.965 87.365 5.87 ;
      RECT 87.135 1.965 87.485 2.315 ;
      RECT 87.16 6.655 87.485 6.98 ;
      RECT 86.045 6.745 87.485 6.915 ;
      RECT 86.045 2.395 86.205 6.915 ;
      RECT 86.36 2.365 86.68 2.685 ;
      RECT 86.045 2.395 86.68 2.565 ;
      RECT 85.31 5.845 85.65 6.195 ;
      RECT 85.395 2.705 85.565 6.195 ;
      RECT 85.32 2.705 85.66 3.055 ;
      RECT 78.925 4.135 85.015 4.325 ;
      RECT 84.845 3.145 85.015 4.325 ;
      RECT 84.825 3.15 85.015 4.325 ;
      RECT 78.925 3.515 79.095 4.325 ;
      RECT 78.87 3.515 79.15 3.885 ;
      RECT 78.94 3.07 79.08 4.325 ;
      RECT 84.755 3.15 85.095 3.5 ;
      RECT 78.75 2.955 79.03 3.325 ;
      RECT 78.46 3.07 79.08 3.21 ;
      RECT 78.46 1.86 78.6 3.21 ;
      RECT 78.4 1.86 78.66 2.18 ;
      RECT 70.935 6.655 71.285 7.005 ;
      RECT 81.72 6.61 82.07 6.96 ;
      RECT 70.935 6.685 82.07 6.885 ;
      RECT 81.36 2.98 81.62 3.3 ;
      RECT 81.42 1.86 81.56 3.3 ;
      RECT 81.36 1.86 81.62 2.18 ;
      RECT 80.36 3.54 80.62 3.86 ;
      RECT 80.36 2.955 80.56 3.86 ;
      RECT 80.3 1.86 80.44 3.49 ;
      RECT 80.3 2.955 80.8 3.325 ;
      RECT 80.24 1.86 80.5 2.18 ;
      RECT 79.88 3.54 80.14 3.86 ;
      RECT 79.94 1.95 80.08 3.86 ;
      RECT 79.64 1.95 80.08 2.18 ;
      RECT 79.64 1.86 79.9 2.18 ;
      RECT 79.4 2.42 79.66 2.74 ;
      RECT 78.82 2.51 79.66 2.65 ;
      RECT 78.82 1.57 78.96 2.65 ;
      RECT 75.48 1.86 75.74 2.18 ;
      RECT 75.48 1.95 76.52 2.09 ;
      RECT 76.38 1.57 76.52 2.09 ;
      RECT 76.38 1.57 78.96 1.71 ;
      RECT 77.67 2.955 77.95 3.325 ;
      RECT 77.74 1.86 77.88 3.325 ;
      RECT 77.68 1.86 77.94 2.18 ;
      RECT 77.32 3.54 77.58 3.86 ;
      RECT 77.38 1.95 77.52 3.86 ;
      RECT 76.96 1.86 77.22 2.18 ;
      RECT 76.96 1.95 77.52 2.09 ;
      RECT 74.99 2.955 75.27 3.325 ;
      RECT 76.96 2.98 77.22 3.3 ;
      RECT 74.64 2.98 75.27 3.3 ;
      RECT 74.64 3.07 77.22 3.21 ;
      RECT 76.43 2.395 76.71 2.765 ;
      RECT 76.43 2.42 76.96 2.74 ;
      RECT 74 2.98 74.26 3.3 ;
      RECT 73.94 2.51 74.08 3.21 ;
      RECT 74.25 2.395 74.53 2.765 ;
      RECT 75.72 2.42 75.98 2.74 ;
      RECT 73.94 2.51 75.98 2.65 ;
      RECT 74.345 1 74.515 2.765 ;
      RECT 74.32 1 74.66 1.34 ;
      RECT 73.52 2.98 73.78 3.3 ;
      RECT 73.58 1.86 73.72 3.3 ;
      RECT 73.52 1.86 73.78 2.18 ;
      RECT 72.55 3.515 72.83 3.885 ;
      RECT 72.56 3.26 72.82 3.885 ;
      RECT 67.8 6.22 68.12 6.545 ;
      RECT 67.83 5.695 68 6.545 ;
      RECT 67.83 5.695 68.005 6.045 ;
      RECT 67.83 5.695 68.805 5.87 ;
      RECT 68.63 1.965 68.805 5.87 ;
      RECT 68.575 1.965 68.925 2.315 ;
      RECT 68.6 6.655 68.925 6.98 ;
      RECT 67.485 6.745 68.925 6.915 ;
      RECT 67.485 2.395 67.645 6.915 ;
      RECT 67.8 2.365 68.12 2.685 ;
      RECT 67.485 2.395 68.12 2.565 ;
      RECT 66.75 5.845 67.09 6.195 ;
      RECT 66.835 2.705 67.005 6.195 ;
      RECT 66.76 2.705 67.1 3.055 ;
      RECT 60.365 4.135 66.455 4.325 ;
      RECT 66.285 3.145 66.455 4.325 ;
      RECT 66.265 3.15 66.455 4.325 ;
      RECT 60.365 3.515 60.535 4.325 ;
      RECT 60.31 3.515 60.59 3.885 ;
      RECT 60.38 3.07 60.52 4.325 ;
      RECT 66.195 3.15 66.535 3.5 ;
      RECT 60.19 2.955 60.47 3.325 ;
      RECT 59.9 3.07 60.52 3.21 ;
      RECT 59.9 1.86 60.04 3.21 ;
      RECT 59.84 1.86 60.1 2.18 ;
      RECT 52.375 6.655 52.725 7.005 ;
      RECT 63.16 6.61 63.51 6.96 ;
      RECT 52.375 6.685 63.51 6.885 ;
      RECT 62.8 2.98 63.06 3.3 ;
      RECT 62.86 1.86 63 3.3 ;
      RECT 62.8 1.86 63.06 2.18 ;
      RECT 61.8 3.54 62.06 3.86 ;
      RECT 61.8 2.955 62 3.86 ;
      RECT 61.74 1.86 61.88 3.49 ;
      RECT 61.74 2.955 62.24 3.325 ;
      RECT 61.68 1.86 61.94 2.18 ;
      RECT 61.32 3.54 61.58 3.86 ;
      RECT 61.38 1.95 61.52 3.86 ;
      RECT 61.08 1.95 61.52 2.18 ;
      RECT 61.08 1.86 61.34 2.18 ;
      RECT 60.84 2.42 61.1 2.74 ;
      RECT 60.26 2.51 61.1 2.65 ;
      RECT 60.26 1.57 60.4 2.65 ;
      RECT 56.92 1.86 57.18 2.18 ;
      RECT 56.92 1.95 57.96 2.09 ;
      RECT 57.82 1.57 57.96 2.09 ;
      RECT 57.82 1.57 60.4 1.71 ;
      RECT 59.11 2.955 59.39 3.325 ;
      RECT 59.18 1.86 59.32 3.325 ;
      RECT 59.12 1.86 59.38 2.18 ;
      RECT 58.76 3.54 59.02 3.86 ;
      RECT 58.82 1.95 58.96 3.86 ;
      RECT 58.4 1.86 58.66 2.18 ;
      RECT 58.4 1.95 58.96 2.09 ;
      RECT 56.43 2.955 56.71 3.325 ;
      RECT 58.4 2.98 58.66 3.3 ;
      RECT 56.08 2.98 56.71 3.3 ;
      RECT 56.08 3.07 58.66 3.21 ;
      RECT 57.87 2.395 58.15 2.765 ;
      RECT 57.87 2.42 58.4 2.74 ;
      RECT 55.44 2.98 55.7 3.3 ;
      RECT 55.38 2.51 55.52 3.21 ;
      RECT 55.69 2.395 55.97 2.765 ;
      RECT 57.16 2.42 57.42 2.74 ;
      RECT 55.38 2.51 57.42 2.65 ;
      RECT 55.785 1 55.955 2.765 ;
      RECT 55.76 1 56.1 1.34 ;
      RECT 54.96 2.98 55.22 3.3 ;
      RECT 55.02 1.86 55.16 3.3 ;
      RECT 54.96 1.86 55.22 2.18 ;
      RECT 53.99 3.515 54.27 3.885 ;
      RECT 54 3.26 54.26 3.885 ;
      RECT 49.24 6.22 49.56 6.545 ;
      RECT 49.27 5.695 49.44 6.545 ;
      RECT 49.27 5.695 49.445 6.045 ;
      RECT 49.27 5.695 50.245 5.87 ;
      RECT 50.07 1.965 50.245 5.87 ;
      RECT 50.015 1.965 50.365 2.315 ;
      RECT 50.04 6.655 50.365 6.98 ;
      RECT 48.925 6.745 50.365 6.915 ;
      RECT 48.925 2.395 49.085 6.915 ;
      RECT 49.24 2.365 49.56 2.685 ;
      RECT 48.925 2.395 49.56 2.565 ;
      RECT 48.19 5.845 48.53 6.195 ;
      RECT 48.275 2.705 48.445 6.195 ;
      RECT 48.2 2.705 48.54 3.055 ;
      RECT 41.805 4.135 47.895 4.325 ;
      RECT 47.725 3.145 47.895 4.325 ;
      RECT 47.705 3.15 47.895 4.325 ;
      RECT 41.805 3.515 41.975 4.325 ;
      RECT 41.75 3.515 42.03 3.885 ;
      RECT 41.82 3.07 41.96 4.325 ;
      RECT 47.635 3.15 47.975 3.5 ;
      RECT 41.63 2.955 41.91 3.325 ;
      RECT 41.34 3.07 41.96 3.21 ;
      RECT 41.34 1.86 41.48 3.21 ;
      RECT 41.28 1.86 41.54 2.18 ;
      RECT 33.86 6.66 34.21 7.01 ;
      RECT 44.6 6.615 44.95 6.965 ;
      RECT 33.86 6.69 44.95 6.89 ;
      RECT 44.24 2.98 44.5 3.3 ;
      RECT 44.3 1.86 44.44 3.3 ;
      RECT 44.24 1.86 44.5 2.18 ;
      RECT 43.24 3.54 43.5 3.86 ;
      RECT 43.24 2.955 43.44 3.86 ;
      RECT 43.18 1.86 43.32 3.49 ;
      RECT 43.18 2.955 43.68 3.325 ;
      RECT 43.12 1.86 43.38 2.18 ;
      RECT 42.76 3.54 43.02 3.86 ;
      RECT 42.82 1.95 42.96 3.86 ;
      RECT 42.52 1.95 42.96 2.18 ;
      RECT 42.52 1.86 42.78 2.18 ;
      RECT 42.28 2.42 42.54 2.74 ;
      RECT 41.7 2.51 42.54 2.65 ;
      RECT 41.7 1.57 41.84 2.65 ;
      RECT 38.36 1.86 38.62 2.18 ;
      RECT 38.36 1.95 39.4 2.09 ;
      RECT 39.26 1.57 39.4 2.09 ;
      RECT 39.26 1.57 41.84 1.71 ;
      RECT 40.55 2.955 40.83 3.325 ;
      RECT 40.62 1.86 40.76 3.325 ;
      RECT 40.56 1.86 40.82 2.18 ;
      RECT 40.2 3.54 40.46 3.86 ;
      RECT 40.26 1.95 40.4 3.86 ;
      RECT 39.84 1.86 40.1 2.18 ;
      RECT 39.84 1.95 40.4 2.09 ;
      RECT 37.87 2.955 38.15 3.325 ;
      RECT 39.84 2.98 40.1 3.3 ;
      RECT 37.52 2.98 38.15 3.3 ;
      RECT 37.52 3.07 40.1 3.21 ;
      RECT 39.31 2.395 39.59 2.765 ;
      RECT 39.31 2.42 39.84 2.74 ;
      RECT 36.88 2.98 37.14 3.3 ;
      RECT 36.82 2.51 36.96 3.21 ;
      RECT 37.13 2.395 37.41 2.765 ;
      RECT 38.6 2.42 38.86 2.74 ;
      RECT 36.82 2.51 38.86 2.65 ;
      RECT 37.225 1 37.395 2.765 ;
      RECT 37.2 1 37.54 1.34 ;
      RECT 36.4 2.98 36.66 3.3 ;
      RECT 36.46 1.86 36.6 3.3 ;
      RECT 36.4 1.86 36.66 2.18 ;
      RECT 35.43 3.515 35.71 3.885 ;
      RECT 35.44 3.26 35.7 3.885 ;
      RECT 30.68 6.22 31 6.545 ;
      RECT 30.71 5.695 30.88 6.545 ;
      RECT 30.71 5.695 30.885 6.045 ;
      RECT 30.71 5.695 31.685 5.87 ;
      RECT 31.51 1.965 31.685 5.87 ;
      RECT 31.455 1.965 31.805 2.315 ;
      RECT 31.48 6.655 31.805 6.98 ;
      RECT 30.365 6.745 31.805 6.915 ;
      RECT 30.365 2.395 30.525 6.915 ;
      RECT 30.68 2.365 31 2.685 ;
      RECT 30.365 2.395 31 2.565 ;
      RECT 29.63 5.845 29.97 6.195 ;
      RECT 29.715 2.705 29.885 6.195 ;
      RECT 29.64 2.705 29.98 3.055 ;
      RECT 23.245 4.135 29.335 4.325 ;
      RECT 29.165 3.145 29.335 4.325 ;
      RECT 29.145 3.15 29.335 4.325 ;
      RECT 23.245 3.515 23.415 4.325 ;
      RECT 23.19 3.515 23.47 3.885 ;
      RECT 23.26 3.07 23.4 4.325 ;
      RECT 29.075 3.15 29.415 3.5 ;
      RECT 23.07 2.955 23.35 3.325 ;
      RECT 22.78 3.07 23.4 3.21 ;
      RECT 22.78 1.86 22.92 3.21 ;
      RECT 22.72 1.86 22.98 2.18 ;
      RECT 15.3 6.655 15.65 7.005 ;
      RECT 26.045 6.61 26.395 6.96 ;
      RECT 15.3 6.685 26.395 6.885 ;
      RECT 25.68 2.98 25.94 3.3 ;
      RECT 25.74 1.86 25.88 3.3 ;
      RECT 25.68 1.86 25.94 2.18 ;
      RECT 24.68 3.54 24.94 3.86 ;
      RECT 24.68 2.955 24.88 3.86 ;
      RECT 24.62 1.86 24.76 3.49 ;
      RECT 24.62 2.955 25.12 3.325 ;
      RECT 24.56 1.86 24.82 2.18 ;
      RECT 24.2 3.54 24.46 3.86 ;
      RECT 24.26 1.95 24.4 3.86 ;
      RECT 23.96 1.95 24.4 2.18 ;
      RECT 23.96 1.86 24.22 2.18 ;
      RECT 23.72 2.42 23.98 2.74 ;
      RECT 23.14 2.51 23.98 2.65 ;
      RECT 23.14 1.57 23.28 2.65 ;
      RECT 19.8 1.86 20.06 2.18 ;
      RECT 19.8 1.95 20.84 2.09 ;
      RECT 20.7 1.57 20.84 2.09 ;
      RECT 20.7 1.57 23.28 1.71 ;
      RECT 21.99 2.955 22.27 3.325 ;
      RECT 22.06 1.86 22.2 3.325 ;
      RECT 22 1.86 22.26 2.18 ;
      RECT 21.64 3.54 21.9 3.86 ;
      RECT 21.7 1.95 21.84 3.86 ;
      RECT 21.28 1.86 21.54 2.18 ;
      RECT 21.28 1.95 21.84 2.09 ;
      RECT 19.31 2.955 19.59 3.325 ;
      RECT 21.28 2.98 21.54 3.3 ;
      RECT 18.96 2.98 19.59 3.3 ;
      RECT 18.96 3.07 21.54 3.21 ;
      RECT 20.75 2.395 21.03 2.765 ;
      RECT 20.75 2.42 21.28 2.74 ;
      RECT 18.32 2.98 18.58 3.3 ;
      RECT 18.26 2.51 18.4 3.21 ;
      RECT 18.57 2.395 18.85 2.765 ;
      RECT 20.04 2.42 20.3 2.74 ;
      RECT 18.26 2.51 20.3 2.65 ;
      RECT 18.665 1 18.835 2.765 ;
      RECT 18.64 1 18.98 1.34 ;
      RECT 17.84 2.98 18.1 3.3 ;
      RECT 17.9 1.86 18.04 3.3 ;
      RECT 17.84 1.86 18.1 2.18 ;
      RECT 16.87 3.515 17.15 3.885 ;
      RECT 16.88 3.26 17.14 3.885 ;
      RECT 12.12 6.22 12.44 6.545 ;
      RECT 12.15 5.695 12.32 6.545 ;
      RECT 12.15 5.695 12.325 6.045 ;
      RECT 12.15 5.695 13.125 5.87 ;
      RECT 12.95 1.965 13.125 5.87 ;
      RECT 12.895 1.965 13.245 2.315 ;
      RECT 12.92 6.655 13.245 6.98 ;
      RECT 11.805 6.745 13.245 6.915 ;
      RECT 11.805 2.395 11.965 6.915 ;
      RECT 12.12 2.365 12.44 2.685 ;
      RECT 11.805 2.395 12.44 2.565 ;
      RECT 11.07 5.845 11.41 6.195 ;
      RECT 11.155 2.705 11.325 6.195 ;
      RECT 11.08 2.705 11.42 3.055 ;
      RECT 4.685 4.135 10.775 4.325 ;
      RECT 10.605 3.145 10.775 4.325 ;
      RECT 10.585 3.15 10.775 4.325 ;
      RECT 4.685 3.515 4.855 4.325 ;
      RECT 4.63 3.515 4.91 3.885 ;
      RECT 4.7 3.07 4.84 4.325 ;
      RECT 10.515 3.15 10.855 3.5 ;
      RECT 4.51 2.955 4.79 3.325 ;
      RECT 4.22 3.07 4.84 3.21 ;
      RECT 4.22 1.86 4.36 3.21 ;
      RECT 4.16 1.86 4.42 2.18 ;
      RECT -3.965 6.995 -3.675 7.345 ;
      RECT -3.965 7.055 -2.775 7.225 ;
      RECT -2.945 6.685 -2.775 7.225 ;
      RECT 7.485 6.605 7.835 6.955 ;
      RECT -2.945 6.685 7.835 6.855 ;
      RECT 7.12 2.98 7.38 3.3 ;
      RECT 7.18 1.86 7.32 3.3 ;
      RECT 7.12 1.86 7.38 2.18 ;
      RECT 6.12 3.54 6.38 3.86 ;
      RECT 6.12 2.955 6.32 3.86 ;
      RECT 6.06 1.86 6.2 3.49 ;
      RECT 6.06 2.955 6.56 3.325 ;
      RECT 6 1.86 6.26 2.18 ;
      RECT 5.64 3.54 5.9 3.86 ;
      RECT 5.7 1.95 5.84 3.86 ;
      RECT 5.4 1.95 5.84 2.18 ;
      RECT 5.4 1.86 5.66 2.18 ;
      RECT 5.16 2.42 5.42 2.74 ;
      RECT 4.58 2.51 5.42 2.65 ;
      RECT 4.58 1.57 4.72 2.65 ;
      RECT 1.24 1.86 1.5 2.18 ;
      RECT 1.24 1.95 2.28 2.09 ;
      RECT 2.14 1.57 2.28 2.09 ;
      RECT 2.14 1.57 4.72 1.71 ;
      RECT 3.43 2.955 3.71 3.325 ;
      RECT 3.5 1.86 3.64 3.325 ;
      RECT 3.44 1.86 3.7 2.18 ;
      RECT 3.08 3.54 3.34 3.86 ;
      RECT 3.14 1.95 3.28 3.86 ;
      RECT 2.72 1.86 2.98 2.18 ;
      RECT 2.72 1.95 3.28 2.09 ;
      RECT 0.75 2.955 1.03 3.325 ;
      RECT 2.72 2.98 2.98 3.3 ;
      RECT 0.4 2.98 1.03 3.3 ;
      RECT 0.4 3.07 2.98 3.21 ;
      RECT 2.19 2.395 2.47 2.765 ;
      RECT 2.19 2.42 2.72 2.74 ;
      RECT -0.24 2.98 0.02 3.3 ;
      RECT -0.3 2.51 -0.16 3.21 ;
      RECT 0.01 2.395 0.29 2.765 ;
      RECT 1.48 2.42 1.74 2.74 ;
      RECT -0.3 2.51 1.74 2.65 ;
      RECT 0.105 1 0.275 2.765 ;
      RECT 0.08 1 0.42 1.34 ;
      RECT -0.72 2.98 -0.46 3.3 ;
      RECT -0.66 1.86 -0.52 3.3 ;
      RECT -0.72 1.86 -0.46 2.18 ;
      RECT -1.69 3.515 -1.41 3.885 ;
      RECT -1.68 3.26 -1.42 3.885 ;
      RECT 82.79 1.835 83.07 2.205 ;
      RECT 81.83 3.515 82.11 3.885 ;
      RECT 81.05 7.055 81.425 7.425 ;
      RECT 80.83 3.515 81.11 3.885 ;
      RECT 73.03 2.395 73.31 2.765 ;
      RECT 64.23 1.835 64.51 2.205 ;
      RECT 63.27 3.515 63.55 3.885 ;
      RECT 62.49 7.055 62.865 7.425 ;
      RECT 62.27 3.515 62.55 3.885 ;
      RECT 54.47 2.395 54.75 2.765 ;
      RECT 45.67 1.835 45.95 2.205 ;
      RECT 44.71 3.515 44.99 3.885 ;
      RECT 43.93 7.055 44.305 7.425 ;
      RECT 43.71 3.515 43.99 3.885 ;
      RECT 35.91 2.395 36.19 2.765 ;
      RECT 27.11 1.835 27.39 2.205 ;
      RECT 26.15 3.515 26.43 3.885 ;
      RECT 25.37 7.055 25.745 7.425 ;
      RECT 25.15 3.515 25.43 3.885 ;
      RECT 17.35 2.395 17.63 2.765 ;
      RECT 8.55 1.835 8.83 2.205 ;
      RECT 7.59 3.515 7.87 3.885 ;
      RECT 6.81 7.055 7.185 7.425 ;
      RECT 6.59 3.515 6.87 3.885 ;
      RECT -1.21 2.395 -0.93 2.765 ;
    LAYER via1 ;
      RECT 89.62 7.375 89.77 7.525 ;
      RECT 87.25 6.74 87.4 6.89 ;
      RECT 87.235 2.065 87.385 2.215 ;
      RECT 86.445 2.45 86.595 2.6 ;
      RECT 86.445 6.325 86.595 6.475 ;
      RECT 85.42 2.805 85.57 2.955 ;
      RECT 85.41 5.945 85.56 6.095 ;
      RECT 84.855 3.25 85.005 3.4 ;
      RECT 82.855 1.945 83.005 2.095 ;
      RECT 81.895 3.625 82.045 3.775 ;
      RECT 81.82 6.71 81.97 6.86 ;
      RECT 81.415 1.945 81.565 2.095 ;
      RECT 81.415 3.065 81.565 3.215 ;
      RECT 81.16 7.165 81.31 7.315 ;
      RECT 80.895 3.625 81.045 3.775 ;
      RECT 80.415 3.625 80.565 3.775 ;
      RECT 80.295 1.945 80.445 2.095 ;
      RECT 79.935 3.625 80.085 3.775 ;
      RECT 79.695 1.945 79.845 2.095 ;
      RECT 79.455 2.505 79.605 2.655 ;
      RECT 78.935 3.625 79.085 3.775 ;
      RECT 78.455 1.945 78.605 2.095 ;
      RECT 77.735 1.945 77.885 2.095 ;
      RECT 77.735 3.065 77.885 3.215 ;
      RECT 77.375 3.625 77.525 3.775 ;
      RECT 77.015 1.945 77.165 2.095 ;
      RECT 77.015 3.065 77.165 3.215 ;
      RECT 76.755 2.505 76.905 2.655 ;
      RECT 75.775 2.505 75.925 2.655 ;
      RECT 75.535 1.945 75.685 2.095 ;
      RECT 74.695 3.065 74.845 3.215 ;
      RECT 74.415 1.095 74.565 1.245 ;
      RECT 74.055 3.065 74.205 3.215 ;
      RECT 73.575 1.945 73.725 2.095 ;
      RECT 73.575 3.065 73.725 3.215 ;
      RECT 73.095 2.505 73.245 2.655 ;
      RECT 72.615 3.345 72.765 3.495 ;
      RECT 71.035 6.755 71.185 6.905 ;
      RECT 68.69 6.74 68.84 6.89 ;
      RECT 68.675 2.065 68.825 2.215 ;
      RECT 67.885 2.45 68.035 2.6 ;
      RECT 67.885 6.325 68.035 6.475 ;
      RECT 66.86 2.805 67.01 2.955 ;
      RECT 66.85 5.945 67 6.095 ;
      RECT 66.295 3.25 66.445 3.4 ;
      RECT 64.295 1.945 64.445 2.095 ;
      RECT 63.335 3.625 63.485 3.775 ;
      RECT 63.26 6.71 63.41 6.86 ;
      RECT 62.855 1.945 63.005 2.095 ;
      RECT 62.855 3.065 63.005 3.215 ;
      RECT 62.6 7.165 62.75 7.315 ;
      RECT 62.335 3.625 62.485 3.775 ;
      RECT 61.855 3.625 62.005 3.775 ;
      RECT 61.735 1.945 61.885 2.095 ;
      RECT 61.375 3.625 61.525 3.775 ;
      RECT 61.135 1.945 61.285 2.095 ;
      RECT 60.895 2.505 61.045 2.655 ;
      RECT 60.375 3.625 60.525 3.775 ;
      RECT 59.895 1.945 60.045 2.095 ;
      RECT 59.175 1.945 59.325 2.095 ;
      RECT 59.175 3.065 59.325 3.215 ;
      RECT 58.815 3.625 58.965 3.775 ;
      RECT 58.455 1.945 58.605 2.095 ;
      RECT 58.455 3.065 58.605 3.215 ;
      RECT 58.195 2.505 58.345 2.655 ;
      RECT 57.215 2.505 57.365 2.655 ;
      RECT 56.975 1.945 57.125 2.095 ;
      RECT 56.135 3.065 56.285 3.215 ;
      RECT 55.855 1.095 56.005 1.245 ;
      RECT 55.495 3.065 55.645 3.215 ;
      RECT 55.015 1.945 55.165 2.095 ;
      RECT 55.015 3.065 55.165 3.215 ;
      RECT 54.535 2.505 54.685 2.655 ;
      RECT 54.055 3.345 54.205 3.495 ;
      RECT 52.475 6.755 52.625 6.905 ;
      RECT 50.13 6.74 50.28 6.89 ;
      RECT 50.115 2.065 50.265 2.215 ;
      RECT 49.325 2.45 49.475 2.6 ;
      RECT 49.325 6.325 49.475 6.475 ;
      RECT 48.3 2.805 48.45 2.955 ;
      RECT 48.29 5.945 48.44 6.095 ;
      RECT 47.735 3.25 47.885 3.4 ;
      RECT 45.735 1.945 45.885 2.095 ;
      RECT 44.775 3.625 44.925 3.775 ;
      RECT 44.7 6.715 44.85 6.865 ;
      RECT 44.295 1.945 44.445 2.095 ;
      RECT 44.295 3.065 44.445 3.215 ;
      RECT 44.04 7.165 44.19 7.315 ;
      RECT 43.775 3.625 43.925 3.775 ;
      RECT 43.295 3.625 43.445 3.775 ;
      RECT 43.175 1.945 43.325 2.095 ;
      RECT 42.815 3.625 42.965 3.775 ;
      RECT 42.575 1.945 42.725 2.095 ;
      RECT 42.335 2.505 42.485 2.655 ;
      RECT 41.815 3.625 41.965 3.775 ;
      RECT 41.335 1.945 41.485 2.095 ;
      RECT 40.615 1.945 40.765 2.095 ;
      RECT 40.615 3.065 40.765 3.215 ;
      RECT 40.255 3.625 40.405 3.775 ;
      RECT 39.895 1.945 40.045 2.095 ;
      RECT 39.895 3.065 40.045 3.215 ;
      RECT 39.635 2.505 39.785 2.655 ;
      RECT 38.655 2.505 38.805 2.655 ;
      RECT 38.415 1.945 38.565 2.095 ;
      RECT 37.575 3.065 37.725 3.215 ;
      RECT 37.295 1.095 37.445 1.245 ;
      RECT 36.935 3.065 37.085 3.215 ;
      RECT 36.455 1.945 36.605 2.095 ;
      RECT 36.455 3.065 36.605 3.215 ;
      RECT 35.975 2.505 36.125 2.655 ;
      RECT 35.495 3.345 35.645 3.495 ;
      RECT 33.96 6.76 34.11 6.91 ;
      RECT 31.57 6.74 31.72 6.89 ;
      RECT 31.555 2.065 31.705 2.215 ;
      RECT 30.765 2.45 30.915 2.6 ;
      RECT 30.765 6.325 30.915 6.475 ;
      RECT 29.74 2.805 29.89 2.955 ;
      RECT 29.73 5.945 29.88 6.095 ;
      RECT 29.175 3.25 29.325 3.4 ;
      RECT 27.175 1.945 27.325 2.095 ;
      RECT 26.215 3.625 26.365 3.775 ;
      RECT 26.145 6.71 26.295 6.86 ;
      RECT 25.735 1.945 25.885 2.095 ;
      RECT 25.735 3.065 25.885 3.215 ;
      RECT 25.48 7.165 25.63 7.315 ;
      RECT 25.215 3.625 25.365 3.775 ;
      RECT 24.735 3.625 24.885 3.775 ;
      RECT 24.615 1.945 24.765 2.095 ;
      RECT 24.255 3.625 24.405 3.775 ;
      RECT 24.015 1.945 24.165 2.095 ;
      RECT 23.775 2.505 23.925 2.655 ;
      RECT 23.255 3.625 23.405 3.775 ;
      RECT 22.775 1.945 22.925 2.095 ;
      RECT 22.055 1.945 22.205 2.095 ;
      RECT 22.055 3.065 22.205 3.215 ;
      RECT 21.695 3.625 21.845 3.775 ;
      RECT 21.335 1.945 21.485 2.095 ;
      RECT 21.335 3.065 21.485 3.215 ;
      RECT 21.075 2.505 21.225 2.655 ;
      RECT 20.095 2.505 20.245 2.655 ;
      RECT 19.855 1.945 20.005 2.095 ;
      RECT 19.015 3.065 19.165 3.215 ;
      RECT 18.735 1.095 18.885 1.245 ;
      RECT 18.375 3.065 18.525 3.215 ;
      RECT 17.895 1.945 18.045 2.095 ;
      RECT 17.895 3.065 18.045 3.215 ;
      RECT 17.415 2.505 17.565 2.655 ;
      RECT 16.935 3.345 17.085 3.495 ;
      RECT 15.4 6.755 15.55 6.905 ;
      RECT 13.01 6.74 13.16 6.89 ;
      RECT 12.995 2.065 13.145 2.215 ;
      RECT 12.205 2.45 12.355 2.6 ;
      RECT 12.205 6.325 12.355 6.475 ;
      RECT 11.18 2.805 11.33 2.955 ;
      RECT 11.17 5.945 11.32 6.095 ;
      RECT 10.615 3.25 10.765 3.4 ;
      RECT 8.615 1.945 8.765 2.095 ;
      RECT 7.655 3.625 7.805 3.775 ;
      RECT 7.585 6.705 7.735 6.855 ;
      RECT 7.175 1.945 7.325 2.095 ;
      RECT 7.175 3.065 7.325 3.215 ;
      RECT 6.92 7.165 7.07 7.315 ;
      RECT 6.655 3.625 6.805 3.775 ;
      RECT 6.175 3.625 6.325 3.775 ;
      RECT 6.055 1.945 6.205 2.095 ;
      RECT 5.695 3.625 5.845 3.775 ;
      RECT 5.455 1.945 5.605 2.095 ;
      RECT 5.215 2.505 5.365 2.655 ;
      RECT 4.695 3.625 4.845 3.775 ;
      RECT 4.215 1.945 4.365 2.095 ;
      RECT 3.495 1.945 3.645 2.095 ;
      RECT 3.495 3.065 3.645 3.215 ;
      RECT 3.135 3.625 3.285 3.775 ;
      RECT 2.775 1.945 2.925 2.095 ;
      RECT 2.775 3.065 2.925 3.215 ;
      RECT 2.515 2.505 2.665 2.655 ;
      RECT 1.535 2.505 1.685 2.655 ;
      RECT 1.295 1.945 1.445 2.095 ;
      RECT 0.455 3.065 0.605 3.215 ;
      RECT 0.175 1.095 0.325 1.245 ;
      RECT -0.185 3.065 -0.035 3.215 ;
      RECT -0.665 1.945 -0.515 2.095 ;
      RECT -0.665 3.065 -0.515 3.215 ;
      RECT -1.145 2.505 -0.995 2.655 ;
      RECT -1.625 3.345 -1.475 3.495 ;
      RECT -3.895 7.095 -3.745 7.245 ;
      RECT -4.27 6.355 -4.12 6.505 ;
    LAYER met1 ;
      RECT 72.275 0 84.235 1.74 ;
      RECT 53.715 0 65.675 1.74 ;
      RECT 35.155 0 47.115 1.74 ;
      RECT 16.595 0 28.555 1.74 ;
      RECT -1.965 0 9.995 1.74 ;
      RECT 72.275 0 84.32 1.585 ;
      RECT 53.715 0 65.76 1.585 ;
      RECT 35.155 0 47.2 1.585 ;
      RECT 16.595 0 28.64 1.585 ;
      RECT -1.965 0 10.08 1.585 ;
      RECT -5.465 0 90.09 0.305 ;
      RECT 71.53 4.145 73.995 4.75 ;
      RECT 52.97 4.145 55.435 4.75 ;
      RECT 34.41 4.145 36.875 4.75 ;
      RECT 15.85 4.145 18.315 4.75 ;
      RECT -5.46 4.145 -0.245 4.75 ;
      RECT 72.275 4.135 90.09 4.745 ;
      RECT 53.715 4.135 71.53 4.745 ;
      RECT 35.155 4.135 52.97 4.745 ;
      RECT 16.595 4.135 34.41 4.745 ;
      RECT -1.965 4.135 15.85 4.745 ;
      RECT 72.275 3.98 84.235 4.745 ;
      RECT 53.715 3.98 65.675 4.745 ;
      RECT 35.155 3.98 47.115 4.745 ;
      RECT 16.595 3.98 28.555 4.745 ;
      RECT -1.965 3.98 9.995 4.745 ;
      RECT -5.465 8.575 90.09 8.88 ;
      RECT 80.28 6.315 80.45 8.88 ;
      RECT 61.72 6.315 61.89 8.88 ;
      RECT 43.16 6.315 43.33 8.88 ;
      RECT 24.6 6.315 24.77 8.88 ;
      RECT 6.04 6.315 6.21 8.88 ;
      RECT 80.715 6.285 81.005 6.515 ;
      RECT 62.155 6.285 62.445 6.515 ;
      RECT 43.595 6.285 43.885 6.515 ;
      RECT 25.035 6.285 25.325 6.515 ;
      RECT 6.475 6.285 6.765 6.515 ;
      RECT 80.28 6.315 81.005 6.485 ;
      RECT 61.72 6.315 62.445 6.485 ;
      RECT 43.16 6.315 43.885 6.485 ;
      RECT 24.6 6.315 25.325 6.485 ;
      RECT 6.04 6.315 6.765 6.485 ;
      RECT 89.49 7.765 89.78 7.995 ;
      RECT 89.55 6.285 89.72 7.995 ;
      RECT 89.52 7.275 89.87 7.625 ;
      RECT 89.49 6.285 89.78 6.515 ;
      RECT 89.49 2.365 89.78 2.595 ;
      RECT 89.55 0.885 89.72 2.595 ;
      RECT 89.49 0.885 89.78 1.115 ;
      RECT 89.08 2.735 89.41 2.965 ;
      RECT 89.08 2.765 89.58 2.935 ;
      RECT 89.08 2.395 89.27 2.965 ;
      RECT 88.5 2.365 88.79 2.595 ;
      RECT 88.5 2.395 89.27 2.565 ;
      RECT 88.56 0.885 88.73 2.595 ;
      RECT 88.5 0.885 88.79 1.115 ;
      RECT 88.5 7.765 88.79 7.995 ;
      RECT 88.56 6.285 88.73 7.995 ;
      RECT 88.5 6.285 88.79 6.515 ;
      RECT 88.5 6.325 89.35 6.485 ;
      RECT 89.18 5.915 89.35 6.485 ;
      RECT 88.5 6.32 88.89 6.485 ;
      RECT 89.12 5.915 89.41 6.145 ;
      RECT 89.12 5.945 89.58 6.115 ;
      RECT 88.13 2.735 88.42 2.965 ;
      RECT 88.13 2.765 88.59 2.935 ;
      RECT 88.19 1.655 88.355 2.965 ;
      RECT 86.705 1.625 86.995 1.855 ;
      RECT 86.705 1.655 88.355 1.825 ;
      RECT 86.765 0.885 86.935 1.855 ;
      RECT 86.705 0.885 86.995 1.115 ;
      RECT 86.705 7.765 86.995 7.995 ;
      RECT 86.765 7.025 86.935 7.995 ;
      RECT 86.765 7.12 88.355 7.29 ;
      RECT 88.185 5.915 88.355 7.29 ;
      RECT 86.705 7.025 86.995 7.255 ;
      RECT 88.13 5.915 88.42 6.145 ;
      RECT 88.13 5.945 88.59 6.115 ;
      RECT 84.755 3.15 85.095 3.5 ;
      RECT 84.845 2.025 85.015 3.5 ;
      RECT 87.135 1.965 87.485 2.315 ;
      RECT 84.845 2.025 87.485 2.195 ;
      RECT 87.16 6.655 87.485 6.98 ;
      RECT 81.72 6.61 82.07 6.96 ;
      RECT 87.135 6.655 87.485 6.885 ;
      RECT 81.52 6.655 82.07 6.885 ;
      RECT 81.35 6.685 87.485 6.855 ;
      RECT 86.36 2.365 86.68 2.685 ;
      RECT 86.33 2.365 86.68 2.595 ;
      RECT 86.16 2.395 86.68 2.565 ;
      RECT 86.36 6.255 86.68 6.545 ;
      RECT 86.33 6.285 86.68 6.515 ;
      RECT 86.16 6.315 86.68 6.485 ;
      RECT 85.32 2.705 85.66 3.055 ;
      RECT 85.32 2.765 85.795 2.935 ;
      RECT 85.31 5.845 85.65 6.195 ;
      RECT 79.72 5.915 80.01 6.145 ;
      RECT 79.72 5.945 85.795 6.115 ;
      RECT 81.81 3.57 82.13 3.83 ;
      RECT 83.1 2.745 83.24 3.605 ;
      RECT 81.9 3.465 83.24 3.605 ;
      RECT 81.9 3.025 82.04 3.83 ;
      RECT 81.825 3.025 82.115 3.255 ;
      RECT 83.025 2.745 83.315 2.975 ;
      RECT 82.545 3.025 82.835 3.255 ;
      RECT 82.74 1.95 82.88 3.21 ;
      RECT 82.77 1.89 83.09 2.15 ;
      RECT 79.37 2.45 79.69 2.71 ;
      RECT 82.065 2.465 82.355 2.695 ;
      RECT 79.46 2.37 82.28 2.51 ;
      RECT 81.33 1.89 81.65 2.15 ;
      RECT 81.825 1.905 82.115 2.135 ;
      RECT 81.33 1.95 82.115 2.09 ;
      RECT 81.33 3.01 81.65 3.27 ;
      RECT 81.33 2.79 81.56 3.27 ;
      RECT 80.825 2.745 81.115 2.975 ;
      RECT 80.825 2.79 81.56 2.93 ;
      RECT 81.09 7.765 81.38 7.995 ;
      RECT 81.15 7.025 81.32 7.995 ;
      RECT 81.05 7.055 81.43 7.425 ;
      RECT 81.09 7.025 81.38 7.425 ;
      RECT 79.85 3.57 80.17 3.83 ;
      RECT 79.385 3.585 79.675 3.815 ;
      RECT 79.385 3.63 80.17 3.77 ;
      RECT 78.145 2.465 78.435 2.695 ;
      RECT 78.145 2.51 79.08 2.65 ;
      RECT 78.94 1.95 79.08 2.65 ;
      RECT 79.61 1.89 79.93 2.15 ;
      RECT 79.385 1.905 79.93 2.135 ;
      RECT 78.94 1.95 79.93 2.09 ;
      RECT 77.29 3.57 77.61 3.83 ;
      RECT 77.29 3.63 78.36 3.77 ;
      RECT 78.22 3.07 78.36 3.77 ;
      RECT 79.385 3.025 79.675 3.255 ;
      RECT 78.22 3.07 79.675 3.21 ;
      RECT 77.65 1.89 77.97 2.15 ;
      RECT 77.425 1.905 77.97 2.135 ;
      RECT 76.67 2.45 76.99 2.71 ;
      RECT 77.665 2.465 77.955 2.695 ;
      RECT 76.425 2.465 76.99 2.695 ;
      RECT 76.425 2.51 77.955 2.65 ;
      RECT 75.945 3.025 76.235 3.255 ;
      RECT 76.14 1.95 76.28 3.21 ;
      RECT 76.93 1.89 77.25 2.15 ;
      RECT 75.945 1.905 76.235 2.135 ;
      RECT 75.945 1.95 77.25 2.09 ;
      RECT 75.54 3.465 76.64 3.605 ;
      RECT 76.425 3.305 76.715 3.535 ;
      RECT 75.465 3.305 75.755 3.535 ;
      RECT 75.705 2.37 75.995 2.74 ;
      RECT 74.94 2.37 75.995 2.51 ;
      RECT 75.45 1.89 75.77 2.15 ;
      RECT 73.49 1.89 73.81 2.15 ;
      RECT 73.49 1.95 75.77 2.09 ;
      RECT 74.61 3.01 74.93 3.27 ;
      RECT 74.61 3.01 75.44 3.15 ;
      RECT 75.225 2.745 75.44 3.15 ;
      RECT 75.225 2.745 75.515 2.975 ;
      RECT 73.01 2.45 73.33 2.71 ;
      RECT 74.42 2.465 74.71 2.695 ;
      RECT 73.01 2.465 73.555 2.695 ;
      RECT 73.01 2.55 73.96 2.69 ;
      RECT 73.82 2.37 73.96 2.69 ;
      RECT 74.32 2.465 74.71 2.65 ;
      RECT 73.82 2.37 74.46 2.51 ;
      RECT 72.53 3.26 72.85 3.675 ;
      RECT 72.61 1.905 72.765 3.675 ;
      RECT 72.545 1.905 72.835 2.135 ;
      RECT 70.93 7.765 71.22 7.995 ;
      RECT 70.99 6.285 71.16 7.995 ;
      RECT 70.935 6.655 71.285 7.005 ;
      RECT 70.93 6.285 71.22 6.515 ;
      RECT 70.93 2.365 71.22 2.595 ;
      RECT 70.99 0.885 71.16 2.595 ;
      RECT 70.93 0.885 71.22 1.115 ;
      RECT 70.52 2.735 70.85 2.965 ;
      RECT 70.52 2.765 71.02 2.935 ;
      RECT 70.52 2.395 70.71 2.965 ;
      RECT 69.94 2.365 70.23 2.595 ;
      RECT 69.94 2.395 70.71 2.565 ;
      RECT 70 0.885 70.17 2.595 ;
      RECT 69.94 0.885 70.23 1.115 ;
      RECT 69.94 7.765 70.23 7.995 ;
      RECT 70 6.285 70.17 7.995 ;
      RECT 69.94 6.285 70.23 6.515 ;
      RECT 69.94 6.325 70.79 6.485 ;
      RECT 70.62 5.915 70.79 6.485 ;
      RECT 69.94 6.32 70.33 6.485 ;
      RECT 70.56 5.915 70.85 6.145 ;
      RECT 70.56 5.945 71.02 6.115 ;
      RECT 69.57 2.735 69.86 2.965 ;
      RECT 69.57 2.765 70.03 2.935 ;
      RECT 69.63 1.655 69.795 2.965 ;
      RECT 68.145 1.625 68.435 1.855 ;
      RECT 68.145 1.655 69.795 1.825 ;
      RECT 68.205 0.885 68.375 1.855 ;
      RECT 68.145 0.885 68.435 1.115 ;
      RECT 68.145 7.765 68.435 7.995 ;
      RECT 68.205 7.025 68.375 7.995 ;
      RECT 68.205 7.12 69.795 7.29 ;
      RECT 69.625 5.915 69.795 7.29 ;
      RECT 68.145 7.025 68.435 7.255 ;
      RECT 69.57 5.915 69.86 6.145 ;
      RECT 69.57 5.945 70.03 6.115 ;
      RECT 66.195 3.15 66.535 3.5 ;
      RECT 66.285 2.025 66.455 3.5 ;
      RECT 68.575 1.965 68.925 2.315 ;
      RECT 66.285 2.025 68.925 2.195 ;
      RECT 68.6 6.655 68.925 6.98 ;
      RECT 63.16 6.61 63.51 6.96 ;
      RECT 68.575 6.655 68.925 6.885 ;
      RECT 62.96 6.655 63.51 6.885 ;
      RECT 62.79 6.685 68.925 6.855 ;
      RECT 67.8 2.365 68.12 2.685 ;
      RECT 67.77 2.365 68.12 2.595 ;
      RECT 67.6 2.395 68.12 2.565 ;
      RECT 67.8 6.255 68.12 6.545 ;
      RECT 67.77 6.285 68.12 6.515 ;
      RECT 67.6 6.315 68.12 6.485 ;
      RECT 66.76 2.705 67.1 3.055 ;
      RECT 66.76 2.765 67.235 2.935 ;
      RECT 66.75 5.845 67.09 6.195 ;
      RECT 61.16 5.915 61.45 6.145 ;
      RECT 61.16 5.945 67.235 6.115 ;
      RECT 63.25 3.57 63.57 3.83 ;
      RECT 64.54 2.745 64.68 3.605 ;
      RECT 63.34 3.465 64.68 3.605 ;
      RECT 63.34 3.025 63.48 3.83 ;
      RECT 63.265 3.025 63.555 3.255 ;
      RECT 64.465 2.745 64.755 2.975 ;
      RECT 63.985 3.025 64.275 3.255 ;
      RECT 64.18 1.95 64.32 3.21 ;
      RECT 64.21 1.89 64.53 2.15 ;
      RECT 60.81 2.45 61.13 2.71 ;
      RECT 63.505 2.465 63.795 2.695 ;
      RECT 60.9 2.37 63.72 2.51 ;
      RECT 62.77 1.89 63.09 2.15 ;
      RECT 63.265 1.905 63.555 2.135 ;
      RECT 62.77 1.95 63.555 2.09 ;
      RECT 62.77 3.01 63.09 3.27 ;
      RECT 62.77 2.79 63 3.27 ;
      RECT 62.265 2.745 62.555 2.975 ;
      RECT 62.265 2.79 63 2.93 ;
      RECT 62.53 7.765 62.82 7.995 ;
      RECT 62.59 7.025 62.76 7.995 ;
      RECT 62.49 7.055 62.87 7.425 ;
      RECT 62.53 7.025 62.82 7.425 ;
      RECT 61.29 3.57 61.61 3.83 ;
      RECT 60.825 3.585 61.115 3.815 ;
      RECT 60.825 3.63 61.61 3.77 ;
      RECT 59.585 2.465 59.875 2.695 ;
      RECT 59.585 2.51 60.52 2.65 ;
      RECT 60.38 1.95 60.52 2.65 ;
      RECT 61.05 1.89 61.37 2.15 ;
      RECT 60.825 1.905 61.37 2.135 ;
      RECT 60.38 1.95 61.37 2.09 ;
      RECT 58.73 3.57 59.05 3.83 ;
      RECT 58.73 3.63 59.8 3.77 ;
      RECT 59.66 3.07 59.8 3.77 ;
      RECT 60.825 3.025 61.115 3.255 ;
      RECT 59.66 3.07 61.115 3.21 ;
      RECT 59.09 1.89 59.41 2.15 ;
      RECT 58.865 1.905 59.41 2.135 ;
      RECT 58.11 2.45 58.43 2.71 ;
      RECT 59.105 2.465 59.395 2.695 ;
      RECT 57.865 2.465 58.43 2.695 ;
      RECT 57.865 2.51 59.395 2.65 ;
      RECT 57.385 3.025 57.675 3.255 ;
      RECT 57.58 1.95 57.72 3.21 ;
      RECT 58.37 1.89 58.69 2.15 ;
      RECT 57.385 1.905 57.675 2.135 ;
      RECT 57.385 1.95 58.69 2.09 ;
      RECT 56.98 3.465 58.08 3.605 ;
      RECT 57.865 3.305 58.155 3.535 ;
      RECT 56.905 3.305 57.195 3.535 ;
      RECT 57.145 2.37 57.435 2.74 ;
      RECT 56.38 2.37 57.435 2.51 ;
      RECT 56.89 1.89 57.21 2.15 ;
      RECT 54.93 1.89 55.25 2.15 ;
      RECT 54.93 1.95 57.21 2.09 ;
      RECT 56.05 3.01 56.37 3.27 ;
      RECT 56.05 3.01 56.88 3.15 ;
      RECT 56.665 2.745 56.88 3.15 ;
      RECT 56.665 2.745 56.955 2.975 ;
      RECT 54.45 2.45 54.77 2.71 ;
      RECT 55.86 2.465 56.15 2.695 ;
      RECT 54.45 2.465 54.995 2.695 ;
      RECT 54.45 2.55 55.4 2.69 ;
      RECT 55.26 2.37 55.4 2.69 ;
      RECT 55.76 2.465 56.15 2.65 ;
      RECT 55.26 2.37 55.9 2.51 ;
      RECT 53.97 3.26 54.29 3.675 ;
      RECT 54.05 1.905 54.205 3.675 ;
      RECT 53.985 1.905 54.275 2.135 ;
      RECT 52.37 7.765 52.66 7.995 ;
      RECT 52.43 6.285 52.6 7.995 ;
      RECT 52.375 6.655 52.725 7.005 ;
      RECT 52.37 6.285 52.66 6.515 ;
      RECT 52.37 2.365 52.66 2.595 ;
      RECT 52.43 0.885 52.6 2.595 ;
      RECT 52.37 0.885 52.66 1.115 ;
      RECT 51.96 2.735 52.29 2.965 ;
      RECT 51.96 2.765 52.46 2.935 ;
      RECT 51.96 2.395 52.15 2.965 ;
      RECT 51.38 2.365 51.67 2.595 ;
      RECT 51.38 2.395 52.15 2.565 ;
      RECT 51.44 0.885 51.61 2.595 ;
      RECT 51.38 0.885 51.67 1.115 ;
      RECT 51.38 7.765 51.67 7.995 ;
      RECT 51.44 6.285 51.61 7.995 ;
      RECT 51.38 6.285 51.67 6.515 ;
      RECT 51.38 6.325 52.23 6.485 ;
      RECT 52.06 5.915 52.23 6.485 ;
      RECT 51.38 6.32 51.77 6.485 ;
      RECT 52 5.915 52.29 6.145 ;
      RECT 52 5.945 52.46 6.115 ;
      RECT 51.01 2.735 51.3 2.965 ;
      RECT 51.01 2.765 51.47 2.935 ;
      RECT 51.07 1.655 51.235 2.965 ;
      RECT 49.585 1.625 49.875 1.855 ;
      RECT 49.585 1.655 51.235 1.825 ;
      RECT 49.645 0.885 49.815 1.855 ;
      RECT 49.585 0.885 49.875 1.115 ;
      RECT 49.585 7.765 49.875 7.995 ;
      RECT 49.645 7.025 49.815 7.995 ;
      RECT 49.645 7.12 51.235 7.29 ;
      RECT 51.065 5.915 51.235 7.29 ;
      RECT 49.585 7.025 49.875 7.255 ;
      RECT 51.01 5.915 51.3 6.145 ;
      RECT 51.01 5.945 51.47 6.115 ;
      RECT 47.635 3.15 47.975 3.5 ;
      RECT 47.725 2.025 47.895 3.5 ;
      RECT 50.015 1.965 50.365 2.315 ;
      RECT 47.725 2.025 50.365 2.195 ;
      RECT 50.04 6.655 50.365 6.98 ;
      RECT 44.6 6.615 44.95 6.965 ;
      RECT 50.015 6.655 50.365 6.885 ;
      RECT 44.4 6.655 44.95 6.885 ;
      RECT 44.23 6.685 50.365 6.855 ;
      RECT 49.24 2.365 49.56 2.685 ;
      RECT 49.21 2.365 49.56 2.595 ;
      RECT 49.04 2.395 49.56 2.565 ;
      RECT 49.24 6.255 49.56 6.545 ;
      RECT 49.21 6.285 49.56 6.515 ;
      RECT 49.04 6.315 49.56 6.485 ;
      RECT 48.2 2.705 48.54 3.055 ;
      RECT 48.2 2.765 48.675 2.935 ;
      RECT 48.19 5.845 48.53 6.195 ;
      RECT 42.6 5.915 42.89 6.145 ;
      RECT 42.6 5.945 48.675 6.115 ;
      RECT 44.69 3.57 45.01 3.83 ;
      RECT 45.98 2.745 46.12 3.605 ;
      RECT 44.78 3.465 46.12 3.605 ;
      RECT 44.78 3.025 44.92 3.83 ;
      RECT 44.705 3.025 44.995 3.255 ;
      RECT 45.905 2.745 46.195 2.975 ;
      RECT 45.425 3.025 45.715 3.255 ;
      RECT 45.62 1.95 45.76 3.21 ;
      RECT 45.65 1.89 45.97 2.15 ;
      RECT 42.25 2.45 42.57 2.71 ;
      RECT 44.945 2.465 45.235 2.695 ;
      RECT 42.34 2.37 45.16 2.51 ;
      RECT 44.21 1.89 44.53 2.15 ;
      RECT 44.705 1.905 44.995 2.135 ;
      RECT 44.21 1.95 44.995 2.09 ;
      RECT 44.21 3.01 44.53 3.27 ;
      RECT 44.21 2.79 44.44 3.27 ;
      RECT 43.705 2.745 43.995 2.975 ;
      RECT 43.705 2.79 44.44 2.93 ;
      RECT 43.97 7.765 44.26 7.995 ;
      RECT 44.03 7.025 44.2 7.995 ;
      RECT 43.93 7.055 44.31 7.425 ;
      RECT 43.97 7.025 44.26 7.425 ;
      RECT 42.73 3.57 43.05 3.83 ;
      RECT 42.265 3.585 42.555 3.815 ;
      RECT 42.265 3.63 43.05 3.77 ;
      RECT 41.025 2.465 41.315 2.695 ;
      RECT 41.025 2.51 41.96 2.65 ;
      RECT 41.82 1.95 41.96 2.65 ;
      RECT 42.49 1.89 42.81 2.15 ;
      RECT 42.265 1.905 42.81 2.135 ;
      RECT 41.82 1.95 42.81 2.09 ;
      RECT 40.17 3.57 40.49 3.83 ;
      RECT 40.17 3.63 41.24 3.77 ;
      RECT 41.1 3.07 41.24 3.77 ;
      RECT 42.265 3.025 42.555 3.255 ;
      RECT 41.1 3.07 42.555 3.21 ;
      RECT 40.53 1.89 40.85 2.15 ;
      RECT 40.305 1.905 40.85 2.135 ;
      RECT 39.55 2.45 39.87 2.71 ;
      RECT 40.545 2.465 40.835 2.695 ;
      RECT 39.305 2.465 39.87 2.695 ;
      RECT 39.305 2.51 40.835 2.65 ;
      RECT 38.825 3.025 39.115 3.255 ;
      RECT 39.02 1.95 39.16 3.21 ;
      RECT 39.81 1.89 40.13 2.15 ;
      RECT 38.825 1.905 39.115 2.135 ;
      RECT 38.825 1.95 40.13 2.09 ;
      RECT 38.42 3.465 39.52 3.605 ;
      RECT 39.305 3.305 39.595 3.535 ;
      RECT 38.345 3.305 38.635 3.535 ;
      RECT 38.585 2.37 38.875 2.74 ;
      RECT 37.82 2.37 38.875 2.51 ;
      RECT 38.33 1.89 38.65 2.15 ;
      RECT 36.37 1.89 36.69 2.15 ;
      RECT 36.37 1.95 38.65 2.09 ;
      RECT 37.49 3.01 37.81 3.27 ;
      RECT 37.49 3.01 38.32 3.15 ;
      RECT 38.105 2.745 38.32 3.15 ;
      RECT 38.105 2.745 38.395 2.975 ;
      RECT 35.89 2.45 36.21 2.71 ;
      RECT 37.3 2.465 37.59 2.695 ;
      RECT 35.89 2.465 36.435 2.695 ;
      RECT 35.89 2.55 36.84 2.69 ;
      RECT 36.7 2.37 36.84 2.69 ;
      RECT 37.2 2.465 37.59 2.65 ;
      RECT 36.7 2.37 37.34 2.51 ;
      RECT 35.41 3.26 35.73 3.675 ;
      RECT 35.49 1.905 35.645 3.675 ;
      RECT 35.425 1.905 35.715 2.135 ;
      RECT 33.81 7.765 34.1 7.995 ;
      RECT 33.87 6.285 34.04 7.995 ;
      RECT 33.855 6.66 34.21 7.015 ;
      RECT 33.81 6.285 34.1 6.515 ;
      RECT 33.81 2.365 34.1 2.595 ;
      RECT 33.87 0.885 34.04 2.595 ;
      RECT 33.81 0.885 34.1 1.115 ;
      RECT 33.4 2.735 33.73 2.965 ;
      RECT 33.4 2.765 33.9 2.935 ;
      RECT 33.4 2.395 33.59 2.965 ;
      RECT 32.82 2.365 33.11 2.595 ;
      RECT 32.82 2.395 33.59 2.565 ;
      RECT 32.88 0.885 33.05 2.595 ;
      RECT 32.82 0.885 33.11 1.115 ;
      RECT 32.82 7.765 33.11 7.995 ;
      RECT 32.88 6.285 33.05 7.995 ;
      RECT 32.82 6.285 33.11 6.515 ;
      RECT 32.82 6.325 33.67 6.485 ;
      RECT 33.5 5.915 33.67 6.485 ;
      RECT 32.82 6.32 33.21 6.485 ;
      RECT 33.44 5.915 33.73 6.145 ;
      RECT 33.44 5.945 33.9 6.115 ;
      RECT 32.45 2.735 32.74 2.965 ;
      RECT 32.45 2.765 32.91 2.935 ;
      RECT 32.51 1.655 32.675 2.965 ;
      RECT 31.025 1.625 31.315 1.855 ;
      RECT 31.025 1.655 32.675 1.825 ;
      RECT 31.085 0.885 31.255 1.855 ;
      RECT 31.025 0.885 31.315 1.115 ;
      RECT 31.025 7.765 31.315 7.995 ;
      RECT 31.085 7.025 31.255 7.995 ;
      RECT 31.085 7.12 32.675 7.29 ;
      RECT 32.505 5.915 32.675 7.29 ;
      RECT 31.025 7.025 31.315 7.255 ;
      RECT 32.45 5.915 32.74 6.145 ;
      RECT 32.45 5.945 32.91 6.115 ;
      RECT 29.075 3.15 29.415 3.5 ;
      RECT 29.165 2.025 29.335 3.5 ;
      RECT 31.455 1.965 31.805 2.315 ;
      RECT 29.165 2.025 31.805 2.195 ;
      RECT 31.48 6.655 31.805 6.98 ;
      RECT 26.045 6.61 26.395 6.96 ;
      RECT 31.455 6.655 31.805 6.885 ;
      RECT 25.84 6.655 26.395 6.885 ;
      RECT 25.67 6.685 31.805 6.855 ;
      RECT 30.68 2.365 31 2.685 ;
      RECT 30.65 2.365 31 2.595 ;
      RECT 30.48 2.395 31 2.565 ;
      RECT 30.68 6.255 31 6.545 ;
      RECT 30.65 6.285 31 6.515 ;
      RECT 30.48 6.315 31 6.485 ;
      RECT 29.64 2.705 29.98 3.055 ;
      RECT 29.64 2.765 30.115 2.935 ;
      RECT 29.63 5.845 29.97 6.195 ;
      RECT 24.04 5.915 24.33 6.145 ;
      RECT 24.04 5.945 30.115 6.115 ;
      RECT 26.13 3.57 26.45 3.83 ;
      RECT 27.42 2.745 27.56 3.605 ;
      RECT 26.22 3.465 27.56 3.605 ;
      RECT 26.22 3.025 26.36 3.83 ;
      RECT 26.145 3.025 26.435 3.255 ;
      RECT 27.345 2.745 27.635 2.975 ;
      RECT 26.865 3.025 27.155 3.255 ;
      RECT 27.06 1.95 27.2 3.21 ;
      RECT 27.09 1.89 27.41 2.15 ;
      RECT 23.69 2.45 24.01 2.71 ;
      RECT 26.385 2.465 26.675 2.695 ;
      RECT 23.78 2.37 26.6 2.51 ;
      RECT 25.65 1.89 25.97 2.15 ;
      RECT 26.145 1.905 26.435 2.135 ;
      RECT 25.65 1.95 26.435 2.09 ;
      RECT 25.65 3.01 25.97 3.27 ;
      RECT 25.65 2.79 25.88 3.27 ;
      RECT 25.145 2.745 25.435 2.975 ;
      RECT 25.145 2.79 25.88 2.93 ;
      RECT 25.41 7.765 25.7 7.995 ;
      RECT 25.47 7.025 25.64 7.995 ;
      RECT 25.37 7.055 25.75 7.425 ;
      RECT 25.41 7.025 25.7 7.425 ;
      RECT 24.17 3.57 24.49 3.83 ;
      RECT 23.705 3.585 23.995 3.815 ;
      RECT 23.705 3.63 24.49 3.77 ;
      RECT 22.465 2.465 22.755 2.695 ;
      RECT 22.465 2.51 23.4 2.65 ;
      RECT 23.26 1.95 23.4 2.65 ;
      RECT 23.93 1.89 24.25 2.15 ;
      RECT 23.705 1.905 24.25 2.135 ;
      RECT 23.26 1.95 24.25 2.09 ;
      RECT 21.61 3.57 21.93 3.83 ;
      RECT 21.61 3.63 22.68 3.77 ;
      RECT 22.54 3.07 22.68 3.77 ;
      RECT 23.705 3.025 23.995 3.255 ;
      RECT 22.54 3.07 23.995 3.21 ;
      RECT 21.97 1.89 22.29 2.15 ;
      RECT 21.745 1.905 22.29 2.135 ;
      RECT 20.99 2.45 21.31 2.71 ;
      RECT 21.985 2.465 22.275 2.695 ;
      RECT 20.745 2.465 21.31 2.695 ;
      RECT 20.745 2.51 22.275 2.65 ;
      RECT 20.265 3.025 20.555 3.255 ;
      RECT 20.46 1.95 20.6 3.21 ;
      RECT 21.25 1.89 21.57 2.15 ;
      RECT 20.265 1.905 20.555 2.135 ;
      RECT 20.265 1.95 21.57 2.09 ;
      RECT 19.86 3.465 20.96 3.605 ;
      RECT 20.745 3.305 21.035 3.535 ;
      RECT 19.785 3.305 20.075 3.535 ;
      RECT 20.025 2.37 20.315 2.74 ;
      RECT 19.26 2.37 20.315 2.51 ;
      RECT 19.77 1.89 20.09 2.15 ;
      RECT 17.81 1.89 18.13 2.15 ;
      RECT 17.81 1.95 20.09 2.09 ;
      RECT 18.93 3.01 19.25 3.27 ;
      RECT 18.93 3.01 19.76 3.15 ;
      RECT 19.545 2.745 19.76 3.15 ;
      RECT 19.545 2.745 19.835 2.975 ;
      RECT 17.33 2.45 17.65 2.71 ;
      RECT 18.74 2.465 19.03 2.695 ;
      RECT 17.33 2.465 17.875 2.695 ;
      RECT 17.33 2.55 18.28 2.69 ;
      RECT 18.14 2.37 18.28 2.69 ;
      RECT 18.64 2.465 19.03 2.65 ;
      RECT 18.14 2.37 18.78 2.51 ;
      RECT 16.85 3.26 17.17 3.675 ;
      RECT 16.93 1.905 17.085 3.675 ;
      RECT 16.865 1.905 17.155 2.135 ;
      RECT 15.25 7.765 15.54 7.995 ;
      RECT 15.31 6.285 15.48 7.995 ;
      RECT 15.3 6.655 15.65 7.005 ;
      RECT 15.25 6.285 15.54 6.515 ;
      RECT 15.25 2.365 15.54 2.595 ;
      RECT 15.31 0.885 15.48 2.595 ;
      RECT 15.25 0.885 15.54 1.115 ;
      RECT 14.84 2.735 15.17 2.965 ;
      RECT 14.84 2.765 15.34 2.935 ;
      RECT 14.84 2.395 15.03 2.965 ;
      RECT 14.26 2.365 14.55 2.595 ;
      RECT 14.26 2.395 15.03 2.565 ;
      RECT 14.32 0.885 14.49 2.595 ;
      RECT 14.26 0.885 14.55 1.115 ;
      RECT 14.26 7.765 14.55 7.995 ;
      RECT 14.32 6.285 14.49 7.995 ;
      RECT 14.26 6.285 14.55 6.515 ;
      RECT 14.26 6.325 15.11 6.485 ;
      RECT 14.94 5.915 15.11 6.485 ;
      RECT 14.26 6.32 14.65 6.485 ;
      RECT 14.88 5.915 15.17 6.145 ;
      RECT 14.88 5.945 15.34 6.115 ;
      RECT 13.89 2.735 14.18 2.965 ;
      RECT 13.89 2.765 14.35 2.935 ;
      RECT 13.95 1.655 14.115 2.965 ;
      RECT 12.465 1.625 12.755 1.855 ;
      RECT 12.465 1.655 14.115 1.825 ;
      RECT 12.525 0.885 12.695 1.855 ;
      RECT 12.465 0.885 12.755 1.115 ;
      RECT 12.465 7.765 12.755 7.995 ;
      RECT 12.525 7.025 12.695 7.995 ;
      RECT 12.525 7.12 14.115 7.29 ;
      RECT 13.945 5.915 14.115 7.29 ;
      RECT 12.465 7.025 12.755 7.255 ;
      RECT 13.89 5.915 14.18 6.145 ;
      RECT 13.89 5.945 14.35 6.115 ;
      RECT 10.515 3.15 10.855 3.5 ;
      RECT 10.605 2.025 10.775 3.5 ;
      RECT 12.895 1.965 13.245 2.315 ;
      RECT 10.605 2.025 13.245 2.195 ;
      RECT 12.92 6.655 13.245 6.98 ;
      RECT 7.485 6.605 7.835 6.955 ;
      RECT 12.895 6.655 13.245 6.885 ;
      RECT 7.28 6.655 7.835 6.885 ;
      RECT 7.11 6.685 13.245 6.855 ;
      RECT 12.12 2.365 12.44 2.685 ;
      RECT 12.09 2.365 12.44 2.595 ;
      RECT 11.92 2.395 12.44 2.565 ;
      RECT 12.12 6.255 12.44 6.545 ;
      RECT 12.09 6.285 12.44 6.515 ;
      RECT 11.92 6.315 12.44 6.485 ;
      RECT 11.08 2.705 11.42 3.055 ;
      RECT 11.08 2.765 11.555 2.935 ;
      RECT 11.07 5.845 11.41 6.195 ;
      RECT 5.48 5.915 5.77 6.145 ;
      RECT 5.48 5.945 11.555 6.115 ;
      RECT 7.57 3.57 7.89 3.83 ;
      RECT 8.86 2.745 9 3.605 ;
      RECT 7.66 3.465 9 3.605 ;
      RECT 7.66 3.025 7.8 3.83 ;
      RECT 7.585 3.025 7.875 3.255 ;
      RECT 8.785 2.745 9.075 2.975 ;
      RECT 8.305 3.025 8.595 3.255 ;
      RECT 8.5 1.95 8.64 3.21 ;
      RECT 8.53 1.89 8.85 2.15 ;
      RECT 5.13 2.45 5.45 2.71 ;
      RECT 7.825 2.465 8.115 2.695 ;
      RECT 5.22 2.37 8.04 2.51 ;
      RECT 7.09 1.89 7.41 2.15 ;
      RECT 7.585 1.905 7.875 2.135 ;
      RECT 7.09 1.95 7.875 2.09 ;
      RECT 7.09 3.01 7.41 3.27 ;
      RECT 7.09 2.79 7.32 3.27 ;
      RECT 6.585 2.745 6.875 2.975 ;
      RECT 6.585 2.79 7.32 2.93 ;
      RECT 6.85 7.765 7.14 7.995 ;
      RECT 6.91 7.025 7.08 7.995 ;
      RECT 6.81 7.055 7.19 7.425 ;
      RECT 6.85 7.025 7.14 7.425 ;
      RECT 5.61 3.57 5.93 3.83 ;
      RECT 5.145 3.585 5.435 3.815 ;
      RECT 5.145 3.63 5.93 3.77 ;
      RECT 3.905 2.465 4.195 2.695 ;
      RECT 3.905 2.51 4.84 2.65 ;
      RECT 4.7 1.95 4.84 2.65 ;
      RECT 5.37 1.89 5.69 2.15 ;
      RECT 5.145 1.905 5.69 2.135 ;
      RECT 4.7 1.95 5.69 2.09 ;
      RECT 3.05 3.57 3.37 3.83 ;
      RECT 3.05 3.63 4.12 3.77 ;
      RECT 3.98 3.07 4.12 3.77 ;
      RECT 5.145 3.025 5.435 3.255 ;
      RECT 3.98 3.07 5.435 3.21 ;
      RECT 3.41 1.89 3.73 2.15 ;
      RECT 3.185 1.905 3.73 2.135 ;
      RECT 2.43 2.45 2.75 2.71 ;
      RECT 3.425 2.465 3.715 2.695 ;
      RECT 2.185 2.465 2.75 2.695 ;
      RECT 2.185 2.51 3.715 2.65 ;
      RECT 1.705 3.025 1.995 3.255 ;
      RECT 1.9 1.95 2.04 3.21 ;
      RECT 2.69 1.89 3.01 2.15 ;
      RECT 1.705 1.905 1.995 2.135 ;
      RECT 1.705 1.95 3.01 2.09 ;
      RECT 1.3 3.465 2.4 3.605 ;
      RECT 2.185 3.305 2.475 3.535 ;
      RECT 1.225 3.305 1.515 3.535 ;
      RECT 1.465 2.37 1.755 2.74 ;
      RECT 0.7 2.37 1.755 2.51 ;
      RECT 1.21 1.89 1.53 2.15 ;
      RECT -0.75 1.89 -0.43 2.15 ;
      RECT -0.75 1.95 1.53 2.09 ;
      RECT 0.37 3.01 0.69 3.27 ;
      RECT 0.37 3.01 1.2 3.15 ;
      RECT 0.985 2.745 1.2 3.15 ;
      RECT 0.985 2.745 1.275 2.975 ;
      RECT -1.23 2.45 -0.91 2.71 ;
      RECT 0.18 2.465 0.47 2.695 ;
      RECT -1.23 2.465 -0.685 2.695 ;
      RECT -1.23 2.55 -0.28 2.69 ;
      RECT -0.42 2.37 -0.28 2.69 ;
      RECT 0.08 2.465 0.47 2.65 ;
      RECT -0.42 2.37 0.22 2.51 ;
      RECT -1.71 3.26 -1.39 3.675 ;
      RECT -1.63 1.905 -1.475 3.675 ;
      RECT -1.695 1.905 -1.405 2.135 ;
      RECT -3.535 6.655 -3.245 6.885 ;
      RECT -3.705 6.685 -3.245 6.855 ;
      RECT -3.965 7.765 -3.675 7.995 ;
      RECT -3.905 7.025 -3.735 7.995 ;
      RECT -3.995 7.025 -3.645 7.315 ;
      RECT -4.37 6.285 -4.02 6.575 ;
      RECT -4.51 6.315 -4.02 6.485 ;
      RECT -5.365 5.905 -5.025 6.165 ;
      RECT -5.365 5.945 -4.875 6.115 ;
      RECT 80.81 3.57 81.13 3.83 ;
      RECT 80.21 1.89 80.89 2.15 ;
      RECT 80.33 3.57 80.65 3.83 ;
      RECT 78.85 3.57 79.17 3.83 ;
      RECT 78.37 1.89 78.69 2.15 ;
      RECT 77.65 3.01 77.97 3.27 ;
      RECT 76.93 3.01 77.25 3.27 ;
      RECT 73.97 3.01 74.29 3.27 ;
      RECT 73.49 3.01 73.81 3.27 ;
      RECT 62.25 3.57 62.57 3.83 ;
      RECT 61.65 1.89 62.33 2.15 ;
      RECT 61.77 3.57 62.09 3.83 ;
      RECT 60.29 3.57 60.61 3.83 ;
      RECT 59.81 1.89 60.13 2.15 ;
      RECT 59.09 3.01 59.41 3.27 ;
      RECT 58.37 3.01 58.69 3.27 ;
      RECT 55.41 3.01 55.73 3.27 ;
      RECT 54.93 3.01 55.25 3.27 ;
      RECT 43.69 3.57 44.01 3.83 ;
      RECT 43.09 1.89 43.77 2.15 ;
      RECT 43.21 3.57 43.53 3.83 ;
      RECT 41.73 3.57 42.05 3.83 ;
      RECT 41.25 1.89 41.57 2.15 ;
      RECT 40.53 3.01 40.85 3.27 ;
      RECT 39.81 3.01 40.13 3.27 ;
      RECT 36.85 3.01 37.17 3.27 ;
      RECT 36.37 3.01 36.69 3.27 ;
      RECT 25.13 3.57 25.45 3.83 ;
      RECT 24.53 1.89 25.21 2.15 ;
      RECT 24.65 3.57 24.97 3.83 ;
      RECT 23.17 3.57 23.49 3.83 ;
      RECT 22.69 1.89 23.01 2.15 ;
      RECT 21.97 3.01 22.29 3.27 ;
      RECT 21.25 3.01 21.57 3.27 ;
      RECT 18.29 3.01 18.61 3.27 ;
      RECT 17.81 3.01 18.13 3.27 ;
      RECT 6.57 3.57 6.89 3.83 ;
      RECT 5.97 1.89 6.65 2.15 ;
      RECT 6.09 3.57 6.41 3.83 ;
      RECT 4.61 3.57 4.93 3.83 ;
      RECT 4.13 1.89 4.45 2.15 ;
      RECT 3.41 3.01 3.73 3.27 ;
      RECT 2.69 3.01 3.01 3.27 ;
      RECT -0.27 3.01 0.05 3.27 ;
      RECT -0.75 3.01 -0.43 3.27 ;
    LAYER mcon ;
      RECT 89.55 0.915 89.72 1.085 ;
      RECT 89.55 2.395 89.72 2.565 ;
      RECT 89.55 6.315 89.72 6.485 ;
      RECT 89.55 7.795 89.72 7.965 ;
      RECT 89.2 0.105 89.37 0.275 ;
      RECT 89.2 4.165 89.37 4.335 ;
      RECT 89.2 4.545 89.37 4.715 ;
      RECT 89.2 8.605 89.37 8.775 ;
      RECT 89.18 2.765 89.35 2.935 ;
      RECT 89.18 5.945 89.35 6.115 ;
      RECT 88.56 0.915 88.73 1.085 ;
      RECT 88.56 2.395 88.73 2.565 ;
      RECT 88.56 6.315 88.73 6.485 ;
      RECT 88.56 7.795 88.73 7.965 ;
      RECT 88.21 0.105 88.38 0.275 ;
      RECT 88.21 4.165 88.38 4.335 ;
      RECT 88.21 4.545 88.38 4.715 ;
      RECT 88.21 8.605 88.38 8.775 ;
      RECT 88.19 2.765 88.36 2.935 ;
      RECT 88.19 5.945 88.36 6.115 ;
      RECT 87.505 0.105 87.675 0.275 ;
      RECT 87.505 4.165 87.675 4.335 ;
      RECT 87.505 4.545 87.675 4.715 ;
      RECT 87.505 8.605 87.675 8.775 ;
      RECT 87.195 2.025 87.365 2.195 ;
      RECT 87.195 6.685 87.365 6.855 ;
      RECT 86.825 0.105 86.995 0.275 ;
      RECT 86.825 8.605 86.995 8.775 ;
      RECT 86.765 0.915 86.935 1.085 ;
      RECT 86.765 1.655 86.935 1.825 ;
      RECT 86.765 7.055 86.935 7.225 ;
      RECT 86.765 7.795 86.935 7.965 ;
      RECT 86.39 2.395 86.56 2.565 ;
      RECT 86.39 6.315 86.56 6.485 ;
      RECT 86.145 0.105 86.315 0.275 ;
      RECT 86.145 8.605 86.315 8.775 ;
      RECT 85.465 0.105 85.635 0.275 ;
      RECT 85.465 8.605 85.635 8.775 ;
      RECT 85.395 2.765 85.565 2.935 ;
      RECT 85.395 5.945 85.565 6.115 ;
      RECT 83.92 1.415 84.09 1.585 ;
      RECT 83.92 4.135 84.09 4.305 ;
      RECT 83.46 1.415 83.63 1.585 ;
      RECT 83.46 4.135 83.63 4.305 ;
      RECT 83.085 2.775 83.255 2.945 ;
      RECT 83 1.415 83.17 1.585 ;
      RECT 83 4.135 83.17 4.305 ;
      RECT 82.845 1.935 83.015 2.105 ;
      RECT 82.605 3.055 82.775 3.225 ;
      RECT 82.54 1.415 82.71 1.585 ;
      RECT 82.54 4.135 82.71 4.305 ;
      RECT 82.125 2.495 82.295 2.665 ;
      RECT 82.08 1.415 82.25 1.585 ;
      RECT 82.08 4.135 82.25 4.305 ;
      RECT 81.89 4.545 82.06 4.715 ;
      RECT 81.89 8.605 82.06 8.775 ;
      RECT 81.885 1.935 82.055 2.105 ;
      RECT 81.885 3.055 82.055 3.225 ;
      RECT 81.885 3.615 82.055 3.785 ;
      RECT 81.62 1.415 81.79 1.585 ;
      RECT 81.62 4.135 81.79 4.305 ;
      RECT 81.58 6.685 81.75 6.855 ;
      RECT 81.405 3.055 81.575 3.225 ;
      RECT 81.21 8.605 81.38 8.775 ;
      RECT 81.16 1.415 81.33 1.585 ;
      RECT 81.16 4.135 81.33 4.305 ;
      RECT 81.15 7.055 81.32 7.225 ;
      RECT 81.15 7.795 81.32 7.965 ;
      RECT 80.885 2.775 81.055 2.945 ;
      RECT 80.885 3.615 81.055 3.785 ;
      RECT 80.775 6.315 80.945 6.485 ;
      RECT 80.7 1.415 80.87 1.585 ;
      RECT 80.7 4.135 80.87 4.305 ;
      RECT 80.53 8.605 80.7 8.775 ;
      RECT 80.405 1.935 80.575 2.105 ;
      RECT 80.405 3.615 80.575 3.785 ;
      RECT 80.24 1.415 80.41 1.585 ;
      RECT 80.24 4.135 80.41 4.305 ;
      RECT 79.85 8.605 80.02 8.775 ;
      RECT 79.78 1.415 79.95 1.585 ;
      RECT 79.78 4.135 79.95 4.305 ;
      RECT 79.78 5.945 79.95 6.115 ;
      RECT 79.445 1.935 79.615 2.105 ;
      RECT 79.445 2.495 79.615 2.665 ;
      RECT 79.445 3.055 79.615 3.225 ;
      RECT 79.445 3.615 79.615 3.785 ;
      RECT 79.32 1.415 79.49 1.585 ;
      RECT 79.32 4.135 79.49 4.305 ;
      RECT 78.925 3.615 79.095 3.785 ;
      RECT 78.86 1.415 79.03 1.585 ;
      RECT 78.86 4.135 79.03 4.305 ;
      RECT 78.445 1.935 78.615 2.105 ;
      RECT 78.4 1.415 78.57 1.585 ;
      RECT 78.4 4.135 78.57 4.305 ;
      RECT 78.205 2.495 78.375 2.665 ;
      RECT 77.94 1.415 78.11 1.585 ;
      RECT 77.94 4.135 78.11 4.305 ;
      RECT 77.725 2.495 77.895 2.665 ;
      RECT 77.725 3.055 77.895 3.225 ;
      RECT 77.485 1.935 77.655 2.105 ;
      RECT 77.48 1.415 77.65 1.585 ;
      RECT 77.48 4.135 77.65 4.305 ;
      RECT 77.02 1.415 77.19 1.585 ;
      RECT 77.02 4.135 77.19 4.305 ;
      RECT 77.005 3.055 77.175 3.225 ;
      RECT 76.56 1.415 76.73 1.585 ;
      RECT 76.56 4.135 76.73 4.305 ;
      RECT 76.485 2.495 76.655 2.665 ;
      RECT 76.485 3.335 76.655 3.505 ;
      RECT 76.1 1.415 76.27 1.585 ;
      RECT 76.1 4.135 76.27 4.305 ;
      RECT 76.005 1.935 76.175 2.105 ;
      RECT 76.005 3.055 76.175 3.225 ;
      RECT 75.765 2.495 75.935 2.665 ;
      RECT 75.64 1.415 75.81 1.585 ;
      RECT 75.64 4.135 75.81 4.305 ;
      RECT 75.525 3.335 75.695 3.505 ;
      RECT 75.285 2.775 75.455 2.945 ;
      RECT 75.18 1.415 75.35 1.585 ;
      RECT 75.18 4.135 75.35 4.305 ;
      RECT 74.72 1.415 74.89 1.585 ;
      RECT 74.72 4.135 74.89 4.305 ;
      RECT 74.48 2.495 74.65 2.665 ;
      RECT 74.26 1.415 74.43 1.585 ;
      RECT 74.26 4.135 74.43 4.305 ;
      RECT 74.045 3.055 74.215 3.225 ;
      RECT 73.8 1.415 73.97 1.585 ;
      RECT 73.8 4.135 73.97 4.305 ;
      RECT 73.565 1.935 73.735 2.105 ;
      RECT 73.565 3.055 73.735 3.225 ;
      RECT 73.34 1.415 73.51 1.585 ;
      RECT 73.34 4.135 73.51 4.305 ;
      RECT 73.325 2.495 73.495 2.665 ;
      RECT 72.88 1.415 73.05 1.585 ;
      RECT 72.88 4.135 73.05 4.305 ;
      RECT 72.605 1.935 72.775 2.105 ;
      RECT 72.605 3.475 72.775 3.645 ;
      RECT 72.42 1.415 72.59 1.585 ;
      RECT 72.42 4.135 72.59 4.305 ;
      RECT 70.99 0.915 71.16 1.085 ;
      RECT 70.99 2.395 71.16 2.565 ;
      RECT 70.99 6.315 71.16 6.485 ;
      RECT 70.99 7.795 71.16 7.965 ;
      RECT 70.64 0.105 70.81 0.275 ;
      RECT 70.64 4.165 70.81 4.335 ;
      RECT 70.64 4.545 70.81 4.715 ;
      RECT 70.64 8.605 70.81 8.775 ;
      RECT 70.62 2.765 70.79 2.935 ;
      RECT 70.62 5.945 70.79 6.115 ;
      RECT 70 0.915 70.17 1.085 ;
      RECT 70 2.395 70.17 2.565 ;
      RECT 70 6.315 70.17 6.485 ;
      RECT 70 7.795 70.17 7.965 ;
      RECT 69.65 0.105 69.82 0.275 ;
      RECT 69.65 4.165 69.82 4.335 ;
      RECT 69.65 4.545 69.82 4.715 ;
      RECT 69.65 8.605 69.82 8.775 ;
      RECT 69.63 2.765 69.8 2.935 ;
      RECT 69.63 5.945 69.8 6.115 ;
      RECT 68.945 0.105 69.115 0.275 ;
      RECT 68.945 4.165 69.115 4.335 ;
      RECT 68.945 4.545 69.115 4.715 ;
      RECT 68.945 8.605 69.115 8.775 ;
      RECT 68.635 2.025 68.805 2.195 ;
      RECT 68.635 6.685 68.805 6.855 ;
      RECT 68.265 0.105 68.435 0.275 ;
      RECT 68.265 8.605 68.435 8.775 ;
      RECT 68.205 0.915 68.375 1.085 ;
      RECT 68.205 1.655 68.375 1.825 ;
      RECT 68.205 7.055 68.375 7.225 ;
      RECT 68.205 7.795 68.375 7.965 ;
      RECT 67.83 2.395 68 2.565 ;
      RECT 67.83 6.315 68 6.485 ;
      RECT 67.585 0.105 67.755 0.275 ;
      RECT 67.585 8.605 67.755 8.775 ;
      RECT 66.905 0.105 67.075 0.275 ;
      RECT 66.905 8.605 67.075 8.775 ;
      RECT 66.835 2.765 67.005 2.935 ;
      RECT 66.835 5.945 67.005 6.115 ;
      RECT 65.36 1.415 65.53 1.585 ;
      RECT 65.36 4.135 65.53 4.305 ;
      RECT 64.9 1.415 65.07 1.585 ;
      RECT 64.9 4.135 65.07 4.305 ;
      RECT 64.525 2.775 64.695 2.945 ;
      RECT 64.44 1.415 64.61 1.585 ;
      RECT 64.44 4.135 64.61 4.305 ;
      RECT 64.285 1.935 64.455 2.105 ;
      RECT 64.045 3.055 64.215 3.225 ;
      RECT 63.98 1.415 64.15 1.585 ;
      RECT 63.98 4.135 64.15 4.305 ;
      RECT 63.565 2.495 63.735 2.665 ;
      RECT 63.52 1.415 63.69 1.585 ;
      RECT 63.52 4.135 63.69 4.305 ;
      RECT 63.33 4.545 63.5 4.715 ;
      RECT 63.33 8.605 63.5 8.775 ;
      RECT 63.325 1.935 63.495 2.105 ;
      RECT 63.325 3.055 63.495 3.225 ;
      RECT 63.325 3.615 63.495 3.785 ;
      RECT 63.06 1.415 63.23 1.585 ;
      RECT 63.06 4.135 63.23 4.305 ;
      RECT 63.02 6.685 63.19 6.855 ;
      RECT 62.845 3.055 63.015 3.225 ;
      RECT 62.65 8.605 62.82 8.775 ;
      RECT 62.6 1.415 62.77 1.585 ;
      RECT 62.6 4.135 62.77 4.305 ;
      RECT 62.59 7.055 62.76 7.225 ;
      RECT 62.59 7.795 62.76 7.965 ;
      RECT 62.325 2.775 62.495 2.945 ;
      RECT 62.325 3.615 62.495 3.785 ;
      RECT 62.215 6.315 62.385 6.485 ;
      RECT 62.14 1.415 62.31 1.585 ;
      RECT 62.14 4.135 62.31 4.305 ;
      RECT 61.97 8.605 62.14 8.775 ;
      RECT 61.845 1.935 62.015 2.105 ;
      RECT 61.845 3.615 62.015 3.785 ;
      RECT 61.68 1.415 61.85 1.585 ;
      RECT 61.68 4.135 61.85 4.305 ;
      RECT 61.29 8.605 61.46 8.775 ;
      RECT 61.22 1.415 61.39 1.585 ;
      RECT 61.22 4.135 61.39 4.305 ;
      RECT 61.22 5.945 61.39 6.115 ;
      RECT 60.885 1.935 61.055 2.105 ;
      RECT 60.885 2.495 61.055 2.665 ;
      RECT 60.885 3.055 61.055 3.225 ;
      RECT 60.885 3.615 61.055 3.785 ;
      RECT 60.76 1.415 60.93 1.585 ;
      RECT 60.76 4.135 60.93 4.305 ;
      RECT 60.365 3.615 60.535 3.785 ;
      RECT 60.3 1.415 60.47 1.585 ;
      RECT 60.3 4.135 60.47 4.305 ;
      RECT 59.885 1.935 60.055 2.105 ;
      RECT 59.84 1.415 60.01 1.585 ;
      RECT 59.84 4.135 60.01 4.305 ;
      RECT 59.645 2.495 59.815 2.665 ;
      RECT 59.38 1.415 59.55 1.585 ;
      RECT 59.38 4.135 59.55 4.305 ;
      RECT 59.165 2.495 59.335 2.665 ;
      RECT 59.165 3.055 59.335 3.225 ;
      RECT 58.925 1.935 59.095 2.105 ;
      RECT 58.92 1.415 59.09 1.585 ;
      RECT 58.92 4.135 59.09 4.305 ;
      RECT 58.46 1.415 58.63 1.585 ;
      RECT 58.46 4.135 58.63 4.305 ;
      RECT 58.445 3.055 58.615 3.225 ;
      RECT 58 1.415 58.17 1.585 ;
      RECT 58 4.135 58.17 4.305 ;
      RECT 57.925 2.495 58.095 2.665 ;
      RECT 57.925 3.335 58.095 3.505 ;
      RECT 57.54 1.415 57.71 1.585 ;
      RECT 57.54 4.135 57.71 4.305 ;
      RECT 57.445 1.935 57.615 2.105 ;
      RECT 57.445 3.055 57.615 3.225 ;
      RECT 57.205 2.495 57.375 2.665 ;
      RECT 57.08 1.415 57.25 1.585 ;
      RECT 57.08 4.135 57.25 4.305 ;
      RECT 56.965 3.335 57.135 3.505 ;
      RECT 56.725 2.775 56.895 2.945 ;
      RECT 56.62 1.415 56.79 1.585 ;
      RECT 56.62 4.135 56.79 4.305 ;
      RECT 56.16 1.415 56.33 1.585 ;
      RECT 56.16 4.135 56.33 4.305 ;
      RECT 55.92 2.495 56.09 2.665 ;
      RECT 55.7 1.415 55.87 1.585 ;
      RECT 55.7 4.135 55.87 4.305 ;
      RECT 55.485 3.055 55.655 3.225 ;
      RECT 55.24 1.415 55.41 1.585 ;
      RECT 55.24 4.135 55.41 4.305 ;
      RECT 55.005 1.935 55.175 2.105 ;
      RECT 55.005 3.055 55.175 3.225 ;
      RECT 54.78 1.415 54.95 1.585 ;
      RECT 54.78 4.135 54.95 4.305 ;
      RECT 54.765 2.495 54.935 2.665 ;
      RECT 54.32 1.415 54.49 1.585 ;
      RECT 54.32 4.135 54.49 4.305 ;
      RECT 54.045 1.935 54.215 2.105 ;
      RECT 54.045 3.475 54.215 3.645 ;
      RECT 53.86 1.415 54.03 1.585 ;
      RECT 53.86 4.135 54.03 4.305 ;
      RECT 52.43 0.915 52.6 1.085 ;
      RECT 52.43 2.395 52.6 2.565 ;
      RECT 52.43 6.315 52.6 6.485 ;
      RECT 52.43 7.795 52.6 7.965 ;
      RECT 52.08 0.105 52.25 0.275 ;
      RECT 52.08 4.165 52.25 4.335 ;
      RECT 52.08 4.545 52.25 4.715 ;
      RECT 52.08 8.605 52.25 8.775 ;
      RECT 52.06 2.765 52.23 2.935 ;
      RECT 52.06 5.945 52.23 6.115 ;
      RECT 51.44 0.915 51.61 1.085 ;
      RECT 51.44 2.395 51.61 2.565 ;
      RECT 51.44 6.315 51.61 6.485 ;
      RECT 51.44 7.795 51.61 7.965 ;
      RECT 51.09 0.105 51.26 0.275 ;
      RECT 51.09 4.165 51.26 4.335 ;
      RECT 51.09 4.545 51.26 4.715 ;
      RECT 51.09 8.605 51.26 8.775 ;
      RECT 51.07 2.765 51.24 2.935 ;
      RECT 51.07 5.945 51.24 6.115 ;
      RECT 50.385 0.105 50.555 0.275 ;
      RECT 50.385 4.165 50.555 4.335 ;
      RECT 50.385 4.545 50.555 4.715 ;
      RECT 50.385 8.605 50.555 8.775 ;
      RECT 50.075 2.025 50.245 2.195 ;
      RECT 50.075 6.685 50.245 6.855 ;
      RECT 49.705 0.105 49.875 0.275 ;
      RECT 49.705 8.605 49.875 8.775 ;
      RECT 49.645 0.915 49.815 1.085 ;
      RECT 49.645 1.655 49.815 1.825 ;
      RECT 49.645 7.055 49.815 7.225 ;
      RECT 49.645 7.795 49.815 7.965 ;
      RECT 49.27 2.395 49.44 2.565 ;
      RECT 49.27 6.315 49.44 6.485 ;
      RECT 49.025 0.105 49.195 0.275 ;
      RECT 49.025 8.605 49.195 8.775 ;
      RECT 48.345 0.105 48.515 0.275 ;
      RECT 48.345 8.605 48.515 8.775 ;
      RECT 48.275 2.765 48.445 2.935 ;
      RECT 48.275 5.945 48.445 6.115 ;
      RECT 46.8 1.415 46.97 1.585 ;
      RECT 46.8 4.135 46.97 4.305 ;
      RECT 46.34 1.415 46.51 1.585 ;
      RECT 46.34 4.135 46.51 4.305 ;
      RECT 45.965 2.775 46.135 2.945 ;
      RECT 45.88 1.415 46.05 1.585 ;
      RECT 45.88 4.135 46.05 4.305 ;
      RECT 45.725 1.935 45.895 2.105 ;
      RECT 45.485 3.055 45.655 3.225 ;
      RECT 45.42 1.415 45.59 1.585 ;
      RECT 45.42 4.135 45.59 4.305 ;
      RECT 45.005 2.495 45.175 2.665 ;
      RECT 44.96 1.415 45.13 1.585 ;
      RECT 44.96 4.135 45.13 4.305 ;
      RECT 44.77 4.545 44.94 4.715 ;
      RECT 44.77 8.605 44.94 8.775 ;
      RECT 44.765 1.935 44.935 2.105 ;
      RECT 44.765 3.055 44.935 3.225 ;
      RECT 44.765 3.615 44.935 3.785 ;
      RECT 44.5 1.415 44.67 1.585 ;
      RECT 44.5 4.135 44.67 4.305 ;
      RECT 44.46 6.685 44.63 6.855 ;
      RECT 44.285 3.055 44.455 3.225 ;
      RECT 44.09 8.605 44.26 8.775 ;
      RECT 44.04 1.415 44.21 1.585 ;
      RECT 44.04 4.135 44.21 4.305 ;
      RECT 44.03 7.055 44.2 7.225 ;
      RECT 44.03 7.795 44.2 7.965 ;
      RECT 43.765 2.775 43.935 2.945 ;
      RECT 43.765 3.615 43.935 3.785 ;
      RECT 43.655 6.315 43.825 6.485 ;
      RECT 43.58 1.415 43.75 1.585 ;
      RECT 43.58 4.135 43.75 4.305 ;
      RECT 43.41 8.605 43.58 8.775 ;
      RECT 43.285 1.935 43.455 2.105 ;
      RECT 43.285 3.615 43.455 3.785 ;
      RECT 43.12 1.415 43.29 1.585 ;
      RECT 43.12 4.135 43.29 4.305 ;
      RECT 42.73 8.605 42.9 8.775 ;
      RECT 42.66 1.415 42.83 1.585 ;
      RECT 42.66 4.135 42.83 4.305 ;
      RECT 42.66 5.945 42.83 6.115 ;
      RECT 42.325 1.935 42.495 2.105 ;
      RECT 42.325 2.495 42.495 2.665 ;
      RECT 42.325 3.055 42.495 3.225 ;
      RECT 42.325 3.615 42.495 3.785 ;
      RECT 42.2 1.415 42.37 1.585 ;
      RECT 42.2 4.135 42.37 4.305 ;
      RECT 41.805 3.615 41.975 3.785 ;
      RECT 41.74 1.415 41.91 1.585 ;
      RECT 41.74 4.135 41.91 4.305 ;
      RECT 41.325 1.935 41.495 2.105 ;
      RECT 41.28 1.415 41.45 1.585 ;
      RECT 41.28 4.135 41.45 4.305 ;
      RECT 41.085 2.495 41.255 2.665 ;
      RECT 40.82 1.415 40.99 1.585 ;
      RECT 40.82 4.135 40.99 4.305 ;
      RECT 40.605 2.495 40.775 2.665 ;
      RECT 40.605 3.055 40.775 3.225 ;
      RECT 40.365 1.935 40.535 2.105 ;
      RECT 40.36 1.415 40.53 1.585 ;
      RECT 40.36 4.135 40.53 4.305 ;
      RECT 39.9 1.415 40.07 1.585 ;
      RECT 39.9 4.135 40.07 4.305 ;
      RECT 39.885 3.055 40.055 3.225 ;
      RECT 39.44 1.415 39.61 1.585 ;
      RECT 39.44 4.135 39.61 4.305 ;
      RECT 39.365 2.495 39.535 2.665 ;
      RECT 39.365 3.335 39.535 3.505 ;
      RECT 38.98 1.415 39.15 1.585 ;
      RECT 38.98 4.135 39.15 4.305 ;
      RECT 38.885 1.935 39.055 2.105 ;
      RECT 38.885 3.055 39.055 3.225 ;
      RECT 38.645 2.495 38.815 2.665 ;
      RECT 38.52 1.415 38.69 1.585 ;
      RECT 38.52 4.135 38.69 4.305 ;
      RECT 38.405 3.335 38.575 3.505 ;
      RECT 38.165 2.775 38.335 2.945 ;
      RECT 38.06 1.415 38.23 1.585 ;
      RECT 38.06 4.135 38.23 4.305 ;
      RECT 37.6 1.415 37.77 1.585 ;
      RECT 37.6 4.135 37.77 4.305 ;
      RECT 37.36 2.495 37.53 2.665 ;
      RECT 37.14 1.415 37.31 1.585 ;
      RECT 37.14 4.135 37.31 4.305 ;
      RECT 36.925 3.055 37.095 3.225 ;
      RECT 36.68 1.415 36.85 1.585 ;
      RECT 36.68 4.135 36.85 4.305 ;
      RECT 36.445 1.935 36.615 2.105 ;
      RECT 36.445 3.055 36.615 3.225 ;
      RECT 36.22 1.415 36.39 1.585 ;
      RECT 36.22 4.135 36.39 4.305 ;
      RECT 36.205 2.495 36.375 2.665 ;
      RECT 35.76 1.415 35.93 1.585 ;
      RECT 35.76 4.135 35.93 4.305 ;
      RECT 35.485 1.935 35.655 2.105 ;
      RECT 35.485 3.475 35.655 3.645 ;
      RECT 35.3 1.415 35.47 1.585 ;
      RECT 35.3 4.135 35.47 4.305 ;
      RECT 33.87 0.915 34.04 1.085 ;
      RECT 33.87 2.395 34.04 2.565 ;
      RECT 33.87 6.315 34.04 6.485 ;
      RECT 33.87 7.795 34.04 7.965 ;
      RECT 33.52 0.105 33.69 0.275 ;
      RECT 33.52 4.165 33.69 4.335 ;
      RECT 33.52 4.545 33.69 4.715 ;
      RECT 33.52 8.605 33.69 8.775 ;
      RECT 33.5 2.765 33.67 2.935 ;
      RECT 33.5 5.945 33.67 6.115 ;
      RECT 32.88 0.915 33.05 1.085 ;
      RECT 32.88 2.395 33.05 2.565 ;
      RECT 32.88 6.315 33.05 6.485 ;
      RECT 32.88 7.795 33.05 7.965 ;
      RECT 32.53 0.105 32.7 0.275 ;
      RECT 32.53 4.165 32.7 4.335 ;
      RECT 32.53 4.545 32.7 4.715 ;
      RECT 32.53 8.605 32.7 8.775 ;
      RECT 32.51 2.765 32.68 2.935 ;
      RECT 32.51 5.945 32.68 6.115 ;
      RECT 31.825 0.105 31.995 0.275 ;
      RECT 31.825 4.165 31.995 4.335 ;
      RECT 31.825 4.545 31.995 4.715 ;
      RECT 31.825 8.605 31.995 8.775 ;
      RECT 31.515 2.025 31.685 2.195 ;
      RECT 31.515 6.685 31.685 6.855 ;
      RECT 31.145 0.105 31.315 0.275 ;
      RECT 31.145 8.605 31.315 8.775 ;
      RECT 31.085 0.915 31.255 1.085 ;
      RECT 31.085 1.655 31.255 1.825 ;
      RECT 31.085 7.055 31.255 7.225 ;
      RECT 31.085 7.795 31.255 7.965 ;
      RECT 30.71 2.395 30.88 2.565 ;
      RECT 30.71 6.315 30.88 6.485 ;
      RECT 30.465 0.105 30.635 0.275 ;
      RECT 30.465 8.605 30.635 8.775 ;
      RECT 29.785 0.105 29.955 0.275 ;
      RECT 29.785 8.605 29.955 8.775 ;
      RECT 29.715 2.765 29.885 2.935 ;
      RECT 29.715 5.945 29.885 6.115 ;
      RECT 28.24 1.415 28.41 1.585 ;
      RECT 28.24 4.135 28.41 4.305 ;
      RECT 27.78 1.415 27.95 1.585 ;
      RECT 27.78 4.135 27.95 4.305 ;
      RECT 27.405 2.775 27.575 2.945 ;
      RECT 27.32 1.415 27.49 1.585 ;
      RECT 27.32 4.135 27.49 4.305 ;
      RECT 27.165 1.935 27.335 2.105 ;
      RECT 26.925 3.055 27.095 3.225 ;
      RECT 26.86 1.415 27.03 1.585 ;
      RECT 26.86 4.135 27.03 4.305 ;
      RECT 26.445 2.495 26.615 2.665 ;
      RECT 26.4 1.415 26.57 1.585 ;
      RECT 26.4 4.135 26.57 4.305 ;
      RECT 26.21 4.545 26.38 4.715 ;
      RECT 26.21 8.605 26.38 8.775 ;
      RECT 26.205 1.935 26.375 2.105 ;
      RECT 26.205 3.055 26.375 3.225 ;
      RECT 26.205 3.615 26.375 3.785 ;
      RECT 25.94 1.415 26.11 1.585 ;
      RECT 25.94 4.135 26.11 4.305 ;
      RECT 25.9 6.685 26.07 6.855 ;
      RECT 25.725 3.055 25.895 3.225 ;
      RECT 25.53 8.605 25.7 8.775 ;
      RECT 25.48 1.415 25.65 1.585 ;
      RECT 25.48 4.135 25.65 4.305 ;
      RECT 25.47 7.055 25.64 7.225 ;
      RECT 25.47 7.795 25.64 7.965 ;
      RECT 25.205 2.775 25.375 2.945 ;
      RECT 25.205 3.615 25.375 3.785 ;
      RECT 25.095 6.315 25.265 6.485 ;
      RECT 25.02 1.415 25.19 1.585 ;
      RECT 25.02 4.135 25.19 4.305 ;
      RECT 24.85 8.605 25.02 8.775 ;
      RECT 24.725 1.935 24.895 2.105 ;
      RECT 24.725 3.615 24.895 3.785 ;
      RECT 24.56 1.415 24.73 1.585 ;
      RECT 24.56 4.135 24.73 4.305 ;
      RECT 24.17 8.605 24.34 8.775 ;
      RECT 24.1 1.415 24.27 1.585 ;
      RECT 24.1 4.135 24.27 4.305 ;
      RECT 24.1 5.945 24.27 6.115 ;
      RECT 23.765 1.935 23.935 2.105 ;
      RECT 23.765 2.495 23.935 2.665 ;
      RECT 23.765 3.055 23.935 3.225 ;
      RECT 23.765 3.615 23.935 3.785 ;
      RECT 23.64 1.415 23.81 1.585 ;
      RECT 23.64 4.135 23.81 4.305 ;
      RECT 23.245 3.615 23.415 3.785 ;
      RECT 23.18 1.415 23.35 1.585 ;
      RECT 23.18 4.135 23.35 4.305 ;
      RECT 22.765 1.935 22.935 2.105 ;
      RECT 22.72 1.415 22.89 1.585 ;
      RECT 22.72 4.135 22.89 4.305 ;
      RECT 22.525 2.495 22.695 2.665 ;
      RECT 22.26 1.415 22.43 1.585 ;
      RECT 22.26 4.135 22.43 4.305 ;
      RECT 22.045 2.495 22.215 2.665 ;
      RECT 22.045 3.055 22.215 3.225 ;
      RECT 21.805 1.935 21.975 2.105 ;
      RECT 21.8 1.415 21.97 1.585 ;
      RECT 21.8 4.135 21.97 4.305 ;
      RECT 21.34 1.415 21.51 1.585 ;
      RECT 21.34 4.135 21.51 4.305 ;
      RECT 21.325 3.055 21.495 3.225 ;
      RECT 20.88 1.415 21.05 1.585 ;
      RECT 20.88 4.135 21.05 4.305 ;
      RECT 20.805 2.495 20.975 2.665 ;
      RECT 20.805 3.335 20.975 3.505 ;
      RECT 20.42 1.415 20.59 1.585 ;
      RECT 20.42 4.135 20.59 4.305 ;
      RECT 20.325 1.935 20.495 2.105 ;
      RECT 20.325 3.055 20.495 3.225 ;
      RECT 20.085 2.495 20.255 2.665 ;
      RECT 19.96 1.415 20.13 1.585 ;
      RECT 19.96 4.135 20.13 4.305 ;
      RECT 19.845 3.335 20.015 3.505 ;
      RECT 19.605 2.775 19.775 2.945 ;
      RECT 19.5 1.415 19.67 1.585 ;
      RECT 19.5 4.135 19.67 4.305 ;
      RECT 19.04 1.415 19.21 1.585 ;
      RECT 19.04 4.135 19.21 4.305 ;
      RECT 18.8 2.495 18.97 2.665 ;
      RECT 18.58 1.415 18.75 1.585 ;
      RECT 18.58 4.135 18.75 4.305 ;
      RECT 18.365 3.055 18.535 3.225 ;
      RECT 18.12 1.415 18.29 1.585 ;
      RECT 18.12 4.135 18.29 4.305 ;
      RECT 17.885 1.935 18.055 2.105 ;
      RECT 17.885 3.055 18.055 3.225 ;
      RECT 17.66 1.415 17.83 1.585 ;
      RECT 17.66 4.135 17.83 4.305 ;
      RECT 17.645 2.495 17.815 2.665 ;
      RECT 17.2 1.415 17.37 1.585 ;
      RECT 17.2 4.135 17.37 4.305 ;
      RECT 16.925 1.935 17.095 2.105 ;
      RECT 16.925 3.475 17.095 3.645 ;
      RECT 16.74 1.415 16.91 1.585 ;
      RECT 16.74 4.135 16.91 4.305 ;
      RECT 15.31 0.915 15.48 1.085 ;
      RECT 15.31 2.395 15.48 2.565 ;
      RECT 15.31 6.315 15.48 6.485 ;
      RECT 15.31 7.795 15.48 7.965 ;
      RECT 14.96 0.105 15.13 0.275 ;
      RECT 14.96 4.165 15.13 4.335 ;
      RECT 14.96 4.545 15.13 4.715 ;
      RECT 14.96 8.605 15.13 8.775 ;
      RECT 14.94 2.765 15.11 2.935 ;
      RECT 14.94 5.945 15.11 6.115 ;
      RECT 14.32 0.915 14.49 1.085 ;
      RECT 14.32 2.395 14.49 2.565 ;
      RECT 14.32 6.315 14.49 6.485 ;
      RECT 14.32 7.795 14.49 7.965 ;
      RECT 13.97 0.105 14.14 0.275 ;
      RECT 13.97 4.165 14.14 4.335 ;
      RECT 13.97 4.545 14.14 4.715 ;
      RECT 13.97 8.605 14.14 8.775 ;
      RECT 13.95 2.765 14.12 2.935 ;
      RECT 13.95 5.945 14.12 6.115 ;
      RECT 13.265 0.105 13.435 0.275 ;
      RECT 13.265 4.165 13.435 4.335 ;
      RECT 13.265 4.545 13.435 4.715 ;
      RECT 13.265 8.605 13.435 8.775 ;
      RECT 12.955 2.025 13.125 2.195 ;
      RECT 12.955 6.685 13.125 6.855 ;
      RECT 12.585 0.105 12.755 0.275 ;
      RECT 12.585 8.605 12.755 8.775 ;
      RECT 12.525 0.915 12.695 1.085 ;
      RECT 12.525 1.655 12.695 1.825 ;
      RECT 12.525 7.055 12.695 7.225 ;
      RECT 12.525 7.795 12.695 7.965 ;
      RECT 12.15 2.395 12.32 2.565 ;
      RECT 12.15 6.315 12.32 6.485 ;
      RECT 11.905 0.105 12.075 0.275 ;
      RECT 11.905 8.605 12.075 8.775 ;
      RECT 11.225 0.105 11.395 0.275 ;
      RECT 11.225 8.605 11.395 8.775 ;
      RECT 11.155 2.765 11.325 2.935 ;
      RECT 11.155 5.945 11.325 6.115 ;
      RECT 9.68 1.415 9.85 1.585 ;
      RECT 9.68 4.135 9.85 4.305 ;
      RECT 9.22 1.415 9.39 1.585 ;
      RECT 9.22 4.135 9.39 4.305 ;
      RECT 8.845 2.775 9.015 2.945 ;
      RECT 8.76 1.415 8.93 1.585 ;
      RECT 8.76 4.135 8.93 4.305 ;
      RECT 8.605 1.935 8.775 2.105 ;
      RECT 8.365 3.055 8.535 3.225 ;
      RECT 8.3 1.415 8.47 1.585 ;
      RECT 8.3 4.135 8.47 4.305 ;
      RECT 7.885 2.495 8.055 2.665 ;
      RECT 7.84 1.415 8.01 1.585 ;
      RECT 7.84 4.135 8.01 4.305 ;
      RECT 7.65 4.545 7.82 4.715 ;
      RECT 7.65 8.605 7.82 8.775 ;
      RECT 7.645 1.935 7.815 2.105 ;
      RECT 7.645 3.055 7.815 3.225 ;
      RECT 7.645 3.615 7.815 3.785 ;
      RECT 7.38 1.415 7.55 1.585 ;
      RECT 7.38 4.135 7.55 4.305 ;
      RECT 7.34 6.685 7.51 6.855 ;
      RECT 7.165 3.055 7.335 3.225 ;
      RECT 6.97 8.605 7.14 8.775 ;
      RECT 6.92 1.415 7.09 1.585 ;
      RECT 6.92 4.135 7.09 4.305 ;
      RECT 6.91 7.055 7.08 7.225 ;
      RECT 6.91 7.795 7.08 7.965 ;
      RECT 6.645 2.775 6.815 2.945 ;
      RECT 6.645 3.615 6.815 3.785 ;
      RECT 6.535 6.315 6.705 6.485 ;
      RECT 6.46 1.415 6.63 1.585 ;
      RECT 6.46 4.135 6.63 4.305 ;
      RECT 6.29 8.605 6.46 8.775 ;
      RECT 6.165 1.935 6.335 2.105 ;
      RECT 6.165 3.615 6.335 3.785 ;
      RECT 6 1.415 6.17 1.585 ;
      RECT 6 4.135 6.17 4.305 ;
      RECT 5.61 8.605 5.78 8.775 ;
      RECT 5.54 1.415 5.71 1.585 ;
      RECT 5.54 4.135 5.71 4.305 ;
      RECT 5.54 5.945 5.71 6.115 ;
      RECT 5.205 1.935 5.375 2.105 ;
      RECT 5.205 2.495 5.375 2.665 ;
      RECT 5.205 3.055 5.375 3.225 ;
      RECT 5.205 3.615 5.375 3.785 ;
      RECT 5.08 1.415 5.25 1.585 ;
      RECT 5.08 4.135 5.25 4.305 ;
      RECT 4.685 3.615 4.855 3.785 ;
      RECT 4.62 1.415 4.79 1.585 ;
      RECT 4.62 4.135 4.79 4.305 ;
      RECT 4.205 1.935 4.375 2.105 ;
      RECT 4.16 1.415 4.33 1.585 ;
      RECT 4.16 4.135 4.33 4.305 ;
      RECT 3.965 2.495 4.135 2.665 ;
      RECT 3.7 1.415 3.87 1.585 ;
      RECT 3.7 4.135 3.87 4.305 ;
      RECT 3.485 2.495 3.655 2.665 ;
      RECT 3.485 3.055 3.655 3.225 ;
      RECT 3.245 1.935 3.415 2.105 ;
      RECT 3.24 1.415 3.41 1.585 ;
      RECT 3.24 4.135 3.41 4.305 ;
      RECT 2.78 1.415 2.95 1.585 ;
      RECT 2.78 4.135 2.95 4.305 ;
      RECT 2.765 3.055 2.935 3.225 ;
      RECT 2.32 1.415 2.49 1.585 ;
      RECT 2.32 4.135 2.49 4.305 ;
      RECT 2.245 2.495 2.415 2.665 ;
      RECT 2.245 3.335 2.415 3.505 ;
      RECT 1.86 1.415 2.03 1.585 ;
      RECT 1.86 4.135 2.03 4.305 ;
      RECT 1.765 1.935 1.935 2.105 ;
      RECT 1.765 3.055 1.935 3.225 ;
      RECT 1.525 2.495 1.695 2.665 ;
      RECT 1.4 1.415 1.57 1.585 ;
      RECT 1.4 4.135 1.57 4.305 ;
      RECT 1.285 3.335 1.455 3.505 ;
      RECT 1.045 2.775 1.215 2.945 ;
      RECT 0.94 1.415 1.11 1.585 ;
      RECT 0.94 4.135 1.11 4.305 ;
      RECT 0.48 1.415 0.65 1.585 ;
      RECT 0.48 4.135 0.65 4.305 ;
      RECT 0.24 2.495 0.41 2.665 ;
      RECT 0.02 1.415 0.19 1.585 ;
      RECT 0.02 4.135 0.19 4.305 ;
      RECT -0.195 3.055 -0.025 3.225 ;
      RECT -0.44 1.415 -0.27 1.585 ;
      RECT -0.44 4.135 -0.27 4.305 ;
      RECT -0.675 1.935 -0.505 2.105 ;
      RECT -0.675 3.055 -0.505 3.225 ;
      RECT -0.9 1.415 -0.73 1.585 ;
      RECT -0.9 4.135 -0.73 4.305 ;
      RECT -0.915 2.495 -0.745 2.665 ;
      RECT -1.36 1.415 -1.19 1.585 ;
      RECT -1.36 4.135 -1.19 4.305 ;
      RECT -1.635 1.935 -1.465 2.105 ;
      RECT -1.635 3.475 -1.465 3.645 ;
      RECT -1.82 1.415 -1.65 1.585 ;
      RECT -1.82 4.135 -1.65 4.305 ;
      RECT -3.165 4.545 -2.995 4.715 ;
      RECT -3.165 8.605 -2.995 8.775 ;
      RECT -3.475 6.685 -3.305 6.855 ;
      RECT -3.845 8.605 -3.675 8.775 ;
      RECT -3.905 7.055 -3.735 7.225 ;
      RECT -3.905 7.795 -3.735 7.965 ;
      RECT -4.28 6.315 -4.11 6.485 ;
      RECT -4.525 8.605 -4.355 8.775 ;
      RECT -5.205 8.605 -5.035 8.775 ;
      RECT -5.275 5.945 -5.105 6.115 ;
    LAYER li ;
      RECT 83.325 0 83.495 2.085 ;
      RECT 82.365 0 82.535 2.085 ;
      RECT 81.405 0 81.575 2.085 ;
      RECT 80.885 0 81.055 2.085 ;
      RECT 79.925 0 80.095 2.085 ;
      RECT 78.925 0 79.095 2.085 ;
      RECT 77.965 0 78.135 2.085 ;
      RECT 76.485 0 76.655 2.085 ;
      RECT 74.565 0 74.735 2.085 ;
      RECT 73.085 0 73.255 2.085 ;
      RECT 64.765 0 64.935 2.085 ;
      RECT 63.805 0 63.975 2.085 ;
      RECT 62.845 0 63.015 2.085 ;
      RECT 62.325 0 62.495 2.085 ;
      RECT 61.365 0 61.535 2.085 ;
      RECT 60.365 0 60.535 2.085 ;
      RECT 59.405 0 59.575 2.085 ;
      RECT 57.925 0 58.095 2.085 ;
      RECT 56.005 0 56.175 2.085 ;
      RECT 54.525 0 54.695 2.085 ;
      RECT 46.205 0 46.375 2.085 ;
      RECT 45.245 0 45.415 2.085 ;
      RECT 44.285 0 44.455 2.085 ;
      RECT 43.765 0 43.935 2.085 ;
      RECT 42.805 0 42.975 2.085 ;
      RECT 41.805 0 41.975 2.085 ;
      RECT 40.845 0 41.015 2.085 ;
      RECT 39.365 0 39.535 2.085 ;
      RECT 37.445 0 37.615 2.085 ;
      RECT 35.965 0 36.135 2.085 ;
      RECT 27.645 0 27.815 2.085 ;
      RECT 26.685 0 26.855 2.085 ;
      RECT 25.725 0 25.895 2.085 ;
      RECT 25.205 0 25.375 2.085 ;
      RECT 24.245 0 24.415 2.085 ;
      RECT 23.245 0 23.415 2.085 ;
      RECT 22.285 0 22.455 2.085 ;
      RECT 20.805 0 20.975 2.085 ;
      RECT 18.885 0 19.055 2.085 ;
      RECT 17.405 0 17.575 2.085 ;
      RECT 9.085 0 9.255 2.085 ;
      RECT 8.125 0 8.295 2.085 ;
      RECT 7.165 0 7.335 2.085 ;
      RECT 6.645 0 6.815 2.085 ;
      RECT 5.685 0 5.855 2.085 ;
      RECT 4.685 0 4.855 2.085 ;
      RECT 3.725 0 3.895 2.085 ;
      RECT 2.245 0 2.415 2.085 ;
      RECT 0.325 0 0.495 2.085 ;
      RECT -1.155 0 -0.985 2.085 ;
      RECT 80.605 0 80.8 1.595 ;
      RECT 76.93 0 77.125 1.595 ;
      RECT 74.565 0 74.825 1.595 ;
      RECT 62.045 0 62.24 1.595 ;
      RECT 58.37 0 58.565 1.595 ;
      RECT 56.005 0 56.265 1.595 ;
      RECT 43.485 0 43.68 1.595 ;
      RECT 39.81 0 40.005 1.595 ;
      RECT 37.445 0 37.705 1.595 ;
      RECT 24.925 0 25.12 1.595 ;
      RECT 21.25 0 21.445 1.595 ;
      RECT 18.885 0 19.145 1.595 ;
      RECT 6.365 0 6.56 1.595 ;
      RECT 2.69 0 2.885 1.595 ;
      RECT 0.325 0 0.585 1.595 ;
      RECT 72.275 0 84.32 1.585 ;
      RECT 53.715 0 65.76 1.585 ;
      RECT 35.155 0 47.2 1.585 ;
      RECT 16.595 0 28.64 1.585 ;
      RECT -1.965 0 10.08 1.585 ;
      RECT 89.12 0 89.29 0.935 ;
      RECT 88.13 0 88.3 0.935 ;
      RECT 85.385 0 85.555 0.935 ;
      RECT 70.56 0 70.73 0.935 ;
      RECT 69.57 0 69.74 0.935 ;
      RECT 66.825 0 66.995 0.935 ;
      RECT 52 0 52.17 0.935 ;
      RECT 51.01 0 51.18 0.935 ;
      RECT 48.265 0 48.435 0.935 ;
      RECT 33.44 0 33.61 0.935 ;
      RECT 32.45 0 32.62 0.935 ;
      RECT 29.705 0 29.875 0.935 ;
      RECT 14.88 0 15.05 0.935 ;
      RECT 13.89 0 14.06 0.935 ;
      RECT 11.145 0 11.315 0.935 ;
      RECT -5.465 0 90.09 0.305 ;
      RECT -3.475 4.145 -3.305 8.305 ;
      RECT 89.12 3.405 89.29 5.475 ;
      RECT 88.13 3.405 88.3 5.475 ;
      RECT 85.385 3.405 85.555 5.475 ;
      RECT 79.77 4.135 79.94 5.475 ;
      RECT 70.56 3.405 70.73 5.475 ;
      RECT 69.57 3.405 69.74 5.475 ;
      RECT 66.825 3.405 66.995 5.475 ;
      RECT 61.21 4.135 61.38 5.475 ;
      RECT 52 3.405 52.17 5.475 ;
      RECT 51.01 3.405 51.18 5.475 ;
      RECT 48.265 3.405 48.435 5.475 ;
      RECT 42.65 4.135 42.82 5.475 ;
      RECT 33.44 3.405 33.61 5.475 ;
      RECT 32.45 3.405 32.62 5.475 ;
      RECT 29.705 3.405 29.875 5.475 ;
      RECT 24.09 4.135 24.26 5.475 ;
      RECT 14.88 3.405 15.05 5.475 ;
      RECT 13.89 3.405 14.06 5.475 ;
      RECT 11.145 3.405 11.315 5.475 ;
      RECT 5.53 4.135 5.7 5.475 ;
      RECT -5.285 4.145 -5.115 5.475 ;
      RECT 71.53 4.145 73.995 4.75 ;
      RECT 52.97 4.145 55.435 4.75 ;
      RECT 34.41 4.145 36.875 4.75 ;
      RECT 15.85 4.145 18.315 4.75 ;
      RECT -5.46 4.145 -0.245 4.75 ;
      RECT 72.275 4.135 90.09 4.745 ;
      RECT 53.715 4.135 71.53 4.745 ;
      RECT 35.155 4.135 52.97 4.745 ;
      RECT 16.595 4.135 34.41 4.745 ;
      RECT -1.965 4.135 15.85 4.745 ;
      RECT 82.365 3.635 82.535 4.745 ;
      RECT 79.925 3.635 80.095 4.745 ;
      RECT 77.965 3.635 78.135 4.745 ;
      RECT 77.005 3.635 77.175 4.745 ;
      RECT 75.045 3.635 75.215 4.745 ;
      RECT 74.045 3.635 74.215 4.745 ;
      RECT 73.085 3.635 73.255 4.75 ;
      RECT 63.805 3.635 63.975 4.745 ;
      RECT 61.365 3.635 61.535 4.745 ;
      RECT 59.405 3.635 59.575 4.745 ;
      RECT 58.445 3.635 58.615 4.745 ;
      RECT 56.485 3.635 56.655 4.745 ;
      RECT 55.485 3.635 55.655 4.745 ;
      RECT 54.525 3.635 54.695 4.75 ;
      RECT 45.245 3.635 45.415 4.745 ;
      RECT 42.805 3.635 42.975 4.745 ;
      RECT 40.845 3.635 41.015 4.745 ;
      RECT 39.885 3.635 40.055 4.745 ;
      RECT 37.925 3.635 38.095 4.745 ;
      RECT 36.925 3.635 37.095 4.745 ;
      RECT 35.965 3.635 36.135 4.75 ;
      RECT 26.685 3.635 26.855 4.745 ;
      RECT 24.245 3.635 24.415 4.745 ;
      RECT 22.285 3.635 22.455 4.745 ;
      RECT 21.325 3.635 21.495 4.745 ;
      RECT 19.365 3.635 19.535 4.745 ;
      RECT 18.365 3.635 18.535 4.745 ;
      RECT 17.405 3.635 17.575 4.75 ;
      RECT 8.125 3.635 8.295 4.745 ;
      RECT 5.685 3.635 5.855 4.745 ;
      RECT 3.725 3.635 3.895 4.745 ;
      RECT 2.765 3.635 2.935 4.745 ;
      RECT 0.805 3.635 0.975 4.745 ;
      RECT -0.195 3.635 -0.025 4.745 ;
      RECT -1.155 3.635 -0.985 4.75 ;
      RECT -5.465 8.575 90.09 8.88 ;
      RECT 89.12 7.945 89.29 8.88 ;
      RECT 88.13 7.945 88.3 8.88 ;
      RECT 85.385 7.945 85.555 8.88 ;
      RECT 79.77 7.945 79.94 8.88 ;
      RECT 70.56 7.945 70.73 8.88 ;
      RECT 69.57 7.945 69.74 8.88 ;
      RECT 66.825 7.945 66.995 8.88 ;
      RECT 61.21 7.945 61.38 8.88 ;
      RECT 52 7.945 52.17 8.88 ;
      RECT 51.01 7.945 51.18 8.88 ;
      RECT 48.265 7.945 48.435 8.88 ;
      RECT 42.65 7.945 42.82 8.88 ;
      RECT 33.44 7.945 33.61 8.88 ;
      RECT 32.45 7.945 32.62 8.88 ;
      RECT 29.705 7.945 29.875 8.88 ;
      RECT 24.09 7.945 24.26 8.88 ;
      RECT 14.88 7.945 15.05 8.88 ;
      RECT 13.89 7.945 14.06 8.88 ;
      RECT 11.145 7.945 11.315 8.88 ;
      RECT 5.53 7.945 5.7 8.88 ;
      RECT -5.285 7.945 -5.115 8.88 ;
      RECT 89.18 1.74 89.35 2.935 ;
      RECT 89.18 1.74 89.645 1.91 ;
      RECT 89.18 6.97 89.645 7.14 ;
      RECT 89.18 5.945 89.35 7.14 ;
      RECT 88.19 1.74 88.36 2.935 ;
      RECT 88.19 1.74 88.655 1.91 ;
      RECT 88.19 6.97 88.655 7.14 ;
      RECT 88.19 5.945 88.36 7.14 ;
      RECT 86.335 2.635 86.505 3.865 ;
      RECT 86.39 0.855 86.56 2.805 ;
      RECT 86.335 0.575 86.505 1.025 ;
      RECT 86.335 7.855 86.505 8.305 ;
      RECT 86.39 6.075 86.56 8.025 ;
      RECT 86.335 5.015 86.505 6.245 ;
      RECT 85.815 0.575 85.985 3.865 ;
      RECT 85.815 2.075 86.22 2.405 ;
      RECT 85.815 1.235 86.22 1.565 ;
      RECT 85.815 5.015 85.985 8.305 ;
      RECT 85.815 7.315 86.22 7.645 ;
      RECT 85.815 6.475 86.22 6.805 ;
      RECT 82.605 3.225 83.575 3.395 ;
      RECT 82.605 3.055 82.775 3.395 ;
      RECT 82.125 2.495 82.295 2.825 ;
      RECT 82.125 2.575 82.855 2.745 ;
      RECT 81.765 3.615 82.055 3.785 ;
      RECT 81.765 2.575 81.935 3.785 ;
      RECT 81.765 3.055 82.055 3.225 ;
      RECT 81.565 2.575 81.935 2.745 ;
      RECT 80.885 2.675 81.055 2.945 ;
      RECT 80.645 2.675 81.055 2.845 ;
      RECT 80.565 2.575 80.895 2.745 ;
      RECT 80.405 3.615 81.055 3.785 ;
      RECT 80.885 3.145 81.055 3.785 ;
      RECT 80.765 3.225 81.055 3.785 ;
      RECT 80.72 7.855 80.89 8.305 ;
      RECT 80.775 6.075 80.945 8.025 ;
      RECT 80.72 5.015 80.89 6.245 ;
      RECT 80.2 5.015 80.37 8.305 ;
      RECT 80.2 7.315 80.605 7.645 ;
      RECT 80.2 6.475 80.605 6.805 ;
      RECT 79.445 2.915 79.615 3.225 ;
      RECT 79.445 2.915 80.335 3.085 ;
      RECT 80.165 2.495 80.335 3.085 ;
      RECT 79.445 2.575 79.935 2.745 ;
      RECT 79.445 2.495 79.615 2.745 ;
      RECT 77.405 3.225 77.895 3.395 ;
      RECT 78.565 2.575 78.735 3.225 ;
      RECT 77.725 3.055 78.735 3.225 ;
      RECT 78.685 2.495 78.855 2.825 ;
      RECT 77.485 1.835 77.655 2.105 ;
      RECT 76.925 1.835 77.655 2.005 ;
      RECT 77.005 2.575 77.175 3.225 ;
      RECT 77.005 2.575 77.495 2.745 ;
      RECT 76.165 2.575 76.655 2.745 ;
      RECT 76.485 2.495 76.655 2.745 ;
      RECT 76.005 1.835 76.175 2.105 ;
      RECT 75.445 1.835 76.175 2.005 ;
      RECT 75.525 3.225 75.695 3.505 ;
      RECT 74.485 3.225 75.775 3.395 ;
      RECT 74.48 2.575 75.055 2.745 ;
      RECT 74.48 2.495 74.65 2.745 ;
      RECT 73.565 1.835 73.735 2.105 ;
      RECT 73.565 1.835 74.295 2.005 ;
      RECT 73.925 3.055 74.215 3.225 ;
      RECT 73.925 2.575 74.095 3.225 ;
      RECT 73.725 2.575 74.095 2.745 ;
      RECT 73.565 3.055 73.735 3.475 ;
      RECT 72.945 3.14 73.735 3.31 ;
      RECT 72.945 2.915 73.115 3.31 ;
      RECT 72.845 2.495 73.015 3.085 ;
      RECT 72.605 2.575 73.015 2.845 ;
      RECT 70.62 1.74 70.79 2.935 ;
      RECT 70.62 1.74 71.085 1.91 ;
      RECT 70.62 6.97 71.085 7.14 ;
      RECT 70.62 5.945 70.79 7.14 ;
      RECT 69.63 1.74 69.8 2.935 ;
      RECT 69.63 1.74 70.095 1.91 ;
      RECT 69.63 6.97 70.095 7.14 ;
      RECT 69.63 5.945 69.8 7.14 ;
      RECT 67.775 2.635 67.945 3.865 ;
      RECT 67.83 0.855 68 2.805 ;
      RECT 67.775 0.575 67.945 1.025 ;
      RECT 67.775 7.855 67.945 8.305 ;
      RECT 67.83 6.075 68 8.025 ;
      RECT 67.775 5.015 67.945 6.245 ;
      RECT 67.255 0.575 67.425 3.865 ;
      RECT 67.255 2.075 67.66 2.405 ;
      RECT 67.255 1.235 67.66 1.565 ;
      RECT 67.255 5.015 67.425 8.305 ;
      RECT 67.255 7.315 67.66 7.645 ;
      RECT 67.255 6.475 67.66 6.805 ;
      RECT 64.045 3.225 65.015 3.395 ;
      RECT 64.045 3.055 64.215 3.395 ;
      RECT 63.565 2.495 63.735 2.825 ;
      RECT 63.565 2.575 64.295 2.745 ;
      RECT 63.205 3.615 63.495 3.785 ;
      RECT 63.205 2.575 63.375 3.785 ;
      RECT 63.205 3.055 63.495 3.225 ;
      RECT 63.005 2.575 63.375 2.745 ;
      RECT 62.325 2.675 62.495 2.945 ;
      RECT 62.085 2.675 62.495 2.845 ;
      RECT 62.005 2.575 62.335 2.745 ;
      RECT 61.845 3.615 62.495 3.785 ;
      RECT 62.325 3.145 62.495 3.785 ;
      RECT 62.205 3.225 62.495 3.785 ;
      RECT 62.16 7.855 62.33 8.305 ;
      RECT 62.215 6.075 62.385 8.025 ;
      RECT 62.16 5.015 62.33 6.245 ;
      RECT 61.64 5.015 61.81 8.305 ;
      RECT 61.64 7.315 62.045 7.645 ;
      RECT 61.64 6.475 62.045 6.805 ;
      RECT 60.885 2.915 61.055 3.225 ;
      RECT 60.885 2.915 61.775 3.085 ;
      RECT 61.605 2.495 61.775 3.085 ;
      RECT 60.885 2.575 61.375 2.745 ;
      RECT 60.885 2.495 61.055 2.745 ;
      RECT 58.845 3.225 59.335 3.395 ;
      RECT 60.005 2.575 60.175 3.225 ;
      RECT 59.165 3.055 60.175 3.225 ;
      RECT 60.125 2.495 60.295 2.825 ;
      RECT 58.925 1.835 59.095 2.105 ;
      RECT 58.365 1.835 59.095 2.005 ;
      RECT 58.445 2.575 58.615 3.225 ;
      RECT 58.445 2.575 58.935 2.745 ;
      RECT 57.605 2.575 58.095 2.745 ;
      RECT 57.925 2.495 58.095 2.745 ;
      RECT 57.445 1.835 57.615 2.105 ;
      RECT 56.885 1.835 57.615 2.005 ;
      RECT 56.965 3.225 57.135 3.505 ;
      RECT 55.925 3.225 57.215 3.395 ;
      RECT 55.92 2.575 56.495 2.745 ;
      RECT 55.92 2.495 56.09 2.745 ;
      RECT 55.005 1.835 55.175 2.105 ;
      RECT 55.005 1.835 55.735 2.005 ;
      RECT 55.365 3.055 55.655 3.225 ;
      RECT 55.365 2.575 55.535 3.225 ;
      RECT 55.165 2.575 55.535 2.745 ;
      RECT 55.005 3.055 55.175 3.475 ;
      RECT 54.385 3.14 55.175 3.31 ;
      RECT 54.385 2.915 54.555 3.31 ;
      RECT 54.285 2.495 54.455 3.085 ;
      RECT 54.045 2.575 54.455 2.845 ;
      RECT 52.06 1.74 52.23 2.935 ;
      RECT 52.06 1.74 52.525 1.91 ;
      RECT 52.06 6.97 52.525 7.14 ;
      RECT 52.06 5.945 52.23 7.14 ;
      RECT 51.07 1.74 51.24 2.935 ;
      RECT 51.07 1.74 51.535 1.91 ;
      RECT 51.07 6.97 51.535 7.14 ;
      RECT 51.07 5.945 51.24 7.14 ;
      RECT 49.215 2.635 49.385 3.865 ;
      RECT 49.27 0.855 49.44 2.805 ;
      RECT 49.215 0.575 49.385 1.025 ;
      RECT 49.215 7.855 49.385 8.305 ;
      RECT 49.27 6.075 49.44 8.025 ;
      RECT 49.215 5.015 49.385 6.245 ;
      RECT 48.695 0.575 48.865 3.865 ;
      RECT 48.695 2.075 49.1 2.405 ;
      RECT 48.695 1.235 49.1 1.565 ;
      RECT 48.695 5.015 48.865 8.305 ;
      RECT 48.695 7.315 49.1 7.645 ;
      RECT 48.695 6.475 49.1 6.805 ;
      RECT 45.485 3.225 46.455 3.395 ;
      RECT 45.485 3.055 45.655 3.395 ;
      RECT 45.005 2.495 45.175 2.825 ;
      RECT 45.005 2.575 45.735 2.745 ;
      RECT 44.645 3.615 44.935 3.785 ;
      RECT 44.645 2.575 44.815 3.785 ;
      RECT 44.645 3.055 44.935 3.225 ;
      RECT 44.445 2.575 44.815 2.745 ;
      RECT 43.765 2.675 43.935 2.945 ;
      RECT 43.525 2.675 43.935 2.845 ;
      RECT 43.445 2.575 43.775 2.745 ;
      RECT 43.285 3.615 43.935 3.785 ;
      RECT 43.765 3.145 43.935 3.785 ;
      RECT 43.645 3.225 43.935 3.785 ;
      RECT 43.6 7.855 43.77 8.305 ;
      RECT 43.655 6.075 43.825 8.025 ;
      RECT 43.6 5.015 43.77 6.245 ;
      RECT 43.08 5.015 43.25 8.305 ;
      RECT 43.08 7.315 43.485 7.645 ;
      RECT 43.08 6.475 43.485 6.805 ;
      RECT 42.325 2.915 42.495 3.225 ;
      RECT 42.325 2.915 43.215 3.085 ;
      RECT 43.045 2.495 43.215 3.085 ;
      RECT 42.325 2.575 42.815 2.745 ;
      RECT 42.325 2.495 42.495 2.745 ;
      RECT 40.285 3.225 40.775 3.395 ;
      RECT 41.445 2.575 41.615 3.225 ;
      RECT 40.605 3.055 41.615 3.225 ;
      RECT 41.565 2.495 41.735 2.825 ;
      RECT 40.365 1.835 40.535 2.105 ;
      RECT 39.805 1.835 40.535 2.005 ;
      RECT 39.885 2.575 40.055 3.225 ;
      RECT 39.885 2.575 40.375 2.745 ;
      RECT 39.045 2.575 39.535 2.745 ;
      RECT 39.365 2.495 39.535 2.745 ;
      RECT 38.885 1.835 39.055 2.105 ;
      RECT 38.325 1.835 39.055 2.005 ;
      RECT 38.405 3.225 38.575 3.505 ;
      RECT 37.365 3.225 38.655 3.395 ;
      RECT 37.36 2.575 37.935 2.745 ;
      RECT 37.36 2.495 37.53 2.745 ;
      RECT 36.445 1.835 36.615 2.105 ;
      RECT 36.445 1.835 37.175 2.005 ;
      RECT 36.805 3.055 37.095 3.225 ;
      RECT 36.805 2.575 36.975 3.225 ;
      RECT 36.605 2.575 36.975 2.745 ;
      RECT 36.445 3.055 36.615 3.475 ;
      RECT 35.825 3.14 36.615 3.31 ;
      RECT 35.825 2.915 35.995 3.31 ;
      RECT 35.725 2.495 35.895 3.085 ;
      RECT 35.485 2.575 35.895 2.845 ;
      RECT 33.5 1.74 33.67 2.935 ;
      RECT 33.5 1.74 33.965 1.91 ;
      RECT 33.5 6.97 33.965 7.14 ;
      RECT 33.5 5.945 33.67 7.14 ;
      RECT 32.51 1.74 32.68 2.935 ;
      RECT 32.51 1.74 32.975 1.91 ;
      RECT 32.51 6.97 32.975 7.14 ;
      RECT 32.51 5.945 32.68 7.14 ;
      RECT 30.655 2.635 30.825 3.865 ;
      RECT 30.71 0.855 30.88 2.805 ;
      RECT 30.655 0.575 30.825 1.025 ;
      RECT 30.655 7.855 30.825 8.305 ;
      RECT 30.71 6.075 30.88 8.025 ;
      RECT 30.655 5.015 30.825 6.245 ;
      RECT 30.135 0.575 30.305 3.865 ;
      RECT 30.135 2.075 30.54 2.405 ;
      RECT 30.135 1.235 30.54 1.565 ;
      RECT 30.135 5.015 30.305 8.305 ;
      RECT 30.135 7.315 30.54 7.645 ;
      RECT 30.135 6.475 30.54 6.805 ;
      RECT 26.925 3.225 27.895 3.395 ;
      RECT 26.925 3.055 27.095 3.395 ;
      RECT 26.445 2.495 26.615 2.825 ;
      RECT 26.445 2.575 27.175 2.745 ;
      RECT 26.085 3.615 26.375 3.785 ;
      RECT 26.085 2.575 26.255 3.785 ;
      RECT 26.085 3.055 26.375 3.225 ;
      RECT 25.885 2.575 26.255 2.745 ;
      RECT 25.205 2.675 25.375 2.945 ;
      RECT 24.965 2.675 25.375 2.845 ;
      RECT 24.885 2.575 25.215 2.745 ;
      RECT 24.725 3.615 25.375 3.785 ;
      RECT 25.205 3.145 25.375 3.785 ;
      RECT 25.085 3.225 25.375 3.785 ;
      RECT 25.04 7.855 25.21 8.305 ;
      RECT 25.095 6.075 25.265 8.025 ;
      RECT 25.04 5.015 25.21 6.245 ;
      RECT 24.52 5.015 24.69 8.305 ;
      RECT 24.52 7.315 24.925 7.645 ;
      RECT 24.52 6.475 24.925 6.805 ;
      RECT 23.765 2.915 23.935 3.225 ;
      RECT 23.765 2.915 24.655 3.085 ;
      RECT 24.485 2.495 24.655 3.085 ;
      RECT 23.765 2.575 24.255 2.745 ;
      RECT 23.765 2.495 23.935 2.745 ;
      RECT 21.725 3.225 22.215 3.395 ;
      RECT 22.885 2.575 23.055 3.225 ;
      RECT 22.045 3.055 23.055 3.225 ;
      RECT 23.005 2.495 23.175 2.825 ;
      RECT 21.805 1.835 21.975 2.105 ;
      RECT 21.245 1.835 21.975 2.005 ;
      RECT 21.325 2.575 21.495 3.225 ;
      RECT 21.325 2.575 21.815 2.745 ;
      RECT 20.485 2.575 20.975 2.745 ;
      RECT 20.805 2.495 20.975 2.745 ;
      RECT 20.325 1.835 20.495 2.105 ;
      RECT 19.765 1.835 20.495 2.005 ;
      RECT 19.845 3.225 20.015 3.505 ;
      RECT 18.805 3.225 20.095 3.395 ;
      RECT 18.8 2.575 19.375 2.745 ;
      RECT 18.8 2.495 18.97 2.745 ;
      RECT 17.885 1.835 18.055 2.105 ;
      RECT 17.885 1.835 18.615 2.005 ;
      RECT 18.245 3.055 18.535 3.225 ;
      RECT 18.245 2.575 18.415 3.225 ;
      RECT 18.045 2.575 18.415 2.745 ;
      RECT 17.885 3.055 18.055 3.475 ;
      RECT 17.265 3.14 18.055 3.31 ;
      RECT 17.265 2.915 17.435 3.31 ;
      RECT 17.165 2.495 17.335 3.085 ;
      RECT 16.925 2.575 17.335 2.845 ;
      RECT 14.94 1.74 15.11 2.935 ;
      RECT 14.94 1.74 15.405 1.91 ;
      RECT 14.94 6.97 15.405 7.14 ;
      RECT 14.94 5.945 15.11 7.14 ;
      RECT 13.95 1.74 14.12 2.935 ;
      RECT 13.95 1.74 14.415 1.91 ;
      RECT 13.95 6.97 14.415 7.14 ;
      RECT 13.95 5.945 14.12 7.14 ;
      RECT 12.095 2.635 12.265 3.865 ;
      RECT 12.15 0.855 12.32 2.805 ;
      RECT 12.095 0.575 12.265 1.025 ;
      RECT 12.095 7.855 12.265 8.305 ;
      RECT 12.15 6.075 12.32 8.025 ;
      RECT 12.095 5.015 12.265 6.245 ;
      RECT 11.575 0.575 11.745 3.865 ;
      RECT 11.575 2.075 11.98 2.405 ;
      RECT 11.575 1.235 11.98 1.565 ;
      RECT 11.575 5.015 11.745 8.305 ;
      RECT 11.575 7.315 11.98 7.645 ;
      RECT 11.575 6.475 11.98 6.805 ;
      RECT 8.365 3.225 9.335 3.395 ;
      RECT 8.365 3.055 8.535 3.395 ;
      RECT 7.885 2.495 8.055 2.825 ;
      RECT 7.885 2.575 8.615 2.745 ;
      RECT 7.525 3.615 7.815 3.785 ;
      RECT 7.525 2.575 7.695 3.785 ;
      RECT 7.525 3.055 7.815 3.225 ;
      RECT 7.325 2.575 7.695 2.745 ;
      RECT 6.645 2.675 6.815 2.945 ;
      RECT 6.405 2.675 6.815 2.845 ;
      RECT 6.325 2.575 6.655 2.745 ;
      RECT 6.165 3.615 6.815 3.785 ;
      RECT 6.645 3.145 6.815 3.785 ;
      RECT 6.525 3.225 6.815 3.785 ;
      RECT 6.48 7.855 6.65 8.305 ;
      RECT 6.535 6.075 6.705 8.025 ;
      RECT 6.48 5.015 6.65 6.245 ;
      RECT 5.96 5.015 6.13 8.305 ;
      RECT 5.96 7.315 6.365 7.645 ;
      RECT 5.96 6.475 6.365 6.805 ;
      RECT 5.205 2.915 5.375 3.225 ;
      RECT 5.205 2.915 6.095 3.085 ;
      RECT 5.925 2.495 6.095 3.085 ;
      RECT 5.205 2.575 5.695 2.745 ;
      RECT 5.205 2.495 5.375 2.745 ;
      RECT 3.165 3.225 3.655 3.395 ;
      RECT 4.325 2.575 4.495 3.225 ;
      RECT 3.485 3.055 4.495 3.225 ;
      RECT 4.445 2.495 4.615 2.825 ;
      RECT 3.245 1.835 3.415 2.105 ;
      RECT 2.685 1.835 3.415 2.005 ;
      RECT 2.765 2.575 2.935 3.225 ;
      RECT 2.765 2.575 3.255 2.745 ;
      RECT 1.925 2.575 2.415 2.745 ;
      RECT 2.245 2.495 2.415 2.745 ;
      RECT 1.765 1.835 1.935 2.105 ;
      RECT 1.205 1.835 1.935 2.005 ;
      RECT 1.285 3.225 1.455 3.505 ;
      RECT 0.245 3.225 1.535 3.395 ;
      RECT 0.24 2.575 0.815 2.745 ;
      RECT 0.24 2.495 0.41 2.745 ;
      RECT -0.675 1.835 -0.505 2.105 ;
      RECT -0.675 1.835 0.055 2.005 ;
      RECT -0.315 3.055 -0.025 3.225 ;
      RECT -0.315 2.575 -0.145 3.225 ;
      RECT -0.515 2.575 -0.145 2.745 ;
      RECT -0.675 3.055 -0.505 3.475 ;
      RECT -1.295 3.14 -0.505 3.31 ;
      RECT -1.295 2.915 -1.125 3.31 ;
      RECT -1.395 2.495 -1.225 3.085 ;
      RECT -1.635 2.575 -1.225 2.845 ;
      RECT -4.335 7.855 -4.165 8.305 ;
      RECT -4.28 6.075 -4.11 8.025 ;
      RECT -4.335 5.015 -4.165 6.245 ;
      RECT -4.855 5.015 -4.685 8.305 ;
      RECT -4.855 7.315 -4.45 7.645 ;
      RECT -4.855 6.475 -4.45 6.805 ;
      RECT 89.55 0.575 89.72 1.085 ;
      RECT 89.55 2.395 89.72 3.865 ;
      RECT 89.55 5.015 89.72 6.485 ;
      RECT 89.55 7.795 89.72 8.305 ;
      RECT 88.56 0.575 88.73 1.085 ;
      RECT 88.56 2.395 88.73 3.865 ;
      RECT 88.56 5.015 88.73 6.485 ;
      RECT 88.56 7.795 88.73 8.305 ;
      RECT 87.195 0.575 87.365 3.865 ;
      RECT 87.195 5.015 87.365 8.305 ;
      RECT 86.765 0.575 86.935 1.085 ;
      RECT 86.765 1.655 86.935 3.865 ;
      RECT 86.765 5.015 86.935 7.225 ;
      RECT 86.765 7.795 86.935 8.305 ;
      RECT 85.395 1.66 85.565 2.935 ;
      RECT 85.395 5.945 85.565 7.22 ;
      RECT 83.085 2.495 83.255 2.945 ;
      RECT 82.845 1.755 83.015 2.105 ;
      RECT 81.885 1.755 82.055 2.105 ;
      RECT 81.58 5.015 81.75 8.305 ;
      RECT 81.405 3.055 81.575 3.475 ;
      RECT 81.15 5.015 81.32 7.225 ;
      RECT 81.15 7.795 81.32 8.305 ;
      RECT 80.405 1.755 80.575 2.105 ;
      RECT 79.78 5.945 79.95 7.22 ;
      RECT 79.445 1.755 79.615 2.105 ;
      RECT 79.445 3.485 79.615 3.815 ;
      RECT 78.925 3.145 79.095 3.785 ;
      RECT 78.445 1.755 78.615 2.105 ;
      RECT 78.205 2.495 78.375 2.825 ;
      RECT 77.725 2.495 77.895 2.825 ;
      RECT 76.485 3.145 76.655 3.505 ;
      RECT 76.005 3.055 76.175 3.475 ;
      RECT 75.765 2.495 75.935 2.825 ;
      RECT 75.285 2.495 75.455 2.945 ;
      RECT 73.325 2.495 73.495 2.825 ;
      RECT 72.605 1.755 72.775 2.105 ;
      RECT 72.605 3.285 72.775 3.645 ;
      RECT 70.99 0.575 71.16 1.085 ;
      RECT 70.99 2.395 71.16 3.865 ;
      RECT 70.99 5.015 71.16 6.485 ;
      RECT 70.99 7.795 71.16 8.305 ;
      RECT 70 0.575 70.17 1.085 ;
      RECT 70 2.395 70.17 3.865 ;
      RECT 70 5.015 70.17 6.485 ;
      RECT 70 7.795 70.17 8.305 ;
      RECT 68.635 0.575 68.805 3.865 ;
      RECT 68.635 5.015 68.805 8.305 ;
      RECT 68.205 0.575 68.375 1.085 ;
      RECT 68.205 1.655 68.375 3.865 ;
      RECT 68.205 5.015 68.375 7.225 ;
      RECT 68.205 7.795 68.375 8.305 ;
      RECT 66.835 1.66 67.005 2.935 ;
      RECT 66.835 5.945 67.005 7.22 ;
      RECT 64.525 2.495 64.695 2.945 ;
      RECT 64.285 1.755 64.455 2.105 ;
      RECT 63.325 1.755 63.495 2.105 ;
      RECT 63.02 5.015 63.19 8.305 ;
      RECT 62.845 3.055 63.015 3.475 ;
      RECT 62.59 5.015 62.76 7.225 ;
      RECT 62.59 7.795 62.76 8.305 ;
      RECT 61.845 1.755 62.015 2.105 ;
      RECT 61.22 5.945 61.39 7.22 ;
      RECT 60.885 1.755 61.055 2.105 ;
      RECT 60.885 3.485 61.055 3.815 ;
      RECT 60.365 3.145 60.535 3.785 ;
      RECT 59.885 1.755 60.055 2.105 ;
      RECT 59.645 2.495 59.815 2.825 ;
      RECT 59.165 2.495 59.335 2.825 ;
      RECT 57.925 3.145 58.095 3.505 ;
      RECT 57.445 3.055 57.615 3.475 ;
      RECT 57.205 2.495 57.375 2.825 ;
      RECT 56.725 2.495 56.895 2.945 ;
      RECT 54.765 2.495 54.935 2.825 ;
      RECT 54.045 1.755 54.215 2.105 ;
      RECT 54.045 3.285 54.215 3.645 ;
      RECT 52.43 0.575 52.6 1.085 ;
      RECT 52.43 2.395 52.6 3.865 ;
      RECT 52.43 5.015 52.6 6.485 ;
      RECT 52.43 7.795 52.6 8.305 ;
      RECT 51.44 0.575 51.61 1.085 ;
      RECT 51.44 2.395 51.61 3.865 ;
      RECT 51.44 5.015 51.61 6.485 ;
      RECT 51.44 7.795 51.61 8.305 ;
      RECT 50.075 0.575 50.245 3.865 ;
      RECT 50.075 5.015 50.245 8.305 ;
      RECT 49.645 0.575 49.815 1.085 ;
      RECT 49.645 1.655 49.815 3.865 ;
      RECT 49.645 5.015 49.815 7.225 ;
      RECT 49.645 7.795 49.815 8.305 ;
      RECT 48.275 1.66 48.445 2.935 ;
      RECT 48.275 5.945 48.445 7.22 ;
      RECT 45.965 2.495 46.135 2.945 ;
      RECT 45.725 1.755 45.895 2.105 ;
      RECT 44.765 1.755 44.935 2.105 ;
      RECT 44.46 5.015 44.63 8.305 ;
      RECT 44.285 3.055 44.455 3.475 ;
      RECT 44.03 5.015 44.2 7.225 ;
      RECT 44.03 7.795 44.2 8.305 ;
      RECT 43.285 1.755 43.455 2.105 ;
      RECT 42.66 5.945 42.83 7.22 ;
      RECT 42.325 1.755 42.495 2.105 ;
      RECT 42.325 3.485 42.495 3.815 ;
      RECT 41.805 3.145 41.975 3.785 ;
      RECT 41.325 1.755 41.495 2.105 ;
      RECT 41.085 2.495 41.255 2.825 ;
      RECT 40.605 2.495 40.775 2.825 ;
      RECT 39.365 3.145 39.535 3.505 ;
      RECT 38.885 3.055 39.055 3.475 ;
      RECT 38.645 2.495 38.815 2.825 ;
      RECT 38.165 2.495 38.335 2.945 ;
      RECT 36.205 2.495 36.375 2.825 ;
      RECT 35.485 1.755 35.655 2.105 ;
      RECT 35.485 3.285 35.655 3.645 ;
      RECT 33.87 0.575 34.04 1.085 ;
      RECT 33.87 2.395 34.04 3.865 ;
      RECT 33.87 5.015 34.04 6.485 ;
      RECT 33.87 7.795 34.04 8.305 ;
      RECT 32.88 0.575 33.05 1.085 ;
      RECT 32.88 2.395 33.05 3.865 ;
      RECT 32.88 5.015 33.05 6.485 ;
      RECT 32.88 7.795 33.05 8.305 ;
      RECT 31.515 0.575 31.685 3.865 ;
      RECT 31.515 5.015 31.685 8.305 ;
      RECT 31.085 0.575 31.255 1.085 ;
      RECT 31.085 1.655 31.255 3.865 ;
      RECT 31.085 5.015 31.255 7.225 ;
      RECT 31.085 7.795 31.255 8.305 ;
      RECT 29.715 1.66 29.885 2.935 ;
      RECT 29.715 5.945 29.885 7.22 ;
      RECT 27.405 2.495 27.575 2.945 ;
      RECT 27.165 1.755 27.335 2.105 ;
      RECT 26.205 1.755 26.375 2.105 ;
      RECT 25.9 5.015 26.07 8.305 ;
      RECT 25.725 3.055 25.895 3.475 ;
      RECT 25.47 5.015 25.64 7.225 ;
      RECT 25.47 7.795 25.64 8.305 ;
      RECT 24.725 1.755 24.895 2.105 ;
      RECT 24.1 5.945 24.27 7.22 ;
      RECT 23.765 1.755 23.935 2.105 ;
      RECT 23.765 3.485 23.935 3.815 ;
      RECT 23.245 3.145 23.415 3.785 ;
      RECT 22.765 1.755 22.935 2.105 ;
      RECT 22.525 2.495 22.695 2.825 ;
      RECT 22.045 2.495 22.215 2.825 ;
      RECT 20.805 3.145 20.975 3.505 ;
      RECT 20.325 3.055 20.495 3.475 ;
      RECT 20.085 2.495 20.255 2.825 ;
      RECT 19.605 2.495 19.775 2.945 ;
      RECT 17.645 2.495 17.815 2.825 ;
      RECT 16.925 1.755 17.095 2.105 ;
      RECT 16.925 3.285 17.095 3.645 ;
      RECT 15.31 0.575 15.48 1.085 ;
      RECT 15.31 2.395 15.48 3.865 ;
      RECT 15.31 5.015 15.48 6.485 ;
      RECT 15.31 7.795 15.48 8.305 ;
      RECT 14.32 0.575 14.49 1.085 ;
      RECT 14.32 2.395 14.49 3.865 ;
      RECT 14.32 5.015 14.49 6.485 ;
      RECT 14.32 7.795 14.49 8.305 ;
      RECT 12.955 0.575 13.125 3.865 ;
      RECT 12.955 5.015 13.125 8.305 ;
      RECT 12.525 0.575 12.695 1.085 ;
      RECT 12.525 1.655 12.695 3.865 ;
      RECT 12.525 5.015 12.695 7.225 ;
      RECT 12.525 7.795 12.695 8.305 ;
      RECT 11.155 1.66 11.325 2.935 ;
      RECT 11.155 5.945 11.325 7.22 ;
      RECT 8.845 2.495 9.015 2.945 ;
      RECT 8.605 1.755 8.775 2.105 ;
      RECT 7.645 1.755 7.815 2.105 ;
      RECT 7.34 5.015 7.51 8.305 ;
      RECT 7.165 3.055 7.335 3.475 ;
      RECT 6.91 5.015 7.08 7.225 ;
      RECT 6.91 7.795 7.08 8.305 ;
      RECT 6.165 1.755 6.335 2.105 ;
      RECT 5.54 5.945 5.71 7.22 ;
      RECT 5.205 1.755 5.375 2.105 ;
      RECT 5.205 3.485 5.375 3.815 ;
      RECT 4.685 3.145 4.855 3.785 ;
      RECT 4.205 1.755 4.375 2.105 ;
      RECT 3.965 2.495 4.135 2.825 ;
      RECT 3.485 2.495 3.655 2.825 ;
      RECT 2.245 3.145 2.415 3.505 ;
      RECT 1.765 3.055 1.935 3.475 ;
      RECT 1.525 2.495 1.695 2.825 ;
      RECT 1.045 2.495 1.215 2.945 ;
      RECT -0.915 2.495 -0.745 2.825 ;
      RECT -1.635 1.755 -1.465 2.105 ;
      RECT -1.635 3.285 -1.465 3.645 ;
      RECT -3.905 5.015 -3.735 7.225 ;
      RECT -3.905 7.795 -3.735 8.305 ;
      RECT -5.275 5.945 -5.105 7.22 ;
  END
END sky130_osu_ring_oscillator_mpr2et_8_b0r2

MACRO sky130_osu_ring_oscillator_mpr2xa_8_b0r1
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 2.8 -0.005 ;
  SIZE 79.1 BY 8.88 ;
  SYMMETRY X Y R90 ;
  SITE CoreSite ;
  OBS
    LAYER met4 ;
      RECT 63.94 2.98 64.27 3.31 ;
      RECT 63.955 2.505 64.27 3.31 ;
      RECT 66.1 2.49 66.43 2.845 ;
      RECT 63.955 2.505 66.43 2.805 ;
      RECT 48.68 2.98 49.01 3.31 ;
      RECT 48.695 2.505 49.01 3.31 ;
      RECT 50.84 2.49 51.17 2.845 ;
      RECT 48.695 2.505 51.17 2.805 ;
      RECT 33.42 2.98 33.75 3.31 ;
      RECT 33.435 2.505 33.75 3.31 ;
      RECT 35.58 2.49 35.91 2.845 ;
      RECT 33.435 2.505 35.91 2.805 ;
      RECT 18.16 2.98 18.49 3.31 ;
      RECT 18.175 2.505 18.49 3.31 ;
      RECT 20.32 2.49 20.65 2.845 ;
      RECT 18.175 2.505 20.65 2.805 ;
      RECT 2.9 2.98 3.23 3.31 ;
      RECT 2.915 2.505 3.23 3.31 ;
      RECT 5.06 2.49 5.39 2.845 ;
      RECT 2.915 2.505 5.39 2.805 ;
    LAYER via3 ;
      RECT 66.165 2.58 66.365 2.78 ;
      RECT 64.005 3.045 64.205 3.245 ;
      RECT 50.905 2.58 51.105 2.78 ;
      RECT 48.745 3.045 48.945 3.245 ;
      RECT 35.645 2.58 35.845 2.78 ;
      RECT 33.485 3.045 33.685 3.245 ;
      RECT 20.385 2.58 20.585 2.78 ;
      RECT 18.225 3.045 18.425 3.245 ;
      RECT 5.125 2.58 5.325 2.78 ;
      RECT 2.965 3.045 3.165 3.245 ;
    LAYER met3 ;
      RECT 67.26 7.06 67.63 7.43 ;
      RECT 67.295 4.48 67.595 7.43 ;
      RECT 65.855 4.48 67.595 4.78 ;
      RECT 63.06 4.26 66.155 4.56 ;
      RECT 65.855 2.52 66.155 4.78 ;
      RECT 63.06 2.98 63.36 4.56 ;
      RECT 66.58 3.515 66.91 3.87 ;
      RECT 64.675 3.555 66.91 3.855 ;
      RECT 64.675 2.42 64.975 3.855 ;
      RECT 62.755 2.98 63.485 3.31 ;
      RECT 65.65 2.525 66.43 2.87 ;
      RECT 66.125 2.49 66.43 2.87 ;
      RECT 64.66 2.42 64.99 2.75 ;
      RECT 63.945 2.42 64.265 3.335 ;
      RECT 63.945 2.42 64.275 2.955 ;
      RECT 52 7.06 52.37 7.43 ;
      RECT 52.035 4.48 52.335 7.43 ;
      RECT 50.595 4.48 52.335 4.78 ;
      RECT 47.8 4.26 50.895 4.56 ;
      RECT 50.595 2.52 50.895 4.78 ;
      RECT 47.8 2.98 48.1 4.56 ;
      RECT 51.32 3.515 51.65 3.87 ;
      RECT 49.415 3.555 51.65 3.855 ;
      RECT 49.415 2.42 49.715 3.855 ;
      RECT 47.495 2.98 48.225 3.31 ;
      RECT 50.39 2.525 51.17 2.87 ;
      RECT 50.865 2.49 51.17 2.87 ;
      RECT 49.4 2.42 49.73 2.75 ;
      RECT 48.685 2.42 49.005 3.335 ;
      RECT 48.685 2.42 49.015 2.955 ;
      RECT 36.74 7.06 37.11 7.43 ;
      RECT 36.775 4.48 37.075 7.43 ;
      RECT 35.335 4.48 37.075 4.78 ;
      RECT 32.54 4.26 35.635 4.56 ;
      RECT 35.335 2.52 35.635 4.78 ;
      RECT 32.54 2.98 32.84 4.56 ;
      RECT 36.06 3.515 36.39 3.87 ;
      RECT 34.155 3.555 36.39 3.855 ;
      RECT 34.155 2.42 34.455 3.855 ;
      RECT 32.235 2.98 32.965 3.31 ;
      RECT 35.13 2.525 35.91 2.87 ;
      RECT 35.605 2.49 35.91 2.87 ;
      RECT 34.14 2.42 34.47 2.75 ;
      RECT 33.425 2.42 33.745 3.335 ;
      RECT 33.425 2.42 33.755 2.955 ;
      RECT 21.48 7.06 21.85 7.43 ;
      RECT 21.515 4.48 21.815 7.43 ;
      RECT 20.075 4.48 21.815 4.78 ;
      RECT 17.28 4.26 20.375 4.56 ;
      RECT 20.075 2.52 20.375 4.78 ;
      RECT 17.28 2.98 17.58 4.56 ;
      RECT 20.8 3.515 21.13 3.87 ;
      RECT 18.895 3.555 21.13 3.855 ;
      RECT 18.895 2.42 19.195 3.855 ;
      RECT 16.975 2.98 17.705 3.31 ;
      RECT 19.87 2.525 20.65 2.87 ;
      RECT 20.345 2.49 20.65 2.87 ;
      RECT 18.88 2.42 19.21 2.75 ;
      RECT 18.165 2.42 18.485 3.335 ;
      RECT 18.165 2.42 18.495 2.955 ;
      RECT 6.22 7.06 6.59 7.43 ;
      RECT 6.255 4.48 6.555 7.43 ;
      RECT 4.815 4.48 6.555 4.78 ;
      RECT 2.02 4.26 5.115 4.56 ;
      RECT 4.815 2.52 5.115 4.78 ;
      RECT 2.02 2.98 2.32 4.56 ;
      RECT 5.54 3.515 5.87 3.87 ;
      RECT 3.635 3.555 5.87 3.855 ;
      RECT 3.635 2.42 3.935 3.855 ;
      RECT 1.715 2.98 2.445 3.31 ;
      RECT 4.61 2.525 5.39 2.87 ;
      RECT 5.085 2.49 5.39 2.87 ;
      RECT 3.62 2.42 3.95 2.75 ;
      RECT 2.905 2.42 3.225 3.335 ;
      RECT 2.905 2.42 3.235 2.955 ;
      RECT 69.5 1.86 70.23 2.19 ;
      RECT 67.81 1.875 68.54 2.205 ;
      RECT 66.775 1.86 67.505 2.21 ;
      RECT 65.225 1.885 65.955 2.215 ;
      RECT 62.62 1.86 63.35 2.19 ;
      RECT 54.24 1.86 54.97 2.19 ;
      RECT 52.55 1.875 53.28 2.205 ;
      RECT 51.515 1.86 52.245 2.21 ;
      RECT 49.965 1.885 50.695 2.215 ;
      RECT 47.36 1.86 48.09 2.19 ;
      RECT 38.98 1.86 39.71 2.19 ;
      RECT 37.29 1.875 38.02 2.205 ;
      RECT 36.255 1.86 36.985 2.21 ;
      RECT 34.705 1.885 35.435 2.215 ;
      RECT 32.1 1.86 32.83 2.19 ;
      RECT 23.72 1.86 24.45 2.19 ;
      RECT 22.03 1.875 22.76 2.205 ;
      RECT 20.995 1.86 21.725 2.21 ;
      RECT 19.445 1.885 20.175 2.215 ;
      RECT 16.84 1.86 17.57 2.19 ;
      RECT 8.46 1.86 9.19 2.19 ;
      RECT 6.77 1.875 7.5 2.205 ;
      RECT 5.735 1.86 6.465 2.21 ;
      RECT 4.185 1.885 4.915 2.215 ;
      RECT 1.58 1.86 2.31 2.19 ;
    LAYER via2 ;
      RECT 69.735 1.925 69.935 2.125 ;
      RECT 67.875 1.94 68.075 2.14 ;
      RECT 67.345 7.145 67.545 7.345 ;
      RECT 66.855 1.945 67.055 2.145 ;
      RECT 66.645 3.58 66.845 3.78 ;
      RECT 66.165 2.58 66.365 2.78 ;
      RECT 65.415 1.95 65.615 2.15 ;
      RECT 64.725 2.485 64.925 2.685 ;
      RECT 64.01 2.485 64.21 2.685 ;
      RECT 63.045 3.045 63.245 3.245 ;
      RECT 62.805 1.925 63.005 2.125 ;
      RECT 54.475 1.925 54.675 2.125 ;
      RECT 52.615 1.94 52.815 2.14 ;
      RECT 52.085 7.145 52.285 7.345 ;
      RECT 51.595 1.945 51.795 2.145 ;
      RECT 51.385 3.58 51.585 3.78 ;
      RECT 50.905 2.58 51.105 2.78 ;
      RECT 50.155 1.95 50.355 2.15 ;
      RECT 49.465 2.485 49.665 2.685 ;
      RECT 48.75 2.485 48.95 2.685 ;
      RECT 47.785 3.045 47.985 3.245 ;
      RECT 47.545 1.925 47.745 2.125 ;
      RECT 39.215 1.925 39.415 2.125 ;
      RECT 37.355 1.94 37.555 2.14 ;
      RECT 36.825 7.145 37.025 7.345 ;
      RECT 36.335 1.945 36.535 2.145 ;
      RECT 36.125 3.58 36.325 3.78 ;
      RECT 35.645 2.58 35.845 2.78 ;
      RECT 34.895 1.95 35.095 2.15 ;
      RECT 34.205 2.485 34.405 2.685 ;
      RECT 33.49 2.485 33.69 2.685 ;
      RECT 32.525 3.045 32.725 3.245 ;
      RECT 32.285 1.925 32.485 2.125 ;
      RECT 23.955 1.925 24.155 2.125 ;
      RECT 22.095 1.94 22.295 2.14 ;
      RECT 21.565 7.145 21.765 7.345 ;
      RECT 21.075 1.945 21.275 2.145 ;
      RECT 20.865 3.58 21.065 3.78 ;
      RECT 20.385 2.58 20.585 2.78 ;
      RECT 19.635 1.95 19.835 2.15 ;
      RECT 18.945 2.485 19.145 2.685 ;
      RECT 18.23 2.485 18.43 2.685 ;
      RECT 17.265 3.045 17.465 3.245 ;
      RECT 17.025 1.925 17.225 2.125 ;
      RECT 8.695 1.925 8.895 2.125 ;
      RECT 6.835 1.94 7.035 2.14 ;
      RECT 6.305 7.145 6.505 7.345 ;
      RECT 5.815 1.945 6.015 2.145 ;
      RECT 5.605 3.58 5.805 3.78 ;
      RECT 5.125 2.58 5.325 2.78 ;
      RECT 4.375 1.95 4.575 2.15 ;
      RECT 3.685 2.485 3.885 2.685 ;
      RECT 2.97 2.485 3.17 2.685 ;
      RECT 2.005 3.045 2.205 3.245 ;
      RECT 1.765 1.925 1.965 2.125 ;
    LAYER met2 ;
      RECT -1.57 8.405 75.93 8.575 ;
      RECT 75.76 7.28 75.93 8.575 ;
      RECT -1.57 6.26 -1.4 8.575 ;
      RECT 75.73 7.28 76.08 7.63 ;
      RECT -1.63 6.26 -1.34 6.61 ;
      RECT 72.57 6.225 72.89 6.55 ;
      RECT 72.6 5.7 72.77 6.55 ;
      RECT 72.6 5.7 72.775 6.05 ;
      RECT 72.6 5.7 73.575 5.875 ;
      RECT 73.4 1.97 73.575 5.875 ;
      RECT 73.345 1.97 73.695 2.32 ;
      RECT 73.37 6.66 73.695 6.985 ;
      RECT 72.255 6.75 73.695 6.92 ;
      RECT 72.255 2.4 72.415 6.92 ;
      RECT 72.57 2.37 72.89 2.69 ;
      RECT 72.255 2.4 72.89 2.57 ;
      RECT 71.525 5.865 71.865 6.215 ;
      RECT 71.605 2.71 71.775 6.215 ;
      RECT 71.525 2.71 71.865 3.06 ;
      RECT 69.705 3.545 69.965 3.865 ;
      RECT 69.765 1.84 69.905 3.865 ;
      RECT 70.965 2.705 71.305 3.055 ;
      RECT 70.34 2.775 71.305 2.975 ;
      RECT 70.34 1.945 70.54 2.975 ;
      RECT 69.59 2.4 69.905 2.77 ;
      RECT 71.055 2.7 71.225 3.055 ;
      RECT 69.66 1.955 69.905 2.77 ;
      RECT 69.695 1.84 69.975 2.21 ;
      RECT 69.695 1.945 70.54 2.145 ;
      RECT 69.015 2.425 69.275 2.745 ;
      RECT 68.355 2.515 69.275 2.655 ;
      RECT 68.355 1.575 68.495 2.655 ;
      RECT 64.815 1.865 65.075 2.185 ;
      RECT 64.995 1.575 65.135 2.095 ;
      RECT 64.995 1.575 68.495 1.715 ;
      RECT 60.445 6.66 60.795 7.01 ;
      RECT 67.93 6.615 68.28 6.965 ;
      RECT 60.445 6.69 68.28 6.89 ;
      RECT 67.845 3.265 68.105 3.585 ;
      RECT 67.905 1.855 68.045 3.585 ;
      RECT 67.835 1.855 68.115 2.225 ;
      RECT 65.235 4.015 67.67 4.155 ;
      RECT 67.53 2.705 67.67 4.155 ;
      RECT 65.235 3.635 65.375 4.155 ;
      RECT 64.935 3.635 65.375 3.865 ;
      RECT 62.595 3.635 65.375 3.775 ;
      RECT 64.935 3.545 65.195 3.865 ;
      RECT 62.595 3.355 62.735 3.775 ;
      RECT 62.085 3.265 62.345 3.585 ;
      RECT 62.085 3.355 62.735 3.495 ;
      RECT 62.145 1.865 62.285 3.585 ;
      RECT 67.47 2.705 67.73 3.025 ;
      RECT 62.085 1.865 62.345 2.185 ;
      RECT 67.095 3.545 67.355 3.865 ;
      RECT 67.155 1.955 67.295 3.865 ;
      RECT 66.815 1.955 67.295 2.23 ;
      RECT 66.615 1.86 67.095 2.205 ;
      RECT 66.605 3.495 66.885 3.865 ;
      RECT 66.675 2.4 66.815 3.865 ;
      RECT 66.615 2.4 66.875 3.025 ;
      RECT 66.605 2.4 66.885 2.77 ;
      RECT 65.535 3.545 65.795 3.865 ;
      RECT 65.535 3.355 65.735 3.865 ;
      RECT 65.34 3.355 65.735 3.495 ;
      RECT 65.34 1.865 65.48 3.495 ;
      RECT 65.34 1.865 65.655 2.235 ;
      RECT 65.28 1.865 65.655 2.185 ;
      RECT 63.005 2.96 63.285 3.33 ;
      RECT 64.455 2.985 64.715 3.305 ;
      RECT 62.835 3.075 64.715 3.215 ;
      RECT 62.835 2.96 63.285 3.215 ;
      RECT 62.775 2.4 63.035 3.025 ;
      RECT 62.765 2.4 63.045 2.77 ;
      RECT 63.845 2.4 64.255 2.77 ;
      RECT 63.255 2.425 63.515 2.745 ;
      RECT 63.255 2.515 64.255 2.655 ;
      RECT 62.765 1.84 63.045 2.21 ;
      RECT 62.765 1.865 63.155 2.185 ;
      RECT 57.31 6.225 57.63 6.55 ;
      RECT 57.34 5.7 57.51 6.55 ;
      RECT 57.34 5.7 57.515 6.05 ;
      RECT 57.34 5.7 58.315 5.875 ;
      RECT 58.14 1.97 58.315 5.875 ;
      RECT 58.085 1.97 58.435 2.32 ;
      RECT 58.11 6.66 58.435 6.985 ;
      RECT 56.995 6.75 58.435 6.92 ;
      RECT 56.995 2.4 57.155 6.92 ;
      RECT 57.31 2.37 57.63 2.69 ;
      RECT 56.995 2.4 57.63 2.57 ;
      RECT 56.265 5.865 56.605 6.215 ;
      RECT 56.345 2.71 56.515 6.215 ;
      RECT 56.265 2.71 56.605 3.06 ;
      RECT 54.445 3.545 54.705 3.865 ;
      RECT 54.505 1.84 54.645 3.865 ;
      RECT 55.705 2.705 56.045 3.055 ;
      RECT 55.08 2.775 56.045 2.975 ;
      RECT 55.08 1.945 55.28 2.975 ;
      RECT 54.33 2.4 54.645 2.77 ;
      RECT 55.795 2.7 55.965 3.055 ;
      RECT 54.4 1.955 54.645 2.77 ;
      RECT 54.435 1.84 54.715 2.21 ;
      RECT 54.435 1.945 55.28 2.145 ;
      RECT 53.755 2.425 54.015 2.745 ;
      RECT 53.095 2.515 54.015 2.655 ;
      RECT 53.095 1.575 53.235 2.655 ;
      RECT 49.555 1.865 49.815 2.185 ;
      RECT 49.735 1.575 49.875 2.095 ;
      RECT 49.735 1.575 53.235 1.715 ;
      RECT 45.185 6.66 45.535 7.01 ;
      RECT 52.675 6.615 53.025 6.965 ;
      RECT 45.185 6.69 53.025 6.89 ;
      RECT 52.585 3.265 52.845 3.585 ;
      RECT 52.645 1.855 52.785 3.585 ;
      RECT 52.575 1.855 52.855 2.225 ;
      RECT 49.975 4.015 52.41 4.155 ;
      RECT 52.27 2.705 52.41 4.155 ;
      RECT 49.975 3.635 50.115 4.155 ;
      RECT 49.675 3.635 50.115 3.865 ;
      RECT 47.335 3.635 50.115 3.775 ;
      RECT 49.675 3.545 49.935 3.865 ;
      RECT 47.335 3.355 47.475 3.775 ;
      RECT 46.825 3.265 47.085 3.585 ;
      RECT 46.825 3.355 47.475 3.495 ;
      RECT 46.885 1.865 47.025 3.585 ;
      RECT 52.21 2.705 52.47 3.025 ;
      RECT 46.825 1.865 47.085 2.185 ;
      RECT 51.835 3.545 52.095 3.865 ;
      RECT 51.895 1.955 52.035 3.865 ;
      RECT 51.555 1.955 52.035 2.23 ;
      RECT 51.355 1.86 51.835 2.205 ;
      RECT 51.345 3.495 51.625 3.865 ;
      RECT 51.415 2.4 51.555 3.865 ;
      RECT 51.355 2.4 51.615 3.025 ;
      RECT 51.345 2.4 51.625 2.77 ;
      RECT 50.275 3.545 50.535 3.865 ;
      RECT 50.275 3.355 50.475 3.865 ;
      RECT 50.08 3.355 50.475 3.495 ;
      RECT 50.08 1.865 50.22 3.495 ;
      RECT 50.08 1.865 50.395 2.235 ;
      RECT 50.02 1.865 50.395 2.185 ;
      RECT 47.745 2.96 48.025 3.33 ;
      RECT 49.195 2.985 49.455 3.305 ;
      RECT 47.575 3.075 49.455 3.215 ;
      RECT 47.575 2.96 48.025 3.215 ;
      RECT 47.515 2.4 47.775 3.025 ;
      RECT 47.505 2.4 47.785 2.77 ;
      RECT 48.585 2.4 48.995 2.77 ;
      RECT 47.995 2.425 48.255 2.745 ;
      RECT 47.995 2.515 48.995 2.655 ;
      RECT 47.505 1.84 47.785 2.21 ;
      RECT 47.505 1.865 47.895 2.185 ;
      RECT 42.05 6.225 42.37 6.55 ;
      RECT 42.08 5.7 42.25 6.55 ;
      RECT 42.08 5.7 42.255 6.05 ;
      RECT 42.08 5.7 43.055 5.875 ;
      RECT 42.88 1.97 43.055 5.875 ;
      RECT 42.825 1.97 43.175 2.32 ;
      RECT 42.85 6.66 43.175 6.985 ;
      RECT 41.735 6.75 43.175 6.92 ;
      RECT 41.735 2.4 41.895 6.92 ;
      RECT 42.05 2.37 42.37 2.69 ;
      RECT 41.735 2.4 42.37 2.57 ;
      RECT 41.005 5.865 41.345 6.215 ;
      RECT 41.085 2.71 41.255 6.215 ;
      RECT 41.005 2.71 41.345 3.06 ;
      RECT 39.185 3.545 39.445 3.865 ;
      RECT 39.245 1.84 39.385 3.865 ;
      RECT 40.445 2.705 40.785 3.055 ;
      RECT 39.82 2.775 40.785 2.975 ;
      RECT 39.82 1.945 40.02 2.975 ;
      RECT 39.07 2.4 39.385 2.77 ;
      RECT 40.535 2.7 40.705 3.055 ;
      RECT 39.14 1.955 39.385 2.77 ;
      RECT 39.175 1.84 39.455 2.21 ;
      RECT 39.175 1.945 40.02 2.145 ;
      RECT 38.495 2.425 38.755 2.745 ;
      RECT 37.835 2.515 38.755 2.655 ;
      RECT 37.835 1.575 37.975 2.655 ;
      RECT 34.295 1.865 34.555 2.185 ;
      RECT 34.475 1.575 34.615 2.095 ;
      RECT 34.475 1.575 37.975 1.715 ;
      RECT 29.97 6.665 30.32 7.015 ;
      RECT 37.41 6.62 37.76 6.97 ;
      RECT 29.97 6.695 37.76 6.895 ;
      RECT 37.325 3.265 37.585 3.585 ;
      RECT 37.385 1.855 37.525 3.585 ;
      RECT 37.315 1.855 37.595 2.225 ;
      RECT 34.715 4.015 37.15 4.155 ;
      RECT 37.01 2.705 37.15 4.155 ;
      RECT 34.715 3.635 34.855 4.155 ;
      RECT 34.415 3.635 34.855 3.865 ;
      RECT 32.075 3.635 34.855 3.775 ;
      RECT 34.415 3.545 34.675 3.865 ;
      RECT 32.075 3.355 32.215 3.775 ;
      RECT 31.565 3.265 31.825 3.585 ;
      RECT 31.565 3.355 32.215 3.495 ;
      RECT 31.625 1.865 31.765 3.585 ;
      RECT 36.95 2.705 37.21 3.025 ;
      RECT 31.565 1.865 31.825 2.185 ;
      RECT 36.575 3.545 36.835 3.865 ;
      RECT 36.635 1.955 36.775 3.865 ;
      RECT 36.295 1.955 36.775 2.23 ;
      RECT 36.095 1.86 36.575 2.205 ;
      RECT 36.085 3.495 36.365 3.865 ;
      RECT 36.155 2.4 36.295 3.865 ;
      RECT 36.095 2.4 36.355 3.025 ;
      RECT 36.085 2.4 36.365 2.77 ;
      RECT 35.015 3.545 35.275 3.865 ;
      RECT 35.015 3.355 35.215 3.865 ;
      RECT 34.82 3.355 35.215 3.495 ;
      RECT 34.82 1.865 34.96 3.495 ;
      RECT 34.82 1.865 35.135 2.235 ;
      RECT 34.76 1.865 35.135 2.185 ;
      RECT 32.485 2.96 32.765 3.33 ;
      RECT 33.935 2.985 34.195 3.305 ;
      RECT 32.315 3.075 34.195 3.215 ;
      RECT 32.315 2.96 32.765 3.215 ;
      RECT 32.255 2.4 32.515 3.025 ;
      RECT 32.245 2.4 32.525 2.77 ;
      RECT 33.325 2.4 33.735 2.77 ;
      RECT 32.735 2.425 32.995 2.745 ;
      RECT 32.735 2.515 33.735 2.655 ;
      RECT 32.245 1.84 32.525 2.21 ;
      RECT 32.245 1.865 32.635 2.185 ;
      RECT 26.79 6.225 27.11 6.55 ;
      RECT 26.82 5.7 26.99 6.55 ;
      RECT 26.82 5.7 26.995 6.05 ;
      RECT 26.82 5.7 27.795 5.875 ;
      RECT 27.62 1.97 27.795 5.875 ;
      RECT 27.565 1.97 27.915 2.32 ;
      RECT 27.59 6.66 27.915 6.985 ;
      RECT 26.475 6.75 27.915 6.92 ;
      RECT 26.475 2.4 26.635 6.92 ;
      RECT 26.79 2.37 27.11 2.69 ;
      RECT 26.475 2.4 27.11 2.57 ;
      RECT 25.745 5.865 26.085 6.215 ;
      RECT 25.825 2.71 25.995 6.215 ;
      RECT 25.745 2.71 26.085 3.06 ;
      RECT 23.925 3.545 24.185 3.865 ;
      RECT 23.985 1.84 24.125 3.865 ;
      RECT 25.185 2.705 25.525 3.055 ;
      RECT 24.56 2.775 25.525 2.975 ;
      RECT 24.56 1.945 24.76 2.975 ;
      RECT 23.81 2.4 24.125 2.77 ;
      RECT 25.275 2.7 25.445 3.055 ;
      RECT 23.88 1.955 24.125 2.77 ;
      RECT 23.915 1.84 24.195 2.21 ;
      RECT 23.915 1.945 24.76 2.145 ;
      RECT 23.235 2.425 23.495 2.745 ;
      RECT 22.575 2.515 23.495 2.655 ;
      RECT 22.575 1.575 22.715 2.655 ;
      RECT 19.035 1.865 19.295 2.185 ;
      RECT 19.215 1.575 19.355 2.095 ;
      RECT 19.215 1.575 22.715 1.715 ;
      RECT 14.71 6.66 15.06 7.01 ;
      RECT 22.15 6.615 22.5 6.965 ;
      RECT 14.71 6.69 22.5 6.89 ;
      RECT 22.065 3.265 22.325 3.585 ;
      RECT 22.125 1.855 22.265 3.585 ;
      RECT 22.055 1.855 22.335 2.225 ;
      RECT 19.455 4.015 21.89 4.155 ;
      RECT 21.75 2.705 21.89 4.155 ;
      RECT 19.455 3.635 19.595 4.155 ;
      RECT 19.155 3.635 19.595 3.865 ;
      RECT 16.815 3.635 19.595 3.775 ;
      RECT 19.155 3.545 19.415 3.865 ;
      RECT 16.815 3.355 16.955 3.775 ;
      RECT 16.305 3.265 16.565 3.585 ;
      RECT 16.305 3.355 16.955 3.495 ;
      RECT 16.365 1.865 16.505 3.585 ;
      RECT 21.69 2.705 21.95 3.025 ;
      RECT 16.305 1.865 16.565 2.185 ;
      RECT 21.315 3.545 21.575 3.865 ;
      RECT 21.375 1.955 21.515 3.865 ;
      RECT 21.035 1.955 21.515 2.23 ;
      RECT 20.835 1.86 21.315 2.205 ;
      RECT 20.825 3.495 21.105 3.865 ;
      RECT 20.895 2.4 21.035 3.865 ;
      RECT 20.835 2.4 21.095 3.025 ;
      RECT 20.825 2.4 21.105 2.77 ;
      RECT 19.755 3.545 20.015 3.865 ;
      RECT 19.755 3.355 19.955 3.865 ;
      RECT 19.56 3.355 19.955 3.495 ;
      RECT 19.56 1.865 19.7 3.495 ;
      RECT 19.56 1.865 19.875 2.235 ;
      RECT 19.5 1.865 19.875 2.185 ;
      RECT 17.225 2.96 17.505 3.33 ;
      RECT 18.675 2.985 18.935 3.305 ;
      RECT 17.055 3.075 18.935 3.215 ;
      RECT 17.055 2.96 17.505 3.215 ;
      RECT 16.995 2.4 17.255 3.025 ;
      RECT 16.985 2.4 17.265 2.77 ;
      RECT 18.065 2.4 18.475 2.77 ;
      RECT 17.475 2.425 17.735 2.745 ;
      RECT 17.475 2.515 18.475 2.655 ;
      RECT 16.985 1.84 17.265 2.21 ;
      RECT 16.985 1.865 17.375 2.185 ;
      RECT 11.53 6.225 11.85 6.55 ;
      RECT 11.56 5.7 11.73 6.55 ;
      RECT 11.56 5.7 11.735 6.05 ;
      RECT 11.56 5.7 12.535 5.875 ;
      RECT 12.36 1.97 12.535 5.875 ;
      RECT 12.305 1.97 12.655 2.32 ;
      RECT 12.33 6.66 12.655 6.985 ;
      RECT 11.215 6.75 12.655 6.92 ;
      RECT 11.215 2.4 11.375 6.92 ;
      RECT 11.53 2.37 11.85 2.69 ;
      RECT 11.215 2.4 11.85 2.57 ;
      RECT 10.485 5.865 10.825 6.215 ;
      RECT 10.565 2.71 10.735 6.215 ;
      RECT 10.485 2.71 10.825 3.06 ;
      RECT 8.665 3.545 8.925 3.865 ;
      RECT 8.725 1.84 8.865 3.865 ;
      RECT 9.925 2.705 10.265 3.055 ;
      RECT 9.3 2.775 10.265 2.975 ;
      RECT 9.3 1.945 9.5 2.975 ;
      RECT 8.55 2.4 8.865 2.77 ;
      RECT 10.015 2.7 10.185 3.055 ;
      RECT 8.62 1.955 8.865 2.77 ;
      RECT 8.655 1.84 8.935 2.21 ;
      RECT 8.655 1.945 9.5 2.145 ;
      RECT 7.975 2.425 8.235 2.745 ;
      RECT 7.315 2.515 8.235 2.655 ;
      RECT 7.315 1.575 7.455 2.655 ;
      RECT 3.775 1.865 4.035 2.185 ;
      RECT 3.955 1.575 4.095 2.095 ;
      RECT 3.955 1.575 7.455 1.715 ;
      RECT -1.255 7 -0.965 7.35 ;
      RECT -1.255 7.07 -0.035 7.24 ;
      RECT -0.205 6.69 -0.035 7.24 ;
      RECT 6.89 6.61 7.24 6.96 ;
      RECT -0.205 6.69 7.24 6.86 ;
      RECT 6.805 3.265 7.065 3.585 ;
      RECT 6.865 1.855 7.005 3.585 ;
      RECT 6.795 1.855 7.075 2.225 ;
      RECT 4.195 4.015 6.63 4.155 ;
      RECT 6.49 2.705 6.63 4.155 ;
      RECT 4.195 3.635 4.335 4.155 ;
      RECT 3.895 3.635 4.335 3.865 ;
      RECT 1.555 3.635 4.335 3.775 ;
      RECT 3.895 3.545 4.155 3.865 ;
      RECT 1.555 3.355 1.695 3.775 ;
      RECT 1.045 3.265 1.305 3.585 ;
      RECT 1.045 3.355 1.695 3.495 ;
      RECT 1.105 1.865 1.245 3.585 ;
      RECT 6.43 2.705 6.69 3.025 ;
      RECT 1.045 1.865 1.305 2.185 ;
      RECT 6.055 3.545 6.315 3.865 ;
      RECT 6.115 1.955 6.255 3.865 ;
      RECT 5.775 1.955 6.255 2.23 ;
      RECT 5.575 1.86 6.055 2.205 ;
      RECT 5.565 3.495 5.845 3.865 ;
      RECT 5.635 2.4 5.775 3.865 ;
      RECT 5.575 2.4 5.835 3.025 ;
      RECT 5.565 2.4 5.845 2.77 ;
      RECT 4.495 3.545 4.755 3.865 ;
      RECT 4.495 3.355 4.695 3.865 ;
      RECT 4.3 3.355 4.695 3.495 ;
      RECT 4.3 1.865 4.44 3.495 ;
      RECT 4.3 1.865 4.615 2.235 ;
      RECT 4.24 1.865 4.615 2.185 ;
      RECT 1.965 2.96 2.245 3.33 ;
      RECT 3.415 2.985 3.675 3.305 ;
      RECT 1.795 3.075 3.675 3.215 ;
      RECT 1.795 2.96 2.245 3.215 ;
      RECT 1.735 2.4 1.995 3.025 ;
      RECT 1.725 2.4 2.005 2.77 ;
      RECT 2.805 2.4 3.215 2.77 ;
      RECT 2.215 2.425 2.475 2.745 ;
      RECT 2.215 2.515 3.215 2.655 ;
      RECT 1.725 1.84 2.005 2.21 ;
      RECT 1.725 1.865 2.115 2.185 ;
      RECT 67.26 7.06 67.63 7.43 ;
      RECT 66.125 2.4 66.405 2.865 ;
      RECT 65.885 1.865 66.165 2.21 ;
      RECT 64.685 2.4 64.965 2.77 ;
      RECT 62.125 1.22 62.495 1.225 ;
      RECT 52 7.06 52.37 7.43 ;
      RECT 50.865 2.4 51.145 2.865 ;
      RECT 50.625 1.865 50.905 2.21 ;
      RECT 49.425 2.4 49.705 2.77 ;
      RECT 46.865 1.22 47.235 1.225 ;
      RECT 36.74 7.06 37.11 7.43 ;
      RECT 35.605 2.4 35.885 2.865 ;
      RECT 35.365 1.865 35.645 2.21 ;
      RECT 34.165 2.4 34.445 2.77 ;
      RECT 31.605 1.22 31.975 1.225 ;
      RECT 21.48 7.06 21.85 7.43 ;
      RECT 20.345 2.4 20.625 2.865 ;
      RECT 20.105 1.865 20.385 2.21 ;
      RECT 18.905 2.4 19.185 2.77 ;
      RECT 16.345 1.22 16.715 1.225 ;
      RECT 6.22 7.06 6.59 7.43 ;
      RECT 5.085 2.4 5.365 2.865 ;
      RECT 4.845 1.865 5.125 2.21 ;
      RECT 3.645 2.4 3.925 2.77 ;
      RECT 1.085 1.22 1.455 1.225 ;
    LAYER via1 ;
      RECT 75.83 7.38 75.98 7.53 ;
      RECT 73.46 6.745 73.61 6.895 ;
      RECT 73.445 2.07 73.595 2.22 ;
      RECT 72.655 2.455 72.805 2.605 ;
      RECT 72.655 6.33 72.805 6.48 ;
      RECT 71.625 2.81 71.775 2.96 ;
      RECT 71.625 5.965 71.775 6.115 ;
      RECT 71.065 2.805 71.215 2.955 ;
      RECT 69.76 1.95 69.91 2.1 ;
      RECT 69.76 3.63 69.91 3.78 ;
      RECT 69.07 2.51 69.22 2.66 ;
      RECT 68.03 6.715 68.18 6.865 ;
      RECT 67.9 1.95 68.05 2.1 ;
      RECT 67.9 3.35 68.05 3.5 ;
      RECT 67.525 2.79 67.675 2.94 ;
      RECT 67.37 7.17 67.52 7.32 ;
      RECT 67.15 3.63 67.3 3.78 ;
      RECT 66.67 1.95 66.82 2.1 ;
      RECT 66.67 2.79 66.82 2.94 ;
      RECT 66.19 2.51 66.34 2.66 ;
      RECT 65.95 1.95 66.1 2.1 ;
      RECT 65.59 3.63 65.74 3.78 ;
      RECT 65.335 1.95 65.485 2.1 ;
      RECT 64.99 3.63 65.14 3.78 ;
      RECT 64.87 1.95 65.02 2.1 ;
      RECT 64.75 2.51 64.9 2.66 ;
      RECT 64.51 3.07 64.66 3.22 ;
      RECT 63.31 2.51 63.46 2.66 ;
      RECT 62.95 1.95 63.1 2.1 ;
      RECT 62.83 2.79 62.98 2.94 ;
      RECT 62.14 1.95 62.29 2.1 ;
      RECT 62.14 3.35 62.29 3.5 ;
      RECT 60.545 6.76 60.695 6.91 ;
      RECT 58.2 6.745 58.35 6.895 ;
      RECT 58.185 2.07 58.335 2.22 ;
      RECT 57.395 2.455 57.545 2.605 ;
      RECT 57.395 6.33 57.545 6.48 ;
      RECT 56.365 2.81 56.515 2.96 ;
      RECT 56.365 5.965 56.515 6.115 ;
      RECT 55.805 2.805 55.955 2.955 ;
      RECT 54.5 1.95 54.65 2.1 ;
      RECT 54.5 3.63 54.65 3.78 ;
      RECT 53.81 2.51 53.96 2.66 ;
      RECT 52.775 6.715 52.925 6.865 ;
      RECT 52.64 1.95 52.79 2.1 ;
      RECT 52.64 3.35 52.79 3.5 ;
      RECT 52.265 2.79 52.415 2.94 ;
      RECT 52.11 7.17 52.26 7.32 ;
      RECT 51.89 3.63 52.04 3.78 ;
      RECT 51.41 1.95 51.56 2.1 ;
      RECT 51.41 2.79 51.56 2.94 ;
      RECT 50.93 2.51 51.08 2.66 ;
      RECT 50.69 1.95 50.84 2.1 ;
      RECT 50.33 3.63 50.48 3.78 ;
      RECT 50.075 1.95 50.225 2.1 ;
      RECT 49.73 3.63 49.88 3.78 ;
      RECT 49.61 1.95 49.76 2.1 ;
      RECT 49.49 2.51 49.64 2.66 ;
      RECT 49.25 3.07 49.4 3.22 ;
      RECT 48.05 2.51 48.2 2.66 ;
      RECT 47.69 1.95 47.84 2.1 ;
      RECT 47.57 2.79 47.72 2.94 ;
      RECT 46.88 1.95 47.03 2.1 ;
      RECT 46.88 3.35 47.03 3.5 ;
      RECT 45.285 6.76 45.435 6.91 ;
      RECT 42.94 6.745 43.09 6.895 ;
      RECT 42.925 2.07 43.075 2.22 ;
      RECT 42.135 2.455 42.285 2.605 ;
      RECT 42.135 6.33 42.285 6.48 ;
      RECT 41.105 2.81 41.255 2.96 ;
      RECT 41.105 5.965 41.255 6.115 ;
      RECT 40.545 2.805 40.695 2.955 ;
      RECT 39.24 1.95 39.39 2.1 ;
      RECT 39.24 3.63 39.39 3.78 ;
      RECT 38.55 2.51 38.7 2.66 ;
      RECT 37.51 6.72 37.66 6.87 ;
      RECT 37.38 1.95 37.53 2.1 ;
      RECT 37.38 3.35 37.53 3.5 ;
      RECT 37.005 2.79 37.155 2.94 ;
      RECT 36.85 7.17 37 7.32 ;
      RECT 36.63 3.63 36.78 3.78 ;
      RECT 36.15 1.95 36.3 2.1 ;
      RECT 36.15 2.79 36.3 2.94 ;
      RECT 35.67 2.51 35.82 2.66 ;
      RECT 35.43 1.95 35.58 2.1 ;
      RECT 35.07 3.63 35.22 3.78 ;
      RECT 34.815 1.95 34.965 2.1 ;
      RECT 34.47 3.63 34.62 3.78 ;
      RECT 34.35 1.95 34.5 2.1 ;
      RECT 34.23 2.51 34.38 2.66 ;
      RECT 33.99 3.07 34.14 3.22 ;
      RECT 32.79 2.51 32.94 2.66 ;
      RECT 32.43 1.95 32.58 2.1 ;
      RECT 32.31 2.79 32.46 2.94 ;
      RECT 31.62 1.95 31.77 2.1 ;
      RECT 31.62 3.35 31.77 3.5 ;
      RECT 30.07 6.765 30.22 6.915 ;
      RECT 27.68 6.745 27.83 6.895 ;
      RECT 27.665 2.07 27.815 2.22 ;
      RECT 26.875 2.455 27.025 2.605 ;
      RECT 26.875 6.33 27.025 6.48 ;
      RECT 25.845 2.81 25.995 2.96 ;
      RECT 25.845 5.965 25.995 6.115 ;
      RECT 25.285 2.805 25.435 2.955 ;
      RECT 23.98 1.95 24.13 2.1 ;
      RECT 23.98 3.63 24.13 3.78 ;
      RECT 23.29 2.51 23.44 2.66 ;
      RECT 22.25 6.715 22.4 6.865 ;
      RECT 22.12 1.95 22.27 2.1 ;
      RECT 22.12 3.35 22.27 3.5 ;
      RECT 21.745 2.79 21.895 2.94 ;
      RECT 21.59 7.17 21.74 7.32 ;
      RECT 21.37 3.63 21.52 3.78 ;
      RECT 20.89 1.95 21.04 2.1 ;
      RECT 20.89 2.79 21.04 2.94 ;
      RECT 20.41 2.51 20.56 2.66 ;
      RECT 20.17 1.95 20.32 2.1 ;
      RECT 19.81 3.63 19.96 3.78 ;
      RECT 19.555 1.95 19.705 2.1 ;
      RECT 19.21 3.63 19.36 3.78 ;
      RECT 19.09 1.95 19.24 2.1 ;
      RECT 18.97 2.51 19.12 2.66 ;
      RECT 18.73 3.07 18.88 3.22 ;
      RECT 17.53 2.51 17.68 2.66 ;
      RECT 17.17 1.95 17.32 2.1 ;
      RECT 17.05 2.79 17.2 2.94 ;
      RECT 16.36 1.95 16.51 2.1 ;
      RECT 16.36 3.35 16.51 3.5 ;
      RECT 14.81 6.76 14.96 6.91 ;
      RECT 12.42 6.745 12.57 6.895 ;
      RECT 12.405 2.07 12.555 2.22 ;
      RECT 11.615 2.455 11.765 2.605 ;
      RECT 11.615 6.33 11.765 6.48 ;
      RECT 10.585 2.81 10.735 2.96 ;
      RECT 10.585 5.965 10.735 6.115 ;
      RECT 10.025 2.805 10.175 2.955 ;
      RECT 8.72 1.95 8.87 2.1 ;
      RECT 8.72 3.63 8.87 3.78 ;
      RECT 8.03 2.51 8.18 2.66 ;
      RECT 6.99 6.71 7.14 6.86 ;
      RECT 6.86 1.95 7.01 2.1 ;
      RECT 6.86 3.35 7.01 3.5 ;
      RECT 6.485 2.79 6.635 2.94 ;
      RECT 6.33 7.17 6.48 7.32 ;
      RECT 6.11 3.63 6.26 3.78 ;
      RECT 5.63 1.95 5.78 2.1 ;
      RECT 5.63 2.79 5.78 2.94 ;
      RECT 5.15 2.51 5.3 2.66 ;
      RECT 4.91 1.95 5.06 2.1 ;
      RECT 4.55 3.63 4.7 3.78 ;
      RECT 4.295 1.95 4.445 2.1 ;
      RECT 3.95 3.63 4.1 3.78 ;
      RECT 3.83 1.95 3.98 2.1 ;
      RECT 3.71 2.51 3.86 2.66 ;
      RECT 3.47 3.07 3.62 3.22 ;
      RECT 2.27 2.51 2.42 2.66 ;
      RECT 1.91 1.95 2.06 2.1 ;
      RECT 1.79 2.79 1.94 2.94 ;
      RECT 1.1 1.95 1.25 2.1 ;
      RECT 1.1 3.35 1.25 3.5 ;
      RECT -1.185 7.1 -1.035 7.25 ;
      RECT -1.56 6.36 -1.41 6.51 ;
    LAYER met1 ;
      RECT 62.28 2.75 62.57 2.98 ;
      RECT 47.02 2.75 47.31 2.98 ;
      RECT 31.76 2.75 32.05 2.98 ;
      RECT 16.5 2.75 16.79 2.98 ;
      RECT 1.24 2.75 1.53 2.98 ;
      RECT 62.355 2.375 62.495 2.98 ;
      RECT 47.095 2.375 47.235 2.98 ;
      RECT 31.835 2.375 31.975 2.98 ;
      RECT 16.575 2.375 16.715 2.98 ;
      RECT 1.315 2.375 1.455 2.98 ;
      RECT 62.355 2.375 62.975 2.515 ;
      RECT 62.835 0.005 62.975 2.515 ;
      RECT 47.095 2.375 47.715 2.515 ;
      RECT 47.575 0.005 47.715 2.515 ;
      RECT 31.835 2.375 32.455 2.515 ;
      RECT 32.315 0.005 32.455 2.515 ;
      RECT 16.575 2.375 17.195 2.515 ;
      RECT 17.055 0.005 17.195 2.515 ;
      RECT 1.315 2.375 1.935 2.515 ;
      RECT 1.795 0.005 1.935 2.515 ;
      RECT 62.595 1.955 62.975 2.215 ;
      RECT 47.335 1.955 47.715 2.215 ;
      RECT 32.075 1.955 32.455 2.215 ;
      RECT 16.815 1.955 17.195 2.215 ;
      RECT 1.555 1.955 1.935 2.215 ;
      RECT 62.775 1.895 63.185 2.155 ;
      RECT 47.515 1.895 47.925 2.155 ;
      RECT 32.255 1.895 32.665 2.155 ;
      RECT 16.995 1.895 17.405 2.155 ;
      RECT 1.735 1.895 2.145 2.155 ;
      RECT 63.48 1.91 63.77 2.14 ;
      RECT 48.22 1.91 48.51 2.14 ;
      RECT 32.96 1.91 33.25 2.14 ;
      RECT 17.7 1.91 17.99 2.14 ;
      RECT 2.44 1.91 2.73 2.14 ;
      RECT 62.595 1.955 63.77 2.095 ;
      RECT 47.335 1.955 48.51 2.095 ;
      RECT 32.075 1.955 33.25 2.095 ;
      RECT 16.815 1.955 17.99 2.095 ;
      RECT 1.555 1.955 2.73 2.095 ;
      RECT 62.775 0.005 63.065 2.155 ;
      RECT 47.515 0.005 47.805 2.155 ;
      RECT 32.255 0.005 32.545 2.155 ;
      RECT 16.995 0.005 17.285 2.155 ;
      RECT 1.735 0.005 2.025 2.155 ;
      RECT 61.79 0.005 70.53 1.745 ;
      RECT 46.53 0.005 55.27 1.745 ;
      RECT 31.27 0.005 40.01 1.745 ;
      RECT 16.01 0.005 24.75 1.745 ;
      RECT 0.75 0.005 9.49 1.745 ;
      RECT -2.75 0.005 76.3 0.31 ;
      RECT -2.75 4.145 76.3 4.75 ;
      RECT 61.79 4.14 76.3 4.75 ;
      RECT 46.53 4.14 61.04 4.75 ;
      RECT 31.27 4.14 45.78 4.75 ;
      RECT 16.01 4.14 30.52 4.75 ;
      RECT 0.75 4.14 15.26 4.75 ;
      RECT 61.79 3.985 70.53 4.75 ;
      RECT 46.53 3.985 55.27 4.75 ;
      RECT 31.27 3.985 40.01 4.75 ;
      RECT 16.01 3.985 24.75 4.75 ;
      RECT 0.75 3.985 9.49 4.75 ;
      RECT -2.75 8.58 76.3 8.885 ;
      RECT 66.76 6.32 66.93 8.885 ;
      RECT 51.5 6.32 51.67 8.885 ;
      RECT 36.24 6.32 36.41 8.885 ;
      RECT 20.98 6.32 21.15 8.885 ;
      RECT 5.72 6.32 5.89 8.885 ;
      RECT 66.925 6.29 67.215 6.52 ;
      RECT 51.665 6.29 51.955 6.52 ;
      RECT 36.405 6.29 36.695 6.52 ;
      RECT 21.145 6.29 21.435 6.52 ;
      RECT 5.885 6.29 6.175 6.52 ;
      RECT 66.755 6.32 67.215 6.49 ;
      RECT 51.495 6.32 51.955 6.49 ;
      RECT 36.235 6.32 36.695 6.49 ;
      RECT 20.975 6.32 21.435 6.49 ;
      RECT 5.715 6.32 6.175 6.49 ;
      RECT 75.7 7.77 75.99 8 ;
      RECT 75.76 6.29 75.93 8 ;
      RECT 75.73 7.28 76.08 7.63 ;
      RECT 75.7 6.29 75.99 6.52 ;
      RECT 75.7 2.37 75.99 2.6 ;
      RECT 75.76 0.89 75.93 2.6 ;
      RECT 75.7 0.89 75.99 1.12 ;
      RECT 75.29 2.74 75.62 2.97 ;
      RECT 75.29 2.77 75.79 2.94 ;
      RECT 75.29 2.4 75.48 2.97 ;
      RECT 74.71 2.37 75 2.6 ;
      RECT 74.71 2.4 75.48 2.57 ;
      RECT 74.77 0.89 74.94 2.6 ;
      RECT 74.71 0.89 75 1.12 ;
      RECT 74.71 7.77 75 8 ;
      RECT 74.77 6.29 74.94 8 ;
      RECT 74.71 6.29 75 6.52 ;
      RECT 74.71 6.33 75.56 6.49 ;
      RECT 75.39 5.92 75.56 6.49 ;
      RECT 74.71 6.325 75.1 6.49 ;
      RECT 75.33 5.92 75.62 6.15 ;
      RECT 75.33 5.95 75.79 6.12 ;
      RECT 74.34 2.74 74.63 2.97 ;
      RECT 74.34 2.77 74.8 2.94 ;
      RECT 74.4 1.66 74.565 2.97 ;
      RECT 72.915 1.63 73.205 1.86 ;
      RECT 72.915 1.66 74.565 1.83 ;
      RECT 72.975 0.89 73.145 1.86 ;
      RECT 72.915 0.89 73.205 1.12 ;
      RECT 72.915 7.77 73.205 8 ;
      RECT 72.975 7.03 73.145 8 ;
      RECT 72.975 7.125 74.565 7.295 ;
      RECT 74.395 5.92 74.565 7.295 ;
      RECT 72.915 7.03 73.205 7.26 ;
      RECT 74.34 5.92 74.63 6.15 ;
      RECT 74.34 5.95 74.8 6.12 ;
      RECT 70.965 2.705 71.305 3.055 ;
      RECT 71.055 2.03 71.225 3.055 ;
      RECT 73.345 1.97 73.695 2.32 ;
      RECT 71.055 2.03 73.695 2.2 ;
      RECT 73.37 6.66 73.695 6.985 ;
      RECT 67.93 6.615 68.28 6.965 ;
      RECT 73.345 6.66 73.695 6.89 ;
      RECT 67.73 6.66 68.28 6.89 ;
      RECT 67.56 6.69 73.695 6.86 ;
      RECT 72.57 2.37 72.89 2.69 ;
      RECT 72.54 2.37 72.89 2.6 ;
      RECT 72.37 2.4 72.89 2.57 ;
      RECT 72.57 6.26 72.89 6.55 ;
      RECT 72.54 6.29 72.89 6.52 ;
      RECT 72.37 6.32 72.89 6.49 ;
      RECT 71.525 2.71 71.865 3.06 ;
      RECT 71.525 2.77 72.005 2.94 ;
      RECT 71.525 5.865 71.865 6.215 ;
      RECT 65.93 5.92 66.22 6.15 ;
      RECT 65.93 5.95 72.005 6.12 ;
      RECT 69.675 1.895 69.995 2.155 ;
      RECT 69.24 1.91 69.53 2.14 ;
      RECT 69.24 1.955 69.995 2.095 ;
      RECT 69.675 3.575 69.995 3.835 ;
      RECT 69.24 3.59 69.53 3.82 ;
      RECT 69.24 3.635 69.995 3.775 ;
      RECT 69 3.03 69.29 3.26 ;
      RECT 69 3.075 69.575 3.215 ;
      RECT 69.435 2.935 69.695 3.075 ;
      RECT 69.48 2.75 69.77 2.98 ;
      RECT 67.635 2.935 68.735 3.075 ;
      RECT 67.44 2.735 67.76 2.995 ;
      RECT 68.52 2.75 68.81 2.98 ;
      RECT 67.44 2.75 67.85 2.995 ;
      RECT 67.815 1.895 68.135 2.155 ;
      RECT 68.28 1.91 68.57 2.14 ;
      RECT 67.815 1.955 68.57 2.095 ;
      RECT 65.115 3.16 67.295 3.3 ;
      RECT 67.155 2.17 67.295 3.3 ;
      RECT 65.115 3.075 66.41 3.3 ;
      RECT 66.12 3.03 66.41 3.3 ;
      RECT 65.115 2.795 65.45 3.3 ;
      RECT 65.16 2.75 65.45 3.3 ;
      RECT 68.04 2.47 68.33 2.7 ;
      RECT 67.155 2.375 68.255 2.515 ;
      RECT 67.08 2.17 67.37 2.42 ;
      RECT 67.3 7.77 67.59 8 ;
      RECT 67.36 7.03 67.53 8 ;
      RECT 67.26 7.06 67.63 7.43 ;
      RECT 67.3 7.03 67.59 7.43 ;
      RECT 67.065 3.575 67.385 3.835 ;
      RECT 67.065 3.59 67.58 3.82 ;
      RECT 65.64 2.47 65.93 2.7 ;
      RECT 65.79 2.075 65.93 2.7 ;
      RECT 65.79 2.075 66.095 2.215 ;
      RECT 66.585 1.895 66.905 2.155 ;
      RECT 65.865 1.895 66.185 2.155 ;
      RECT 66.36 1.91 66.905 2.14 ;
      RECT 65.865 1.955 66.905 2.095 ;
      RECT 65.505 3.575 65.825 3.835 ;
      RECT 65.4 3.59 65.825 3.82 ;
      RECT 63.48 3.03 63.77 3.26 ;
      RECT 63.48 3.03 63.935 3.215 ;
      RECT 63.795 2.555 63.935 3.215 ;
      RECT 63.915 1.955 64.055 2.695 ;
      RECT 64.785 1.895 65.105 2.155 ;
      RECT 63.96 1.91 64.25 2.14 ;
      RECT 63.915 1.955 65.105 2.095 ;
      RECT 64.665 2.455 64.985 2.715 ;
      RECT 64.2 2.47 64.49 2.7 ;
      RECT 64.2 2.515 64.985 2.655 ;
      RECT 64.425 3.015 64.745 3.275 ;
      RECT 64.425 3.03 64.97 3.26 ;
      RECT 63.96 3.59 64.25 3.82 ;
      RECT 63.075 3.47 64.175 3.61 ;
      RECT 63 3.31 63.29 3.54 ;
      RECT 60.44 7.77 60.73 8 ;
      RECT 60.5 6.29 60.67 8 ;
      RECT 60.445 6.66 60.795 7.01 ;
      RECT 60.44 6.29 60.73 6.52 ;
      RECT 60.44 2.37 60.73 2.6 ;
      RECT 60.5 0.89 60.67 2.6 ;
      RECT 60.44 0.89 60.73 1.12 ;
      RECT 60.03 2.74 60.36 2.97 ;
      RECT 60.03 2.77 60.53 2.94 ;
      RECT 60.03 2.4 60.22 2.97 ;
      RECT 59.45 2.37 59.74 2.6 ;
      RECT 59.45 2.4 60.22 2.57 ;
      RECT 59.51 0.89 59.68 2.6 ;
      RECT 59.45 0.89 59.74 1.12 ;
      RECT 59.45 7.77 59.74 8 ;
      RECT 59.51 6.29 59.68 8 ;
      RECT 59.45 6.29 59.74 6.52 ;
      RECT 59.45 6.33 60.3 6.49 ;
      RECT 60.13 5.92 60.3 6.49 ;
      RECT 59.45 6.325 59.84 6.49 ;
      RECT 60.07 5.92 60.36 6.15 ;
      RECT 60.07 5.95 60.53 6.12 ;
      RECT 59.08 2.74 59.37 2.97 ;
      RECT 59.08 2.77 59.54 2.94 ;
      RECT 59.14 1.66 59.305 2.97 ;
      RECT 57.655 1.63 57.945 1.86 ;
      RECT 57.655 1.66 59.305 1.83 ;
      RECT 57.715 0.89 57.885 1.86 ;
      RECT 57.655 0.89 57.945 1.12 ;
      RECT 57.655 7.77 57.945 8 ;
      RECT 57.715 7.03 57.885 8 ;
      RECT 57.715 7.125 59.305 7.295 ;
      RECT 59.135 5.92 59.305 7.295 ;
      RECT 57.655 7.03 57.945 7.26 ;
      RECT 59.08 5.92 59.37 6.15 ;
      RECT 59.08 5.95 59.54 6.12 ;
      RECT 55.705 2.705 56.045 3.055 ;
      RECT 55.795 2.03 55.965 3.055 ;
      RECT 58.085 1.97 58.435 2.32 ;
      RECT 55.795 2.03 58.435 2.2 ;
      RECT 58.11 6.66 58.435 6.985 ;
      RECT 52.675 6.615 53.025 6.965 ;
      RECT 58.085 6.66 58.435 6.89 ;
      RECT 52.47 6.66 53.025 6.89 ;
      RECT 52.3 6.69 58.435 6.86 ;
      RECT 57.31 2.37 57.63 2.69 ;
      RECT 57.28 2.37 57.63 2.6 ;
      RECT 57.11 2.4 57.63 2.57 ;
      RECT 57.31 6.26 57.63 6.55 ;
      RECT 57.28 6.29 57.63 6.52 ;
      RECT 57.11 6.32 57.63 6.49 ;
      RECT 56.265 2.71 56.605 3.06 ;
      RECT 56.265 2.77 56.745 2.94 ;
      RECT 56.265 5.865 56.605 6.215 ;
      RECT 50.67 5.92 50.96 6.15 ;
      RECT 50.67 5.95 56.745 6.12 ;
      RECT 54.415 1.895 54.735 2.155 ;
      RECT 53.98 1.91 54.27 2.14 ;
      RECT 53.98 1.955 54.735 2.095 ;
      RECT 54.415 3.575 54.735 3.835 ;
      RECT 53.98 3.59 54.27 3.82 ;
      RECT 53.98 3.635 54.735 3.775 ;
      RECT 53.74 3.03 54.03 3.26 ;
      RECT 53.74 3.075 54.315 3.215 ;
      RECT 54.175 2.935 54.435 3.075 ;
      RECT 54.22 2.75 54.51 2.98 ;
      RECT 52.375 2.935 53.475 3.075 ;
      RECT 52.18 2.735 52.5 2.995 ;
      RECT 53.26 2.75 53.55 2.98 ;
      RECT 52.18 2.75 52.59 2.995 ;
      RECT 52.555 1.895 52.875 2.155 ;
      RECT 53.02 1.91 53.31 2.14 ;
      RECT 52.555 1.955 53.31 2.095 ;
      RECT 49.855 3.16 52.035 3.3 ;
      RECT 51.895 2.17 52.035 3.3 ;
      RECT 49.855 3.075 51.15 3.3 ;
      RECT 50.86 3.03 51.15 3.3 ;
      RECT 49.855 2.795 50.19 3.3 ;
      RECT 49.9 2.75 50.19 3.3 ;
      RECT 52.78 2.47 53.07 2.7 ;
      RECT 51.895 2.375 52.995 2.515 ;
      RECT 51.82 2.17 52.11 2.42 ;
      RECT 52.04 7.77 52.33 8 ;
      RECT 52.1 7.03 52.27 8 ;
      RECT 52 7.06 52.37 7.43 ;
      RECT 52.04 7.03 52.33 7.43 ;
      RECT 51.805 3.575 52.125 3.835 ;
      RECT 51.805 3.59 52.32 3.82 ;
      RECT 50.38 2.47 50.67 2.7 ;
      RECT 50.53 2.075 50.67 2.7 ;
      RECT 50.53 2.075 50.835 2.215 ;
      RECT 51.325 1.895 51.645 2.155 ;
      RECT 50.605 1.895 50.925 2.155 ;
      RECT 51.1 1.91 51.645 2.14 ;
      RECT 50.605 1.955 51.645 2.095 ;
      RECT 50.245 3.575 50.565 3.835 ;
      RECT 50.14 3.59 50.565 3.82 ;
      RECT 48.22 3.03 48.51 3.26 ;
      RECT 48.22 3.03 48.675 3.215 ;
      RECT 48.535 2.555 48.675 3.215 ;
      RECT 48.655 1.955 48.795 2.695 ;
      RECT 49.525 1.895 49.845 2.155 ;
      RECT 48.7 1.91 48.99 2.14 ;
      RECT 48.655 1.955 49.845 2.095 ;
      RECT 49.405 2.455 49.725 2.715 ;
      RECT 48.94 2.47 49.23 2.7 ;
      RECT 48.94 2.515 49.725 2.655 ;
      RECT 49.165 3.015 49.485 3.275 ;
      RECT 49.165 3.03 49.71 3.26 ;
      RECT 48.7 3.59 48.99 3.82 ;
      RECT 47.815 3.47 48.915 3.61 ;
      RECT 47.74 3.31 48.03 3.54 ;
      RECT 45.18 7.77 45.47 8 ;
      RECT 45.24 6.29 45.41 8 ;
      RECT 45.185 6.66 45.535 7.01 ;
      RECT 45.18 6.29 45.47 6.52 ;
      RECT 45.18 2.37 45.47 2.6 ;
      RECT 45.24 0.89 45.41 2.6 ;
      RECT 45.18 0.89 45.47 1.12 ;
      RECT 44.77 2.74 45.1 2.97 ;
      RECT 44.77 2.77 45.27 2.94 ;
      RECT 44.77 2.4 44.96 2.97 ;
      RECT 44.19 2.37 44.48 2.6 ;
      RECT 44.19 2.4 44.96 2.57 ;
      RECT 44.25 0.89 44.42 2.6 ;
      RECT 44.19 0.89 44.48 1.12 ;
      RECT 44.19 7.77 44.48 8 ;
      RECT 44.25 6.29 44.42 8 ;
      RECT 44.19 6.29 44.48 6.52 ;
      RECT 44.19 6.33 45.04 6.49 ;
      RECT 44.87 5.92 45.04 6.49 ;
      RECT 44.19 6.325 44.58 6.49 ;
      RECT 44.81 5.92 45.1 6.15 ;
      RECT 44.81 5.95 45.27 6.12 ;
      RECT 43.82 2.74 44.11 2.97 ;
      RECT 43.82 2.77 44.28 2.94 ;
      RECT 43.88 1.66 44.045 2.97 ;
      RECT 42.395 1.63 42.685 1.86 ;
      RECT 42.395 1.66 44.045 1.83 ;
      RECT 42.455 0.89 42.625 1.86 ;
      RECT 42.395 0.89 42.685 1.12 ;
      RECT 42.395 7.77 42.685 8 ;
      RECT 42.455 7.03 42.625 8 ;
      RECT 42.455 7.125 44.045 7.295 ;
      RECT 43.875 5.92 44.045 7.295 ;
      RECT 42.395 7.03 42.685 7.26 ;
      RECT 43.82 5.92 44.11 6.15 ;
      RECT 43.82 5.95 44.28 6.12 ;
      RECT 40.445 2.705 40.785 3.055 ;
      RECT 40.535 2.03 40.705 3.055 ;
      RECT 42.825 1.97 43.175 2.32 ;
      RECT 40.535 2.03 43.175 2.2 ;
      RECT 42.85 6.66 43.175 6.985 ;
      RECT 37.41 6.62 37.76 6.97 ;
      RECT 42.825 6.66 43.175 6.89 ;
      RECT 37.21 6.66 37.76 6.89 ;
      RECT 37.04 6.69 43.175 6.86 ;
      RECT 42.05 2.37 42.37 2.69 ;
      RECT 42.02 2.37 42.37 2.6 ;
      RECT 41.85 2.4 42.37 2.57 ;
      RECT 42.05 6.26 42.37 6.55 ;
      RECT 42.02 6.29 42.37 6.52 ;
      RECT 41.85 6.32 42.37 6.49 ;
      RECT 41.005 2.71 41.345 3.06 ;
      RECT 41.005 2.77 41.485 2.94 ;
      RECT 41.005 5.865 41.345 6.215 ;
      RECT 35.41 5.92 35.7 6.15 ;
      RECT 35.41 5.95 41.485 6.12 ;
      RECT 39.155 1.895 39.475 2.155 ;
      RECT 38.72 1.91 39.01 2.14 ;
      RECT 38.72 1.955 39.475 2.095 ;
      RECT 39.155 3.575 39.475 3.835 ;
      RECT 38.72 3.59 39.01 3.82 ;
      RECT 38.72 3.635 39.475 3.775 ;
      RECT 38.48 3.03 38.77 3.26 ;
      RECT 38.48 3.075 39.055 3.215 ;
      RECT 38.915 2.935 39.175 3.075 ;
      RECT 38.96 2.75 39.25 2.98 ;
      RECT 37.115 2.935 38.215 3.075 ;
      RECT 36.92 2.735 37.24 2.995 ;
      RECT 38 2.75 38.29 2.98 ;
      RECT 36.92 2.75 37.33 2.995 ;
      RECT 37.295 1.895 37.615 2.155 ;
      RECT 37.76 1.91 38.05 2.14 ;
      RECT 37.295 1.955 38.05 2.095 ;
      RECT 34.595 3.16 36.775 3.3 ;
      RECT 36.635 2.17 36.775 3.3 ;
      RECT 34.595 3.075 35.89 3.3 ;
      RECT 35.6 3.03 35.89 3.3 ;
      RECT 34.595 2.795 34.93 3.3 ;
      RECT 34.64 2.75 34.93 3.3 ;
      RECT 37.52 2.47 37.81 2.7 ;
      RECT 36.635 2.375 37.735 2.515 ;
      RECT 36.56 2.17 36.85 2.42 ;
      RECT 36.78 7.77 37.07 8 ;
      RECT 36.84 7.03 37.01 8 ;
      RECT 36.74 7.06 37.11 7.43 ;
      RECT 36.78 7.03 37.07 7.43 ;
      RECT 36.545 3.575 36.865 3.835 ;
      RECT 36.545 3.59 37.06 3.82 ;
      RECT 35.12 2.47 35.41 2.7 ;
      RECT 35.27 2.075 35.41 2.7 ;
      RECT 35.27 2.075 35.575 2.215 ;
      RECT 36.065 1.895 36.385 2.155 ;
      RECT 35.345 1.895 35.665 2.155 ;
      RECT 35.84 1.91 36.385 2.14 ;
      RECT 35.345 1.955 36.385 2.095 ;
      RECT 34.985 3.575 35.305 3.835 ;
      RECT 34.88 3.59 35.305 3.82 ;
      RECT 32.96 3.03 33.25 3.26 ;
      RECT 32.96 3.03 33.415 3.215 ;
      RECT 33.275 2.555 33.415 3.215 ;
      RECT 33.395 1.955 33.535 2.695 ;
      RECT 34.265 1.895 34.585 2.155 ;
      RECT 33.44 1.91 33.73 2.14 ;
      RECT 33.395 1.955 34.585 2.095 ;
      RECT 34.145 2.455 34.465 2.715 ;
      RECT 33.68 2.47 33.97 2.7 ;
      RECT 33.68 2.515 34.465 2.655 ;
      RECT 33.905 3.015 34.225 3.275 ;
      RECT 33.905 3.03 34.45 3.26 ;
      RECT 33.44 3.59 33.73 3.82 ;
      RECT 32.555 3.47 33.655 3.61 ;
      RECT 32.48 3.31 32.77 3.54 ;
      RECT 29.92 7.77 30.21 8 ;
      RECT 29.98 6.29 30.15 8 ;
      RECT 29.965 6.665 30.32 7.02 ;
      RECT 29.92 6.29 30.21 6.52 ;
      RECT 29.92 2.37 30.21 2.6 ;
      RECT 29.98 0.89 30.15 2.6 ;
      RECT 29.92 0.89 30.21 1.12 ;
      RECT 29.51 2.74 29.84 2.97 ;
      RECT 29.51 2.77 30.01 2.94 ;
      RECT 29.51 2.4 29.7 2.97 ;
      RECT 28.93 2.37 29.22 2.6 ;
      RECT 28.93 2.4 29.7 2.57 ;
      RECT 28.99 0.89 29.16 2.6 ;
      RECT 28.93 0.89 29.22 1.12 ;
      RECT 28.93 7.77 29.22 8 ;
      RECT 28.99 6.29 29.16 8 ;
      RECT 28.93 6.29 29.22 6.52 ;
      RECT 28.93 6.33 29.78 6.49 ;
      RECT 29.61 5.92 29.78 6.49 ;
      RECT 28.93 6.325 29.32 6.49 ;
      RECT 29.55 5.92 29.84 6.15 ;
      RECT 29.55 5.95 30.01 6.12 ;
      RECT 28.56 2.74 28.85 2.97 ;
      RECT 28.56 2.77 29.02 2.94 ;
      RECT 28.62 1.66 28.785 2.97 ;
      RECT 27.135 1.63 27.425 1.86 ;
      RECT 27.135 1.66 28.785 1.83 ;
      RECT 27.195 0.89 27.365 1.86 ;
      RECT 27.135 0.89 27.425 1.12 ;
      RECT 27.135 7.77 27.425 8 ;
      RECT 27.195 7.03 27.365 8 ;
      RECT 27.195 7.125 28.785 7.295 ;
      RECT 28.615 5.92 28.785 7.295 ;
      RECT 27.135 7.03 27.425 7.26 ;
      RECT 28.56 5.92 28.85 6.15 ;
      RECT 28.56 5.95 29.02 6.12 ;
      RECT 25.185 2.705 25.525 3.055 ;
      RECT 25.275 2.03 25.445 3.055 ;
      RECT 27.565 1.97 27.915 2.32 ;
      RECT 25.275 2.03 27.915 2.2 ;
      RECT 27.59 6.66 27.915 6.985 ;
      RECT 22.15 6.615 22.5 6.965 ;
      RECT 27.565 6.66 27.915 6.89 ;
      RECT 21.95 6.66 22.5 6.89 ;
      RECT 21.78 6.69 27.915 6.86 ;
      RECT 26.79 2.37 27.11 2.69 ;
      RECT 26.76 2.37 27.11 2.6 ;
      RECT 26.59 2.4 27.11 2.57 ;
      RECT 26.79 6.26 27.11 6.55 ;
      RECT 26.76 6.29 27.11 6.52 ;
      RECT 26.59 6.32 27.11 6.49 ;
      RECT 25.745 2.71 26.085 3.06 ;
      RECT 25.745 2.77 26.225 2.94 ;
      RECT 25.745 5.865 26.085 6.215 ;
      RECT 20.15 5.92 20.44 6.15 ;
      RECT 20.15 5.95 26.225 6.12 ;
      RECT 23.895 1.895 24.215 2.155 ;
      RECT 23.46 1.91 23.75 2.14 ;
      RECT 23.46 1.955 24.215 2.095 ;
      RECT 23.895 3.575 24.215 3.835 ;
      RECT 23.46 3.59 23.75 3.82 ;
      RECT 23.46 3.635 24.215 3.775 ;
      RECT 23.22 3.03 23.51 3.26 ;
      RECT 23.22 3.075 23.795 3.215 ;
      RECT 23.655 2.935 23.915 3.075 ;
      RECT 23.7 2.75 23.99 2.98 ;
      RECT 21.855 2.935 22.955 3.075 ;
      RECT 21.66 2.735 21.98 2.995 ;
      RECT 22.74 2.75 23.03 2.98 ;
      RECT 21.66 2.75 22.07 2.995 ;
      RECT 22.035 1.895 22.355 2.155 ;
      RECT 22.5 1.91 22.79 2.14 ;
      RECT 22.035 1.955 22.79 2.095 ;
      RECT 19.335 3.16 21.515 3.3 ;
      RECT 21.375 2.17 21.515 3.3 ;
      RECT 19.335 3.075 20.63 3.3 ;
      RECT 20.34 3.03 20.63 3.3 ;
      RECT 19.335 2.795 19.67 3.3 ;
      RECT 19.38 2.75 19.67 3.3 ;
      RECT 22.26 2.47 22.55 2.7 ;
      RECT 21.375 2.375 22.475 2.515 ;
      RECT 21.3 2.17 21.59 2.42 ;
      RECT 21.52 7.77 21.81 8 ;
      RECT 21.58 7.03 21.75 8 ;
      RECT 21.48 7.06 21.85 7.43 ;
      RECT 21.52 7.03 21.81 7.43 ;
      RECT 21.285 3.575 21.605 3.835 ;
      RECT 21.285 3.59 21.8 3.82 ;
      RECT 19.86 2.47 20.15 2.7 ;
      RECT 20.01 2.075 20.15 2.7 ;
      RECT 20.01 2.075 20.315 2.215 ;
      RECT 20.805 1.895 21.125 2.155 ;
      RECT 20.085 1.895 20.405 2.155 ;
      RECT 20.58 1.91 21.125 2.14 ;
      RECT 20.085 1.955 21.125 2.095 ;
      RECT 19.725 3.575 20.045 3.835 ;
      RECT 19.62 3.59 20.045 3.82 ;
      RECT 17.7 3.03 17.99 3.26 ;
      RECT 17.7 3.03 18.155 3.215 ;
      RECT 18.015 2.555 18.155 3.215 ;
      RECT 18.135 1.955 18.275 2.695 ;
      RECT 19.005 1.895 19.325 2.155 ;
      RECT 18.18 1.91 18.47 2.14 ;
      RECT 18.135 1.955 19.325 2.095 ;
      RECT 18.885 2.455 19.205 2.715 ;
      RECT 18.42 2.47 18.71 2.7 ;
      RECT 18.42 2.515 19.205 2.655 ;
      RECT 18.645 3.015 18.965 3.275 ;
      RECT 18.645 3.03 19.19 3.26 ;
      RECT 18.18 3.59 18.47 3.82 ;
      RECT 17.295 3.47 18.395 3.61 ;
      RECT 17.22 3.31 17.51 3.54 ;
      RECT 14.66 7.77 14.95 8 ;
      RECT 14.72 6.29 14.89 8 ;
      RECT 14.71 6.66 15.06 7.01 ;
      RECT 14.66 6.29 14.95 6.52 ;
      RECT 14.66 2.37 14.95 2.6 ;
      RECT 14.72 0.89 14.89 2.6 ;
      RECT 14.66 0.89 14.95 1.12 ;
      RECT 14.25 2.74 14.58 2.97 ;
      RECT 14.25 2.77 14.75 2.94 ;
      RECT 14.25 2.4 14.44 2.97 ;
      RECT 13.67 2.37 13.96 2.6 ;
      RECT 13.67 2.4 14.44 2.57 ;
      RECT 13.73 0.89 13.9 2.6 ;
      RECT 13.67 0.89 13.96 1.12 ;
      RECT 13.67 7.77 13.96 8 ;
      RECT 13.73 6.29 13.9 8 ;
      RECT 13.67 6.29 13.96 6.52 ;
      RECT 13.67 6.33 14.52 6.49 ;
      RECT 14.35 5.92 14.52 6.49 ;
      RECT 13.67 6.325 14.06 6.49 ;
      RECT 14.29 5.92 14.58 6.15 ;
      RECT 14.29 5.95 14.75 6.12 ;
      RECT 13.3 2.74 13.59 2.97 ;
      RECT 13.3 2.77 13.76 2.94 ;
      RECT 13.36 1.66 13.525 2.97 ;
      RECT 11.875 1.63 12.165 1.86 ;
      RECT 11.875 1.66 13.525 1.83 ;
      RECT 11.935 0.89 12.105 1.86 ;
      RECT 11.875 0.89 12.165 1.12 ;
      RECT 11.875 7.77 12.165 8 ;
      RECT 11.935 7.03 12.105 8 ;
      RECT 11.935 7.125 13.525 7.295 ;
      RECT 13.355 5.92 13.525 7.295 ;
      RECT 11.875 7.03 12.165 7.26 ;
      RECT 13.3 5.92 13.59 6.15 ;
      RECT 13.3 5.95 13.76 6.12 ;
      RECT 9.925 2.705 10.265 3.055 ;
      RECT 10.015 2.03 10.185 3.055 ;
      RECT 12.305 1.97 12.655 2.32 ;
      RECT 10.015 2.03 12.655 2.2 ;
      RECT 12.33 6.66 12.655 6.985 ;
      RECT 6.89 6.61 7.24 6.96 ;
      RECT 12.305 6.66 12.655 6.89 ;
      RECT 6.69 6.66 7.24 6.89 ;
      RECT 6.52 6.69 12.655 6.86 ;
      RECT 11.53 2.37 11.85 2.69 ;
      RECT 11.5 2.37 11.85 2.6 ;
      RECT 11.33 2.4 11.85 2.57 ;
      RECT 11.53 6.26 11.85 6.55 ;
      RECT 11.5 6.29 11.85 6.52 ;
      RECT 11.33 6.32 11.85 6.49 ;
      RECT 10.485 2.71 10.825 3.06 ;
      RECT 10.485 2.77 10.965 2.94 ;
      RECT 10.485 5.865 10.825 6.215 ;
      RECT 4.89 5.92 5.18 6.15 ;
      RECT 4.89 5.95 10.965 6.12 ;
      RECT 8.635 1.895 8.955 2.155 ;
      RECT 8.2 1.91 8.49 2.14 ;
      RECT 8.2 1.955 8.955 2.095 ;
      RECT 8.635 3.575 8.955 3.835 ;
      RECT 8.2 3.59 8.49 3.82 ;
      RECT 8.2 3.635 8.955 3.775 ;
      RECT 7.96 3.03 8.25 3.26 ;
      RECT 7.96 3.075 8.535 3.215 ;
      RECT 8.395 2.935 8.655 3.075 ;
      RECT 8.44 2.75 8.73 2.98 ;
      RECT 6.595 2.935 7.695 3.075 ;
      RECT 6.4 2.735 6.72 2.995 ;
      RECT 7.48 2.75 7.77 2.98 ;
      RECT 6.4 2.75 6.81 2.995 ;
      RECT 6.775 1.895 7.095 2.155 ;
      RECT 7.24 1.91 7.53 2.14 ;
      RECT 6.775 1.955 7.53 2.095 ;
      RECT 4.075 3.16 6.255 3.3 ;
      RECT 6.115 2.17 6.255 3.3 ;
      RECT 4.075 3.075 5.37 3.3 ;
      RECT 5.08 3.03 5.37 3.3 ;
      RECT 4.075 2.795 4.41 3.3 ;
      RECT 4.12 2.75 4.41 3.3 ;
      RECT 7 2.47 7.29 2.7 ;
      RECT 6.115 2.375 7.215 2.515 ;
      RECT 6.04 2.17 6.33 2.42 ;
      RECT 6.26 7.77 6.55 8 ;
      RECT 6.32 7.03 6.49 8 ;
      RECT 6.22 7.06 6.59 7.43 ;
      RECT 6.26 7.03 6.55 7.43 ;
      RECT 6.025 3.575 6.345 3.835 ;
      RECT 6.025 3.59 6.54 3.82 ;
      RECT 4.6 2.47 4.89 2.7 ;
      RECT 4.75 2.075 4.89 2.7 ;
      RECT 4.75 2.075 5.055 2.215 ;
      RECT 5.545 1.895 5.865 2.155 ;
      RECT 4.825 1.895 5.145 2.155 ;
      RECT 5.32 1.91 5.865 2.14 ;
      RECT 4.825 1.955 5.865 2.095 ;
      RECT 4.465 3.575 4.785 3.835 ;
      RECT 4.36 3.59 4.785 3.82 ;
      RECT 2.44 3.03 2.73 3.26 ;
      RECT 2.44 3.03 2.895 3.215 ;
      RECT 2.755 2.555 2.895 3.215 ;
      RECT 2.875 1.955 3.015 2.695 ;
      RECT 3.745 1.895 4.065 2.155 ;
      RECT 2.92 1.91 3.21 2.14 ;
      RECT 2.875 1.955 4.065 2.095 ;
      RECT 3.625 2.455 3.945 2.715 ;
      RECT 3.16 2.47 3.45 2.7 ;
      RECT 3.16 2.515 3.945 2.655 ;
      RECT 3.385 3.015 3.705 3.275 ;
      RECT 3.385 3.03 3.93 3.26 ;
      RECT 2.92 3.59 3.21 3.82 ;
      RECT 2.035 3.47 3.135 3.61 ;
      RECT 1.96 3.31 2.25 3.54 ;
      RECT -0.825 6.66 -0.535 6.89 ;
      RECT -0.995 6.69 -0.535 6.86 ;
      RECT -1.255 7.77 -0.965 8 ;
      RECT -1.195 7.03 -1.025 8 ;
      RECT -1.285 7.03 -0.935 7.32 ;
      RECT -1.66 6.29 -1.31 6.58 ;
      RECT -1.8 6.32 -1.31 6.49 ;
      RECT -2.625 5.92 -2.335 6.15 ;
      RECT -2.625 5.95 -2.165 6.12 ;
      RECT 68.985 2.455 69.305 2.715 ;
      RECT 67.815 3.295 68.135 3.555 ;
      RECT 66.585 2.735 66.905 2.995 ;
      RECT 66.105 2.455 66.425 2.715 ;
      RECT 65.25 1.895 65.65 2.155 ;
      RECT 64.905 3.575 65.225 3.835 ;
      RECT 63.225 2.455 63.545 2.715 ;
      RECT 62.745 2.735 63.065 2.995 ;
      RECT 62.055 1.895 62.375 2.155 ;
      RECT 62.055 3.295 62.375 3.555 ;
      RECT 53.725 2.455 54.045 2.715 ;
      RECT 52.555 3.295 52.875 3.555 ;
      RECT 51.325 2.735 51.645 2.995 ;
      RECT 50.845 2.455 51.165 2.715 ;
      RECT 49.99 1.895 50.39 2.155 ;
      RECT 49.645 3.575 49.965 3.835 ;
      RECT 47.965 2.455 48.285 2.715 ;
      RECT 47.485 2.735 47.805 2.995 ;
      RECT 46.795 1.895 47.115 2.155 ;
      RECT 46.795 3.295 47.115 3.555 ;
      RECT 38.465 2.455 38.785 2.715 ;
      RECT 37.295 3.295 37.615 3.555 ;
      RECT 36.065 2.735 36.385 2.995 ;
      RECT 35.585 2.455 35.905 2.715 ;
      RECT 34.73 1.895 35.13 2.155 ;
      RECT 34.385 3.575 34.705 3.835 ;
      RECT 32.705 2.455 33.025 2.715 ;
      RECT 32.225 2.735 32.545 2.995 ;
      RECT 31.535 1.895 31.855 2.155 ;
      RECT 31.535 3.295 31.855 3.555 ;
      RECT 23.205 2.455 23.525 2.715 ;
      RECT 22.035 3.295 22.355 3.555 ;
      RECT 20.805 2.735 21.125 2.995 ;
      RECT 20.325 2.455 20.645 2.715 ;
      RECT 19.47 1.895 19.87 2.155 ;
      RECT 19.125 3.575 19.445 3.835 ;
      RECT 17.445 2.455 17.765 2.715 ;
      RECT 16.965 2.735 17.285 2.995 ;
      RECT 16.275 1.895 16.595 2.155 ;
      RECT 16.275 3.295 16.595 3.555 ;
      RECT 7.945 2.455 8.265 2.715 ;
      RECT 6.775 3.295 7.095 3.555 ;
      RECT 5.545 2.735 5.865 2.995 ;
      RECT 5.065 2.455 5.385 2.715 ;
      RECT 4.21 1.895 4.61 2.155 ;
      RECT 3.865 3.575 4.185 3.835 ;
      RECT 2.185 2.455 2.505 2.715 ;
      RECT 1.705 2.735 2.025 2.995 ;
      RECT 1.015 1.895 1.335 2.155 ;
      RECT 1.015 3.295 1.335 3.555 ;
    LAYER mcon ;
      RECT 75.76 0.92 75.93 1.09 ;
      RECT 75.76 2.4 75.93 2.57 ;
      RECT 75.76 6.32 75.93 6.49 ;
      RECT 75.76 7.8 75.93 7.97 ;
      RECT 75.41 0.11 75.58 0.28 ;
      RECT 75.41 4.17 75.58 4.34 ;
      RECT 75.41 4.55 75.58 4.72 ;
      RECT 75.41 8.61 75.58 8.78 ;
      RECT 75.39 2.77 75.56 2.94 ;
      RECT 75.39 5.95 75.56 6.12 ;
      RECT 74.77 0.92 74.94 1.09 ;
      RECT 74.77 2.4 74.94 2.57 ;
      RECT 74.77 6.32 74.94 6.49 ;
      RECT 74.77 7.8 74.94 7.97 ;
      RECT 74.42 0.11 74.59 0.28 ;
      RECT 74.42 4.17 74.59 4.34 ;
      RECT 74.42 4.55 74.59 4.72 ;
      RECT 74.42 8.61 74.59 8.78 ;
      RECT 74.4 2.77 74.57 2.94 ;
      RECT 74.4 5.95 74.57 6.12 ;
      RECT 73.715 0.11 73.885 0.28 ;
      RECT 73.715 4.17 73.885 4.34 ;
      RECT 73.715 4.55 73.885 4.72 ;
      RECT 73.715 8.61 73.885 8.78 ;
      RECT 73.405 2.03 73.575 2.2 ;
      RECT 73.405 6.69 73.575 6.86 ;
      RECT 73.035 0.11 73.205 0.28 ;
      RECT 73.035 8.61 73.205 8.78 ;
      RECT 72.975 0.92 73.145 1.09 ;
      RECT 72.975 1.66 73.145 1.83 ;
      RECT 72.975 7.06 73.145 7.23 ;
      RECT 72.975 7.8 73.145 7.97 ;
      RECT 72.6 2.4 72.77 2.57 ;
      RECT 72.6 6.32 72.77 6.49 ;
      RECT 72.355 0.11 72.525 0.28 ;
      RECT 72.355 8.61 72.525 8.78 ;
      RECT 71.675 0.11 71.845 0.28 ;
      RECT 71.675 8.61 71.845 8.78 ;
      RECT 71.605 2.77 71.775 2.94 ;
      RECT 71.605 5.95 71.775 6.12 ;
      RECT 70.215 1.42 70.385 1.59 ;
      RECT 70.215 4.14 70.385 4.31 ;
      RECT 69.755 1.42 69.925 1.59 ;
      RECT 69.755 4.14 69.925 4.31 ;
      RECT 69.54 2.78 69.71 2.95 ;
      RECT 69.3 1.94 69.47 2.11 ;
      RECT 69.3 3.62 69.47 3.79 ;
      RECT 69.295 1.42 69.465 1.59 ;
      RECT 69.295 4.14 69.465 4.31 ;
      RECT 69.06 2.5 69.23 2.67 ;
      RECT 69.06 3.06 69.23 3.23 ;
      RECT 68.835 1.42 69.005 1.59 ;
      RECT 68.835 4.14 69.005 4.31 ;
      RECT 68.58 2.78 68.75 2.95 ;
      RECT 68.375 1.42 68.545 1.59 ;
      RECT 68.375 4.14 68.545 4.31 ;
      RECT 68.34 1.94 68.51 2.11 ;
      RECT 68.1 2.5 68.27 2.67 ;
      RECT 68.1 4.55 68.27 4.72 ;
      RECT 68.1 8.61 68.27 8.78 ;
      RECT 67.915 1.42 68.085 1.59 ;
      RECT 67.915 4.14 68.085 4.31 ;
      RECT 67.89 3.34 68.06 3.51 ;
      RECT 67.79 6.69 67.96 6.86 ;
      RECT 67.62 2.78 67.79 2.95 ;
      RECT 67.455 1.42 67.625 1.59 ;
      RECT 67.455 4.14 67.625 4.31 ;
      RECT 67.42 8.61 67.59 8.78 ;
      RECT 67.36 7.06 67.53 7.23 ;
      RECT 67.36 7.8 67.53 7.97 ;
      RECT 67.35 3.62 67.52 3.79 ;
      RECT 67.14 2.2 67.31 2.37 ;
      RECT 66.995 1.42 67.165 1.59 ;
      RECT 66.995 4.14 67.165 4.31 ;
      RECT 66.985 6.32 67.155 6.49 ;
      RECT 66.74 8.61 66.91 8.78 ;
      RECT 66.66 2.78 66.83 2.95 ;
      RECT 66.535 1.42 66.705 1.59 ;
      RECT 66.535 4.14 66.705 4.31 ;
      RECT 66.42 1.94 66.59 2.11 ;
      RECT 66.18 2.5 66.35 2.67 ;
      RECT 66.18 3.06 66.35 3.23 ;
      RECT 66.075 1.42 66.245 1.59 ;
      RECT 66.075 4.14 66.245 4.31 ;
      RECT 66.06 8.61 66.23 8.78 ;
      RECT 65.99 5.95 66.16 6.12 ;
      RECT 65.7 2.5 65.87 2.67 ;
      RECT 65.615 1.42 65.785 1.59 ;
      RECT 65.615 4.14 65.785 4.31 ;
      RECT 65.46 3.62 65.63 3.79 ;
      RECT 65.42 1.94 65.59 2.11 ;
      RECT 65.22 2.78 65.39 2.95 ;
      RECT 65.155 1.42 65.325 1.59 ;
      RECT 65.155 4.14 65.325 4.31 ;
      RECT 64.98 3.62 65.15 3.79 ;
      RECT 64.74 3.06 64.91 3.23 ;
      RECT 64.695 1.42 64.865 1.59 ;
      RECT 64.695 4.14 64.865 4.31 ;
      RECT 64.26 2.5 64.43 2.67 ;
      RECT 64.235 1.42 64.405 1.59 ;
      RECT 64.235 4.14 64.405 4.31 ;
      RECT 64.02 1.94 64.19 2.11 ;
      RECT 64.02 3.62 64.19 3.79 ;
      RECT 63.775 1.42 63.945 1.59 ;
      RECT 63.775 4.14 63.945 4.31 ;
      RECT 63.54 1.94 63.71 2.11 ;
      RECT 63.54 3.06 63.71 3.23 ;
      RECT 63.315 1.42 63.485 1.59 ;
      RECT 63.315 4.14 63.485 4.31 ;
      RECT 63.3 2.5 63.47 2.67 ;
      RECT 63.06 3.34 63.23 3.51 ;
      RECT 62.855 1.42 63.025 1.59 ;
      RECT 62.855 4.14 63.025 4.31 ;
      RECT 62.82 2.78 62.99 2.95 ;
      RECT 62.395 1.42 62.565 1.59 ;
      RECT 62.395 4.14 62.565 4.31 ;
      RECT 62.34 2.78 62.51 2.95 ;
      RECT 62.13 1.94 62.3 2.11 ;
      RECT 62.13 3.34 62.3 3.51 ;
      RECT 61.935 1.42 62.105 1.59 ;
      RECT 61.935 4.14 62.105 4.31 ;
      RECT 60.5 0.92 60.67 1.09 ;
      RECT 60.5 2.4 60.67 2.57 ;
      RECT 60.5 6.32 60.67 6.49 ;
      RECT 60.5 7.8 60.67 7.97 ;
      RECT 60.15 0.11 60.32 0.28 ;
      RECT 60.15 4.17 60.32 4.34 ;
      RECT 60.15 4.55 60.32 4.72 ;
      RECT 60.15 8.61 60.32 8.78 ;
      RECT 60.13 2.77 60.3 2.94 ;
      RECT 60.13 5.95 60.3 6.12 ;
      RECT 59.51 0.92 59.68 1.09 ;
      RECT 59.51 2.4 59.68 2.57 ;
      RECT 59.51 6.32 59.68 6.49 ;
      RECT 59.51 7.8 59.68 7.97 ;
      RECT 59.16 0.11 59.33 0.28 ;
      RECT 59.16 4.17 59.33 4.34 ;
      RECT 59.16 4.55 59.33 4.72 ;
      RECT 59.16 8.61 59.33 8.78 ;
      RECT 59.14 2.77 59.31 2.94 ;
      RECT 59.14 5.95 59.31 6.12 ;
      RECT 58.455 0.11 58.625 0.28 ;
      RECT 58.455 4.17 58.625 4.34 ;
      RECT 58.455 4.55 58.625 4.72 ;
      RECT 58.455 8.61 58.625 8.78 ;
      RECT 58.145 2.03 58.315 2.2 ;
      RECT 58.145 6.69 58.315 6.86 ;
      RECT 57.775 0.11 57.945 0.28 ;
      RECT 57.775 8.61 57.945 8.78 ;
      RECT 57.715 0.92 57.885 1.09 ;
      RECT 57.715 1.66 57.885 1.83 ;
      RECT 57.715 7.06 57.885 7.23 ;
      RECT 57.715 7.8 57.885 7.97 ;
      RECT 57.34 2.4 57.51 2.57 ;
      RECT 57.34 6.32 57.51 6.49 ;
      RECT 57.095 0.11 57.265 0.28 ;
      RECT 57.095 8.61 57.265 8.78 ;
      RECT 56.415 0.11 56.585 0.28 ;
      RECT 56.415 8.61 56.585 8.78 ;
      RECT 56.345 2.77 56.515 2.94 ;
      RECT 56.345 5.95 56.515 6.12 ;
      RECT 54.955 1.42 55.125 1.59 ;
      RECT 54.955 4.14 55.125 4.31 ;
      RECT 54.495 1.42 54.665 1.59 ;
      RECT 54.495 4.14 54.665 4.31 ;
      RECT 54.28 2.78 54.45 2.95 ;
      RECT 54.04 1.94 54.21 2.11 ;
      RECT 54.04 3.62 54.21 3.79 ;
      RECT 54.035 1.42 54.205 1.59 ;
      RECT 54.035 4.14 54.205 4.31 ;
      RECT 53.8 2.5 53.97 2.67 ;
      RECT 53.8 3.06 53.97 3.23 ;
      RECT 53.575 1.42 53.745 1.59 ;
      RECT 53.575 4.14 53.745 4.31 ;
      RECT 53.32 2.78 53.49 2.95 ;
      RECT 53.115 1.42 53.285 1.59 ;
      RECT 53.115 4.14 53.285 4.31 ;
      RECT 53.08 1.94 53.25 2.11 ;
      RECT 52.84 2.5 53.01 2.67 ;
      RECT 52.84 4.55 53.01 4.72 ;
      RECT 52.84 8.61 53.01 8.78 ;
      RECT 52.655 1.42 52.825 1.59 ;
      RECT 52.655 4.14 52.825 4.31 ;
      RECT 52.63 3.34 52.8 3.51 ;
      RECT 52.53 6.69 52.7 6.86 ;
      RECT 52.36 2.78 52.53 2.95 ;
      RECT 52.195 1.42 52.365 1.59 ;
      RECT 52.195 4.14 52.365 4.31 ;
      RECT 52.16 8.61 52.33 8.78 ;
      RECT 52.1 7.06 52.27 7.23 ;
      RECT 52.1 7.8 52.27 7.97 ;
      RECT 52.09 3.62 52.26 3.79 ;
      RECT 51.88 2.2 52.05 2.37 ;
      RECT 51.735 1.42 51.905 1.59 ;
      RECT 51.735 4.14 51.905 4.31 ;
      RECT 51.725 6.32 51.895 6.49 ;
      RECT 51.48 8.61 51.65 8.78 ;
      RECT 51.4 2.78 51.57 2.95 ;
      RECT 51.275 1.42 51.445 1.59 ;
      RECT 51.275 4.14 51.445 4.31 ;
      RECT 51.16 1.94 51.33 2.11 ;
      RECT 50.92 2.5 51.09 2.67 ;
      RECT 50.92 3.06 51.09 3.23 ;
      RECT 50.815 1.42 50.985 1.59 ;
      RECT 50.815 4.14 50.985 4.31 ;
      RECT 50.8 8.61 50.97 8.78 ;
      RECT 50.73 5.95 50.9 6.12 ;
      RECT 50.44 2.5 50.61 2.67 ;
      RECT 50.355 1.42 50.525 1.59 ;
      RECT 50.355 4.14 50.525 4.31 ;
      RECT 50.2 3.62 50.37 3.79 ;
      RECT 50.16 1.94 50.33 2.11 ;
      RECT 49.96 2.78 50.13 2.95 ;
      RECT 49.895 1.42 50.065 1.59 ;
      RECT 49.895 4.14 50.065 4.31 ;
      RECT 49.72 3.62 49.89 3.79 ;
      RECT 49.48 3.06 49.65 3.23 ;
      RECT 49.435 1.42 49.605 1.59 ;
      RECT 49.435 4.14 49.605 4.31 ;
      RECT 49 2.5 49.17 2.67 ;
      RECT 48.975 1.42 49.145 1.59 ;
      RECT 48.975 4.14 49.145 4.31 ;
      RECT 48.76 1.94 48.93 2.11 ;
      RECT 48.76 3.62 48.93 3.79 ;
      RECT 48.515 1.42 48.685 1.59 ;
      RECT 48.515 4.14 48.685 4.31 ;
      RECT 48.28 1.94 48.45 2.11 ;
      RECT 48.28 3.06 48.45 3.23 ;
      RECT 48.055 1.42 48.225 1.59 ;
      RECT 48.055 4.14 48.225 4.31 ;
      RECT 48.04 2.5 48.21 2.67 ;
      RECT 47.8 3.34 47.97 3.51 ;
      RECT 47.595 1.42 47.765 1.59 ;
      RECT 47.595 4.14 47.765 4.31 ;
      RECT 47.56 2.78 47.73 2.95 ;
      RECT 47.135 1.42 47.305 1.59 ;
      RECT 47.135 4.14 47.305 4.31 ;
      RECT 47.08 2.78 47.25 2.95 ;
      RECT 46.87 1.94 47.04 2.11 ;
      RECT 46.87 3.34 47.04 3.51 ;
      RECT 46.675 1.42 46.845 1.59 ;
      RECT 46.675 4.14 46.845 4.31 ;
      RECT 45.24 0.92 45.41 1.09 ;
      RECT 45.24 2.4 45.41 2.57 ;
      RECT 45.24 6.32 45.41 6.49 ;
      RECT 45.24 7.8 45.41 7.97 ;
      RECT 44.89 0.11 45.06 0.28 ;
      RECT 44.89 4.17 45.06 4.34 ;
      RECT 44.89 4.55 45.06 4.72 ;
      RECT 44.89 8.61 45.06 8.78 ;
      RECT 44.87 2.77 45.04 2.94 ;
      RECT 44.87 5.95 45.04 6.12 ;
      RECT 44.25 0.92 44.42 1.09 ;
      RECT 44.25 2.4 44.42 2.57 ;
      RECT 44.25 6.32 44.42 6.49 ;
      RECT 44.25 7.8 44.42 7.97 ;
      RECT 43.9 0.11 44.07 0.28 ;
      RECT 43.9 4.17 44.07 4.34 ;
      RECT 43.9 4.55 44.07 4.72 ;
      RECT 43.9 8.61 44.07 8.78 ;
      RECT 43.88 2.77 44.05 2.94 ;
      RECT 43.88 5.95 44.05 6.12 ;
      RECT 43.195 0.11 43.365 0.28 ;
      RECT 43.195 4.17 43.365 4.34 ;
      RECT 43.195 4.55 43.365 4.72 ;
      RECT 43.195 8.61 43.365 8.78 ;
      RECT 42.885 2.03 43.055 2.2 ;
      RECT 42.885 6.69 43.055 6.86 ;
      RECT 42.515 0.11 42.685 0.28 ;
      RECT 42.515 8.61 42.685 8.78 ;
      RECT 42.455 0.92 42.625 1.09 ;
      RECT 42.455 1.66 42.625 1.83 ;
      RECT 42.455 7.06 42.625 7.23 ;
      RECT 42.455 7.8 42.625 7.97 ;
      RECT 42.08 2.4 42.25 2.57 ;
      RECT 42.08 6.32 42.25 6.49 ;
      RECT 41.835 0.11 42.005 0.28 ;
      RECT 41.835 8.61 42.005 8.78 ;
      RECT 41.155 0.11 41.325 0.28 ;
      RECT 41.155 8.61 41.325 8.78 ;
      RECT 41.085 2.77 41.255 2.94 ;
      RECT 41.085 5.95 41.255 6.12 ;
      RECT 39.695 1.42 39.865 1.59 ;
      RECT 39.695 4.14 39.865 4.31 ;
      RECT 39.235 1.42 39.405 1.59 ;
      RECT 39.235 4.14 39.405 4.31 ;
      RECT 39.02 2.78 39.19 2.95 ;
      RECT 38.78 1.94 38.95 2.11 ;
      RECT 38.78 3.62 38.95 3.79 ;
      RECT 38.775 1.42 38.945 1.59 ;
      RECT 38.775 4.14 38.945 4.31 ;
      RECT 38.54 2.5 38.71 2.67 ;
      RECT 38.54 3.06 38.71 3.23 ;
      RECT 38.315 1.42 38.485 1.59 ;
      RECT 38.315 4.14 38.485 4.31 ;
      RECT 38.06 2.78 38.23 2.95 ;
      RECT 37.855 1.42 38.025 1.59 ;
      RECT 37.855 4.14 38.025 4.31 ;
      RECT 37.82 1.94 37.99 2.11 ;
      RECT 37.58 2.5 37.75 2.67 ;
      RECT 37.58 4.55 37.75 4.72 ;
      RECT 37.58 8.61 37.75 8.78 ;
      RECT 37.395 1.42 37.565 1.59 ;
      RECT 37.395 4.14 37.565 4.31 ;
      RECT 37.37 3.34 37.54 3.51 ;
      RECT 37.27 6.69 37.44 6.86 ;
      RECT 37.1 2.78 37.27 2.95 ;
      RECT 36.935 1.42 37.105 1.59 ;
      RECT 36.935 4.14 37.105 4.31 ;
      RECT 36.9 8.61 37.07 8.78 ;
      RECT 36.84 7.06 37.01 7.23 ;
      RECT 36.84 7.8 37.01 7.97 ;
      RECT 36.83 3.62 37 3.79 ;
      RECT 36.62 2.2 36.79 2.37 ;
      RECT 36.475 1.42 36.645 1.59 ;
      RECT 36.475 4.14 36.645 4.31 ;
      RECT 36.465 6.32 36.635 6.49 ;
      RECT 36.22 8.61 36.39 8.78 ;
      RECT 36.14 2.78 36.31 2.95 ;
      RECT 36.015 1.42 36.185 1.59 ;
      RECT 36.015 4.14 36.185 4.31 ;
      RECT 35.9 1.94 36.07 2.11 ;
      RECT 35.66 2.5 35.83 2.67 ;
      RECT 35.66 3.06 35.83 3.23 ;
      RECT 35.555 1.42 35.725 1.59 ;
      RECT 35.555 4.14 35.725 4.31 ;
      RECT 35.54 8.61 35.71 8.78 ;
      RECT 35.47 5.95 35.64 6.12 ;
      RECT 35.18 2.5 35.35 2.67 ;
      RECT 35.095 1.42 35.265 1.59 ;
      RECT 35.095 4.14 35.265 4.31 ;
      RECT 34.94 3.62 35.11 3.79 ;
      RECT 34.9 1.94 35.07 2.11 ;
      RECT 34.7 2.78 34.87 2.95 ;
      RECT 34.635 1.42 34.805 1.59 ;
      RECT 34.635 4.14 34.805 4.31 ;
      RECT 34.46 3.62 34.63 3.79 ;
      RECT 34.22 3.06 34.39 3.23 ;
      RECT 34.175 1.42 34.345 1.59 ;
      RECT 34.175 4.14 34.345 4.31 ;
      RECT 33.74 2.5 33.91 2.67 ;
      RECT 33.715 1.42 33.885 1.59 ;
      RECT 33.715 4.14 33.885 4.31 ;
      RECT 33.5 1.94 33.67 2.11 ;
      RECT 33.5 3.62 33.67 3.79 ;
      RECT 33.255 1.42 33.425 1.59 ;
      RECT 33.255 4.14 33.425 4.31 ;
      RECT 33.02 1.94 33.19 2.11 ;
      RECT 33.02 3.06 33.19 3.23 ;
      RECT 32.795 1.42 32.965 1.59 ;
      RECT 32.795 4.14 32.965 4.31 ;
      RECT 32.78 2.5 32.95 2.67 ;
      RECT 32.54 3.34 32.71 3.51 ;
      RECT 32.335 1.42 32.505 1.59 ;
      RECT 32.335 4.14 32.505 4.31 ;
      RECT 32.3 2.78 32.47 2.95 ;
      RECT 31.875 1.42 32.045 1.59 ;
      RECT 31.875 4.14 32.045 4.31 ;
      RECT 31.82 2.78 31.99 2.95 ;
      RECT 31.61 1.94 31.78 2.11 ;
      RECT 31.61 3.34 31.78 3.51 ;
      RECT 31.415 1.42 31.585 1.59 ;
      RECT 31.415 4.14 31.585 4.31 ;
      RECT 29.98 0.92 30.15 1.09 ;
      RECT 29.98 2.4 30.15 2.57 ;
      RECT 29.98 6.32 30.15 6.49 ;
      RECT 29.98 7.8 30.15 7.97 ;
      RECT 29.63 0.11 29.8 0.28 ;
      RECT 29.63 4.17 29.8 4.34 ;
      RECT 29.63 4.55 29.8 4.72 ;
      RECT 29.63 8.61 29.8 8.78 ;
      RECT 29.61 2.77 29.78 2.94 ;
      RECT 29.61 5.95 29.78 6.12 ;
      RECT 28.99 0.92 29.16 1.09 ;
      RECT 28.99 2.4 29.16 2.57 ;
      RECT 28.99 6.32 29.16 6.49 ;
      RECT 28.99 7.8 29.16 7.97 ;
      RECT 28.64 0.11 28.81 0.28 ;
      RECT 28.64 4.17 28.81 4.34 ;
      RECT 28.64 4.55 28.81 4.72 ;
      RECT 28.64 8.61 28.81 8.78 ;
      RECT 28.62 2.77 28.79 2.94 ;
      RECT 28.62 5.95 28.79 6.12 ;
      RECT 27.935 0.11 28.105 0.28 ;
      RECT 27.935 4.17 28.105 4.34 ;
      RECT 27.935 4.55 28.105 4.72 ;
      RECT 27.935 8.61 28.105 8.78 ;
      RECT 27.625 2.03 27.795 2.2 ;
      RECT 27.625 6.69 27.795 6.86 ;
      RECT 27.255 0.11 27.425 0.28 ;
      RECT 27.255 8.61 27.425 8.78 ;
      RECT 27.195 0.92 27.365 1.09 ;
      RECT 27.195 1.66 27.365 1.83 ;
      RECT 27.195 7.06 27.365 7.23 ;
      RECT 27.195 7.8 27.365 7.97 ;
      RECT 26.82 2.4 26.99 2.57 ;
      RECT 26.82 6.32 26.99 6.49 ;
      RECT 26.575 0.11 26.745 0.28 ;
      RECT 26.575 8.61 26.745 8.78 ;
      RECT 25.895 0.11 26.065 0.28 ;
      RECT 25.895 8.61 26.065 8.78 ;
      RECT 25.825 2.77 25.995 2.94 ;
      RECT 25.825 5.95 25.995 6.12 ;
      RECT 24.435 1.42 24.605 1.59 ;
      RECT 24.435 4.14 24.605 4.31 ;
      RECT 23.975 1.42 24.145 1.59 ;
      RECT 23.975 4.14 24.145 4.31 ;
      RECT 23.76 2.78 23.93 2.95 ;
      RECT 23.52 1.94 23.69 2.11 ;
      RECT 23.52 3.62 23.69 3.79 ;
      RECT 23.515 1.42 23.685 1.59 ;
      RECT 23.515 4.14 23.685 4.31 ;
      RECT 23.28 2.5 23.45 2.67 ;
      RECT 23.28 3.06 23.45 3.23 ;
      RECT 23.055 1.42 23.225 1.59 ;
      RECT 23.055 4.14 23.225 4.31 ;
      RECT 22.8 2.78 22.97 2.95 ;
      RECT 22.595 1.42 22.765 1.59 ;
      RECT 22.595 4.14 22.765 4.31 ;
      RECT 22.56 1.94 22.73 2.11 ;
      RECT 22.32 2.5 22.49 2.67 ;
      RECT 22.32 4.55 22.49 4.72 ;
      RECT 22.32 8.61 22.49 8.78 ;
      RECT 22.135 1.42 22.305 1.59 ;
      RECT 22.135 4.14 22.305 4.31 ;
      RECT 22.11 3.34 22.28 3.51 ;
      RECT 22.01 6.69 22.18 6.86 ;
      RECT 21.84 2.78 22.01 2.95 ;
      RECT 21.675 1.42 21.845 1.59 ;
      RECT 21.675 4.14 21.845 4.31 ;
      RECT 21.64 8.61 21.81 8.78 ;
      RECT 21.58 7.06 21.75 7.23 ;
      RECT 21.58 7.8 21.75 7.97 ;
      RECT 21.57 3.62 21.74 3.79 ;
      RECT 21.36 2.2 21.53 2.37 ;
      RECT 21.215 1.42 21.385 1.59 ;
      RECT 21.215 4.14 21.385 4.31 ;
      RECT 21.205 6.32 21.375 6.49 ;
      RECT 20.96 8.61 21.13 8.78 ;
      RECT 20.88 2.78 21.05 2.95 ;
      RECT 20.755 1.42 20.925 1.59 ;
      RECT 20.755 4.14 20.925 4.31 ;
      RECT 20.64 1.94 20.81 2.11 ;
      RECT 20.4 2.5 20.57 2.67 ;
      RECT 20.4 3.06 20.57 3.23 ;
      RECT 20.295 1.42 20.465 1.59 ;
      RECT 20.295 4.14 20.465 4.31 ;
      RECT 20.28 8.61 20.45 8.78 ;
      RECT 20.21 5.95 20.38 6.12 ;
      RECT 19.92 2.5 20.09 2.67 ;
      RECT 19.835 1.42 20.005 1.59 ;
      RECT 19.835 4.14 20.005 4.31 ;
      RECT 19.68 3.62 19.85 3.79 ;
      RECT 19.64 1.94 19.81 2.11 ;
      RECT 19.44 2.78 19.61 2.95 ;
      RECT 19.375 1.42 19.545 1.59 ;
      RECT 19.375 4.14 19.545 4.31 ;
      RECT 19.2 3.62 19.37 3.79 ;
      RECT 18.96 3.06 19.13 3.23 ;
      RECT 18.915 1.42 19.085 1.59 ;
      RECT 18.915 4.14 19.085 4.31 ;
      RECT 18.48 2.5 18.65 2.67 ;
      RECT 18.455 1.42 18.625 1.59 ;
      RECT 18.455 4.14 18.625 4.31 ;
      RECT 18.24 1.94 18.41 2.11 ;
      RECT 18.24 3.62 18.41 3.79 ;
      RECT 17.995 1.42 18.165 1.59 ;
      RECT 17.995 4.14 18.165 4.31 ;
      RECT 17.76 1.94 17.93 2.11 ;
      RECT 17.76 3.06 17.93 3.23 ;
      RECT 17.535 1.42 17.705 1.59 ;
      RECT 17.535 4.14 17.705 4.31 ;
      RECT 17.52 2.5 17.69 2.67 ;
      RECT 17.28 3.34 17.45 3.51 ;
      RECT 17.075 1.42 17.245 1.59 ;
      RECT 17.075 4.14 17.245 4.31 ;
      RECT 17.04 2.78 17.21 2.95 ;
      RECT 16.615 1.42 16.785 1.59 ;
      RECT 16.615 4.14 16.785 4.31 ;
      RECT 16.56 2.78 16.73 2.95 ;
      RECT 16.35 1.94 16.52 2.11 ;
      RECT 16.35 3.34 16.52 3.51 ;
      RECT 16.155 1.42 16.325 1.59 ;
      RECT 16.155 4.14 16.325 4.31 ;
      RECT 14.72 0.92 14.89 1.09 ;
      RECT 14.72 2.4 14.89 2.57 ;
      RECT 14.72 6.32 14.89 6.49 ;
      RECT 14.72 7.8 14.89 7.97 ;
      RECT 14.37 0.11 14.54 0.28 ;
      RECT 14.37 4.17 14.54 4.34 ;
      RECT 14.37 4.55 14.54 4.72 ;
      RECT 14.37 8.61 14.54 8.78 ;
      RECT 14.35 2.77 14.52 2.94 ;
      RECT 14.35 5.95 14.52 6.12 ;
      RECT 13.73 0.92 13.9 1.09 ;
      RECT 13.73 2.4 13.9 2.57 ;
      RECT 13.73 6.32 13.9 6.49 ;
      RECT 13.73 7.8 13.9 7.97 ;
      RECT 13.38 0.11 13.55 0.28 ;
      RECT 13.38 4.17 13.55 4.34 ;
      RECT 13.38 4.55 13.55 4.72 ;
      RECT 13.38 8.61 13.55 8.78 ;
      RECT 13.36 2.77 13.53 2.94 ;
      RECT 13.36 5.95 13.53 6.12 ;
      RECT 12.675 0.11 12.845 0.28 ;
      RECT 12.675 4.17 12.845 4.34 ;
      RECT 12.675 4.55 12.845 4.72 ;
      RECT 12.675 8.61 12.845 8.78 ;
      RECT 12.365 2.03 12.535 2.2 ;
      RECT 12.365 6.69 12.535 6.86 ;
      RECT 11.995 0.11 12.165 0.28 ;
      RECT 11.995 8.61 12.165 8.78 ;
      RECT 11.935 0.92 12.105 1.09 ;
      RECT 11.935 1.66 12.105 1.83 ;
      RECT 11.935 7.06 12.105 7.23 ;
      RECT 11.935 7.8 12.105 7.97 ;
      RECT 11.56 2.4 11.73 2.57 ;
      RECT 11.56 6.32 11.73 6.49 ;
      RECT 11.315 0.11 11.485 0.28 ;
      RECT 11.315 8.61 11.485 8.78 ;
      RECT 10.635 0.11 10.805 0.28 ;
      RECT 10.635 8.61 10.805 8.78 ;
      RECT 10.565 2.77 10.735 2.94 ;
      RECT 10.565 5.95 10.735 6.12 ;
      RECT 9.175 1.42 9.345 1.59 ;
      RECT 9.175 4.14 9.345 4.31 ;
      RECT 8.715 1.42 8.885 1.59 ;
      RECT 8.715 4.14 8.885 4.31 ;
      RECT 8.5 2.78 8.67 2.95 ;
      RECT 8.26 1.94 8.43 2.11 ;
      RECT 8.26 3.62 8.43 3.79 ;
      RECT 8.255 1.42 8.425 1.59 ;
      RECT 8.255 4.14 8.425 4.31 ;
      RECT 8.02 2.5 8.19 2.67 ;
      RECT 8.02 3.06 8.19 3.23 ;
      RECT 7.795 1.42 7.965 1.59 ;
      RECT 7.795 4.14 7.965 4.31 ;
      RECT 7.54 2.78 7.71 2.95 ;
      RECT 7.335 1.42 7.505 1.59 ;
      RECT 7.335 4.14 7.505 4.31 ;
      RECT 7.3 1.94 7.47 2.11 ;
      RECT 7.06 2.5 7.23 2.67 ;
      RECT 7.06 4.55 7.23 4.72 ;
      RECT 7.06 8.61 7.23 8.78 ;
      RECT 6.875 1.42 7.045 1.59 ;
      RECT 6.875 4.14 7.045 4.31 ;
      RECT 6.85 3.34 7.02 3.51 ;
      RECT 6.75 6.69 6.92 6.86 ;
      RECT 6.58 2.78 6.75 2.95 ;
      RECT 6.415 1.42 6.585 1.59 ;
      RECT 6.415 4.14 6.585 4.31 ;
      RECT 6.38 8.61 6.55 8.78 ;
      RECT 6.32 7.06 6.49 7.23 ;
      RECT 6.32 7.8 6.49 7.97 ;
      RECT 6.31 3.62 6.48 3.79 ;
      RECT 6.1 2.2 6.27 2.37 ;
      RECT 5.955 1.42 6.125 1.59 ;
      RECT 5.955 4.14 6.125 4.31 ;
      RECT 5.945 6.32 6.115 6.49 ;
      RECT 5.7 8.61 5.87 8.78 ;
      RECT 5.62 2.78 5.79 2.95 ;
      RECT 5.495 1.42 5.665 1.59 ;
      RECT 5.495 4.14 5.665 4.31 ;
      RECT 5.38 1.94 5.55 2.11 ;
      RECT 5.14 2.5 5.31 2.67 ;
      RECT 5.14 3.06 5.31 3.23 ;
      RECT 5.035 1.42 5.205 1.59 ;
      RECT 5.035 4.14 5.205 4.31 ;
      RECT 5.02 8.61 5.19 8.78 ;
      RECT 4.95 5.95 5.12 6.12 ;
      RECT 4.66 2.5 4.83 2.67 ;
      RECT 4.575 1.42 4.745 1.59 ;
      RECT 4.575 4.14 4.745 4.31 ;
      RECT 4.42 3.62 4.59 3.79 ;
      RECT 4.38 1.94 4.55 2.11 ;
      RECT 4.18 2.78 4.35 2.95 ;
      RECT 4.115 1.42 4.285 1.59 ;
      RECT 4.115 4.14 4.285 4.31 ;
      RECT 3.94 3.62 4.11 3.79 ;
      RECT 3.7 3.06 3.87 3.23 ;
      RECT 3.655 1.42 3.825 1.59 ;
      RECT 3.655 4.14 3.825 4.31 ;
      RECT 3.22 2.5 3.39 2.67 ;
      RECT 3.195 1.42 3.365 1.59 ;
      RECT 3.195 4.14 3.365 4.31 ;
      RECT 2.98 1.94 3.15 2.11 ;
      RECT 2.98 3.62 3.15 3.79 ;
      RECT 2.735 1.42 2.905 1.59 ;
      RECT 2.735 4.14 2.905 4.31 ;
      RECT 2.5 1.94 2.67 2.11 ;
      RECT 2.5 3.06 2.67 3.23 ;
      RECT 2.275 1.42 2.445 1.59 ;
      RECT 2.275 4.14 2.445 4.31 ;
      RECT 2.26 2.5 2.43 2.67 ;
      RECT 2.02 3.34 2.19 3.51 ;
      RECT 1.815 1.42 1.985 1.59 ;
      RECT 1.815 4.14 1.985 4.31 ;
      RECT 1.78 2.78 1.95 2.95 ;
      RECT 1.355 1.42 1.525 1.59 ;
      RECT 1.355 4.14 1.525 4.31 ;
      RECT 1.3 2.78 1.47 2.95 ;
      RECT 1.09 1.94 1.26 2.11 ;
      RECT 1.09 3.34 1.26 3.51 ;
      RECT 0.895 1.42 1.065 1.59 ;
      RECT 0.895 4.14 1.065 4.31 ;
      RECT -0.455 4.55 -0.285 4.72 ;
      RECT -0.455 8.61 -0.285 8.78 ;
      RECT -0.765 6.69 -0.595 6.86 ;
      RECT -1.135 8.61 -0.965 8.78 ;
      RECT -1.195 7.06 -1.025 7.23 ;
      RECT -1.195 7.8 -1.025 7.97 ;
      RECT -1.57 6.32 -1.4 6.49 ;
      RECT -1.815 8.61 -1.645 8.78 ;
      RECT -2.495 8.61 -2.325 8.78 ;
      RECT -2.565 5.95 -2.395 6.12 ;
    LAYER li ;
      RECT 69.76 0.005 69.93 2.09 ;
      RECT 68.82 0.005 68.99 2.09 ;
      RECT 67.86 0.005 68.03 2.09 ;
      RECT 65.94 0.005 66.11 2.09 ;
      RECT 64.98 0.005 65.15 2.09 ;
      RECT 63.06 0.005 63.23 2.09 ;
      RECT 54.5 0.005 54.67 2.09 ;
      RECT 53.56 0.005 53.73 2.09 ;
      RECT 52.6 0.005 52.77 2.09 ;
      RECT 50.68 0.005 50.85 2.09 ;
      RECT 49.72 0.005 49.89 2.09 ;
      RECT 47.8 0.005 47.97 2.09 ;
      RECT 39.24 0.005 39.41 2.09 ;
      RECT 38.3 0.005 38.47 2.09 ;
      RECT 37.34 0.005 37.51 2.09 ;
      RECT 35.42 0.005 35.59 2.09 ;
      RECT 34.46 0.005 34.63 2.09 ;
      RECT 32.54 0.005 32.71 2.09 ;
      RECT 23.98 0.005 24.15 2.09 ;
      RECT 23.04 0.005 23.21 2.09 ;
      RECT 22.08 0.005 22.25 2.09 ;
      RECT 20.16 0.005 20.33 2.09 ;
      RECT 19.2 0.005 19.37 2.09 ;
      RECT 17.28 0.005 17.45 2.09 ;
      RECT 8.72 0.005 8.89 2.09 ;
      RECT 7.78 0.005 7.95 2.09 ;
      RECT 6.82 0.005 6.99 2.09 ;
      RECT 4.9 0.005 5.07 2.09 ;
      RECT 3.94 0.005 4.11 2.09 ;
      RECT 2.02 0.005 2.19 2.09 ;
      RECT 66.815 0.005 67.01 1.6 ;
      RECT 63.06 0.005 63.335 1.6 ;
      RECT 51.555 0.005 51.75 1.6 ;
      RECT 47.8 0.005 48.075 1.6 ;
      RECT 36.295 0.005 36.49 1.6 ;
      RECT 32.54 0.005 32.815 1.6 ;
      RECT 21.035 0.005 21.23 1.6 ;
      RECT 17.28 0.005 17.555 1.6 ;
      RECT 5.775 0.005 5.97 1.6 ;
      RECT 2.02 0.005 2.295 1.6 ;
      RECT 61.79 0.005 70.53 1.59 ;
      RECT 46.53 0.005 55.27 1.59 ;
      RECT 31.27 0.005 40.01 1.59 ;
      RECT 16.01 0.005 24.75 1.59 ;
      RECT 0.75 0.005 9.49 1.59 ;
      RECT 75.33 0.005 75.5 0.94 ;
      RECT 74.34 0.005 74.51 0.94 ;
      RECT 71.595 0.005 71.765 0.94 ;
      RECT 60.07 0.005 60.24 0.94 ;
      RECT 59.08 0.005 59.25 0.94 ;
      RECT 56.335 0.005 56.505 0.94 ;
      RECT 44.81 0.005 44.98 0.94 ;
      RECT 43.82 0.005 43.99 0.94 ;
      RECT 41.075 0.005 41.245 0.94 ;
      RECT 29.55 0.005 29.72 0.94 ;
      RECT 28.56 0.005 28.73 0.94 ;
      RECT 25.815 0.005 25.985 0.94 ;
      RECT 14.29 0.005 14.46 0.94 ;
      RECT 13.3 0.005 13.47 0.94 ;
      RECT 10.555 0.005 10.725 0.94 ;
      RECT -2.75 0.005 76.3 0.31 ;
      RECT -0.765 4.145 -0.595 8.31 ;
      RECT 75.33 3.41 75.5 5.48 ;
      RECT 74.34 3.41 74.51 5.48 ;
      RECT 71.595 3.41 71.765 5.48 ;
      RECT 65.98 4.14 66.15 5.48 ;
      RECT 60.07 3.41 60.24 5.48 ;
      RECT 59.08 3.41 59.25 5.48 ;
      RECT 56.335 3.41 56.505 5.48 ;
      RECT 50.72 4.14 50.89 5.48 ;
      RECT 44.81 3.41 44.98 5.48 ;
      RECT 43.82 3.41 43.99 5.48 ;
      RECT 41.075 3.41 41.245 5.48 ;
      RECT 35.46 4.14 35.63 5.48 ;
      RECT 29.55 3.41 29.72 5.48 ;
      RECT 28.56 3.41 28.73 5.48 ;
      RECT 25.815 3.41 25.985 5.48 ;
      RECT 20.2 4.14 20.37 5.48 ;
      RECT 14.29 3.41 14.46 5.48 ;
      RECT 13.3 3.41 13.47 5.48 ;
      RECT 10.555 3.41 10.725 5.48 ;
      RECT 4.94 4.14 5.11 5.48 ;
      RECT -2.575 4.145 -2.405 5.48 ;
      RECT -2.75 4.145 76.3 4.75 ;
      RECT 61.79 4.14 76.3 4.75 ;
      RECT 46.53 4.14 61.04 4.75 ;
      RECT 31.27 4.14 45.78 4.75 ;
      RECT 16.01 4.14 30.52 4.75 ;
      RECT 0.75 4.14 15.26 4.75 ;
      RECT 68.82 3.64 68.99 4.75 ;
      RECT 66.9 3.64 67.07 4.75 ;
      RECT 65.96 3.64 66.13 4.75 ;
      RECT 64.5 3.64 64.67 4.75 ;
      RECT 62.58 3.64 62.75 4.75 ;
      RECT 53.56 3.64 53.73 4.75 ;
      RECT 51.64 3.64 51.81 4.75 ;
      RECT 50.7 3.64 50.87 4.75 ;
      RECT 49.24 3.64 49.41 4.75 ;
      RECT 47.32 3.64 47.49 4.75 ;
      RECT 38.3 3.64 38.47 4.75 ;
      RECT 36.38 3.64 36.55 4.75 ;
      RECT 35.44 3.64 35.61 4.75 ;
      RECT 33.98 3.64 34.15 4.75 ;
      RECT 32.06 3.64 32.23 4.75 ;
      RECT 23.04 3.64 23.21 4.75 ;
      RECT 21.12 3.64 21.29 4.75 ;
      RECT 20.18 3.64 20.35 4.75 ;
      RECT 18.72 3.64 18.89 4.75 ;
      RECT 16.8 3.64 16.97 4.75 ;
      RECT 7.78 3.64 7.95 4.75 ;
      RECT 5.86 3.64 6.03 4.75 ;
      RECT 4.92 3.64 5.09 4.75 ;
      RECT 3.46 3.64 3.63 4.75 ;
      RECT 1.54 3.64 1.71 4.75 ;
      RECT -2.75 8.58 76.3 8.885 ;
      RECT 75.33 7.95 75.5 8.885 ;
      RECT 74.34 7.95 74.51 8.885 ;
      RECT 71.595 7.95 71.765 8.885 ;
      RECT 65.98 7.95 66.15 8.885 ;
      RECT 60.07 7.95 60.24 8.885 ;
      RECT 59.08 7.95 59.25 8.885 ;
      RECT 56.335 7.95 56.505 8.885 ;
      RECT 50.72 7.95 50.89 8.885 ;
      RECT 44.81 7.95 44.98 8.885 ;
      RECT 43.82 7.95 43.99 8.885 ;
      RECT 41.075 7.95 41.245 8.885 ;
      RECT 35.46 7.95 35.63 8.885 ;
      RECT 29.55 7.95 29.72 8.885 ;
      RECT 28.56 7.95 28.73 8.885 ;
      RECT 25.815 7.95 25.985 8.885 ;
      RECT 20.2 7.95 20.37 8.885 ;
      RECT 14.29 7.95 14.46 8.885 ;
      RECT 13.3 7.95 13.47 8.885 ;
      RECT 10.555 7.95 10.725 8.885 ;
      RECT 4.94 7.95 5.11 8.885 ;
      RECT -2.575 7.95 -2.405 8.885 ;
      RECT 75.39 1.745 75.56 2.94 ;
      RECT 75.39 1.745 75.855 1.915 ;
      RECT 75.39 6.975 75.855 7.145 ;
      RECT 75.39 5.95 75.56 7.145 ;
      RECT 74.4 1.745 74.57 2.94 ;
      RECT 74.4 1.745 74.865 1.915 ;
      RECT 74.4 6.975 74.865 7.145 ;
      RECT 74.4 5.95 74.57 7.145 ;
      RECT 72.545 2.64 72.715 3.87 ;
      RECT 72.6 0.86 72.77 2.81 ;
      RECT 72.545 0.58 72.715 1.03 ;
      RECT 72.545 7.86 72.715 8.31 ;
      RECT 72.6 6.08 72.77 8.03 ;
      RECT 72.545 5.02 72.715 6.25 ;
      RECT 72.025 0.58 72.195 3.87 ;
      RECT 72.025 2.08 72.43 2.41 ;
      RECT 72.025 1.24 72.43 1.57 ;
      RECT 72.025 5.02 72.195 8.31 ;
      RECT 72.025 7.32 72.43 7.65 ;
      RECT 72.025 6.48 72.43 6.81 ;
      RECT 69.3 3.62 69.815 3.79 ;
      RECT 69.645 3.23 69.815 3.79 ;
      RECT 69.75 3.15 69.92 3.48 ;
      RECT 69.54 2.54 69.815 2.95 ;
      RECT 69.42 2.54 69.815 2.75 ;
      RECT 67.89 3.15 68.06 3.51 ;
      RECT 67.89 3.23 69.23 3.4 ;
      RECT 69.06 3.06 69.23 3.4 ;
      RECT 67.62 2.58 67.79 2.95 ;
      RECT 67.14 2.58 67.79 2.85 ;
      RECT 67.06 2.58 67.87 2.75 ;
      RECT 66.42 1.82 66.59 2.11 ;
      RECT 66.42 1.82 67.66 1.99 ;
      RECT 67.14 2.16 67.31 2.37 ;
      RECT 66.78 2.16 67.31 2.33 ;
      RECT 66.93 7.86 67.1 8.31 ;
      RECT 66.985 6.08 67.155 8.03 ;
      RECT 66.93 5.02 67.1 6.25 ;
      RECT 66.41 5.02 66.58 8.31 ;
      RECT 66.41 7.32 66.815 7.65 ;
      RECT 66.41 6.48 66.815 6.81 ;
      RECT 66.18 3.23 66.67 3.4 ;
      RECT 66.18 3.06 66.35 3.4 ;
      RECT 65.46 3.23 65.63 3.79 ;
      RECT 65.35 3.23 65.68 3.4 ;
      RECT 65.42 1.84 65.59 2.11 ;
      RECT 65.46 1.76 65.63 2.09 ;
      RECT 65.325 1.84 65.63 2.06 ;
      RECT 63.9 3.23 64.19 3.79 ;
      RECT 64.02 3.15 64.19 3.79 ;
      RECT 63.66 2.58 64.03 2.75 ;
      RECT 63.66 1.94 63.83 2.75 ;
      RECT 63.54 1.94 63.83 2.11 ;
      RECT 60.13 1.745 60.3 2.94 ;
      RECT 60.13 1.745 60.595 1.915 ;
      RECT 60.13 6.975 60.595 7.145 ;
      RECT 60.13 5.95 60.3 7.145 ;
      RECT 59.14 1.745 59.31 2.94 ;
      RECT 59.14 1.745 59.605 1.915 ;
      RECT 59.14 6.975 59.605 7.145 ;
      RECT 59.14 5.95 59.31 7.145 ;
      RECT 57.285 2.64 57.455 3.87 ;
      RECT 57.34 0.86 57.51 2.81 ;
      RECT 57.285 0.58 57.455 1.03 ;
      RECT 57.285 7.86 57.455 8.31 ;
      RECT 57.34 6.08 57.51 8.03 ;
      RECT 57.285 5.02 57.455 6.25 ;
      RECT 56.765 0.58 56.935 3.87 ;
      RECT 56.765 2.08 57.17 2.41 ;
      RECT 56.765 1.24 57.17 1.57 ;
      RECT 56.765 5.02 56.935 8.31 ;
      RECT 56.765 7.32 57.17 7.65 ;
      RECT 56.765 6.48 57.17 6.81 ;
      RECT 54.04 3.62 54.555 3.79 ;
      RECT 54.385 3.23 54.555 3.79 ;
      RECT 54.49 3.15 54.66 3.48 ;
      RECT 54.28 2.54 54.555 2.95 ;
      RECT 54.16 2.54 54.555 2.75 ;
      RECT 52.63 3.15 52.8 3.51 ;
      RECT 52.63 3.23 53.97 3.4 ;
      RECT 53.8 3.06 53.97 3.4 ;
      RECT 52.36 2.58 52.53 2.95 ;
      RECT 51.88 2.58 52.53 2.85 ;
      RECT 51.8 2.58 52.61 2.75 ;
      RECT 51.16 1.82 51.33 2.11 ;
      RECT 51.16 1.82 52.4 1.99 ;
      RECT 51.88 2.16 52.05 2.37 ;
      RECT 51.52 2.16 52.05 2.33 ;
      RECT 51.67 7.86 51.84 8.31 ;
      RECT 51.725 6.08 51.895 8.03 ;
      RECT 51.67 5.02 51.84 6.25 ;
      RECT 51.15 5.02 51.32 8.31 ;
      RECT 51.15 7.32 51.555 7.65 ;
      RECT 51.15 6.48 51.555 6.81 ;
      RECT 50.92 3.23 51.41 3.4 ;
      RECT 50.92 3.06 51.09 3.4 ;
      RECT 50.2 3.23 50.37 3.79 ;
      RECT 50.09 3.23 50.42 3.4 ;
      RECT 50.16 1.84 50.33 2.11 ;
      RECT 50.2 1.76 50.37 2.09 ;
      RECT 50.065 1.84 50.37 2.06 ;
      RECT 48.64 3.23 48.93 3.79 ;
      RECT 48.76 3.15 48.93 3.79 ;
      RECT 48.4 2.58 48.77 2.75 ;
      RECT 48.4 1.94 48.57 2.75 ;
      RECT 48.28 1.94 48.57 2.11 ;
      RECT 44.87 1.745 45.04 2.94 ;
      RECT 44.87 1.745 45.335 1.915 ;
      RECT 44.87 6.975 45.335 7.145 ;
      RECT 44.87 5.95 45.04 7.145 ;
      RECT 43.88 1.745 44.05 2.94 ;
      RECT 43.88 1.745 44.345 1.915 ;
      RECT 43.88 6.975 44.345 7.145 ;
      RECT 43.88 5.95 44.05 7.145 ;
      RECT 42.025 2.64 42.195 3.87 ;
      RECT 42.08 0.86 42.25 2.81 ;
      RECT 42.025 0.58 42.195 1.03 ;
      RECT 42.025 7.86 42.195 8.31 ;
      RECT 42.08 6.08 42.25 8.03 ;
      RECT 42.025 5.02 42.195 6.25 ;
      RECT 41.505 0.58 41.675 3.87 ;
      RECT 41.505 2.08 41.91 2.41 ;
      RECT 41.505 1.24 41.91 1.57 ;
      RECT 41.505 5.02 41.675 8.31 ;
      RECT 41.505 7.32 41.91 7.65 ;
      RECT 41.505 6.48 41.91 6.81 ;
      RECT 38.78 3.62 39.295 3.79 ;
      RECT 39.125 3.23 39.295 3.79 ;
      RECT 39.23 3.15 39.4 3.48 ;
      RECT 39.02 2.54 39.295 2.95 ;
      RECT 38.9 2.54 39.295 2.75 ;
      RECT 37.37 3.15 37.54 3.51 ;
      RECT 37.37 3.23 38.71 3.4 ;
      RECT 38.54 3.06 38.71 3.4 ;
      RECT 37.1 2.58 37.27 2.95 ;
      RECT 36.62 2.58 37.27 2.85 ;
      RECT 36.54 2.58 37.35 2.75 ;
      RECT 35.9 1.82 36.07 2.11 ;
      RECT 35.9 1.82 37.14 1.99 ;
      RECT 36.62 2.16 36.79 2.37 ;
      RECT 36.26 2.16 36.79 2.33 ;
      RECT 36.41 7.86 36.58 8.31 ;
      RECT 36.465 6.08 36.635 8.03 ;
      RECT 36.41 5.02 36.58 6.25 ;
      RECT 35.89 5.02 36.06 8.31 ;
      RECT 35.89 7.32 36.295 7.65 ;
      RECT 35.89 6.48 36.295 6.81 ;
      RECT 35.66 3.23 36.15 3.4 ;
      RECT 35.66 3.06 35.83 3.4 ;
      RECT 34.94 3.23 35.11 3.79 ;
      RECT 34.83 3.23 35.16 3.4 ;
      RECT 34.9 1.84 35.07 2.11 ;
      RECT 34.94 1.76 35.11 2.09 ;
      RECT 34.805 1.84 35.11 2.06 ;
      RECT 33.38 3.23 33.67 3.79 ;
      RECT 33.5 3.15 33.67 3.79 ;
      RECT 33.14 2.58 33.51 2.75 ;
      RECT 33.14 1.94 33.31 2.75 ;
      RECT 33.02 1.94 33.31 2.11 ;
      RECT 29.61 1.745 29.78 2.94 ;
      RECT 29.61 1.745 30.075 1.915 ;
      RECT 29.61 6.975 30.075 7.145 ;
      RECT 29.61 5.95 29.78 7.145 ;
      RECT 28.62 1.745 28.79 2.94 ;
      RECT 28.62 1.745 29.085 1.915 ;
      RECT 28.62 6.975 29.085 7.145 ;
      RECT 28.62 5.95 28.79 7.145 ;
      RECT 26.765 2.64 26.935 3.87 ;
      RECT 26.82 0.86 26.99 2.81 ;
      RECT 26.765 0.58 26.935 1.03 ;
      RECT 26.765 7.86 26.935 8.31 ;
      RECT 26.82 6.08 26.99 8.03 ;
      RECT 26.765 5.02 26.935 6.25 ;
      RECT 26.245 0.58 26.415 3.87 ;
      RECT 26.245 2.08 26.65 2.41 ;
      RECT 26.245 1.24 26.65 1.57 ;
      RECT 26.245 5.02 26.415 8.31 ;
      RECT 26.245 7.32 26.65 7.65 ;
      RECT 26.245 6.48 26.65 6.81 ;
      RECT 23.52 3.62 24.035 3.79 ;
      RECT 23.865 3.23 24.035 3.79 ;
      RECT 23.97 3.15 24.14 3.48 ;
      RECT 23.76 2.54 24.035 2.95 ;
      RECT 23.64 2.54 24.035 2.75 ;
      RECT 22.11 3.15 22.28 3.51 ;
      RECT 22.11 3.23 23.45 3.4 ;
      RECT 23.28 3.06 23.45 3.4 ;
      RECT 21.84 2.58 22.01 2.95 ;
      RECT 21.36 2.58 22.01 2.85 ;
      RECT 21.28 2.58 22.09 2.75 ;
      RECT 20.64 1.82 20.81 2.11 ;
      RECT 20.64 1.82 21.88 1.99 ;
      RECT 21.36 2.16 21.53 2.37 ;
      RECT 21 2.16 21.53 2.33 ;
      RECT 21.15 7.86 21.32 8.31 ;
      RECT 21.205 6.08 21.375 8.03 ;
      RECT 21.15 5.02 21.32 6.25 ;
      RECT 20.63 5.02 20.8 8.31 ;
      RECT 20.63 7.32 21.035 7.65 ;
      RECT 20.63 6.48 21.035 6.81 ;
      RECT 20.4 3.23 20.89 3.4 ;
      RECT 20.4 3.06 20.57 3.4 ;
      RECT 19.68 3.23 19.85 3.79 ;
      RECT 19.57 3.23 19.9 3.4 ;
      RECT 19.64 1.84 19.81 2.11 ;
      RECT 19.68 1.76 19.85 2.09 ;
      RECT 19.545 1.84 19.85 2.06 ;
      RECT 18.12 3.23 18.41 3.79 ;
      RECT 18.24 3.15 18.41 3.79 ;
      RECT 17.88 2.58 18.25 2.75 ;
      RECT 17.88 1.94 18.05 2.75 ;
      RECT 17.76 1.94 18.05 2.11 ;
      RECT 14.35 1.745 14.52 2.94 ;
      RECT 14.35 1.745 14.815 1.915 ;
      RECT 14.35 6.975 14.815 7.145 ;
      RECT 14.35 5.95 14.52 7.145 ;
      RECT 13.36 1.745 13.53 2.94 ;
      RECT 13.36 1.745 13.825 1.915 ;
      RECT 13.36 6.975 13.825 7.145 ;
      RECT 13.36 5.95 13.53 7.145 ;
      RECT 11.505 2.64 11.675 3.87 ;
      RECT 11.56 0.86 11.73 2.81 ;
      RECT 11.505 0.58 11.675 1.03 ;
      RECT 11.505 7.86 11.675 8.31 ;
      RECT 11.56 6.08 11.73 8.03 ;
      RECT 11.505 5.02 11.675 6.25 ;
      RECT 10.985 0.58 11.155 3.87 ;
      RECT 10.985 2.08 11.39 2.41 ;
      RECT 10.985 1.24 11.39 1.57 ;
      RECT 10.985 5.02 11.155 8.31 ;
      RECT 10.985 7.32 11.39 7.65 ;
      RECT 10.985 6.48 11.39 6.81 ;
      RECT 8.26 3.62 8.775 3.79 ;
      RECT 8.605 3.23 8.775 3.79 ;
      RECT 8.71 3.15 8.88 3.48 ;
      RECT 8.5 2.54 8.775 2.95 ;
      RECT 8.38 2.54 8.775 2.75 ;
      RECT 6.85 3.15 7.02 3.51 ;
      RECT 6.85 3.23 8.19 3.4 ;
      RECT 8.02 3.06 8.19 3.4 ;
      RECT 6.58 2.58 6.75 2.95 ;
      RECT 6.1 2.58 6.75 2.85 ;
      RECT 6.02 2.58 6.83 2.75 ;
      RECT 5.38 1.82 5.55 2.11 ;
      RECT 5.38 1.82 6.62 1.99 ;
      RECT 6.1 2.16 6.27 2.37 ;
      RECT 5.74 2.16 6.27 2.33 ;
      RECT 5.89 7.86 6.06 8.31 ;
      RECT 5.945 6.08 6.115 8.03 ;
      RECT 5.89 5.02 6.06 6.25 ;
      RECT 5.37 5.02 5.54 8.31 ;
      RECT 5.37 7.32 5.775 7.65 ;
      RECT 5.37 6.48 5.775 6.81 ;
      RECT 5.14 3.23 5.63 3.4 ;
      RECT 5.14 3.06 5.31 3.4 ;
      RECT 4.42 3.23 4.59 3.79 ;
      RECT 4.31 3.23 4.64 3.4 ;
      RECT 4.38 1.84 4.55 2.11 ;
      RECT 4.42 1.76 4.59 2.09 ;
      RECT 4.285 1.84 4.59 2.06 ;
      RECT 2.86 3.23 3.15 3.79 ;
      RECT 2.98 3.15 3.15 3.79 ;
      RECT 2.62 2.58 2.99 2.75 ;
      RECT 2.62 1.94 2.79 2.75 ;
      RECT 2.5 1.94 2.79 2.11 ;
      RECT -1.625 7.86 -1.455 8.31 ;
      RECT -1.57 6.08 -1.4 8.03 ;
      RECT -1.625 5.02 -1.455 6.25 ;
      RECT -2.145 5.02 -1.975 8.31 ;
      RECT -2.145 7.32 -1.74 7.65 ;
      RECT -2.145 6.48 -1.74 6.81 ;
      RECT 75.76 0.58 75.93 1.09 ;
      RECT 75.76 2.4 75.93 3.87 ;
      RECT 75.76 5.02 75.93 6.49 ;
      RECT 75.76 7.8 75.93 8.31 ;
      RECT 74.77 0.58 74.94 1.09 ;
      RECT 74.77 2.4 74.94 3.87 ;
      RECT 74.77 5.02 74.94 6.49 ;
      RECT 74.77 7.8 74.94 8.31 ;
      RECT 73.405 0.58 73.575 3.87 ;
      RECT 73.405 5.02 73.575 8.31 ;
      RECT 72.975 0.58 73.145 1.09 ;
      RECT 72.975 1.66 73.145 3.87 ;
      RECT 72.975 5.02 73.145 7.23 ;
      RECT 72.975 7.8 73.145 8.31 ;
      RECT 71.605 1.665 71.775 2.94 ;
      RECT 71.605 5.95 71.775 7.225 ;
      RECT 69.3 1.76 69.47 2.11 ;
      RECT 69.06 2.5 69.23 2.83 ;
      RECT 68.58 2.5 68.75 2.95 ;
      RECT 68.34 1.76 68.51 2.11 ;
      RECT 68.1 2.5 68.27 2.83 ;
      RECT 67.79 5.02 67.96 8.31 ;
      RECT 67.36 5.02 67.53 7.23 ;
      RECT 67.36 7.8 67.53 8.31 ;
      RECT 67.35 3.49 67.52 3.82 ;
      RECT 66.66 2.5 66.83 2.95 ;
      RECT 66.18 2.5 66.35 2.83 ;
      RECT 65.99 5.95 66.16 7.225 ;
      RECT 65.7 2.5 65.87 2.83 ;
      RECT 65.22 2.5 65.39 2.95 ;
      RECT 64.98 3.49 65.15 3.82 ;
      RECT 64.74 2.5 64.91 3.23 ;
      RECT 64.26 2.5 64.43 2.83 ;
      RECT 64.02 1.76 64.19 2.11 ;
      RECT 63.54 3.06 63.71 3.48 ;
      RECT 63.3 2.5 63.47 2.83 ;
      RECT 63.06 3.15 63.23 3.51 ;
      RECT 62.82 2.5 62.99 2.95 ;
      RECT 62.34 2.5 62.51 2.95 ;
      RECT 62.13 1.76 62.3 2.11 ;
      RECT 62.13 3.15 62.3 3.51 ;
      RECT 60.5 0.58 60.67 1.09 ;
      RECT 60.5 2.4 60.67 3.87 ;
      RECT 60.5 5.02 60.67 6.49 ;
      RECT 60.5 7.8 60.67 8.31 ;
      RECT 59.51 0.58 59.68 1.09 ;
      RECT 59.51 2.4 59.68 3.87 ;
      RECT 59.51 5.02 59.68 6.49 ;
      RECT 59.51 7.8 59.68 8.31 ;
      RECT 58.145 0.58 58.315 3.87 ;
      RECT 58.145 5.02 58.315 8.31 ;
      RECT 57.715 0.58 57.885 1.09 ;
      RECT 57.715 1.66 57.885 3.87 ;
      RECT 57.715 5.02 57.885 7.23 ;
      RECT 57.715 7.8 57.885 8.31 ;
      RECT 56.345 1.665 56.515 2.94 ;
      RECT 56.345 5.95 56.515 7.225 ;
      RECT 54.04 1.76 54.21 2.11 ;
      RECT 53.8 2.5 53.97 2.83 ;
      RECT 53.32 2.5 53.49 2.95 ;
      RECT 53.08 1.76 53.25 2.11 ;
      RECT 52.84 2.5 53.01 2.83 ;
      RECT 52.53 5.02 52.7 8.31 ;
      RECT 52.1 5.02 52.27 7.23 ;
      RECT 52.1 7.8 52.27 8.31 ;
      RECT 52.09 3.49 52.26 3.82 ;
      RECT 51.4 2.5 51.57 2.95 ;
      RECT 50.92 2.5 51.09 2.83 ;
      RECT 50.73 5.95 50.9 7.225 ;
      RECT 50.44 2.5 50.61 2.83 ;
      RECT 49.96 2.5 50.13 2.95 ;
      RECT 49.72 3.49 49.89 3.82 ;
      RECT 49.48 2.5 49.65 3.23 ;
      RECT 49 2.5 49.17 2.83 ;
      RECT 48.76 1.76 48.93 2.11 ;
      RECT 48.28 3.06 48.45 3.48 ;
      RECT 48.04 2.5 48.21 2.83 ;
      RECT 47.8 3.15 47.97 3.51 ;
      RECT 47.56 2.5 47.73 2.95 ;
      RECT 47.08 2.5 47.25 2.95 ;
      RECT 46.87 1.76 47.04 2.11 ;
      RECT 46.87 3.15 47.04 3.51 ;
      RECT 45.24 0.58 45.41 1.09 ;
      RECT 45.24 2.4 45.41 3.87 ;
      RECT 45.24 5.02 45.41 6.49 ;
      RECT 45.24 7.8 45.41 8.31 ;
      RECT 44.25 0.58 44.42 1.09 ;
      RECT 44.25 2.4 44.42 3.87 ;
      RECT 44.25 5.02 44.42 6.49 ;
      RECT 44.25 7.8 44.42 8.31 ;
      RECT 42.885 0.58 43.055 3.87 ;
      RECT 42.885 5.02 43.055 8.31 ;
      RECT 42.455 0.58 42.625 1.09 ;
      RECT 42.455 1.66 42.625 3.87 ;
      RECT 42.455 5.02 42.625 7.23 ;
      RECT 42.455 7.8 42.625 8.31 ;
      RECT 41.085 1.665 41.255 2.94 ;
      RECT 41.085 5.95 41.255 7.225 ;
      RECT 38.78 1.76 38.95 2.11 ;
      RECT 38.54 2.5 38.71 2.83 ;
      RECT 38.06 2.5 38.23 2.95 ;
      RECT 37.82 1.76 37.99 2.11 ;
      RECT 37.58 2.5 37.75 2.83 ;
      RECT 37.27 5.02 37.44 8.31 ;
      RECT 36.84 5.02 37.01 7.23 ;
      RECT 36.84 7.8 37.01 8.31 ;
      RECT 36.83 3.49 37 3.82 ;
      RECT 36.14 2.5 36.31 2.95 ;
      RECT 35.66 2.5 35.83 2.83 ;
      RECT 35.47 5.95 35.64 7.225 ;
      RECT 35.18 2.5 35.35 2.83 ;
      RECT 34.7 2.5 34.87 2.95 ;
      RECT 34.46 3.49 34.63 3.82 ;
      RECT 34.22 2.5 34.39 3.23 ;
      RECT 33.74 2.5 33.91 2.83 ;
      RECT 33.5 1.76 33.67 2.11 ;
      RECT 33.02 3.06 33.19 3.48 ;
      RECT 32.78 2.5 32.95 2.83 ;
      RECT 32.54 3.15 32.71 3.51 ;
      RECT 32.3 2.5 32.47 2.95 ;
      RECT 31.82 2.5 31.99 2.95 ;
      RECT 31.61 1.76 31.78 2.11 ;
      RECT 31.61 3.15 31.78 3.51 ;
      RECT 29.98 0.58 30.15 1.09 ;
      RECT 29.98 2.4 30.15 3.87 ;
      RECT 29.98 5.02 30.15 6.49 ;
      RECT 29.98 7.8 30.15 8.31 ;
      RECT 28.99 0.58 29.16 1.09 ;
      RECT 28.99 2.4 29.16 3.87 ;
      RECT 28.99 5.02 29.16 6.49 ;
      RECT 28.99 7.8 29.16 8.31 ;
      RECT 27.625 0.58 27.795 3.87 ;
      RECT 27.625 5.02 27.795 8.31 ;
      RECT 27.195 0.58 27.365 1.09 ;
      RECT 27.195 1.66 27.365 3.87 ;
      RECT 27.195 5.02 27.365 7.23 ;
      RECT 27.195 7.8 27.365 8.31 ;
      RECT 25.825 1.665 25.995 2.94 ;
      RECT 25.825 5.95 25.995 7.225 ;
      RECT 23.52 1.76 23.69 2.11 ;
      RECT 23.28 2.5 23.45 2.83 ;
      RECT 22.8 2.5 22.97 2.95 ;
      RECT 22.56 1.76 22.73 2.11 ;
      RECT 22.32 2.5 22.49 2.83 ;
      RECT 22.01 5.02 22.18 8.31 ;
      RECT 21.58 5.02 21.75 7.23 ;
      RECT 21.58 7.8 21.75 8.31 ;
      RECT 21.57 3.49 21.74 3.82 ;
      RECT 20.88 2.5 21.05 2.95 ;
      RECT 20.4 2.5 20.57 2.83 ;
      RECT 20.21 5.95 20.38 7.225 ;
      RECT 19.92 2.5 20.09 2.83 ;
      RECT 19.44 2.5 19.61 2.95 ;
      RECT 19.2 3.49 19.37 3.82 ;
      RECT 18.96 2.5 19.13 3.23 ;
      RECT 18.48 2.5 18.65 2.83 ;
      RECT 18.24 1.76 18.41 2.11 ;
      RECT 17.76 3.06 17.93 3.48 ;
      RECT 17.52 2.5 17.69 2.83 ;
      RECT 17.28 3.15 17.45 3.51 ;
      RECT 17.04 2.5 17.21 2.95 ;
      RECT 16.56 2.5 16.73 2.95 ;
      RECT 16.35 1.76 16.52 2.11 ;
      RECT 16.35 3.15 16.52 3.51 ;
      RECT 14.72 0.58 14.89 1.09 ;
      RECT 14.72 2.4 14.89 3.87 ;
      RECT 14.72 5.02 14.89 6.49 ;
      RECT 14.72 7.8 14.89 8.31 ;
      RECT 13.73 0.58 13.9 1.09 ;
      RECT 13.73 2.4 13.9 3.87 ;
      RECT 13.73 5.02 13.9 6.49 ;
      RECT 13.73 7.8 13.9 8.31 ;
      RECT 12.365 0.58 12.535 3.87 ;
      RECT 12.365 5.02 12.535 8.31 ;
      RECT 11.935 0.58 12.105 1.09 ;
      RECT 11.935 1.66 12.105 3.87 ;
      RECT 11.935 5.02 12.105 7.23 ;
      RECT 11.935 7.8 12.105 8.31 ;
      RECT 10.565 1.665 10.735 2.94 ;
      RECT 10.565 5.95 10.735 7.225 ;
      RECT 8.26 1.76 8.43 2.11 ;
      RECT 8.02 2.5 8.19 2.83 ;
      RECT 7.54 2.5 7.71 2.95 ;
      RECT 7.3 1.76 7.47 2.11 ;
      RECT 7.06 2.5 7.23 2.83 ;
      RECT 6.75 5.02 6.92 8.31 ;
      RECT 6.32 5.02 6.49 7.23 ;
      RECT 6.32 7.8 6.49 8.31 ;
      RECT 6.31 3.49 6.48 3.82 ;
      RECT 5.62 2.5 5.79 2.95 ;
      RECT 5.14 2.5 5.31 2.83 ;
      RECT 4.95 5.95 5.12 7.225 ;
      RECT 4.66 2.5 4.83 2.83 ;
      RECT 4.18 2.5 4.35 2.95 ;
      RECT 3.94 3.49 4.11 3.82 ;
      RECT 3.7 2.5 3.87 3.23 ;
      RECT 3.22 2.5 3.39 2.83 ;
      RECT 2.98 1.76 3.15 2.11 ;
      RECT 2.5 3.06 2.67 3.48 ;
      RECT 2.26 2.5 2.43 2.83 ;
      RECT 2.02 3.15 2.19 3.51 ;
      RECT 1.78 2.5 1.95 2.95 ;
      RECT 1.3 2.5 1.47 2.95 ;
      RECT 1.09 1.76 1.26 2.11 ;
      RECT 1.09 3.15 1.26 3.51 ;
      RECT -1.195 5.02 -1.025 7.23 ;
      RECT -1.195 7.8 -1.025 8.31 ;
      RECT -2.565 5.95 -2.395 7.225 ;
  END
END sky130_osu_ring_oscillator_mpr2xa_8_b0r1

MACRO sky130_osu_ring_oscillator_mpr2xa_8_b0r2
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 2.795 -0.005 ;
  SIZE 79.095 BY 8.88 ;
  SYMMETRY X Y R90 ;
  SITE CoreSite ;
  OBS
    LAYER met4 ;
      RECT 63.94 2.98 64.27 3.31 ;
      RECT 63.955 2.505 64.27 3.31 ;
      RECT 66.1 2.49 66.43 2.845 ;
      RECT 63.955 2.505 66.43 2.805 ;
      RECT 48.68 2.98 49.01 3.31 ;
      RECT 48.695 2.505 49.01 3.31 ;
      RECT 50.84 2.49 51.17 2.845 ;
      RECT 48.695 2.505 51.17 2.805 ;
      RECT 33.42 2.98 33.75 3.31 ;
      RECT 33.435 2.505 33.75 3.31 ;
      RECT 35.58 2.49 35.91 2.845 ;
      RECT 33.435 2.505 35.91 2.805 ;
      RECT 18.16 2.98 18.49 3.31 ;
      RECT 18.175 2.505 18.49 3.31 ;
      RECT 20.32 2.49 20.65 2.845 ;
      RECT 18.175 2.505 20.65 2.805 ;
      RECT 2.9 2.98 3.23 3.31 ;
      RECT 2.915 2.505 3.23 3.31 ;
      RECT 5.06 2.49 5.39 2.845 ;
      RECT 2.915 2.505 5.39 2.805 ;
    LAYER via3 ;
      RECT 66.165 2.58 66.365 2.78 ;
      RECT 64.005 3.045 64.205 3.245 ;
      RECT 50.905 2.58 51.105 2.78 ;
      RECT 48.745 3.045 48.945 3.245 ;
      RECT 35.645 2.58 35.845 2.78 ;
      RECT 33.485 3.045 33.685 3.245 ;
      RECT 20.385 2.58 20.585 2.78 ;
      RECT 18.225 3.045 18.425 3.245 ;
      RECT 5.125 2.58 5.325 2.78 ;
      RECT 2.965 3.045 3.165 3.245 ;
    LAYER met3 ;
      RECT 70.965 1.11 71.305 3.07 ;
      RECT 65.225 1.885 65.955 2.215 ;
      RECT 65.375 1.11 65.675 2.215 ;
      RECT 65.375 1.11 71.305 1.41 ;
      RECT 67.26 7.06 67.63 7.43 ;
      RECT 67.295 4.48 67.595 7.43 ;
      RECT 65.855 4.48 67.595 4.78 ;
      RECT 63.06 4.26 66.155 4.56 ;
      RECT 65.855 2.52 66.155 4.78 ;
      RECT 63.06 2.98 63.36 4.56 ;
      RECT 66.58 3.515 66.91 3.87 ;
      RECT 64.675 3.555 66.91 3.855 ;
      RECT 64.675 2.42 64.975 3.855 ;
      RECT 62.755 2.98 63.485 3.31 ;
      RECT 65.65 2.525 66.43 2.87 ;
      RECT 66.125 2.49 66.43 2.87 ;
      RECT 64.66 2.42 64.99 2.75 ;
      RECT 63.945 2.42 64.265 3.335 ;
      RECT 63.945 2.42 64.275 2.955 ;
      RECT 55.705 1.11 56.045 3.07 ;
      RECT 49.965 1.885 50.695 2.215 ;
      RECT 50.115 1.11 50.415 2.215 ;
      RECT 50.115 1.11 56.045 1.41 ;
      RECT 52 7.06 52.37 7.43 ;
      RECT 52.035 4.48 52.335 7.43 ;
      RECT 50.595 4.48 52.335 4.78 ;
      RECT 47.8 4.26 50.895 4.56 ;
      RECT 50.595 2.52 50.895 4.78 ;
      RECT 47.8 2.98 48.1 4.56 ;
      RECT 51.32 3.515 51.65 3.87 ;
      RECT 49.415 3.555 51.65 3.855 ;
      RECT 49.415 2.42 49.715 3.855 ;
      RECT 47.495 2.98 48.225 3.31 ;
      RECT 50.39 2.525 51.17 2.87 ;
      RECT 50.865 2.49 51.17 2.87 ;
      RECT 49.4 2.42 49.73 2.75 ;
      RECT 48.685 2.42 49.005 3.335 ;
      RECT 48.685 2.42 49.015 2.955 ;
      RECT 40.445 1.11 40.785 3.07 ;
      RECT 34.705 1.885 35.435 2.215 ;
      RECT 34.855 1.11 35.155 2.215 ;
      RECT 34.855 1.11 40.785 1.41 ;
      RECT 36.74 7.06 37.11 7.43 ;
      RECT 36.775 4.48 37.075 7.43 ;
      RECT 35.335 4.48 37.075 4.78 ;
      RECT 32.54 4.26 35.635 4.56 ;
      RECT 35.335 2.52 35.635 4.78 ;
      RECT 32.54 2.98 32.84 4.56 ;
      RECT 36.06 3.515 36.39 3.87 ;
      RECT 34.155 3.555 36.39 3.855 ;
      RECT 34.155 2.42 34.455 3.855 ;
      RECT 32.235 2.98 32.965 3.31 ;
      RECT 35.13 2.525 35.91 2.87 ;
      RECT 35.605 2.49 35.91 2.87 ;
      RECT 34.14 2.42 34.47 2.75 ;
      RECT 33.425 2.42 33.745 3.335 ;
      RECT 33.425 2.42 33.755 2.955 ;
      RECT 25.185 1.11 25.525 3.07 ;
      RECT 19.445 1.885 20.175 2.215 ;
      RECT 19.595 1.11 19.895 2.215 ;
      RECT 19.595 1.11 25.525 1.41 ;
      RECT 21.48 7.06 21.85 7.43 ;
      RECT 21.515 4.48 21.815 7.43 ;
      RECT 20.075 4.48 21.815 4.78 ;
      RECT 17.28 4.26 20.375 4.56 ;
      RECT 20.075 2.52 20.375 4.78 ;
      RECT 17.28 2.98 17.58 4.56 ;
      RECT 20.8 3.515 21.13 3.87 ;
      RECT 18.895 3.555 21.13 3.855 ;
      RECT 18.895 2.42 19.195 3.855 ;
      RECT 16.975 2.98 17.705 3.31 ;
      RECT 19.87 2.525 20.65 2.87 ;
      RECT 20.345 2.49 20.65 2.87 ;
      RECT 18.88 2.42 19.21 2.75 ;
      RECT 18.165 2.42 18.485 3.335 ;
      RECT 18.165 2.42 18.495 2.955 ;
      RECT 9.925 1.11 10.265 3.07 ;
      RECT 4.185 1.885 4.915 2.215 ;
      RECT 4.335 1.11 4.635 2.215 ;
      RECT 4.335 1.11 10.265 1.41 ;
      RECT 6.22 7.06 6.59 7.43 ;
      RECT 6.255 4.48 6.555 7.43 ;
      RECT 4.815 4.48 6.555 4.78 ;
      RECT 2.02 4.26 5.115 4.56 ;
      RECT 4.815 2.52 5.115 4.78 ;
      RECT 2.02 2.98 2.32 4.56 ;
      RECT 5.54 3.515 5.87 3.87 ;
      RECT 3.635 3.555 5.87 3.855 ;
      RECT 3.635 2.42 3.935 3.855 ;
      RECT 1.715 2.98 2.445 3.31 ;
      RECT 4.61 2.525 5.39 2.87 ;
      RECT 5.085 2.49 5.39 2.87 ;
      RECT 3.62 2.42 3.95 2.75 ;
      RECT 2.905 2.42 3.225 3.335 ;
      RECT 2.905 2.42 3.235 2.955 ;
      RECT 69.5 1.86 70.23 2.19 ;
      RECT 67.81 1.875 68.54 2.205 ;
      RECT 66.775 1.86 67.505 2.21 ;
      RECT 62.62 1.86 63.35 2.19 ;
      RECT 54.24 1.86 54.97 2.19 ;
      RECT 52.55 1.875 53.28 2.205 ;
      RECT 51.515 1.86 52.245 2.21 ;
      RECT 47.36 1.86 48.09 2.19 ;
      RECT 38.98 1.86 39.71 2.19 ;
      RECT 37.29 1.875 38.02 2.205 ;
      RECT 36.255 1.86 36.985 2.21 ;
      RECT 32.1 1.86 32.83 2.19 ;
      RECT 23.72 1.86 24.45 2.19 ;
      RECT 22.03 1.875 22.76 2.205 ;
      RECT 20.995 1.86 21.725 2.21 ;
      RECT 16.84 1.86 17.57 2.19 ;
      RECT 8.46 1.86 9.19 2.19 ;
      RECT 6.77 1.875 7.5 2.205 ;
      RECT 5.735 1.86 6.465 2.21 ;
      RECT 1.58 1.86 2.31 2.19 ;
    LAYER via2 ;
      RECT 71.04 2.78 71.24 2.98 ;
      RECT 69.735 1.925 69.935 2.125 ;
      RECT 67.875 1.94 68.075 2.14 ;
      RECT 67.345 7.145 67.545 7.345 ;
      RECT 66.855 1.945 67.055 2.145 ;
      RECT 66.645 3.58 66.845 3.78 ;
      RECT 66.165 2.58 66.365 2.78 ;
      RECT 65.415 1.95 65.615 2.15 ;
      RECT 64.725 2.485 64.925 2.685 ;
      RECT 64.01 2.485 64.21 2.685 ;
      RECT 63.045 3.045 63.245 3.245 ;
      RECT 62.805 1.925 63.005 2.125 ;
      RECT 55.78 2.78 55.98 2.98 ;
      RECT 54.475 1.925 54.675 2.125 ;
      RECT 52.615 1.94 52.815 2.14 ;
      RECT 52.085 7.145 52.285 7.345 ;
      RECT 51.595 1.945 51.795 2.145 ;
      RECT 51.385 3.58 51.585 3.78 ;
      RECT 50.905 2.58 51.105 2.78 ;
      RECT 50.155 1.95 50.355 2.15 ;
      RECT 49.465 2.485 49.665 2.685 ;
      RECT 48.75 2.485 48.95 2.685 ;
      RECT 47.785 3.045 47.985 3.245 ;
      RECT 47.545 1.925 47.745 2.125 ;
      RECT 40.52 2.78 40.72 2.98 ;
      RECT 39.215 1.925 39.415 2.125 ;
      RECT 37.355 1.94 37.555 2.14 ;
      RECT 36.825 7.145 37.025 7.345 ;
      RECT 36.335 1.945 36.535 2.145 ;
      RECT 36.125 3.58 36.325 3.78 ;
      RECT 35.645 2.58 35.845 2.78 ;
      RECT 34.895 1.95 35.095 2.15 ;
      RECT 34.205 2.485 34.405 2.685 ;
      RECT 33.49 2.485 33.69 2.685 ;
      RECT 32.525 3.045 32.725 3.245 ;
      RECT 32.285 1.925 32.485 2.125 ;
      RECT 25.26 2.78 25.46 2.98 ;
      RECT 23.955 1.925 24.155 2.125 ;
      RECT 22.095 1.94 22.295 2.14 ;
      RECT 21.565 7.145 21.765 7.345 ;
      RECT 21.075 1.945 21.275 2.145 ;
      RECT 20.865 3.58 21.065 3.78 ;
      RECT 20.385 2.58 20.585 2.78 ;
      RECT 19.635 1.95 19.835 2.15 ;
      RECT 18.945 2.485 19.145 2.685 ;
      RECT 18.23 2.485 18.43 2.685 ;
      RECT 17.265 3.045 17.465 3.245 ;
      RECT 17.025 1.925 17.225 2.125 ;
      RECT 10 2.78 10.2 2.98 ;
      RECT 8.695 1.925 8.895 2.125 ;
      RECT 6.835 1.94 7.035 2.14 ;
      RECT 6.305 7.145 6.505 7.345 ;
      RECT 5.815 1.945 6.015 2.145 ;
      RECT 5.605 3.58 5.805 3.78 ;
      RECT 5.125 2.58 5.325 2.78 ;
      RECT 4.375 1.95 4.575 2.15 ;
      RECT 3.685 2.485 3.885 2.685 ;
      RECT 2.97 2.485 3.17 2.685 ;
      RECT 2.005 3.045 2.205 3.245 ;
      RECT 1.765 1.925 1.965 2.125 ;
    LAYER met2 ;
      RECT -1.565 8.405 75.93 8.575 ;
      RECT 75.76 7.28 75.93 8.575 ;
      RECT -1.565 6.26 -1.395 8.575 ;
      RECT 75.73 7.28 76.08 7.63 ;
      RECT -1.63 6.26 -1.34 6.61 ;
      RECT 72.57 6.225 72.89 6.55 ;
      RECT 72.6 5.7 72.77 6.55 ;
      RECT 72.6 5.7 72.775 6.05 ;
      RECT 72.6 5.7 73.575 5.875 ;
      RECT 73.4 1.97 73.575 5.875 ;
      RECT 73.345 1.97 73.695 2.32 ;
      RECT 73.37 6.66 73.695 6.985 ;
      RECT 72.255 6.75 73.695 6.92 ;
      RECT 72.255 2.4 72.415 6.92 ;
      RECT 72.57 2.37 72.89 2.69 ;
      RECT 72.255 2.4 72.89 2.57 ;
      RECT 71.525 5.865 71.865 6.215 ;
      RECT 71.605 2.71 71.775 6.215 ;
      RECT 71.525 2.71 71.865 3.06 ;
      RECT 70.995 2.69 71.285 3.07 ;
      RECT 70.965 2.705 71.305 3.055 ;
      RECT 69.705 3.545 69.965 3.865 ;
      RECT 69.765 1.84 69.905 3.865 ;
      RECT 69.59 2.4 69.905 2.77 ;
      RECT 69.66 1.955 69.905 2.77 ;
      RECT 69.695 1.84 69.975 2.21 ;
      RECT 69.015 2.425 69.275 2.745 ;
      RECT 68.355 2.515 69.275 2.655 ;
      RECT 68.355 1.575 68.495 2.655 ;
      RECT 64.815 1.865 65.075 2.185 ;
      RECT 64.995 1.575 65.135 2.095 ;
      RECT 64.995 1.575 68.495 1.715 ;
      RECT 60.445 6.66 60.795 7.01 ;
      RECT 67.93 6.615 68.28 6.965 ;
      RECT 60.445 6.69 68.28 6.89 ;
      RECT 67.845 3.265 68.105 3.585 ;
      RECT 67.905 1.855 68.045 3.585 ;
      RECT 67.835 1.855 68.115 2.225 ;
      RECT 65.235 4.015 67.67 4.155 ;
      RECT 67.53 2.705 67.67 4.155 ;
      RECT 65.235 3.635 65.375 4.155 ;
      RECT 64.935 3.635 65.375 3.865 ;
      RECT 62.595 3.635 65.375 3.775 ;
      RECT 64.935 3.545 65.195 3.865 ;
      RECT 62.595 3.355 62.735 3.775 ;
      RECT 62.085 3.265 62.345 3.585 ;
      RECT 62.085 3.355 62.735 3.495 ;
      RECT 62.145 1.865 62.285 3.585 ;
      RECT 67.47 2.705 67.73 3.025 ;
      RECT 62.085 1.865 62.345 2.185 ;
      RECT 67.095 3.545 67.355 3.865 ;
      RECT 67.155 1.955 67.295 3.865 ;
      RECT 66.815 1.955 67.295 2.23 ;
      RECT 66.615 1.86 67.095 2.205 ;
      RECT 66.605 3.495 66.885 3.865 ;
      RECT 66.675 2.4 66.815 3.865 ;
      RECT 66.615 2.4 66.875 3.025 ;
      RECT 66.605 2.4 66.885 2.77 ;
      RECT 65.535 3.545 65.795 3.865 ;
      RECT 65.535 3.355 65.735 3.865 ;
      RECT 65.34 3.355 65.735 3.495 ;
      RECT 65.34 1.865 65.48 3.495 ;
      RECT 65.34 1.865 65.655 2.235 ;
      RECT 65.28 1.865 65.655 2.185 ;
      RECT 63.005 2.96 63.285 3.33 ;
      RECT 64.455 2.985 64.715 3.305 ;
      RECT 62.835 3.075 64.715 3.215 ;
      RECT 62.835 2.96 63.285 3.215 ;
      RECT 62.775 2.4 63.035 3.025 ;
      RECT 62.765 2.4 63.045 2.77 ;
      RECT 63.845 2.4 64.255 2.77 ;
      RECT 63.255 2.425 63.515 2.745 ;
      RECT 63.255 2.515 64.255 2.655 ;
      RECT 62.765 1.84 63.045 2.21 ;
      RECT 62.765 1.865 63.155 2.185 ;
      RECT 57.31 6.225 57.63 6.55 ;
      RECT 57.34 5.7 57.51 6.55 ;
      RECT 57.34 5.7 57.515 6.05 ;
      RECT 57.34 5.7 58.315 5.875 ;
      RECT 58.14 1.97 58.315 5.875 ;
      RECT 58.085 1.97 58.435 2.32 ;
      RECT 58.11 6.66 58.435 6.985 ;
      RECT 56.995 6.75 58.435 6.92 ;
      RECT 56.995 2.4 57.155 6.92 ;
      RECT 57.31 2.37 57.63 2.69 ;
      RECT 56.995 2.4 57.63 2.57 ;
      RECT 56.265 5.865 56.605 6.215 ;
      RECT 56.345 2.71 56.515 6.215 ;
      RECT 56.265 2.71 56.605 3.06 ;
      RECT 55.735 2.69 56.025 3.07 ;
      RECT 55.705 2.705 56.045 3.055 ;
      RECT 54.445 3.545 54.705 3.865 ;
      RECT 54.505 1.84 54.645 3.865 ;
      RECT 54.33 2.4 54.645 2.77 ;
      RECT 54.4 1.955 54.645 2.77 ;
      RECT 54.435 1.84 54.715 2.21 ;
      RECT 53.755 2.425 54.015 2.745 ;
      RECT 53.095 2.515 54.015 2.655 ;
      RECT 53.095 1.575 53.235 2.655 ;
      RECT 49.555 1.865 49.815 2.185 ;
      RECT 49.735 1.575 49.875 2.095 ;
      RECT 49.735 1.575 53.235 1.715 ;
      RECT 45.185 6.66 45.535 7.01 ;
      RECT 52.675 6.615 53.025 6.965 ;
      RECT 45.185 6.69 53.025 6.89 ;
      RECT 52.585 3.265 52.845 3.585 ;
      RECT 52.645 1.855 52.785 3.585 ;
      RECT 52.575 1.855 52.855 2.225 ;
      RECT 49.975 4.015 52.41 4.155 ;
      RECT 52.27 2.705 52.41 4.155 ;
      RECT 49.975 3.635 50.115 4.155 ;
      RECT 49.675 3.635 50.115 3.865 ;
      RECT 47.335 3.635 50.115 3.775 ;
      RECT 49.675 3.545 49.935 3.865 ;
      RECT 47.335 3.355 47.475 3.775 ;
      RECT 46.825 3.265 47.085 3.585 ;
      RECT 46.825 3.355 47.475 3.495 ;
      RECT 46.885 1.865 47.025 3.585 ;
      RECT 52.21 2.705 52.47 3.025 ;
      RECT 46.825 1.865 47.085 2.185 ;
      RECT 51.835 3.545 52.095 3.865 ;
      RECT 51.895 1.955 52.035 3.865 ;
      RECT 51.555 1.955 52.035 2.23 ;
      RECT 51.355 1.86 51.835 2.205 ;
      RECT 51.345 3.495 51.625 3.865 ;
      RECT 51.415 2.4 51.555 3.865 ;
      RECT 51.355 2.4 51.615 3.025 ;
      RECT 51.345 2.4 51.625 2.77 ;
      RECT 50.275 3.545 50.535 3.865 ;
      RECT 50.275 3.355 50.475 3.865 ;
      RECT 50.08 3.355 50.475 3.495 ;
      RECT 50.08 1.865 50.22 3.495 ;
      RECT 50.08 1.865 50.395 2.235 ;
      RECT 50.02 1.865 50.395 2.185 ;
      RECT 47.745 2.96 48.025 3.33 ;
      RECT 49.195 2.985 49.455 3.305 ;
      RECT 47.575 3.075 49.455 3.215 ;
      RECT 47.575 2.96 48.025 3.215 ;
      RECT 47.515 2.4 47.775 3.025 ;
      RECT 47.505 2.4 47.785 2.77 ;
      RECT 48.585 2.4 48.995 2.77 ;
      RECT 47.995 2.425 48.255 2.745 ;
      RECT 47.995 2.515 48.995 2.655 ;
      RECT 47.505 1.84 47.785 2.21 ;
      RECT 47.505 1.865 47.895 2.185 ;
      RECT 42.05 6.225 42.37 6.55 ;
      RECT 42.08 5.7 42.25 6.55 ;
      RECT 42.08 5.7 42.255 6.05 ;
      RECT 42.08 5.7 43.055 5.875 ;
      RECT 42.88 1.97 43.055 5.875 ;
      RECT 42.825 1.97 43.175 2.32 ;
      RECT 42.85 6.66 43.175 6.985 ;
      RECT 41.735 6.75 43.175 6.92 ;
      RECT 41.735 2.4 41.895 6.92 ;
      RECT 42.05 2.37 42.37 2.69 ;
      RECT 41.735 2.4 42.37 2.57 ;
      RECT 41.005 5.865 41.345 6.215 ;
      RECT 41.085 2.71 41.255 6.215 ;
      RECT 41.005 2.71 41.345 3.06 ;
      RECT 40.475 2.69 40.765 3.07 ;
      RECT 40.445 2.705 40.785 3.055 ;
      RECT 39.185 3.545 39.445 3.865 ;
      RECT 39.245 1.84 39.385 3.865 ;
      RECT 39.07 2.4 39.385 2.77 ;
      RECT 39.14 1.955 39.385 2.77 ;
      RECT 39.175 1.84 39.455 2.21 ;
      RECT 38.495 2.425 38.755 2.745 ;
      RECT 37.835 2.515 38.755 2.655 ;
      RECT 37.835 1.575 37.975 2.655 ;
      RECT 34.295 1.865 34.555 2.185 ;
      RECT 34.475 1.575 34.615 2.095 ;
      RECT 34.475 1.575 37.975 1.715 ;
      RECT 29.97 6.665 30.32 7.015 ;
      RECT 37.41 6.62 37.76 6.97 ;
      RECT 29.97 6.695 37.76 6.895 ;
      RECT 37.325 3.265 37.585 3.585 ;
      RECT 37.385 1.855 37.525 3.585 ;
      RECT 37.315 1.855 37.595 2.225 ;
      RECT 34.715 4.015 37.15 4.155 ;
      RECT 37.01 2.705 37.15 4.155 ;
      RECT 34.715 3.635 34.855 4.155 ;
      RECT 34.415 3.635 34.855 3.865 ;
      RECT 32.075 3.635 34.855 3.775 ;
      RECT 34.415 3.545 34.675 3.865 ;
      RECT 32.075 3.355 32.215 3.775 ;
      RECT 31.565 3.265 31.825 3.585 ;
      RECT 31.565 3.355 32.215 3.495 ;
      RECT 31.625 1.865 31.765 3.585 ;
      RECT 36.95 2.705 37.21 3.025 ;
      RECT 31.565 1.865 31.825 2.185 ;
      RECT 36.575 3.545 36.835 3.865 ;
      RECT 36.635 1.955 36.775 3.865 ;
      RECT 36.295 1.955 36.775 2.23 ;
      RECT 36.095 1.86 36.575 2.205 ;
      RECT 36.085 3.495 36.365 3.865 ;
      RECT 36.155 2.4 36.295 3.865 ;
      RECT 36.095 2.4 36.355 3.025 ;
      RECT 36.085 2.4 36.365 2.77 ;
      RECT 35.015 3.545 35.275 3.865 ;
      RECT 35.015 3.355 35.215 3.865 ;
      RECT 34.82 3.355 35.215 3.495 ;
      RECT 34.82 1.865 34.96 3.495 ;
      RECT 34.82 1.865 35.135 2.235 ;
      RECT 34.76 1.865 35.135 2.185 ;
      RECT 32.485 2.96 32.765 3.33 ;
      RECT 33.935 2.985 34.195 3.305 ;
      RECT 32.315 3.075 34.195 3.215 ;
      RECT 32.315 2.96 32.765 3.215 ;
      RECT 32.255 2.4 32.515 3.025 ;
      RECT 32.245 2.4 32.525 2.77 ;
      RECT 33.325 2.4 33.735 2.77 ;
      RECT 32.735 2.425 32.995 2.745 ;
      RECT 32.735 2.515 33.735 2.655 ;
      RECT 32.245 1.84 32.525 2.21 ;
      RECT 32.245 1.865 32.635 2.185 ;
      RECT 26.79 6.225 27.11 6.55 ;
      RECT 26.82 5.7 26.99 6.55 ;
      RECT 26.82 5.7 26.995 6.05 ;
      RECT 26.82 5.7 27.795 5.875 ;
      RECT 27.62 1.97 27.795 5.875 ;
      RECT 27.565 1.97 27.915 2.32 ;
      RECT 27.59 6.66 27.915 6.985 ;
      RECT 26.475 6.75 27.915 6.92 ;
      RECT 26.475 2.4 26.635 6.92 ;
      RECT 26.79 2.37 27.11 2.69 ;
      RECT 26.475 2.4 27.11 2.57 ;
      RECT 25.745 5.865 26.085 6.215 ;
      RECT 25.825 2.71 25.995 6.215 ;
      RECT 25.745 2.71 26.085 3.06 ;
      RECT 25.215 2.69 25.505 3.07 ;
      RECT 25.185 2.705 25.525 3.055 ;
      RECT 23.925 3.545 24.185 3.865 ;
      RECT 23.985 1.84 24.125 3.865 ;
      RECT 23.81 2.4 24.125 2.77 ;
      RECT 23.88 1.955 24.125 2.77 ;
      RECT 23.915 1.84 24.195 2.21 ;
      RECT 23.235 2.425 23.495 2.745 ;
      RECT 22.575 2.515 23.495 2.655 ;
      RECT 22.575 1.575 22.715 2.655 ;
      RECT 19.035 1.865 19.295 2.185 ;
      RECT 19.215 1.575 19.355 2.095 ;
      RECT 19.215 1.575 22.715 1.715 ;
      RECT 14.71 6.66 15.06 7.01 ;
      RECT 22.15 6.615 22.5 6.965 ;
      RECT 14.71 6.69 22.5 6.89 ;
      RECT 22.065 3.265 22.325 3.585 ;
      RECT 22.125 1.855 22.265 3.585 ;
      RECT 22.055 1.855 22.335 2.225 ;
      RECT 19.455 4.015 21.89 4.155 ;
      RECT 21.75 2.705 21.89 4.155 ;
      RECT 19.455 3.635 19.595 4.155 ;
      RECT 19.155 3.635 19.595 3.865 ;
      RECT 16.815 3.635 19.595 3.775 ;
      RECT 19.155 3.545 19.415 3.865 ;
      RECT 16.815 3.355 16.955 3.775 ;
      RECT 16.305 3.265 16.565 3.585 ;
      RECT 16.305 3.355 16.955 3.495 ;
      RECT 16.365 1.865 16.505 3.585 ;
      RECT 21.69 2.705 21.95 3.025 ;
      RECT 16.305 1.865 16.565 2.185 ;
      RECT 21.315 3.545 21.575 3.865 ;
      RECT 21.375 1.955 21.515 3.865 ;
      RECT 21.035 1.955 21.515 2.23 ;
      RECT 20.835 1.86 21.315 2.205 ;
      RECT 20.825 3.495 21.105 3.865 ;
      RECT 20.895 2.4 21.035 3.865 ;
      RECT 20.835 2.4 21.095 3.025 ;
      RECT 20.825 2.4 21.105 2.77 ;
      RECT 19.755 3.545 20.015 3.865 ;
      RECT 19.755 3.355 19.955 3.865 ;
      RECT 19.56 3.355 19.955 3.495 ;
      RECT 19.56 1.865 19.7 3.495 ;
      RECT 19.56 1.865 19.875 2.235 ;
      RECT 19.5 1.865 19.875 2.185 ;
      RECT 17.225 2.96 17.505 3.33 ;
      RECT 18.675 2.985 18.935 3.305 ;
      RECT 17.055 3.075 18.935 3.215 ;
      RECT 17.055 2.96 17.505 3.215 ;
      RECT 16.995 2.4 17.255 3.025 ;
      RECT 16.985 2.4 17.265 2.77 ;
      RECT 18.065 2.4 18.475 2.77 ;
      RECT 17.475 2.425 17.735 2.745 ;
      RECT 17.475 2.515 18.475 2.655 ;
      RECT 16.985 1.84 17.265 2.21 ;
      RECT 16.985 1.865 17.375 2.185 ;
      RECT 11.53 6.225 11.85 6.55 ;
      RECT 11.56 5.7 11.73 6.55 ;
      RECT 11.56 5.7 11.735 6.05 ;
      RECT 11.56 5.7 12.535 5.875 ;
      RECT 12.36 1.97 12.535 5.875 ;
      RECT 12.305 1.97 12.655 2.32 ;
      RECT 12.33 6.66 12.655 6.985 ;
      RECT 11.215 6.75 12.655 6.92 ;
      RECT 11.215 2.4 11.375 6.92 ;
      RECT 11.53 2.37 11.85 2.69 ;
      RECT 11.215 2.4 11.85 2.57 ;
      RECT 10.485 5.865 10.825 6.215 ;
      RECT 10.565 2.71 10.735 6.215 ;
      RECT 10.485 2.71 10.825 3.06 ;
      RECT 9.955 2.69 10.245 3.07 ;
      RECT 9.925 2.705 10.265 3.055 ;
      RECT 8.665 3.545 8.925 3.865 ;
      RECT 8.725 1.84 8.865 3.865 ;
      RECT 8.55 2.4 8.865 2.77 ;
      RECT 8.62 1.955 8.865 2.77 ;
      RECT 8.655 1.84 8.935 2.21 ;
      RECT 7.975 2.425 8.235 2.745 ;
      RECT 7.315 2.515 8.235 2.655 ;
      RECT 7.315 1.575 7.455 2.655 ;
      RECT 3.775 1.865 4.035 2.185 ;
      RECT 3.955 1.575 4.095 2.095 ;
      RECT 3.955 1.575 7.455 1.715 ;
      RECT -1.255 7 -0.965 7.35 ;
      RECT -1.255 7.055 0 7.225 ;
      RECT -0.17 6.69 0 7.225 ;
      RECT 6.89 6.61 7.24 6.96 ;
      RECT -0.17 6.69 7.24 6.86 ;
      RECT 6.805 3.265 7.065 3.585 ;
      RECT 6.865 1.855 7.005 3.585 ;
      RECT 6.795 1.855 7.075 2.225 ;
      RECT 4.195 4.015 6.63 4.155 ;
      RECT 6.49 2.705 6.63 4.155 ;
      RECT 4.195 3.635 4.335 4.155 ;
      RECT 3.895 3.635 4.335 3.865 ;
      RECT 1.555 3.635 4.335 3.775 ;
      RECT 3.895 3.545 4.155 3.865 ;
      RECT 1.555 3.355 1.695 3.775 ;
      RECT 1.045 3.265 1.305 3.585 ;
      RECT 1.045 3.355 1.695 3.495 ;
      RECT 1.105 1.865 1.245 3.585 ;
      RECT 6.43 2.705 6.69 3.025 ;
      RECT 1.045 1.865 1.305 2.185 ;
      RECT 6.055 3.545 6.315 3.865 ;
      RECT 6.115 1.955 6.255 3.865 ;
      RECT 5.775 1.955 6.255 2.23 ;
      RECT 5.575 1.86 6.055 2.205 ;
      RECT 5.565 3.495 5.845 3.865 ;
      RECT 5.635 2.4 5.775 3.865 ;
      RECT 5.575 2.4 5.835 3.025 ;
      RECT 5.565 2.4 5.845 2.77 ;
      RECT 4.495 3.545 4.755 3.865 ;
      RECT 4.495 3.355 4.695 3.865 ;
      RECT 4.3 3.355 4.695 3.495 ;
      RECT 4.3 1.865 4.44 3.495 ;
      RECT 4.3 1.865 4.615 2.235 ;
      RECT 4.24 1.865 4.615 2.185 ;
      RECT 1.965 2.96 2.245 3.33 ;
      RECT 3.415 2.985 3.675 3.305 ;
      RECT 1.795 3.075 3.675 3.215 ;
      RECT 1.795 2.96 2.245 3.215 ;
      RECT 1.735 2.4 1.995 3.025 ;
      RECT 1.725 2.4 2.005 2.77 ;
      RECT 2.805 2.4 3.215 2.77 ;
      RECT 2.215 2.425 2.475 2.745 ;
      RECT 2.215 2.515 3.215 2.655 ;
      RECT 1.725 1.84 2.005 2.21 ;
      RECT 1.725 1.865 2.115 2.185 ;
      RECT 67.26 7.06 67.63 7.43 ;
      RECT 66.125 2.4 66.405 2.865 ;
      RECT 65.885 1.865 66.165 2.21 ;
      RECT 64.685 2.4 64.965 2.77 ;
      RECT 62.125 1.22 62.495 1.225 ;
      RECT 52 7.06 52.37 7.43 ;
      RECT 50.865 2.4 51.145 2.865 ;
      RECT 50.625 1.865 50.905 2.21 ;
      RECT 49.425 2.4 49.705 2.77 ;
      RECT 46.865 1.22 47.235 1.225 ;
      RECT 36.74 7.06 37.11 7.43 ;
      RECT 35.605 2.4 35.885 2.865 ;
      RECT 35.365 1.865 35.645 2.21 ;
      RECT 34.165 2.4 34.445 2.77 ;
      RECT 31.605 1.22 31.975 1.225 ;
      RECT 21.48 7.06 21.85 7.43 ;
      RECT 20.345 2.4 20.625 2.865 ;
      RECT 20.105 1.865 20.385 2.21 ;
      RECT 18.905 2.4 19.185 2.77 ;
      RECT 16.345 1.22 16.715 1.225 ;
      RECT 6.22 7.06 6.59 7.43 ;
      RECT 5.085 2.4 5.365 2.865 ;
      RECT 4.845 1.865 5.125 2.21 ;
      RECT 3.645 2.4 3.925 2.77 ;
      RECT 1.085 1.22 1.455 1.225 ;
    LAYER via1 ;
      RECT 75.83 7.38 75.98 7.53 ;
      RECT 73.46 6.745 73.61 6.895 ;
      RECT 73.445 2.07 73.595 2.22 ;
      RECT 72.655 2.455 72.805 2.605 ;
      RECT 72.655 6.33 72.805 6.48 ;
      RECT 71.625 2.81 71.775 2.96 ;
      RECT 71.625 5.965 71.775 6.115 ;
      RECT 71.065 2.805 71.215 2.955 ;
      RECT 69.76 1.95 69.91 2.1 ;
      RECT 69.76 3.63 69.91 3.78 ;
      RECT 69.07 2.51 69.22 2.66 ;
      RECT 68.03 6.715 68.18 6.865 ;
      RECT 67.9 1.95 68.05 2.1 ;
      RECT 67.9 3.35 68.05 3.5 ;
      RECT 67.525 2.79 67.675 2.94 ;
      RECT 67.37 7.17 67.52 7.32 ;
      RECT 67.15 3.63 67.3 3.78 ;
      RECT 66.67 1.95 66.82 2.1 ;
      RECT 66.67 2.79 66.82 2.94 ;
      RECT 66.19 2.51 66.34 2.66 ;
      RECT 65.95 1.95 66.1 2.1 ;
      RECT 65.59 3.63 65.74 3.78 ;
      RECT 65.335 1.95 65.485 2.1 ;
      RECT 64.99 3.63 65.14 3.78 ;
      RECT 64.87 1.95 65.02 2.1 ;
      RECT 64.75 2.51 64.9 2.66 ;
      RECT 64.51 3.07 64.66 3.22 ;
      RECT 63.31 2.51 63.46 2.66 ;
      RECT 62.95 1.95 63.1 2.1 ;
      RECT 62.83 2.79 62.98 2.94 ;
      RECT 62.14 1.95 62.29 2.1 ;
      RECT 62.14 3.35 62.29 3.5 ;
      RECT 60.545 6.76 60.695 6.91 ;
      RECT 58.2 6.745 58.35 6.895 ;
      RECT 58.185 2.07 58.335 2.22 ;
      RECT 57.395 2.455 57.545 2.605 ;
      RECT 57.395 6.33 57.545 6.48 ;
      RECT 56.365 2.81 56.515 2.96 ;
      RECT 56.365 5.965 56.515 6.115 ;
      RECT 55.805 2.805 55.955 2.955 ;
      RECT 54.5 1.95 54.65 2.1 ;
      RECT 54.5 3.63 54.65 3.78 ;
      RECT 53.81 2.51 53.96 2.66 ;
      RECT 52.775 6.715 52.925 6.865 ;
      RECT 52.64 1.95 52.79 2.1 ;
      RECT 52.64 3.35 52.79 3.5 ;
      RECT 52.265 2.79 52.415 2.94 ;
      RECT 52.11 7.17 52.26 7.32 ;
      RECT 51.89 3.63 52.04 3.78 ;
      RECT 51.41 1.95 51.56 2.1 ;
      RECT 51.41 2.79 51.56 2.94 ;
      RECT 50.93 2.51 51.08 2.66 ;
      RECT 50.69 1.95 50.84 2.1 ;
      RECT 50.33 3.63 50.48 3.78 ;
      RECT 50.075 1.95 50.225 2.1 ;
      RECT 49.73 3.63 49.88 3.78 ;
      RECT 49.61 1.95 49.76 2.1 ;
      RECT 49.49 2.51 49.64 2.66 ;
      RECT 49.25 3.07 49.4 3.22 ;
      RECT 48.05 2.51 48.2 2.66 ;
      RECT 47.69 1.95 47.84 2.1 ;
      RECT 47.57 2.79 47.72 2.94 ;
      RECT 46.88 1.95 47.03 2.1 ;
      RECT 46.88 3.35 47.03 3.5 ;
      RECT 45.285 6.76 45.435 6.91 ;
      RECT 42.94 6.745 43.09 6.895 ;
      RECT 42.925 2.07 43.075 2.22 ;
      RECT 42.135 2.455 42.285 2.605 ;
      RECT 42.135 6.33 42.285 6.48 ;
      RECT 41.105 2.81 41.255 2.96 ;
      RECT 41.105 5.965 41.255 6.115 ;
      RECT 40.545 2.805 40.695 2.955 ;
      RECT 39.24 1.95 39.39 2.1 ;
      RECT 39.24 3.63 39.39 3.78 ;
      RECT 38.55 2.51 38.7 2.66 ;
      RECT 37.51 6.72 37.66 6.87 ;
      RECT 37.38 1.95 37.53 2.1 ;
      RECT 37.38 3.35 37.53 3.5 ;
      RECT 37.005 2.79 37.155 2.94 ;
      RECT 36.85 7.17 37 7.32 ;
      RECT 36.63 3.63 36.78 3.78 ;
      RECT 36.15 1.95 36.3 2.1 ;
      RECT 36.15 2.79 36.3 2.94 ;
      RECT 35.67 2.51 35.82 2.66 ;
      RECT 35.43 1.95 35.58 2.1 ;
      RECT 35.07 3.63 35.22 3.78 ;
      RECT 34.815 1.95 34.965 2.1 ;
      RECT 34.47 3.63 34.62 3.78 ;
      RECT 34.35 1.95 34.5 2.1 ;
      RECT 34.23 2.51 34.38 2.66 ;
      RECT 33.99 3.07 34.14 3.22 ;
      RECT 32.79 2.51 32.94 2.66 ;
      RECT 32.43 1.95 32.58 2.1 ;
      RECT 32.31 2.79 32.46 2.94 ;
      RECT 31.62 1.95 31.77 2.1 ;
      RECT 31.62 3.35 31.77 3.5 ;
      RECT 30.07 6.765 30.22 6.915 ;
      RECT 27.68 6.745 27.83 6.895 ;
      RECT 27.665 2.07 27.815 2.22 ;
      RECT 26.875 2.455 27.025 2.605 ;
      RECT 26.875 6.33 27.025 6.48 ;
      RECT 25.845 2.81 25.995 2.96 ;
      RECT 25.845 5.965 25.995 6.115 ;
      RECT 25.285 2.805 25.435 2.955 ;
      RECT 23.98 1.95 24.13 2.1 ;
      RECT 23.98 3.63 24.13 3.78 ;
      RECT 23.29 2.51 23.44 2.66 ;
      RECT 22.25 6.715 22.4 6.865 ;
      RECT 22.12 1.95 22.27 2.1 ;
      RECT 22.12 3.35 22.27 3.5 ;
      RECT 21.745 2.79 21.895 2.94 ;
      RECT 21.59 7.17 21.74 7.32 ;
      RECT 21.37 3.63 21.52 3.78 ;
      RECT 20.89 1.95 21.04 2.1 ;
      RECT 20.89 2.79 21.04 2.94 ;
      RECT 20.41 2.51 20.56 2.66 ;
      RECT 20.17 1.95 20.32 2.1 ;
      RECT 19.81 3.63 19.96 3.78 ;
      RECT 19.555 1.95 19.705 2.1 ;
      RECT 19.21 3.63 19.36 3.78 ;
      RECT 19.09 1.95 19.24 2.1 ;
      RECT 18.97 2.51 19.12 2.66 ;
      RECT 18.73 3.07 18.88 3.22 ;
      RECT 17.53 2.51 17.68 2.66 ;
      RECT 17.17 1.95 17.32 2.1 ;
      RECT 17.05 2.79 17.2 2.94 ;
      RECT 16.36 1.95 16.51 2.1 ;
      RECT 16.36 3.35 16.51 3.5 ;
      RECT 14.81 6.76 14.96 6.91 ;
      RECT 12.42 6.745 12.57 6.895 ;
      RECT 12.405 2.07 12.555 2.22 ;
      RECT 11.615 2.455 11.765 2.605 ;
      RECT 11.615 6.33 11.765 6.48 ;
      RECT 10.585 2.81 10.735 2.96 ;
      RECT 10.585 5.965 10.735 6.115 ;
      RECT 10.025 2.805 10.175 2.955 ;
      RECT 8.72 1.95 8.87 2.1 ;
      RECT 8.72 3.63 8.87 3.78 ;
      RECT 8.03 2.51 8.18 2.66 ;
      RECT 6.99 6.71 7.14 6.86 ;
      RECT 6.86 1.95 7.01 2.1 ;
      RECT 6.86 3.35 7.01 3.5 ;
      RECT 6.485 2.79 6.635 2.94 ;
      RECT 6.33 7.17 6.48 7.32 ;
      RECT 6.11 3.63 6.26 3.78 ;
      RECT 5.63 1.95 5.78 2.1 ;
      RECT 5.63 2.79 5.78 2.94 ;
      RECT 5.15 2.51 5.3 2.66 ;
      RECT 4.91 1.95 5.06 2.1 ;
      RECT 4.55 3.63 4.7 3.78 ;
      RECT 4.295 1.95 4.445 2.1 ;
      RECT 3.95 3.63 4.1 3.78 ;
      RECT 3.83 1.95 3.98 2.1 ;
      RECT 3.71 2.51 3.86 2.66 ;
      RECT 3.47 3.07 3.62 3.22 ;
      RECT 2.27 2.51 2.42 2.66 ;
      RECT 1.91 1.95 2.06 2.1 ;
      RECT 1.79 2.79 1.94 2.94 ;
      RECT 1.1 1.95 1.25 2.1 ;
      RECT 1.1 3.35 1.25 3.5 ;
      RECT -1.185 7.1 -1.035 7.25 ;
      RECT -1.56 6.36 -1.41 6.51 ;
    LAYER met1 ;
      RECT 62.28 2.75 62.57 2.98 ;
      RECT 47.02 2.75 47.31 2.98 ;
      RECT 31.76 2.75 32.05 2.98 ;
      RECT 16.5 2.75 16.79 2.98 ;
      RECT 1.24 2.75 1.53 2.98 ;
      RECT 62.355 2.375 62.495 2.98 ;
      RECT 47.095 2.375 47.235 2.98 ;
      RECT 31.835 2.375 31.975 2.98 ;
      RECT 16.575 2.375 16.715 2.98 ;
      RECT 1.315 2.375 1.455 2.98 ;
      RECT 62.355 2.375 62.975 2.515 ;
      RECT 62.835 0.005 62.975 2.515 ;
      RECT 47.095 2.375 47.715 2.515 ;
      RECT 47.575 0.005 47.715 2.515 ;
      RECT 31.835 2.375 32.455 2.515 ;
      RECT 32.315 0.005 32.455 2.515 ;
      RECT 16.575 2.375 17.195 2.515 ;
      RECT 17.055 0.005 17.195 2.515 ;
      RECT 1.315 2.375 1.935 2.515 ;
      RECT 1.795 0.005 1.935 2.515 ;
      RECT 62.595 1.955 62.975 2.215 ;
      RECT 47.335 1.955 47.715 2.215 ;
      RECT 32.075 1.955 32.455 2.215 ;
      RECT 16.815 1.955 17.195 2.215 ;
      RECT 1.555 1.955 1.935 2.215 ;
      RECT 62.775 1.895 63.185 2.155 ;
      RECT 47.515 1.895 47.925 2.155 ;
      RECT 32.255 1.895 32.665 2.155 ;
      RECT 16.995 1.895 17.405 2.155 ;
      RECT 1.735 1.895 2.145 2.155 ;
      RECT 63.48 1.91 63.77 2.14 ;
      RECT 48.22 1.91 48.51 2.14 ;
      RECT 32.96 1.91 33.25 2.14 ;
      RECT 17.7 1.91 17.99 2.14 ;
      RECT 2.44 1.91 2.73 2.14 ;
      RECT 62.595 1.955 63.77 2.095 ;
      RECT 47.335 1.955 48.51 2.095 ;
      RECT 32.075 1.955 33.25 2.095 ;
      RECT 16.815 1.955 17.99 2.095 ;
      RECT 1.555 1.955 2.73 2.095 ;
      RECT 62.775 0.005 63.065 2.155 ;
      RECT 47.515 0.005 47.805 2.155 ;
      RECT 32.255 0.005 32.545 2.155 ;
      RECT 16.995 0.005 17.285 2.155 ;
      RECT 1.735 0.005 2.025 2.155 ;
      RECT 61.79 0.005 70.53 1.745 ;
      RECT 46.53 0.005 55.27 1.745 ;
      RECT 31.27 0.005 40.01 1.745 ;
      RECT 16.01 0.005 24.75 1.745 ;
      RECT 0.75 0.005 9.49 1.745 ;
      RECT -2.75 0.005 76.3 0.31 ;
      RECT -2.75 4.145 76.3 4.75 ;
      RECT 61.79 4.14 76.3 4.75 ;
      RECT 46.53 4.14 61.04 4.75 ;
      RECT 31.27 4.14 45.78 4.75 ;
      RECT 16.01 4.14 30.52 4.75 ;
      RECT 0.75 4.14 15.26 4.75 ;
      RECT 61.79 3.985 70.53 4.75 ;
      RECT 46.53 3.985 55.27 4.75 ;
      RECT 31.27 3.985 40.01 4.75 ;
      RECT 16.01 3.985 24.75 4.75 ;
      RECT 0.75 3.985 9.49 4.75 ;
      RECT -2.75 8.58 76.3 8.885 ;
      RECT 66.76 6.32 66.93 8.885 ;
      RECT 51.5 6.32 51.67 8.885 ;
      RECT 36.24 6.32 36.41 8.885 ;
      RECT 20.98 6.32 21.15 8.885 ;
      RECT 5.72 6.32 5.89 8.885 ;
      RECT 66.925 6.29 67.215 6.52 ;
      RECT 51.665 6.29 51.955 6.52 ;
      RECT 36.405 6.29 36.695 6.52 ;
      RECT 21.145 6.29 21.435 6.52 ;
      RECT 5.885 6.29 6.175 6.52 ;
      RECT 66.755 6.32 67.215 6.49 ;
      RECT 51.495 6.32 51.955 6.49 ;
      RECT 36.235 6.32 36.695 6.49 ;
      RECT 20.975 6.32 21.435 6.49 ;
      RECT 5.715 6.32 6.175 6.49 ;
      RECT 75.7 7.77 75.99 8 ;
      RECT 75.76 6.29 75.93 8 ;
      RECT 75.73 7.28 76.08 7.63 ;
      RECT 75.7 6.29 75.99 6.52 ;
      RECT 75.7 2.37 75.99 2.6 ;
      RECT 75.76 0.89 75.93 2.6 ;
      RECT 75.7 0.89 75.99 1.12 ;
      RECT 75.29 2.74 75.62 2.97 ;
      RECT 75.29 2.77 75.79 2.94 ;
      RECT 75.29 2.4 75.48 2.97 ;
      RECT 74.71 2.37 75 2.6 ;
      RECT 74.71 2.4 75.48 2.57 ;
      RECT 74.77 0.89 74.94 2.6 ;
      RECT 74.71 0.89 75 1.12 ;
      RECT 74.71 7.77 75 8 ;
      RECT 74.77 6.29 74.94 8 ;
      RECT 74.71 6.29 75 6.52 ;
      RECT 74.71 6.33 75.56 6.49 ;
      RECT 75.39 5.92 75.56 6.49 ;
      RECT 74.71 6.325 75.1 6.49 ;
      RECT 75.33 5.92 75.62 6.15 ;
      RECT 75.33 5.95 75.79 6.12 ;
      RECT 74.34 2.74 74.63 2.97 ;
      RECT 74.34 2.77 74.8 2.94 ;
      RECT 74.4 1.66 74.565 2.97 ;
      RECT 72.915 1.63 73.205 1.86 ;
      RECT 72.915 1.66 74.565 1.83 ;
      RECT 72.975 0.89 73.145 1.86 ;
      RECT 72.915 0.89 73.205 1.12 ;
      RECT 72.915 7.77 73.205 8 ;
      RECT 72.975 7.03 73.145 8 ;
      RECT 72.975 7.125 74.565 7.295 ;
      RECT 74.395 5.92 74.565 7.295 ;
      RECT 72.915 7.03 73.205 7.26 ;
      RECT 74.34 5.92 74.63 6.15 ;
      RECT 74.34 5.95 74.8 6.12 ;
      RECT 70.965 2.705 71.305 3.055 ;
      RECT 71.055 2.03 71.225 3.055 ;
      RECT 73.345 1.97 73.695 2.32 ;
      RECT 71.055 2.03 73.695 2.2 ;
      RECT 73.37 6.66 73.695 6.985 ;
      RECT 67.93 6.615 68.28 6.965 ;
      RECT 73.345 6.66 73.695 6.89 ;
      RECT 67.73 6.66 68.28 6.89 ;
      RECT 67.56 6.69 73.695 6.86 ;
      RECT 72.57 2.37 72.89 2.69 ;
      RECT 72.54 2.37 72.89 2.6 ;
      RECT 72.37 2.4 72.89 2.57 ;
      RECT 72.57 6.26 72.89 6.55 ;
      RECT 72.54 6.29 72.89 6.52 ;
      RECT 72.37 6.32 72.89 6.49 ;
      RECT 71.525 2.71 71.865 3.06 ;
      RECT 71.525 2.77 72.005 2.94 ;
      RECT 71.525 5.865 71.865 6.215 ;
      RECT 65.93 5.92 66.22 6.15 ;
      RECT 65.93 5.95 72.005 6.12 ;
      RECT 69.675 1.895 69.995 2.155 ;
      RECT 69.24 1.91 69.53 2.14 ;
      RECT 69.24 1.955 69.995 2.095 ;
      RECT 69.675 3.575 69.995 3.835 ;
      RECT 69.24 3.59 69.53 3.82 ;
      RECT 69.24 3.635 69.995 3.775 ;
      RECT 69 3.03 69.29 3.26 ;
      RECT 69 3.075 69.575 3.215 ;
      RECT 69.435 2.935 69.695 3.075 ;
      RECT 69.48 2.75 69.77 2.98 ;
      RECT 67.635 2.935 68.735 3.075 ;
      RECT 67.44 2.735 67.76 2.995 ;
      RECT 68.52 2.75 68.81 2.98 ;
      RECT 67.44 2.75 67.85 2.995 ;
      RECT 67.815 1.895 68.135 2.155 ;
      RECT 68.28 1.91 68.57 2.14 ;
      RECT 67.815 1.955 68.57 2.095 ;
      RECT 65.115 3.16 67.295 3.3 ;
      RECT 67.155 2.17 67.295 3.3 ;
      RECT 65.115 3.075 66.41 3.3 ;
      RECT 66.12 3.03 66.41 3.3 ;
      RECT 65.115 2.795 65.45 3.3 ;
      RECT 65.16 2.75 65.45 3.3 ;
      RECT 68.04 2.47 68.33 2.7 ;
      RECT 67.155 2.375 68.255 2.515 ;
      RECT 67.08 2.17 67.37 2.42 ;
      RECT 67.3 7.77 67.59 8 ;
      RECT 67.36 7.03 67.53 8 ;
      RECT 67.26 7.06 67.63 7.43 ;
      RECT 67.3 7.03 67.59 7.43 ;
      RECT 67.065 3.575 67.385 3.835 ;
      RECT 67.065 3.59 67.58 3.82 ;
      RECT 65.64 2.47 65.93 2.7 ;
      RECT 65.79 2.075 65.93 2.7 ;
      RECT 65.79 2.075 66.095 2.215 ;
      RECT 66.585 1.895 66.905 2.155 ;
      RECT 65.865 1.895 66.185 2.155 ;
      RECT 66.36 1.91 66.905 2.14 ;
      RECT 65.865 1.955 66.905 2.095 ;
      RECT 65.505 3.575 65.825 3.835 ;
      RECT 65.4 3.59 65.825 3.82 ;
      RECT 63.48 3.03 63.77 3.26 ;
      RECT 63.48 3.03 63.935 3.215 ;
      RECT 63.795 2.555 63.935 3.215 ;
      RECT 63.915 1.955 64.055 2.695 ;
      RECT 64.785 1.895 65.105 2.155 ;
      RECT 63.96 1.91 64.25 2.14 ;
      RECT 63.915 1.955 65.105 2.095 ;
      RECT 64.665 2.455 64.985 2.715 ;
      RECT 64.2 2.47 64.49 2.7 ;
      RECT 64.2 2.515 64.985 2.655 ;
      RECT 64.425 3.015 64.745 3.275 ;
      RECT 64.425 3.03 64.97 3.26 ;
      RECT 63.96 3.59 64.25 3.82 ;
      RECT 63.075 3.47 64.175 3.61 ;
      RECT 63 3.31 63.29 3.54 ;
      RECT 60.44 7.77 60.73 8 ;
      RECT 60.5 6.29 60.67 8 ;
      RECT 60.445 6.66 60.795 7.01 ;
      RECT 60.44 6.29 60.73 6.52 ;
      RECT 60.44 2.37 60.73 2.6 ;
      RECT 60.5 0.89 60.67 2.6 ;
      RECT 60.44 0.89 60.73 1.12 ;
      RECT 60.03 2.74 60.36 2.97 ;
      RECT 60.03 2.77 60.53 2.94 ;
      RECT 60.03 2.4 60.22 2.97 ;
      RECT 59.45 2.37 59.74 2.6 ;
      RECT 59.45 2.4 60.22 2.57 ;
      RECT 59.51 0.89 59.68 2.6 ;
      RECT 59.45 0.89 59.74 1.12 ;
      RECT 59.45 7.77 59.74 8 ;
      RECT 59.51 6.29 59.68 8 ;
      RECT 59.45 6.29 59.74 6.52 ;
      RECT 59.45 6.33 60.3 6.49 ;
      RECT 60.13 5.92 60.3 6.49 ;
      RECT 59.45 6.325 59.84 6.49 ;
      RECT 60.07 5.92 60.36 6.15 ;
      RECT 60.07 5.95 60.53 6.12 ;
      RECT 59.08 2.74 59.37 2.97 ;
      RECT 59.08 2.77 59.54 2.94 ;
      RECT 59.14 1.66 59.305 2.97 ;
      RECT 57.655 1.63 57.945 1.86 ;
      RECT 57.655 1.66 59.305 1.83 ;
      RECT 57.715 0.89 57.885 1.86 ;
      RECT 57.655 0.89 57.945 1.12 ;
      RECT 57.655 7.77 57.945 8 ;
      RECT 57.715 7.03 57.885 8 ;
      RECT 57.715 7.125 59.305 7.295 ;
      RECT 59.135 5.92 59.305 7.295 ;
      RECT 57.655 7.03 57.945 7.26 ;
      RECT 59.08 5.92 59.37 6.15 ;
      RECT 59.08 5.95 59.54 6.12 ;
      RECT 55.705 2.705 56.045 3.055 ;
      RECT 55.795 2.03 55.965 3.055 ;
      RECT 58.085 1.97 58.435 2.32 ;
      RECT 55.795 2.03 58.435 2.2 ;
      RECT 58.11 6.66 58.435 6.985 ;
      RECT 52.675 6.615 53.025 6.965 ;
      RECT 58.085 6.66 58.435 6.89 ;
      RECT 52.47 6.66 53.025 6.89 ;
      RECT 52.3 6.69 58.435 6.86 ;
      RECT 57.31 2.37 57.63 2.69 ;
      RECT 57.28 2.37 57.63 2.6 ;
      RECT 57.11 2.4 57.63 2.57 ;
      RECT 57.31 6.26 57.63 6.55 ;
      RECT 57.28 6.29 57.63 6.52 ;
      RECT 57.11 6.32 57.63 6.49 ;
      RECT 56.265 2.71 56.605 3.06 ;
      RECT 56.265 2.77 56.745 2.94 ;
      RECT 56.265 5.865 56.605 6.215 ;
      RECT 50.67 5.92 50.96 6.15 ;
      RECT 50.67 5.95 56.745 6.12 ;
      RECT 54.415 1.895 54.735 2.155 ;
      RECT 53.98 1.91 54.27 2.14 ;
      RECT 53.98 1.955 54.735 2.095 ;
      RECT 54.415 3.575 54.735 3.835 ;
      RECT 53.98 3.59 54.27 3.82 ;
      RECT 53.98 3.635 54.735 3.775 ;
      RECT 53.74 3.03 54.03 3.26 ;
      RECT 53.74 3.075 54.315 3.215 ;
      RECT 54.175 2.935 54.435 3.075 ;
      RECT 54.22 2.75 54.51 2.98 ;
      RECT 52.375 2.935 53.475 3.075 ;
      RECT 52.18 2.735 52.5 2.995 ;
      RECT 53.26 2.75 53.55 2.98 ;
      RECT 52.18 2.75 52.59 2.995 ;
      RECT 52.555 1.895 52.875 2.155 ;
      RECT 53.02 1.91 53.31 2.14 ;
      RECT 52.555 1.955 53.31 2.095 ;
      RECT 49.855 3.16 52.035 3.3 ;
      RECT 51.895 2.17 52.035 3.3 ;
      RECT 49.855 3.075 51.15 3.3 ;
      RECT 50.86 3.03 51.15 3.3 ;
      RECT 49.855 2.795 50.19 3.3 ;
      RECT 49.9 2.75 50.19 3.3 ;
      RECT 52.78 2.47 53.07 2.7 ;
      RECT 51.895 2.375 52.995 2.515 ;
      RECT 51.82 2.17 52.11 2.42 ;
      RECT 52.04 7.77 52.33 8 ;
      RECT 52.1 7.03 52.27 8 ;
      RECT 52 7.06 52.37 7.43 ;
      RECT 52.04 7.03 52.33 7.43 ;
      RECT 51.805 3.575 52.125 3.835 ;
      RECT 51.805 3.59 52.32 3.82 ;
      RECT 50.38 2.47 50.67 2.7 ;
      RECT 50.53 2.075 50.67 2.7 ;
      RECT 50.53 2.075 50.835 2.215 ;
      RECT 51.325 1.895 51.645 2.155 ;
      RECT 50.605 1.895 50.925 2.155 ;
      RECT 51.1 1.91 51.645 2.14 ;
      RECT 50.605 1.955 51.645 2.095 ;
      RECT 50.245 3.575 50.565 3.835 ;
      RECT 50.14 3.59 50.565 3.82 ;
      RECT 48.22 3.03 48.51 3.26 ;
      RECT 48.22 3.03 48.675 3.215 ;
      RECT 48.535 2.555 48.675 3.215 ;
      RECT 48.655 1.955 48.795 2.695 ;
      RECT 49.525 1.895 49.845 2.155 ;
      RECT 48.7 1.91 48.99 2.14 ;
      RECT 48.655 1.955 49.845 2.095 ;
      RECT 49.405 2.455 49.725 2.715 ;
      RECT 48.94 2.47 49.23 2.7 ;
      RECT 48.94 2.515 49.725 2.655 ;
      RECT 49.165 3.015 49.485 3.275 ;
      RECT 49.165 3.03 49.71 3.26 ;
      RECT 48.7 3.59 48.99 3.82 ;
      RECT 47.815 3.47 48.915 3.61 ;
      RECT 47.74 3.31 48.03 3.54 ;
      RECT 45.18 7.77 45.47 8 ;
      RECT 45.24 6.29 45.41 8 ;
      RECT 45.185 6.66 45.535 7.01 ;
      RECT 45.18 6.29 45.47 6.52 ;
      RECT 45.18 2.37 45.47 2.6 ;
      RECT 45.24 0.89 45.41 2.6 ;
      RECT 45.18 0.89 45.47 1.12 ;
      RECT 44.77 2.74 45.1 2.97 ;
      RECT 44.77 2.77 45.27 2.94 ;
      RECT 44.77 2.4 44.96 2.97 ;
      RECT 44.19 2.37 44.48 2.6 ;
      RECT 44.19 2.4 44.96 2.57 ;
      RECT 44.25 0.89 44.42 2.6 ;
      RECT 44.19 0.89 44.48 1.12 ;
      RECT 44.19 7.77 44.48 8 ;
      RECT 44.25 6.29 44.42 8 ;
      RECT 44.19 6.29 44.48 6.52 ;
      RECT 44.19 6.33 45.04 6.49 ;
      RECT 44.87 5.92 45.04 6.49 ;
      RECT 44.19 6.325 44.58 6.49 ;
      RECT 44.81 5.92 45.1 6.15 ;
      RECT 44.81 5.95 45.27 6.12 ;
      RECT 43.82 2.74 44.11 2.97 ;
      RECT 43.82 2.77 44.28 2.94 ;
      RECT 43.88 1.66 44.045 2.97 ;
      RECT 42.395 1.63 42.685 1.86 ;
      RECT 42.395 1.66 44.045 1.83 ;
      RECT 42.455 0.89 42.625 1.86 ;
      RECT 42.395 0.89 42.685 1.12 ;
      RECT 42.395 7.77 42.685 8 ;
      RECT 42.455 7.03 42.625 8 ;
      RECT 42.455 7.125 44.045 7.295 ;
      RECT 43.875 5.92 44.045 7.295 ;
      RECT 42.395 7.03 42.685 7.26 ;
      RECT 43.82 5.92 44.11 6.15 ;
      RECT 43.82 5.95 44.28 6.12 ;
      RECT 40.445 2.705 40.785 3.055 ;
      RECT 40.535 2.03 40.705 3.055 ;
      RECT 42.825 1.97 43.175 2.32 ;
      RECT 40.535 2.03 43.175 2.2 ;
      RECT 42.85 6.66 43.175 6.985 ;
      RECT 37.41 6.62 37.76 6.97 ;
      RECT 42.825 6.66 43.175 6.89 ;
      RECT 37.21 6.66 37.76 6.89 ;
      RECT 37.04 6.69 43.175 6.86 ;
      RECT 42.05 2.37 42.37 2.69 ;
      RECT 42.02 2.37 42.37 2.6 ;
      RECT 41.85 2.4 42.37 2.57 ;
      RECT 42.05 6.26 42.37 6.55 ;
      RECT 42.02 6.29 42.37 6.52 ;
      RECT 41.85 6.32 42.37 6.49 ;
      RECT 41.005 2.71 41.345 3.06 ;
      RECT 41.005 2.77 41.485 2.94 ;
      RECT 41.005 5.865 41.345 6.215 ;
      RECT 35.41 5.92 35.7 6.15 ;
      RECT 35.41 5.95 41.485 6.12 ;
      RECT 39.155 1.895 39.475 2.155 ;
      RECT 38.72 1.91 39.01 2.14 ;
      RECT 38.72 1.955 39.475 2.095 ;
      RECT 39.155 3.575 39.475 3.835 ;
      RECT 38.72 3.59 39.01 3.82 ;
      RECT 38.72 3.635 39.475 3.775 ;
      RECT 38.48 3.03 38.77 3.26 ;
      RECT 38.48 3.075 39.055 3.215 ;
      RECT 38.915 2.935 39.175 3.075 ;
      RECT 38.96 2.75 39.25 2.98 ;
      RECT 37.115 2.935 38.215 3.075 ;
      RECT 36.92 2.735 37.24 2.995 ;
      RECT 38 2.75 38.29 2.98 ;
      RECT 36.92 2.75 37.33 2.995 ;
      RECT 37.295 1.895 37.615 2.155 ;
      RECT 37.76 1.91 38.05 2.14 ;
      RECT 37.295 1.955 38.05 2.095 ;
      RECT 34.595 3.16 36.775 3.3 ;
      RECT 36.635 2.17 36.775 3.3 ;
      RECT 34.595 3.075 35.89 3.3 ;
      RECT 35.6 3.03 35.89 3.3 ;
      RECT 34.595 2.795 34.93 3.3 ;
      RECT 34.64 2.75 34.93 3.3 ;
      RECT 37.52 2.47 37.81 2.7 ;
      RECT 36.635 2.375 37.735 2.515 ;
      RECT 36.56 2.17 36.85 2.42 ;
      RECT 36.78 7.77 37.07 8 ;
      RECT 36.84 7.03 37.01 8 ;
      RECT 36.74 7.06 37.11 7.43 ;
      RECT 36.78 7.03 37.07 7.43 ;
      RECT 36.545 3.575 36.865 3.835 ;
      RECT 36.545 3.59 37.06 3.82 ;
      RECT 35.12 2.47 35.41 2.7 ;
      RECT 35.27 2.075 35.41 2.7 ;
      RECT 35.27 2.075 35.575 2.215 ;
      RECT 36.065 1.895 36.385 2.155 ;
      RECT 35.345 1.895 35.665 2.155 ;
      RECT 35.84 1.91 36.385 2.14 ;
      RECT 35.345 1.955 36.385 2.095 ;
      RECT 34.985 3.575 35.305 3.835 ;
      RECT 34.88 3.59 35.305 3.82 ;
      RECT 32.96 3.03 33.25 3.26 ;
      RECT 32.96 3.03 33.415 3.215 ;
      RECT 33.275 2.555 33.415 3.215 ;
      RECT 33.395 1.955 33.535 2.695 ;
      RECT 34.265 1.895 34.585 2.155 ;
      RECT 33.44 1.91 33.73 2.14 ;
      RECT 33.395 1.955 34.585 2.095 ;
      RECT 34.145 2.455 34.465 2.715 ;
      RECT 33.68 2.47 33.97 2.7 ;
      RECT 33.68 2.515 34.465 2.655 ;
      RECT 33.905 3.015 34.225 3.275 ;
      RECT 33.905 3.03 34.45 3.26 ;
      RECT 33.44 3.59 33.73 3.82 ;
      RECT 32.555 3.47 33.655 3.61 ;
      RECT 32.48 3.31 32.77 3.54 ;
      RECT 29.92 7.77 30.21 8 ;
      RECT 29.98 6.29 30.15 8 ;
      RECT 29.965 6.665 30.32 7.02 ;
      RECT 29.92 6.29 30.21 6.52 ;
      RECT 29.92 2.37 30.21 2.6 ;
      RECT 29.98 0.89 30.15 2.6 ;
      RECT 29.92 0.89 30.21 1.12 ;
      RECT 29.51 2.74 29.84 2.97 ;
      RECT 29.51 2.77 30.01 2.94 ;
      RECT 29.51 2.4 29.7 2.97 ;
      RECT 28.93 2.37 29.22 2.6 ;
      RECT 28.93 2.4 29.7 2.57 ;
      RECT 28.99 0.89 29.16 2.6 ;
      RECT 28.93 0.89 29.22 1.12 ;
      RECT 28.93 7.77 29.22 8 ;
      RECT 28.99 6.29 29.16 8 ;
      RECT 28.93 6.29 29.22 6.52 ;
      RECT 28.93 6.33 29.78 6.49 ;
      RECT 29.61 5.92 29.78 6.49 ;
      RECT 28.93 6.325 29.32 6.49 ;
      RECT 29.55 5.92 29.84 6.15 ;
      RECT 29.55 5.95 30.01 6.12 ;
      RECT 28.56 2.74 28.85 2.97 ;
      RECT 28.56 2.77 29.02 2.94 ;
      RECT 28.62 1.66 28.785 2.97 ;
      RECT 27.135 1.63 27.425 1.86 ;
      RECT 27.135 1.66 28.785 1.83 ;
      RECT 27.195 0.89 27.365 1.86 ;
      RECT 27.135 0.89 27.425 1.12 ;
      RECT 27.135 7.77 27.425 8 ;
      RECT 27.195 7.03 27.365 8 ;
      RECT 27.195 7.125 28.785 7.295 ;
      RECT 28.615 5.92 28.785 7.295 ;
      RECT 27.135 7.03 27.425 7.26 ;
      RECT 28.56 5.92 28.85 6.15 ;
      RECT 28.56 5.95 29.02 6.12 ;
      RECT 25.185 2.705 25.525 3.055 ;
      RECT 25.275 2.03 25.445 3.055 ;
      RECT 27.565 1.97 27.915 2.32 ;
      RECT 25.275 2.03 27.915 2.2 ;
      RECT 27.59 6.66 27.915 6.985 ;
      RECT 22.15 6.615 22.5 6.965 ;
      RECT 27.565 6.66 27.915 6.89 ;
      RECT 21.95 6.66 22.5 6.89 ;
      RECT 21.78 6.69 27.915 6.86 ;
      RECT 26.79 2.37 27.11 2.69 ;
      RECT 26.76 2.37 27.11 2.6 ;
      RECT 26.59 2.4 27.11 2.57 ;
      RECT 26.79 6.26 27.11 6.55 ;
      RECT 26.76 6.29 27.11 6.52 ;
      RECT 26.59 6.32 27.11 6.49 ;
      RECT 25.745 2.71 26.085 3.06 ;
      RECT 25.745 2.77 26.225 2.94 ;
      RECT 25.745 5.865 26.085 6.215 ;
      RECT 20.15 5.92 20.44 6.15 ;
      RECT 20.15 5.95 26.225 6.12 ;
      RECT 23.895 1.895 24.215 2.155 ;
      RECT 23.46 1.91 23.75 2.14 ;
      RECT 23.46 1.955 24.215 2.095 ;
      RECT 23.895 3.575 24.215 3.835 ;
      RECT 23.46 3.59 23.75 3.82 ;
      RECT 23.46 3.635 24.215 3.775 ;
      RECT 23.22 3.03 23.51 3.26 ;
      RECT 23.22 3.075 23.795 3.215 ;
      RECT 23.655 2.935 23.915 3.075 ;
      RECT 23.7 2.75 23.99 2.98 ;
      RECT 21.855 2.935 22.955 3.075 ;
      RECT 21.66 2.735 21.98 2.995 ;
      RECT 22.74 2.75 23.03 2.98 ;
      RECT 21.66 2.75 22.07 2.995 ;
      RECT 22.035 1.895 22.355 2.155 ;
      RECT 22.5 1.91 22.79 2.14 ;
      RECT 22.035 1.955 22.79 2.095 ;
      RECT 19.335 3.16 21.515 3.3 ;
      RECT 21.375 2.17 21.515 3.3 ;
      RECT 19.335 3.075 20.63 3.3 ;
      RECT 20.34 3.03 20.63 3.3 ;
      RECT 19.335 2.795 19.67 3.3 ;
      RECT 19.38 2.75 19.67 3.3 ;
      RECT 22.26 2.47 22.55 2.7 ;
      RECT 21.375 2.375 22.475 2.515 ;
      RECT 21.3 2.17 21.59 2.42 ;
      RECT 21.52 7.77 21.81 8 ;
      RECT 21.58 7.03 21.75 8 ;
      RECT 21.48 7.06 21.85 7.43 ;
      RECT 21.52 7.03 21.81 7.43 ;
      RECT 21.285 3.575 21.605 3.835 ;
      RECT 21.285 3.59 21.8 3.82 ;
      RECT 19.86 2.47 20.15 2.7 ;
      RECT 20.01 2.075 20.15 2.7 ;
      RECT 20.01 2.075 20.315 2.215 ;
      RECT 20.805 1.895 21.125 2.155 ;
      RECT 20.085 1.895 20.405 2.155 ;
      RECT 20.58 1.91 21.125 2.14 ;
      RECT 20.085 1.955 21.125 2.095 ;
      RECT 19.725 3.575 20.045 3.835 ;
      RECT 19.62 3.59 20.045 3.82 ;
      RECT 17.7 3.03 17.99 3.26 ;
      RECT 17.7 3.03 18.155 3.215 ;
      RECT 18.015 2.555 18.155 3.215 ;
      RECT 18.135 1.955 18.275 2.695 ;
      RECT 19.005 1.895 19.325 2.155 ;
      RECT 18.18 1.91 18.47 2.14 ;
      RECT 18.135 1.955 19.325 2.095 ;
      RECT 18.885 2.455 19.205 2.715 ;
      RECT 18.42 2.47 18.71 2.7 ;
      RECT 18.42 2.515 19.205 2.655 ;
      RECT 18.645 3.015 18.965 3.275 ;
      RECT 18.645 3.03 19.19 3.26 ;
      RECT 18.18 3.59 18.47 3.82 ;
      RECT 17.295 3.47 18.395 3.61 ;
      RECT 17.22 3.31 17.51 3.54 ;
      RECT 14.66 7.77 14.95 8 ;
      RECT 14.72 6.29 14.89 8 ;
      RECT 14.71 6.66 15.06 7.01 ;
      RECT 14.66 6.29 14.95 6.52 ;
      RECT 14.66 2.37 14.95 2.6 ;
      RECT 14.72 0.89 14.89 2.6 ;
      RECT 14.66 0.89 14.95 1.12 ;
      RECT 14.25 2.74 14.58 2.97 ;
      RECT 14.25 2.77 14.75 2.94 ;
      RECT 14.25 2.4 14.44 2.97 ;
      RECT 13.67 2.37 13.96 2.6 ;
      RECT 13.67 2.4 14.44 2.57 ;
      RECT 13.73 0.89 13.9 2.6 ;
      RECT 13.67 0.89 13.96 1.12 ;
      RECT 13.67 7.77 13.96 8 ;
      RECT 13.73 6.29 13.9 8 ;
      RECT 13.67 6.29 13.96 6.52 ;
      RECT 13.67 6.33 14.52 6.49 ;
      RECT 14.35 5.92 14.52 6.49 ;
      RECT 13.67 6.325 14.06 6.49 ;
      RECT 14.29 5.92 14.58 6.15 ;
      RECT 14.29 5.95 14.75 6.12 ;
      RECT 13.3 2.74 13.59 2.97 ;
      RECT 13.3 2.77 13.76 2.94 ;
      RECT 13.36 1.66 13.525 2.97 ;
      RECT 11.875 1.63 12.165 1.86 ;
      RECT 11.875 1.66 13.525 1.83 ;
      RECT 11.935 0.89 12.105 1.86 ;
      RECT 11.875 0.89 12.165 1.12 ;
      RECT 11.875 7.77 12.165 8 ;
      RECT 11.935 7.03 12.105 8 ;
      RECT 11.935 7.125 13.525 7.295 ;
      RECT 13.355 5.92 13.525 7.295 ;
      RECT 11.875 7.03 12.165 7.26 ;
      RECT 13.3 5.92 13.59 6.15 ;
      RECT 13.3 5.95 13.76 6.12 ;
      RECT 9.925 2.705 10.265 3.055 ;
      RECT 10.015 2.03 10.185 3.055 ;
      RECT 12.305 1.97 12.655 2.32 ;
      RECT 10.015 2.03 12.655 2.2 ;
      RECT 12.33 6.66 12.655 6.985 ;
      RECT 6.89 6.61 7.24 6.96 ;
      RECT 12.305 6.66 12.655 6.89 ;
      RECT 6.69 6.66 7.24 6.89 ;
      RECT 6.52 6.69 12.655 6.86 ;
      RECT 11.53 2.37 11.85 2.69 ;
      RECT 11.5 2.37 11.85 2.6 ;
      RECT 11.33 2.4 11.85 2.57 ;
      RECT 11.53 6.26 11.85 6.55 ;
      RECT 11.5 6.29 11.85 6.52 ;
      RECT 11.33 6.32 11.85 6.49 ;
      RECT 10.485 2.71 10.825 3.06 ;
      RECT 10.485 2.77 10.965 2.94 ;
      RECT 10.485 5.865 10.825 6.215 ;
      RECT 4.89 5.92 5.18 6.15 ;
      RECT 4.89 5.95 10.965 6.12 ;
      RECT 8.635 1.895 8.955 2.155 ;
      RECT 8.2 1.91 8.49 2.14 ;
      RECT 8.2 1.955 8.955 2.095 ;
      RECT 8.635 3.575 8.955 3.835 ;
      RECT 8.2 3.59 8.49 3.82 ;
      RECT 8.2 3.635 8.955 3.775 ;
      RECT 7.96 3.03 8.25 3.26 ;
      RECT 7.96 3.075 8.535 3.215 ;
      RECT 8.395 2.935 8.655 3.075 ;
      RECT 8.44 2.75 8.73 2.98 ;
      RECT 6.595 2.935 7.695 3.075 ;
      RECT 6.4 2.735 6.72 2.995 ;
      RECT 7.48 2.75 7.77 2.98 ;
      RECT 6.4 2.75 6.81 2.995 ;
      RECT 6.775 1.895 7.095 2.155 ;
      RECT 7.24 1.91 7.53 2.14 ;
      RECT 6.775 1.955 7.53 2.095 ;
      RECT 4.075 3.16 6.255 3.3 ;
      RECT 6.115 2.17 6.255 3.3 ;
      RECT 4.075 3.075 5.37 3.3 ;
      RECT 5.08 3.03 5.37 3.3 ;
      RECT 4.075 2.795 4.41 3.3 ;
      RECT 4.12 2.75 4.41 3.3 ;
      RECT 7 2.47 7.29 2.7 ;
      RECT 6.115 2.375 7.215 2.515 ;
      RECT 6.04 2.17 6.33 2.42 ;
      RECT 6.26 7.77 6.55 8 ;
      RECT 6.32 7.03 6.49 8 ;
      RECT 6.22 7.06 6.59 7.43 ;
      RECT 6.26 7.03 6.55 7.43 ;
      RECT 6.025 3.575 6.345 3.835 ;
      RECT 6.025 3.59 6.54 3.82 ;
      RECT 4.6 2.47 4.89 2.7 ;
      RECT 4.75 2.075 4.89 2.7 ;
      RECT 4.75 2.075 5.055 2.215 ;
      RECT 5.545 1.895 5.865 2.155 ;
      RECT 4.825 1.895 5.145 2.155 ;
      RECT 5.32 1.91 5.865 2.14 ;
      RECT 4.825 1.955 5.865 2.095 ;
      RECT 4.465 3.575 4.785 3.835 ;
      RECT 4.36 3.59 4.785 3.82 ;
      RECT 2.44 3.03 2.73 3.26 ;
      RECT 2.44 3.03 2.895 3.215 ;
      RECT 2.755 2.555 2.895 3.215 ;
      RECT 2.875 1.955 3.015 2.695 ;
      RECT 3.745 1.895 4.065 2.155 ;
      RECT 2.92 1.91 3.21 2.14 ;
      RECT 2.875 1.955 4.065 2.095 ;
      RECT 3.625 2.455 3.945 2.715 ;
      RECT 3.16 2.47 3.45 2.7 ;
      RECT 3.16 2.515 3.945 2.655 ;
      RECT 3.385 3.015 3.705 3.275 ;
      RECT 3.385 3.03 3.93 3.26 ;
      RECT 2.92 3.59 3.21 3.82 ;
      RECT 2.035 3.47 3.135 3.61 ;
      RECT 1.96 3.31 2.25 3.54 ;
      RECT -0.825 6.66 -0.535 6.89 ;
      RECT -0.995 6.69 -0.535 6.86 ;
      RECT -1.255 7.77 -0.965 8 ;
      RECT -1.195 7.03 -1.025 8 ;
      RECT -1.285 7.03 -0.935 7.32 ;
      RECT -1.66 6.29 -1.31 6.58 ;
      RECT -1.8 6.32 -1.31 6.49 ;
      RECT -2.625 5.92 -2.335 6.15 ;
      RECT -2.625 5.95 -2.165 6.12 ;
      RECT 68.985 2.455 69.305 2.715 ;
      RECT 67.815 3.295 68.135 3.555 ;
      RECT 66.585 2.735 66.905 2.995 ;
      RECT 66.105 2.455 66.425 2.715 ;
      RECT 65.25 1.895 65.65 2.155 ;
      RECT 64.905 3.575 65.225 3.835 ;
      RECT 63.225 2.455 63.545 2.715 ;
      RECT 62.745 2.735 63.065 2.995 ;
      RECT 62.055 1.895 62.375 2.155 ;
      RECT 62.055 3.295 62.375 3.555 ;
      RECT 53.725 2.455 54.045 2.715 ;
      RECT 52.555 3.295 52.875 3.555 ;
      RECT 51.325 2.735 51.645 2.995 ;
      RECT 50.845 2.455 51.165 2.715 ;
      RECT 49.99 1.895 50.39 2.155 ;
      RECT 49.645 3.575 49.965 3.835 ;
      RECT 47.965 2.455 48.285 2.715 ;
      RECT 47.485 2.735 47.805 2.995 ;
      RECT 46.795 1.895 47.115 2.155 ;
      RECT 46.795 3.295 47.115 3.555 ;
      RECT 38.465 2.455 38.785 2.715 ;
      RECT 37.295 3.295 37.615 3.555 ;
      RECT 36.065 2.735 36.385 2.995 ;
      RECT 35.585 2.455 35.905 2.715 ;
      RECT 34.73 1.895 35.13 2.155 ;
      RECT 34.385 3.575 34.705 3.835 ;
      RECT 32.705 2.455 33.025 2.715 ;
      RECT 32.225 2.735 32.545 2.995 ;
      RECT 31.535 1.895 31.855 2.155 ;
      RECT 31.535 3.295 31.855 3.555 ;
      RECT 23.205 2.455 23.525 2.715 ;
      RECT 22.035 3.295 22.355 3.555 ;
      RECT 20.805 2.735 21.125 2.995 ;
      RECT 20.325 2.455 20.645 2.715 ;
      RECT 19.47 1.895 19.87 2.155 ;
      RECT 19.125 3.575 19.445 3.835 ;
      RECT 17.445 2.455 17.765 2.715 ;
      RECT 16.965 2.735 17.285 2.995 ;
      RECT 16.275 1.895 16.595 2.155 ;
      RECT 16.275 3.295 16.595 3.555 ;
      RECT 7.945 2.455 8.265 2.715 ;
      RECT 6.775 3.295 7.095 3.555 ;
      RECT 5.545 2.735 5.865 2.995 ;
      RECT 5.065 2.455 5.385 2.715 ;
      RECT 4.21 1.895 4.61 2.155 ;
      RECT 3.865 3.575 4.185 3.835 ;
      RECT 2.185 2.455 2.505 2.715 ;
      RECT 1.705 2.735 2.025 2.995 ;
      RECT 1.015 1.895 1.335 2.155 ;
      RECT 1.015 3.295 1.335 3.555 ;
    LAYER mcon ;
      RECT 75.76 0.92 75.93 1.09 ;
      RECT 75.76 2.4 75.93 2.57 ;
      RECT 75.76 6.32 75.93 6.49 ;
      RECT 75.76 7.8 75.93 7.97 ;
      RECT 75.41 0.11 75.58 0.28 ;
      RECT 75.41 4.17 75.58 4.34 ;
      RECT 75.41 4.55 75.58 4.72 ;
      RECT 75.41 8.61 75.58 8.78 ;
      RECT 75.39 2.77 75.56 2.94 ;
      RECT 75.39 5.95 75.56 6.12 ;
      RECT 74.77 0.92 74.94 1.09 ;
      RECT 74.77 2.4 74.94 2.57 ;
      RECT 74.77 6.32 74.94 6.49 ;
      RECT 74.77 7.8 74.94 7.97 ;
      RECT 74.42 0.11 74.59 0.28 ;
      RECT 74.42 4.17 74.59 4.34 ;
      RECT 74.42 4.55 74.59 4.72 ;
      RECT 74.42 8.61 74.59 8.78 ;
      RECT 74.4 2.77 74.57 2.94 ;
      RECT 74.4 5.95 74.57 6.12 ;
      RECT 73.715 0.11 73.885 0.28 ;
      RECT 73.715 4.17 73.885 4.34 ;
      RECT 73.715 4.55 73.885 4.72 ;
      RECT 73.715 8.61 73.885 8.78 ;
      RECT 73.405 2.03 73.575 2.2 ;
      RECT 73.405 6.69 73.575 6.86 ;
      RECT 73.035 0.11 73.205 0.28 ;
      RECT 73.035 8.61 73.205 8.78 ;
      RECT 72.975 0.92 73.145 1.09 ;
      RECT 72.975 1.66 73.145 1.83 ;
      RECT 72.975 7.06 73.145 7.23 ;
      RECT 72.975 7.8 73.145 7.97 ;
      RECT 72.6 2.4 72.77 2.57 ;
      RECT 72.6 6.32 72.77 6.49 ;
      RECT 72.355 0.11 72.525 0.28 ;
      RECT 72.355 8.61 72.525 8.78 ;
      RECT 71.675 0.11 71.845 0.28 ;
      RECT 71.675 8.61 71.845 8.78 ;
      RECT 71.605 2.77 71.775 2.94 ;
      RECT 71.605 5.95 71.775 6.12 ;
      RECT 70.215 1.42 70.385 1.59 ;
      RECT 70.215 4.14 70.385 4.31 ;
      RECT 69.755 1.42 69.925 1.59 ;
      RECT 69.755 4.14 69.925 4.31 ;
      RECT 69.54 2.78 69.71 2.95 ;
      RECT 69.3 1.94 69.47 2.11 ;
      RECT 69.3 3.62 69.47 3.79 ;
      RECT 69.295 1.42 69.465 1.59 ;
      RECT 69.295 4.14 69.465 4.31 ;
      RECT 69.06 2.5 69.23 2.67 ;
      RECT 69.06 3.06 69.23 3.23 ;
      RECT 68.835 1.42 69.005 1.59 ;
      RECT 68.835 4.14 69.005 4.31 ;
      RECT 68.58 2.78 68.75 2.95 ;
      RECT 68.375 1.42 68.545 1.59 ;
      RECT 68.375 4.14 68.545 4.31 ;
      RECT 68.34 1.94 68.51 2.11 ;
      RECT 68.1 2.5 68.27 2.67 ;
      RECT 68.1 4.55 68.27 4.72 ;
      RECT 68.1 8.61 68.27 8.78 ;
      RECT 67.915 1.42 68.085 1.59 ;
      RECT 67.915 4.14 68.085 4.31 ;
      RECT 67.89 3.34 68.06 3.51 ;
      RECT 67.79 6.69 67.96 6.86 ;
      RECT 67.62 2.78 67.79 2.95 ;
      RECT 67.455 1.42 67.625 1.59 ;
      RECT 67.455 4.14 67.625 4.31 ;
      RECT 67.42 8.61 67.59 8.78 ;
      RECT 67.36 7.06 67.53 7.23 ;
      RECT 67.36 7.8 67.53 7.97 ;
      RECT 67.35 3.62 67.52 3.79 ;
      RECT 67.14 2.2 67.31 2.37 ;
      RECT 66.995 1.42 67.165 1.59 ;
      RECT 66.995 4.14 67.165 4.31 ;
      RECT 66.985 6.32 67.155 6.49 ;
      RECT 66.74 8.61 66.91 8.78 ;
      RECT 66.66 2.78 66.83 2.95 ;
      RECT 66.535 1.42 66.705 1.59 ;
      RECT 66.535 4.14 66.705 4.31 ;
      RECT 66.42 1.94 66.59 2.11 ;
      RECT 66.18 2.5 66.35 2.67 ;
      RECT 66.18 3.06 66.35 3.23 ;
      RECT 66.075 1.42 66.245 1.59 ;
      RECT 66.075 4.14 66.245 4.31 ;
      RECT 66.06 8.61 66.23 8.78 ;
      RECT 65.99 5.95 66.16 6.12 ;
      RECT 65.7 2.5 65.87 2.67 ;
      RECT 65.615 1.42 65.785 1.59 ;
      RECT 65.615 4.14 65.785 4.31 ;
      RECT 65.46 3.62 65.63 3.79 ;
      RECT 65.42 1.94 65.59 2.11 ;
      RECT 65.22 2.78 65.39 2.95 ;
      RECT 65.155 1.42 65.325 1.59 ;
      RECT 65.155 4.14 65.325 4.31 ;
      RECT 64.98 3.62 65.15 3.79 ;
      RECT 64.74 3.06 64.91 3.23 ;
      RECT 64.695 1.42 64.865 1.59 ;
      RECT 64.695 4.14 64.865 4.31 ;
      RECT 64.26 2.5 64.43 2.67 ;
      RECT 64.235 1.42 64.405 1.59 ;
      RECT 64.235 4.14 64.405 4.31 ;
      RECT 64.02 1.94 64.19 2.11 ;
      RECT 64.02 3.62 64.19 3.79 ;
      RECT 63.775 1.42 63.945 1.59 ;
      RECT 63.775 4.14 63.945 4.31 ;
      RECT 63.54 1.94 63.71 2.11 ;
      RECT 63.54 3.06 63.71 3.23 ;
      RECT 63.315 1.42 63.485 1.59 ;
      RECT 63.315 4.14 63.485 4.31 ;
      RECT 63.3 2.5 63.47 2.67 ;
      RECT 63.06 3.34 63.23 3.51 ;
      RECT 62.855 1.42 63.025 1.59 ;
      RECT 62.855 4.14 63.025 4.31 ;
      RECT 62.82 2.78 62.99 2.95 ;
      RECT 62.395 1.42 62.565 1.59 ;
      RECT 62.395 4.14 62.565 4.31 ;
      RECT 62.34 2.78 62.51 2.95 ;
      RECT 62.13 1.94 62.3 2.11 ;
      RECT 62.13 3.34 62.3 3.51 ;
      RECT 61.935 1.42 62.105 1.59 ;
      RECT 61.935 4.14 62.105 4.31 ;
      RECT 60.5 0.92 60.67 1.09 ;
      RECT 60.5 2.4 60.67 2.57 ;
      RECT 60.5 6.32 60.67 6.49 ;
      RECT 60.5 7.8 60.67 7.97 ;
      RECT 60.15 0.11 60.32 0.28 ;
      RECT 60.15 4.17 60.32 4.34 ;
      RECT 60.15 4.55 60.32 4.72 ;
      RECT 60.15 8.61 60.32 8.78 ;
      RECT 60.13 2.77 60.3 2.94 ;
      RECT 60.13 5.95 60.3 6.12 ;
      RECT 59.51 0.92 59.68 1.09 ;
      RECT 59.51 2.4 59.68 2.57 ;
      RECT 59.51 6.32 59.68 6.49 ;
      RECT 59.51 7.8 59.68 7.97 ;
      RECT 59.16 0.11 59.33 0.28 ;
      RECT 59.16 4.17 59.33 4.34 ;
      RECT 59.16 4.55 59.33 4.72 ;
      RECT 59.16 8.61 59.33 8.78 ;
      RECT 59.14 2.77 59.31 2.94 ;
      RECT 59.14 5.95 59.31 6.12 ;
      RECT 58.455 0.11 58.625 0.28 ;
      RECT 58.455 4.17 58.625 4.34 ;
      RECT 58.455 4.55 58.625 4.72 ;
      RECT 58.455 8.61 58.625 8.78 ;
      RECT 58.145 2.03 58.315 2.2 ;
      RECT 58.145 6.69 58.315 6.86 ;
      RECT 57.775 0.11 57.945 0.28 ;
      RECT 57.775 8.61 57.945 8.78 ;
      RECT 57.715 0.92 57.885 1.09 ;
      RECT 57.715 1.66 57.885 1.83 ;
      RECT 57.715 7.06 57.885 7.23 ;
      RECT 57.715 7.8 57.885 7.97 ;
      RECT 57.34 2.4 57.51 2.57 ;
      RECT 57.34 6.32 57.51 6.49 ;
      RECT 57.095 0.11 57.265 0.28 ;
      RECT 57.095 8.61 57.265 8.78 ;
      RECT 56.415 0.11 56.585 0.28 ;
      RECT 56.415 8.61 56.585 8.78 ;
      RECT 56.345 2.77 56.515 2.94 ;
      RECT 56.345 5.95 56.515 6.12 ;
      RECT 54.955 1.42 55.125 1.59 ;
      RECT 54.955 4.14 55.125 4.31 ;
      RECT 54.495 1.42 54.665 1.59 ;
      RECT 54.495 4.14 54.665 4.31 ;
      RECT 54.28 2.78 54.45 2.95 ;
      RECT 54.04 1.94 54.21 2.11 ;
      RECT 54.04 3.62 54.21 3.79 ;
      RECT 54.035 1.42 54.205 1.59 ;
      RECT 54.035 4.14 54.205 4.31 ;
      RECT 53.8 2.5 53.97 2.67 ;
      RECT 53.8 3.06 53.97 3.23 ;
      RECT 53.575 1.42 53.745 1.59 ;
      RECT 53.575 4.14 53.745 4.31 ;
      RECT 53.32 2.78 53.49 2.95 ;
      RECT 53.115 1.42 53.285 1.59 ;
      RECT 53.115 4.14 53.285 4.31 ;
      RECT 53.08 1.94 53.25 2.11 ;
      RECT 52.84 2.5 53.01 2.67 ;
      RECT 52.84 4.55 53.01 4.72 ;
      RECT 52.84 8.61 53.01 8.78 ;
      RECT 52.655 1.42 52.825 1.59 ;
      RECT 52.655 4.14 52.825 4.31 ;
      RECT 52.63 3.34 52.8 3.51 ;
      RECT 52.53 6.69 52.7 6.86 ;
      RECT 52.36 2.78 52.53 2.95 ;
      RECT 52.195 1.42 52.365 1.59 ;
      RECT 52.195 4.14 52.365 4.31 ;
      RECT 52.16 8.61 52.33 8.78 ;
      RECT 52.1 7.06 52.27 7.23 ;
      RECT 52.1 7.8 52.27 7.97 ;
      RECT 52.09 3.62 52.26 3.79 ;
      RECT 51.88 2.2 52.05 2.37 ;
      RECT 51.735 1.42 51.905 1.59 ;
      RECT 51.735 4.14 51.905 4.31 ;
      RECT 51.725 6.32 51.895 6.49 ;
      RECT 51.48 8.61 51.65 8.78 ;
      RECT 51.4 2.78 51.57 2.95 ;
      RECT 51.275 1.42 51.445 1.59 ;
      RECT 51.275 4.14 51.445 4.31 ;
      RECT 51.16 1.94 51.33 2.11 ;
      RECT 50.92 2.5 51.09 2.67 ;
      RECT 50.92 3.06 51.09 3.23 ;
      RECT 50.815 1.42 50.985 1.59 ;
      RECT 50.815 4.14 50.985 4.31 ;
      RECT 50.8 8.61 50.97 8.78 ;
      RECT 50.73 5.95 50.9 6.12 ;
      RECT 50.44 2.5 50.61 2.67 ;
      RECT 50.355 1.42 50.525 1.59 ;
      RECT 50.355 4.14 50.525 4.31 ;
      RECT 50.2 3.62 50.37 3.79 ;
      RECT 50.16 1.94 50.33 2.11 ;
      RECT 49.96 2.78 50.13 2.95 ;
      RECT 49.895 1.42 50.065 1.59 ;
      RECT 49.895 4.14 50.065 4.31 ;
      RECT 49.72 3.62 49.89 3.79 ;
      RECT 49.48 3.06 49.65 3.23 ;
      RECT 49.435 1.42 49.605 1.59 ;
      RECT 49.435 4.14 49.605 4.31 ;
      RECT 49 2.5 49.17 2.67 ;
      RECT 48.975 1.42 49.145 1.59 ;
      RECT 48.975 4.14 49.145 4.31 ;
      RECT 48.76 1.94 48.93 2.11 ;
      RECT 48.76 3.62 48.93 3.79 ;
      RECT 48.515 1.42 48.685 1.59 ;
      RECT 48.515 4.14 48.685 4.31 ;
      RECT 48.28 1.94 48.45 2.11 ;
      RECT 48.28 3.06 48.45 3.23 ;
      RECT 48.055 1.42 48.225 1.59 ;
      RECT 48.055 4.14 48.225 4.31 ;
      RECT 48.04 2.5 48.21 2.67 ;
      RECT 47.8 3.34 47.97 3.51 ;
      RECT 47.595 1.42 47.765 1.59 ;
      RECT 47.595 4.14 47.765 4.31 ;
      RECT 47.56 2.78 47.73 2.95 ;
      RECT 47.135 1.42 47.305 1.59 ;
      RECT 47.135 4.14 47.305 4.31 ;
      RECT 47.08 2.78 47.25 2.95 ;
      RECT 46.87 1.94 47.04 2.11 ;
      RECT 46.87 3.34 47.04 3.51 ;
      RECT 46.675 1.42 46.845 1.59 ;
      RECT 46.675 4.14 46.845 4.31 ;
      RECT 45.24 0.92 45.41 1.09 ;
      RECT 45.24 2.4 45.41 2.57 ;
      RECT 45.24 6.32 45.41 6.49 ;
      RECT 45.24 7.8 45.41 7.97 ;
      RECT 44.89 0.11 45.06 0.28 ;
      RECT 44.89 4.17 45.06 4.34 ;
      RECT 44.89 4.55 45.06 4.72 ;
      RECT 44.89 8.61 45.06 8.78 ;
      RECT 44.87 2.77 45.04 2.94 ;
      RECT 44.87 5.95 45.04 6.12 ;
      RECT 44.25 0.92 44.42 1.09 ;
      RECT 44.25 2.4 44.42 2.57 ;
      RECT 44.25 6.32 44.42 6.49 ;
      RECT 44.25 7.8 44.42 7.97 ;
      RECT 43.9 0.11 44.07 0.28 ;
      RECT 43.9 4.17 44.07 4.34 ;
      RECT 43.9 4.55 44.07 4.72 ;
      RECT 43.9 8.61 44.07 8.78 ;
      RECT 43.88 2.77 44.05 2.94 ;
      RECT 43.88 5.95 44.05 6.12 ;
      RECT 43.195 0.11 43.365 0.28 ;
      RECT 43.195 4.17 43.365 4.34 ;
      RECT 43.195 4.55 43.365 4.72 ;
      RECT 43.195 8.61 43.365 8.78 ;
      RECT 42.885 2.03 43.055 2.2 ;
      RECT 42.885 6.69 43.055 6.86 ;
      RECT 42.515 0.11 42.685 0.28 ;
      RECT 42.515 8.61 42.685 8.78 ;
      RECT 42.455 0.92 42.625 1.09 ;
      RECT 42.455 1.66 42.625 1.83 ;
      RECT 42.455 7.06 42.625 7.23 ;
      RECT 42.455 7.8 42.625 7.97 ;
      RECT 42.08 2.4 42.25 2.57 ;
      RECT 42.08 6.32 42.25 6.49 ;
      RECT 41.835 0.11 42.005 0.28 ;
      RECT 41.835 8.61 42.005 8.78 ;
      RECT 41.155 0.11 41.325 0.28 ;
      RECT 41.155 8.61 41.325 8.78 ;
      RECT 41.085 2.77 41.255 2.94 ;
      RECT 41.085 5.95 41.255 6.12 ;
      RECT 39.695 1.42 39.865 1.59 ;
      RECT 39.695 4.14 39.865 4.31 ;
      RECT 39.235 1.42 39.405 1.59 ;
      RECT 39.235 4.14 39.405 4.31 ;
      RECT 39.02 2.78 39.19 2.95 ;
      RECT 38.78 1.94 38.95 2.11 ;
      RECT 38.78 3.62 38.95 3.79 ;
      RECT 38.775 1.42 38.945 1.59 ;
      RECT 38.775 4.14 38.945 4.31 ;
      RECT 38.54 2.5 38.71 2.67 ;
      RECT 38.54 3.06 38.71 3.23 ;
      RECT 38.315 1.42 38.485 1.59 ;
      RECT 38.315 4.14 38.485 4.31 ;
      RECT 38.06 2.78 38.23 2.95 ;
      RECT 37.855 1.42 38.025 1.59 ;
      RECT 37.855 4.14 38.025 4.31 ;
      RECT 37.82 1.94 37.99 2.11 ;
      RECT 37.58 2.5 37.75 2.67 ;
      RECT 37.58 4.55 37.75 4.72 ;
      RECT 37.58 8.61 37.75 8.78 ;
      RECT 37.395 1.42 37.565 1.59 ;
      RECT 37.395 4.14 37.565 4.31 ;
      RECT 37.37 3.34 37.54 3.51 ;
      RECT 37.27 6.69 37.44 6.86 ;
      RECT 37.1 2.78 37.27 2.95 ;
      RECT 36.935 1.42 37.105 1.59 ;
      RECT 36.935 4.14 37.105 4.31 ;
      RECT 36.9 8.61 37.07 8.78 ;
      RECT 36.84 7.06 37.01 7.23 ;
      RECT 36.84 7.8 37.01 7.97 ;
      RECT 36.83 3.62 37 3.79 ;
      RECT 36.62 2.2 36.79 2.37 ;
      RECT 36.475 1.42 36.645 1.59 ;
      RECT 36.475 4.14 36.645 4.31 ;
      RECT 36.465 6.32 36.635 6.49 ;
      RECT 36.22 8.61 36.39 8.78 ;
      RECT 36.14 2.78 36.31 2.95 ;
      RECT 36.015 1.42 36.185 1.59 ;
      RECT 36.015 4.14 36.185 4.31 ;
      RECT 35.9 1.94 36.07 2.11 ;
      RECT 35.66 2.5 35.83 2.67 ;
      RECT 35.66 3.06 35.83 3.23 ;
      RECT 35.555 1.42 35.725 1.59 ;
      RECT 35.555 4.14 35.725 4.31 ;
      RECT 35.54 8.61 35.71 8.78 ;
      RECT 35.47 5.95 35.64 6.12 ;
      RECT 35.18 2.5 35.35 2.67 ;
      RECT 35.095 1.42 35.265 1.59 ;
      RECT 35.095 4.14 35.265 4.31 ;
      RECT 34.94 3.62 35.11 3.79 ;
      RECT 34.9 1.94 35.07 2.11 ;
      RECT 34.7 2.78 34.87 2.95 ;
      RECT 34.635 1.42 34.805 1.59 ;
      RECT 34.635 4.14 34.805 4.31 ;
      RECT 34.46 3.62 34.63 3.79 ;
      RECT 34.22 3.06 34.39 3.23 ;
      RECT 34.175 1.42 34.345 1.59 ;
      RECT 34.175 4.14 34.345 4.31 ;
      RECT 33.74 2.5 33.91 2.67 ;
      RECT 33.715 1.42 33.885 1.59 ;
      RECT 33.715 4.14 33.885 4.31 ;
      RECT 33.5 1.94 33.67 2.11 ;
      RECT 33.5 3.62 33.67 3.79 ;
      RECT 33.255 1.42 33.425 1.59 ;
      RECT 33.255 4.14 33.425 4.31 ;
      RECT 33.02 1.94 33.19 2.11 ;
      RECT 33.02 3.06 33.19 3.23 ;
      RECT 32.795 1.42 32.965 1.59 ;
      RECT 32.795 4.14 32.965 4.31 ;
      RECT 32.78 2.5 32.95 2.67 ;
      RECT 32.54 3.34 32.71 3.51 ;
      RECT 32.335 1.42 32.505 1.59 ;
      RECT 32.335 4.14 32.505 4.31 ;
      RECT 32.3 2.78 32.47 2.95 ;
      RECT 31.875 1.42 32.045 1.59 ;
      RECT 31.875 4.14 32.045 4.31 ;
      RECT 31.82 2.78 31.99 2.95 ;
      RECT 31.61 1.94 31.78 2.11 ;
      RECT 31.61 3.34 31.78 3.51 ;
      RECT 31.415 1.42 31.585 1.59 ;
      RECT 31.415 4.14 31.585 4.31 ;
      RECT 29.98 0.92 30.15 1.09 ;
      RECT 29.98 2.4 30.15 2.57 ;
      RECT 29.98 6.32 30.15 6.49 ;
      RECT 29.98 7.8 30.15 7.97 ;
      RECT 29.63 0.11 29.8 0.28 ;
      RECT 29.63 4.17 29.8 4.34 ;
      RECT 29.63 4.55 29.8 4.72 ;
      RECT 29.63 8.61 29.8 8.78 ;
      RECT 29.61 2.77 29.78 2.94 ;
      RECT 29.61 5.95 29.78 6.12 ;
      RECT 28.99 0.92 29.16 1.09 ;
      RECT 28.99 2.4 29.16 2.57 ;
      RECT 28.99 6.32 29.16 6.49 ;
      RECT 28.99 7.8 29.16 7.97 ;
      RECT 28.64 0.11 28.81 0.28 ;
      RECT 28.64 4.17 28.81 4.34 ;
      RECT 28.64 4.55 28.81 4.72 ;
      RECT 28.64 8.61 28.81 8.78 ;
      RECT 28.62 2.77 28.79 2.94 ;
      RECT 28.62 5.95 28.79 6.12 ;
      RECT 27.935 0.11 28.105 0.28 ;
      RECT 27.935 4.17 28.105 4.34 ;
      RECT 27.935 4.55 28.105 4.72 ;
      RECT 27.935 8.61 28.105 8.78 ;
      RECT 27.625 2.03 27.795 2.2 ;
      RECT 27.625 6.69 27.795 6.86 ;
      RECT 27.255 0.11 27.425 0.28 ;
      RECT 27.255 8.61 27.425 8.78 ;
      RECT 27.195 0.92 27.365 1.09 ;
      RECT 27.195 1.66 27.365 1.83 ;
      RECT 27.195 7.06 27.365 7.23 ;
      RECT 27.195 7.8 27.365 7.97 ;
      RECT 26.82 2.4 26.99 2.57 ;
      RECT 26.82 6.32 26.99 6.49 ;
      RECT 26.575 0.11 26.745 0.28 ;
      RECT 26.575 8.61 26.745 8.78 ;
      RECT 25.895 0.11 26.065 0.28 ;
      RECT 25.895 8.61 26.065 8.78 ;
      RECT 25.825 2.77 25.995 2.94 ;
      RECT 25.825 5.95 25.995 6.12 ;
      RECT 24.435 1.42 24.605 1.59 ;
      RECT 24.435 4.14 24.605 4.31 ;
      RECT 23.975 1.42 24.145 1.59 ;
      RECT 23.975 4.14 24.145 4.31 ;
      RECT 23.76 2.78 23.93 2.95 ;
      RECT 23.52 1.94 23.69 2.11 ;
      RECT 23.52 3.62 23.69 3.79 ;
      RECT 23.515 1.42 23.685 1.59 ;
      RECT 23.515 4.14 23.685 4.31 ;
      RECT 23.28 2.5 23.45 2.67 ;
      RECT 23.28 3.06 23.45 3.23 ;
      RECT 23.055 1.42 23.225 1.59 ;
      RECT 23.055 4.14 23.225 4.31 ;
      RECT 22.8 2.78 22.97 2.95 ;
      RECT 22.595 1.42 22.765 1.59 ;
      RECT 22.595 4.14 22.765 4.31 ;
      RECT 22.56 1.94 22.73 2.11 ;
      RECT 22.32 2.5 22.49 2.67 ;
      RECT 22.32 4.55 22.49 4.72 ;
      RECT 22.32 8.61 22.49 8.78 ;
      RECT 22.135 1.42 22.305 1.59 ;
      RECT 22.135 4.14 22.305 4.31 ;
      RECT 22.11 3.34 22.28 3.51 ;
      RECT 22.01 6.69 22.18 6.86 ;
      RECT 21.84 2.78 22.01 2.95 ;
      RECT 21.675 1.42 21.845 1.59 ;
      RECT 21.675 4.14 21.845 4.31 ;
      RECT 21.64 8.61 21.81 8.78 ;
      RECT 21.58 7.06 21.75 7.23 ;
      RECT 21.58 7.8 21.75 7.97 ;
      RECT 21.57 3.62 21.74 3.79 ;
      RECT 21.36 2.2 21.53 2.37 ;
      RECT 21.215 1.42 21.385 1.59 ;
      RECT 21.215 4.14 21.385 4.31 ;
      RECT 21.205 6.32 21.375 6.49 ;
      RECT 20.96 8.61 21.13 8.78 ;
      RECT 20.88 2.78 21.05 2.95 ;
      RECT 20.755 1.42 20.925 1.59 ;
      RECT 20.755 4.14 20.925 4.31 ;
      RECT 20.64 1.94 20.81 2.11 ;
      RECT 20.4 2.5 20.57 2.67 ;
      RECT 20.4 3.06 20.57 3.23 ;
      RECT 20.295 1.42 20.465 1.59 ;
      RECT 20.295 4.14 20.465 4.31 ;
      RECT 20.28 8.61 20.45 8.78 ;
      RECT 20.21 5.95 20.38 6.12 ;
      RECT 19.92 2.5 20.09 2.67 ;
      RECT 19.835 1.42 20.005 1.59 ;
      RECT 19.835 4.14 20.005 4.31 ;
      RECT 19.68 3.62 19.85 3.79 ;
      RECT 19.64 1.94 19.81 2.11 ;
      RECT 19.44 2.78 19.61 2.95 ;
      RECT 19.375 1.42 19.545 1.59 ;
      RECT 19.375 4.14 19.545 4.31 ;
      RECT 19.2 3.62 19.37 3.79 ;
      RECT 18.96 3.06 19.13 3.23 ;
      RECT 18.915 1.42 19.085 1.59 ;
      RECT 18.915 4.14 19.085 4.31 ;
      RECT 18.48 2.5 18.65 2.67 ;
      RECT 18.455 1.42 18.625 1.59 ;
      RECT 18.455 4.14 18.625 4.31 ;
      RECT 18.24 1.94 18.41 2.11 ;
      RECT 18.24 3.62 18.41 3.79 ;
      RECT 17.995 1.42 18.165 1.59 ;
      RECT 17.995 4.14 18.165 4.31 ;
      RECT 17.76 1.94 17.93 2.11 ;
      RECT 17.76 3.06 17.93 3.23 ;
      RECT 17.535 1.42 17.705 1.59 ;
      RECT 17.535 4.14 17.705 4.31 ;
      RECT 17.52 2.5 17.69 2.67 ;
      RECT 17.28 3.34 17.45 3.51 ;
      RECT 17.075 1.42 17.245 1.59 ;
      RECT 17.075 4.14 17.245 4.31 ;
      RECT 17.04 2.78 17.21 2.95 ;
      RECT 16.615 1.42 16.785 1.59 ;
      RECT 16.615 4.14 16.785 4.31 ;
      RECT 16.56 2.78 16.73 2.95 ;
      RECT 16.35 1.94 16.52 2.11 ;
      RECT 16.35 3.34 16.52 3.51 ;
      RECT 16.155 1.42 16.325 1.59 ;
      RECT 16.155 4.14 16.325 4.31 ;
      RECT 14.72 0.92 14.89 1.09 ;
      RECT 14.72 2.4 14.89 2.57 ;
      RECT 14.72 6.32 14.89 6.49 ;
      RECT 14.72 7.8 14.89 7.97 ;
      RECT 14.37 0.11 14.54 0.28 ;
      RECT 14.37 4.17 14.54 4.34 ;
      RECT 14.37 4.55 14.54 4.72 ;
      RECT 14.37 8.61 14.54 8.78 ;
      RECT 14.35 2.77 14.52 2.94 ;
      RECT 14.35 5.95 14.52 6.12 ;
      RECT 13.73 0.92 13.9 1.09 ;
      RECT 13.73 2.4 13.9 2.57 ;
      RECT 13.73 6.32 13.9 6.49 ;
      RECT 13.73 7.8 13.9 7.97 ;
      RECT 13.38 0.11 13.55 0.28 ;
      RECT 13.38 4.17 13.55 4.34 ;
      RECT 13.38 4.55 13.55 4.72 ;
      RECT 13.38 8.61 13.55 8.78 ;
      RECT 13.36 2.77 13.53 2.94 ;
      RECT 13.36 5.95 13.53 6.12 ;
      RECT 12.675 0.11 12.845 0.28 ;
      RECT 12.675 4.17 12.845 4.34 ;
      RECT 12.675 4.55 12.845 4.72 ;
      RECT 12.675 8.61 12.845 8.78 ;
      RECT 12.365 2.03 12.535 2.2 ;
      RECT 12.365 6.69 12.535 6.86 ;
      RECT 11.995 0.11 12.165 0.28 ;
      RECT 11.995 8.61 12.165 8.78 ;
      RECT 11.935 0.92 12.105 1.09 ;
      RECT 11.935 1.66 12.105 1.83 ;
      RECT 11.935 7.06 12.105 7.23 ;
      RECT 11.935 7.8 12.105 7.97 ;
      RECT 11.56 2.4 11.73 2.57 ;
      RECT 11.56 6.32 11.73 6.49 ;
      RECT 11.315 0.11 11.485 0.28 ;
      RECT 11.315 8.61 11.485 8.78 ;
      RECT 10.635 0.11 10.805 0.28 ;
      RECT 10.635 8.61 10.805 8.78 ;
      RECT 10.565 2.77 10.735 2.94 ;
      RECT 10.565 5.95 10.735 6.12 ;
      RECT 9.175 1.42 9.345 1.59 ;
      RECT 9.175 4.14 9.345 4.31 ;
      RECT 8.715 1.42 8.885 1.59 ;
      RECT 8.715 4.14 8.885 4.31 ;
      RECT 8.5 2.78 8.67 2.95 ;
      RECT 8.26 1.94 8.43 2.11 ;
      RECT 8.26 3.62 8.43 3.79 ;
      RECT 8.255 1.42 8.425 1.59 ;
      RECT 8.255 4.14 8.425 4.31 ;
      RECT 8.02 2.5 8.19 2.67 ;
      RECT 8.02 3.06 8.19 3.23 ;
      RECT 7.795 1.42 7.965 1.59 ;
      RECT 7.795 4.14 7.965 4.31 ;
      RECT 7.54 2.78 7.71 2.95 ;
      RECT 7.335 1.42 7.505 1.59 ;
      RECT 7.335 4.14 7.505 4.31 ;
      RECT 7.3 1.94 7.47 2.11 ;
      RECT 7.06 2.5 7.23 2.67 ;
      RECT 7.06 4.55 7.23 4.72 ;
      RECT 7.06 8.61 7.23 8.78 ;
      RECT 6.875 1.42 7.045 1.59 ;
      RECT 6.875 4.14 7.045 4.31 ;
      RECT 6.85 3.34 7.02 3.51 ;
      RECT 6.75 6.69 6.92 6.86 ;
      RECT 6.58 2.78 6.75 2.95 ;
      RECT 6.415 1.42 6.585 1.59 ;
      RECT 6.415 4.14 6.585 4.31 ;
      RECT 6.38 8.61 6.55 8.78 ;
      RECT 6.32 7.06 6.49 7.23 ;
      RECT 6.32 7.8 6.49 7.97 ;
      RECT 6.31 3.62 6.48 3.79 ;
      RECT 6.1 2.2 6.27 2.37 ;
      RECT 5.955 1.42 6.125 1.59 ;
      RECT 5.955 4.14 6.125 4.31 ;
      RECT 5.945 6.32 6.115 6.49 ;
      RECT 5.7 8.61 5.87 8.78 ;
      RECT 5.62 2.78 5.79 2.95 ;
      RECT 5.495 1.42 5.665 1.59 ;
      RECT 5.495 4.14 5.665 4.31 ;
      RECT 5.38 1.94 5.55 2.11 ;
      RECT 5.14 2.5 5.31 2.67 ;
      RECT 5.14 3.06 5.31 3.23 ;
      RECT 5.035 1.42 5.205 1.59 ;
      RECT 5.035 4.14 5.205 4.31 ;
      RECT 5.02 8.61 5.19 8.78 ;
      RECT 4.95 5.95 5.12 6.12 ;
      RECT 4.66 2.5 4.83 2.67 ;
      RECT 4.575 1.42 4.745 1.59 ;
      RECT 4.575 4.14 4.745 4.31 ;
      RECT 4.42 3.62 4.59 3.79 ;
      RECT 4.38 1.94 4.55 2.11 ;
      RECT 4.18 2.78 4.35 2.95 ;
      RECT 4.115 1.42 4.285 1.59 ;
      RECT 4.115 4.14 4.285 4.31 ;
      RECT 3.94 3.62 4.11 3.79 ;
      RECT 3.7 3.06 3.87 3.23 ;
      RECT 3.655 1.42 3.825 1.59 ;
      RECT 3.655 4.14 3.825 4.31 ;
      RECT 3.22 2.5 3.39 2.67 ;
      RECT 3.195 1.42 3.365 1.59 ;
      RECT 3.195 4.14 3.365 4.31 ;
      RECT 2.98 1.94 3.15 2.11 ;
      RECT 2.98 3.62 3.15 3.79 ;
      RECT 2.735 1.42 2.905 1.59 ;
      RECT 2.735 4.14 2.905 4.31 ;
      RECT 2.5 1.94 2.67 2.11 ;
      RECT 2.5 3.06 2.67 3.23 ;
      RECT 2.275 1.42 2.445 1.59 ;
      RECT 2.275 4.14 2.445 4.31 ;
      RECT 2.26 2.5 2.43 2.67 ;
      RECT 2.02 3.34 2.19 3.51 ;
      RECT 1.815 1.42 1.985 1.59 ;
      RECT 1.815 4.14 1.985 4.31 ;
      RECT 1.78 2.78 1.95 2.95 ;
      RECT 1.355 1.42 1.525 1.59 ;
      RECT 1.355 4.14 1.525 4.31 ;
      RECT 1.3 2.78 1.47 2.95 ;
      RECT 1.09 1.94 1.26 2.11 ;
      RECT 1.09 3.34 1.26 3.51 ;
      RECT 0.895 1.42 1.065 1.59 ;
      RECT 0.895 4.14 1.065 4.31 ;
      RECT -0.455 4.55 -0.285 4.72 ;
      RECT -0.455 8.61 -0.285 8.78 ;
      RECT -0.765 6.69 -0.595 6.86 ;
      RECT -1.135 8.61 -0.965 8.78 ;
      RECT -1.195 7.06 -1.025 7.23 ;
      RECT -1.195 7.8 -1.025 7.97 ;
      RECT -1.57 6.32 -1.4 6.49 ;
      RECT -1.815 8.61 -1.645 8.78 ;
      RECT -2.495 8.61 -2.325 8.78 ;
      RECT -2.565 5.95 -2.395 6.12 ;
    LAYER li ;
      RECT 69.76 0.005 69.93 2.09 ;
      RECT 68.82 0.005 68.99 2.09 ;
      RECT 67.86 0.005 68.03 2.09 ;
      RECT 65.94 0.005 66.11 2.09 ;
      RECT 64.98 0.005 65.15 2.09 ;
      RECT 63.06 0.005 63.23 2.09 ;
      RECT 54.5 0.005 54.67 2.09 ;
      RECT 53.56 0.005 53.73 2.09 ;
      RECT 52.6 0.005 52.77 2.09 ;
      RECT 50.68 0.005 50.85 2.09 ;
      RECT 49.72 0.005 49.89 2.09 ;
      RECT 47.8 0.005 47.97 2.09 ;
      RECT 39.24 0.005 39.41 2.09 ;
      RECT 38.3 0.005 38.47 2.09 ;
      RECT 37.34 0.005 37.51 2.09 ;
      RECT 35.42 0.005 35.59 2.09 ;
      RECT 34.46 0.005 34.63 2.09 ;
      RECT 32.54 0.005 32.71 2.09 ;
      RECT 23.98 0.005 24.15 2.09 ;
      RECT 23.04 0.005 23.21 2.09 ;
      RECT 22.08 0.005 22.25 2.09 ;
      RECT 20.16 0.005 20.33 2.09 ;
      RECT 19.2 0.005 19.37 2.09 ;
      RECT 17.28 0.005 17.45 2.09 ;
      RECT 8.72 0.005 8.89 2.09 ;
      RECT 7.78 0.005 7.95 2.09 ;
      RECT 6.82 0.005 6.99 2.09 ;
      RECT 4.9 0.005 5.07 2.09 ;
      RECT 3.94 0.005 4.11 2.09 ;
      RECT 2.02 0.005 2.19 2.09 ;
      RECT 66.815 0.005 67.01 1.6 ;
      RECT 63.06 0.005 63.335 1.6 ;
      RECT 51.555 0.005 51.75 1.6 ;
      RECT 47.8 0.005 48.075 1.6 ;
      RECT 36.295 0.005 36.49 1.6 ;
      RECT 32.54 0.005 32.815 1.6 ;
      RECT 21.035 0.005 21.23 1.6 ;
      RECT 17.28 0.005 17.555 1.6 ;
      RECT 5.775 0.005 5.97 1.6 ;
      RECT 2.02 0.005 2.295 1.6 ;
      RECT 61.79 0.005 70.53 1.59 ;
      RECT 46.53 0.005 55.27 1.59 ;
      RECT 31.27 0.005 40.01 1.59 ;
      RECT 16.01 0.005 24.75 1.59 ;
      RECT 0.75 0.005 9.49 1.59 ;
      RECT 75.33 0.005 75.5 0.94 ;
      RECT 74.34 0.005 74.51 0.94 ;
      RECT 71.595 0.005 71.765 0.94 ;
      RECT 60.07 0.005 60.24 0.94 ;
      RECT 59.08 0.005 59.25 0.94 ;
      RECT 56.335 0.005 56.505 0.94 ;
      RECT 44.81 0.005 44.98 0.94 ;
      RECT 43.82 0.005 43.99 0.94 ;
      RECT 41.075 0.005 41.245 0.94 ;
      RECT 29.55 0.005 29.72 0.94 ;
      RECT 28.56 0.005 28.73 0.94 ;
      RECT 25.815 0.005 25.985 0.94 ;
      RECT 14.29 0.005 14.46 0.94 ;
      RECT 13.3 0.005 13.47 0.94 ;
      RECT 10.555 0.005 10.725 0.94 ;
      RECT -2.75 0.005 76.3 0.31 ;
      RECT -0.765 4.145 -0.595 8.31 ;
      RECT 75.33 3.41 75.5 5.48 ;
      RECT 74.34 3.41 74.51 5.48 ;
      RECT 71.595 3.41 71.765 5.48 ;
      RECT 65.98 4.14 66.15 5.48 ;
      RECT 60.07 3.41 60.24 5.48 ;
      RECT 59.08 3.41 59.25 5.48 ;
      RECT 56.335 3.41 56.505 5.48 ;
      RECT 50.72 4.14 50.89 5.48 ;
      RECT 44.81 3.41 44.98 5.48 ;
      RECT 43.82 3.41 43.99 5.48 ;
      RECT 41.075 3.41 41.245 5.48 ;
      RECT 35.46 4.14 35.63 5.48 ;
      RECT 29.55 3.41 29.72 5.48 ;
      RECT 28.56 3.41 28.73 5.48 ;
      RECT 25.815 3.41 25.985 5.48 ;
      RECT 20.2 4.14 20.37 5.48 ;
      RECT 14.29 3.41 14.46 5.48 ;
      RECT 13.3 3.41 13.47 5.48 ;
      RECT 10.555 3.41 10.725 5.48 ;
      RECT 4.94 4.14 5.11 5.48 ;
      RECT -2.575 4.145 -2.405 5.48 ;
      RECT -2.75 4.145 76.3 4.75 ;
      RECT 61.79 4.14 76.3 4.75 ;
      RECT 46.53 4.14 61.04 4.75 ;
      RECT 31.27 4.14 45.78 4.75 ;
      RECT 16.01 4.14 30.52 4.75 ;
      RECT 0.75 4.14 15.26 4.75 ;
      RECT 68.82 3.64 68.99 4.75 ;
      RECT 66.9 3.64 67.07 4.75 ;
      RECT 65.96 3.64 66.13 4.75 ;
      RECT 64.5 3.64 64.67 4.75 ;
      RECT 62.58 3.64 62.75 4.75 ;
      RECT 53.56 3.64 53.73 4.75 ;
      RECT 51.64 3.64 51.81 4.75 ;
      RECT 50.7 3.64 50.87 4.75 ;
      RECT 49.24 3.64 49.41 4.75 ;
      RECT 47.32 3.64 47.49 4.75 ;
      RECT 38.3 3.64 38.47 4.75 ;
      RECT 36.38 3.64 36.55 4.75 ;
      RECT 35.44 3.64 35.61 4.75 ;
      RECT 33.98 3.64 34.15 4.75 ;
      RECT 32.06 3.64 32.23 4.75 ;
      RECT 23.04 3.64 23.21 4.75 ;
      RECT 21.12 3.64 21.29 4.75 ;
      RECT 20.18 3.64 20.35 4.75 ;
      RECT 18.72 3.64 18.89 4.75 ;
      RECT 16.8 3.64 16.97 4.75 ;
      RECT 7.78 3.64 7.95 4.75 ;
      RECT 5.86 3.64 6.03 4.75 ;
      RECT 4.92 3.64 5.09 4.75 ;
      RECT 3.46 3.64 3.63 4.75 ;
      RECT 1.54 3.64 1.71 4.75 ;
      RECT -2.75 8.58 76.3 8.885 ;
      RECT 75.33 7.95 75.5 8.885 ;
      RECT 74.34 7.95 74.51 8.885 ;
      RECT 71.595 7.95 71.765 8.885 ;
      RECT 65.98 7.95 66.15 8.885 ;
      RECT 60.07 7.95 60.24 8.885 ;
      RECT 59.08 7.95 59.25 8.885 ;
      RECT 56.335 7.95 56.505 8.885 ;
      RECT 50.72 7.95 50.89 8.885 ;
      RECT 44.81 7.95 44.98 8.885 ;
      RECT 43.82 7.95 43.99 8.885 ;
      RECT 41.075 7.95 41.245 8.885 ;
      RECT 35.46 7.95 35.63 8.885 ;
      RECT 29.55 7.95 29.72 8.885 ;
      RECT 28.56 7.95 28.73 8.885 ;
      RECT 25.815 7.95 25.985 8.885 ;
      RECT 20.2 7.95 20.37 8.885 ;
      RECT 14.29 7.95 14.46 8.885 ;
      RECT 13.3 7.95 13.47 8.885 ;
      RECT 10.555 7.95 10.725 8.885 ;
      RECT 4.94 7.95 5.11 8.885 ;
      RECT -2.575 7.95 -2.405 8.885 ;
      RECT 75.39 1.745 75.56 2.94 ;
      RECT 75.39 1.745 75.855 1.915 ;
      RECT 75.39 6.975 75.855 7.145 ;
      RECT 75.39 5.95 75.56 7.145 ;
      RECT 74.4 1.745 74.57 2.94 ;
      RECT 74.4 1.745 74.865 1.915 ;
      RECT 74.4 6.975 74.865 7.145 ;
      RECT 74.4 5.95 74.57 7.145 ;
      RECT 72.545 2.64 72.715 3.87 ;
      RECT 72.6 0.86 72.77 2.81 ;
      RECT 72.545 0.58 72.715 1.03 ;
      RECT 72.545 7.86 72.715 8.31 ;
      RECT 72.6 6.08 72.77 8.03 ;
      RECT 72.545 5.02 72.715 6.25 ;
      RECT 72.025 0.58 72.195 3.87 ;
      RECT 72.025 2.08 72.43 2.41 ;
      RECT 72.025 1.24 72.43 1.57 ;
      RECT 72.025 5.02 72.195 8.31 ;
      RECT 72.025 7.32 72.43 7.65 ;
      RECT 72.025 6.48 72.43 6.81 ;
      RECT 69.3 3.62 69.815 3.79 ;
      RECT 69.645 3.23 69.815 3.79 ;
      RECT 69.75 3.15 69.92 3.48 ;
      RECT 69.54 2.54 69.815 2.95 ;
      RECT 69.42 2.54 69.815 2.75 ;
      RECT 67.89 3.15 68.06 3.51 ;
      RECT 67.89 3.23 69.23 3.4 ;
      RECT 69.06 3.06 69.23 3.4 ;
      RECT 67.62 2.58 67.79 2.95 ;
      RECT 67.14 2.58 67.79 2.85 ;
      RECT 67.06 2.58 67.87 2.75 ;
      RECT 66.42 1.82 66.59 2.11 ;
      RECT 66.42 1.82 67.66 1.99 ;
      RECT 67.14 2.16 67.31 2.37 ;
      RECT 66.78 2.16 67.31 2.33 ;
      RECT 66.93 7.86 67.1 8.31 ;
      RECT 66.985 6.08 67.155 8.03 ;
      RECT 66.93 5.02 67.1 6.25 ;
      RECT 66.41 5.02 66.58 8.31 ;
      RECT 66.41 7.32 66.815 7.65 ;
      RECT 66.41 6.48 66.815 6.81 ;
      RECT 66.18 3.23 66.67 3.4 ;
      RECT 66.18 3.06 66.35 3.4 ;
      RECT 65.46 3.23 65.63 3.79 ;
      RECT 65.35 3.23 65.68 3.4 ;
      RECT 65.42 1.84 65.59 2.11 ;
      RECT 65.46 1.76 65.63 2.09 ;
      RECT 65.325 1.84 65.63 2.06 ;
      RECT 63.9 3.23 64.19 3.79 ;
      RECT 64.02 3.15 64.19 3.79 ;
      RECT 63.66 2.58 64.03 2.75 ;
      RECT 63.66 1.94 63.83 2.75 ;
      RECT 63.54 1.94 63.83 2.11 ;
      RECT 60.13 1.745 60.3 2.94 ;
      RECT 60.13 1.745 60.595 1.915 ;
      RECT 60.13 6.975 60.595 7.145 ;
      RECT 60.13 5.95 60.3 7.145 ;
      RECT 59.14 1.745 59.31 2.94 ;
      RECT 59.14 1.745 59.605 1.915 ;
      RECT 59.14 6.975 59.605 7.145 ;
      RECT 59.14 5.95 59.31 7.145 ;
      RECT 57.285 2.64 57.455 3.87 ;
      RECT 57.34 0.86 57.51 2.81 ;
      RECT 57.285 0.58 57.455 1.03 ;
      RECT 57.285 7.86 57.455 8.31 ;
      RECT 57.34 6.08 57.51 8.03 ;
      RECT 57.285 5.02 57.455 6.25 ;
      RECT 56.765 0.58 56.935 3.87 ;
      RECT 56.765 2.08 57.17 2.41 ;
      RECT 56.765 1.24 57.17 1.57 ;
      RECT 56.765 5.02 56.935 8.31 ;
      RECT 56.765 7.32 57.17 7.65 ;
      RECT 56.765 6.48 57.17 6.81 ;
      RECT 54.04 3.62 54.555 3.79 ;
      RECT 54.385 3.23 54.555 3.79 ;
      RECT 54.49 3.15 54.66 3.48 ;
      RECT 54.28 2.54 54.555 2.95 ;
      RECT 54.16 2.54 54.555 2.75 ;
      RECT 52.63 3.15 52.8 3.51 ;
      RECT 52.63 3.23 53.97 3.4 ;
      RECT 53.8 3.06 53.97 3.4 ;
      RECT 52.36 2.58 52.53 2.95 ;
      RECT 51.88 2.58 52.53 2.85 ;
      RECT 51.8 2.58 52.61 2.75 ;
      RECT 51.16 1.82 51.33 2.11 ;
      RECT 51.16 1.82 52.4 1.99 ;
      RECT 51.88 2.16 52.05 2.37 ;
      RECT 51.52 2.16 52.05 2.33 ;
      RECT 51.67 7.86 51.84 8.31 ;
      RECT 51.725 6.08 51.895 8.03 ;
      RECT 51.67 5.02 51.84 6.25 ;
      RECT 51.15 5.02 51.32 8.31 ;
      RECT 51.15 7.32 51.555 7.65 ;
      RECT 51.15 6.48 51.555 6.81 ;
      RECT 50.92 3.23 51.41 3.4 ;
      RECT 50.92 3.06 51.09 3.4 ;
      RECT 50.2 3.23 50.37 3.79 ;
      RECT 50.09 3.23 50.42 3.4 ;
      RECT 50.16 1.84 50.33 2.11 ;
      RECT 50.2 1.76 50.37 2.09 ;
      RECT 50.065 1.84 50.37 2.06 ;
      RECT 48.64 3.23 48.93 3.79 ;
      RECT 48.76 3.15 48.93 3.79 ;
      RECT 48.4 2.58 48.77 2.75 ;
      RECT 48.4 1.94 48.57 2.75 ;
      RECT 48.28 1.94 48.57 2.11 ;
      RECT 44.87 1.745 45.04 2.94 ;
      RECT 44.87 1.745 45.335 1.915 ;
      RECT 44.87 6.975 45.335 7.145 ;
      RECT 44.87 5.95 45.04 7.145 ;
      RECT 43.88 1.745 44.05 2.94 ;
      RECT 43.88 1.745 44.345 1.915 ;
      RECT 43.88 6.975 44.345 7.145 ;
      RECT 43.88 5.95 44.05 7.145 ;
      RECT 42.025 2.64 42.195 3.87 ;
      RECT 42.08 0.86 42.25 2.81 ;
      RECT 42.025 0.58 42.195 1.03 ;
      RECT 42.025 7.86 42.195 8.31 ;
      RECT 42.08 6.08 42.25 8.03 ;
      RECT 42.025 5.02 42.195 6.25 ;
      RECT 41.505 0.58 41.675 3.87 ;
      RECT 41.505 2.08 41.91 2.41 ;
      RECT 41.505 1.24 41.91 1.57 ;
      RECT 41.505 5.02 41.675 8.31 ;
      RECT 41.505 7.32 41.91 7.65 ;
      RECT 41.505 6.48 41.91 6.81 ;
      RECT 38.78 3.62 39.295 3.79 ;
      RECT 39.125 3.23 39.295 3.79 ;
      RECT 39.23 3.15 39.4 3.48 ;
      RECT 39.02 2.54 39.295 2.95 ;
      RECT 38.9 2.54 39.295 2.75 ;
      RECT 37.37 3.15 37.54 3.51 ;
      RECT 37.37 3.23 38.71 3.4 ;
      RECT 38.54 3.06 38.71 3.4 ;
      RECT 37.1 2.58 37.27 2.95 ;
      RECT 36.62 2.58 37.27 2.85 ;
      RECT 36.54 2.58 37.35 2.75 ;
      RECT 35.9 1.82 36.07 2.11 ;
      RECT 35.9 1.82 37.14 1.99 ;
      RECT 36.62 2.16 36.79 2.37 ;
      RECT 36.26 2.16 36.79 2.33 ;
      RECT 36.41 7.86 36.58 8.31 ;
      RECT 36.465 6.08 36.635 8.03 ;
      RECT 36.41 5.02 36.58 6.25 ;
      RECT 35.89 5.02 36.06 8.31 ;
      RECT 35.89 7.32 36.295 7.65 ;
      RECT 35.89 6.48 36.295 6.81 ;
      RECT 35.66 3.23 36.15 3.4 ;
      RECT 35.66 3.06 35.83 3.4 ;
      RECT 34.94 3.23 35.11 3.79 ;
      RECT 34.83 3.23 35.16 3.4 ;
      RECT 34.9 1.84 35.07 2.11 ;
      RECT 34.94 1.76 35.11 2.09 ;
      RECT 34.805 1.84 35.11 2.06 ;
      RECT 33.38 3.23 33.67 3.79 ;
      RECT 33.5 3.15 33.67 3.79 ;
      RECT 33.14 2.58 33.51 2.75 ;
      RECT 33.14 1.94 33.31 2.75 ;
      RECT 33.02 1.94 33.31 2.11 ;
      RECT 29.61 1.745 29.78 2.94 ;
      RECT 29.61 1.745 30.075 1.915 ;
      RECT 29.61 6.975 30.075 7.145 ;
      RECT 29.61 5.95 29.78 7.145 ;
      RECT 28.62 1.745 28.79 2.94 ;
      RECT 28.62 1.745 29.085 1.915 ;
      RECT 28.62 6.975 29.085 7.145 ;
      RECT 28.62 5.95 28.79 7.145 ;
      RECT 26.765 2.64 26.935 3.87 ;
      RECT 26.82 0.86 26.99 2.81 ;
      RECT 26.765 0.58 26.935 1.03 ;
      RECT 26.765 7.86 26.935 8.31 ;
      RECT 26.82 6.08 26.99 8.03 ;
      RECT 26.765 5.02 26.935 6.25 ;
      RECT 26.245 0.58 26.415 3.87 ;
      RECT 26.245 2.08 26.65 2.41 ;
      RECT 26.245 1.24 26.65 1.57 ;
      RECT 26.245 5.02 26.415 8.31 ;
      RECT 26.245 7.32 26.65 7.65 ;
      RECT 26.245 6.48 26.65 6.81 ;
      RECT 23.52 3.62 24.035 3.79 ;
      RECT 23.865 3.23 24.035 3.79 ;
      RECT 23.97 3.15 24.14 3.48 ;
      RECT 23.76 2.54 24.035 2.95 ;
      RECT 23.64 2.54 24.035 2.75 ;
      RECT 22.11 3.15 22.28 3.51 ;
      RECT 22.11 3.23 23.45 3.4 ;
      RECT 23.28 3.06 23.45 3.4 ;
      RECT 21.84 2.58 22.01 2.95 ;
      RECT 21.36 2.58 22.01 2.85 ;
      RECT 21.28 2.58 22.09 2.75 ;
      RECT 20.64 1.82 20.81 2.11 ;
      RECT 20.64 1.82 21.88 1.99 ;
      RECT 21.36 2.16 21.53 2.37 ;
      RECT 21 2.16 21.53 2.33 ;
      RECT 21.15 7.86 21.32 8.31 ;
      RECT 21.205 6.08 21.375 8.03 ;
      RECT 21.15 5.02 21.32 6.25 ;
      RECT 20.63 5.02 20.8 8.31 ;
      RECT 20.63 7.32 21.035 7.65 ;
      RECT 20.63 6.48 21.035 6.81 ;
      RECT 20.4 3.23 20.89 3.4 ;
      RECT 20.4 3.06 20.57 3.4 ;
      RECT 19.68 3.23 19.85 3.79 ;
      RECT 19.57 3.23 19.9 3.4 ;
      RECT 19.64 1.84 19.81 2.11 ;
      RECT 19.68 1.76 19.85 2.09 ;
      RECT 19.545 1.84 19.85 2.06 ;
      RECT 18.12 3.23 18.41 3.79 ;
      RECT 18.24 3.15 18.41 3.79 ;
      RECT 17.88 2.58 18.25 2.75 ;
      RECT 17.88 1.94 18.05 2.75 ;
      RECT 17.76 1.94 18.05 2.11 ;
      RECT 14.35 1.745 14.52 2.94 ;
      RECT 14.35 1.745 14.815 1.915 ;
      RECT 14.35 6.975 14.815 7.145 ;
      RECT 14.35 5.95 14.52 7.145 ;
      RECT 13.36 1.745 13.53 2.94 ;
      RECT 13.36 1.745 13.825 1.915 ;
      RECT 13.36 6.975 13.825 7.145 ;
      RECT 13.36 5.95 13.53 7.145 ;
      RECT 11.505 2.64 11.675 3.87 ;
      RECT 11.56 0.86 11.73 2.81 ;
      RECT 11.505 0.58 11.675 1.03 ;
      RECT 11.505 7.86 11.675 8.31 ;
      RECT 11.56 6.08 11.73 8.03 ;
      RECT 11.505 5.02 11.675 6.25 ;
      RECT 10.985 0.58 11.155 3.87 ;
      RECT 10.985 2.08 11.39 2.41 ;
      RECT 10.985 1.24 11.39 1.57 ;
      RECT 10.985 5.02 11.155 8.31 ;
      RECT 10.985 7.32 11.39 7.65 ;
      RECT 10.985 6.48 11.39 6.81 ;
      RECT 8.26 3.62 8.775 3.79 ;
      RECT 8.605 3.23 8.775 3.79 ;
      RECT 8.71 3.15 8.88 3.48 ;
      RECT 8.5 2.54 8.775 2.95 ;
      RECT 8.38 2.54 8.775 2.75 ;
      RECT 6.85 3.15 7.02 3.51 ;
      RECT 6.85 3.23 8.19 3.4 ;
      RECT 8.02 3.06 8.19 3.4 ;
      RECT 6.58 2.58 6.75 2.95 ;
      RECT 6.1 2.58 6.75 2.85 ;
      RECT 6.02 2.58 6.83 2.75 ;
      RECT 5.38 1.82 5.55 2.11 ;
      RECT 5.38 1.82 6.62 1.99 ;
      RECT 6.1 2.16 6.27 2.37 ;
      RECT 5.74 2.16 6.27 2.33 ;
      RECT 5.89 7.86 6.06 8.31 ;
      RECT 5.945 6.08 6.115 8.03 ;
      RECT 5.89 5.02 6.06 6.25 ;
      RECT 5.37 5.02 5.54 8.31 ;
      RECT 5.37 7.32 5.775 7.65 ;
      RECT 5.37 6.48 5.775 6.81 ;
      RECT 5.14 3.23 5.63 3.4 ;
      RECT 5.14 3.06 5.31 3.4 ;
      RECT 4.42 3.23 4.59 3.79 ;
      RECT 4.31 3.23 4.64 3.4 ;
      RECT 4.38 1.84 4.55 2.11 ;
      RECT 4.42 1.76 4.59 2.09 ;
      RECT 4.285 1.84 4.59 2.06 ;
      RECT 2.86 3.23 3.15 3.79 ;
      RECT 2.98 3.15 3.15 3.79 ;
      RECT 2.62 2.58 2.99 2.75 ;
      RECT 2.62 1.94 2.79 2.75 ;
      RECT 2.5 1.94 2.79 2.11 ;
      RECT -1.625 7.86 -1.455 8.31 ;
      RECT -1.57 6.08 -1.4 8.03 ;
      RECT -1.625 5.02 -1.455 6.25 ;
      RECT -2.145 5.02 -1.975 8.31 ;
      RECT -2.145 7.32 -1.74 7.65 ;
      RECT -2.145 6.48 -1.74 6.81 ;
      RECT 75.76 0.58 75.93 1.09 ;
      RECT 75.76 2.4 75.93 3.87 ;
      RECT 75.76 5.02 75.93 6.49 ;
      RECT 75.76 7.8 75.93 8.31 ;
      RECT 74.77 0.58 74.94 1.09 ;
      RECT 74.77 2.4 74.94 3.87 ;
      RECT 74.77 5.02 74.94 6.49 ;
      RECT 74.77 7.8 74.94 8.31 ;
      RECT 73.405 0.58 73.575 3.87 ;
      RECT 73.405 5.02 73.575 8.31 ;
      RECT 72.975 0.58 73.145 1.09 ;
      RECT 72.975 1.66 73.145 3.87 ;
      RECT 72.975 5.02 73.145 7.23 ;
      RECT 72.975 7.8 73.145 8.31 ;
      RECT 71.605 1.665 71.775 2.94 ;
      RECT 71.605 5.95 71.775 7.225 ;
      RECT 69.3 1.76 69.47 2.11 ;
      RECT 69.06 2.5 69.23 2.83 ;
      RECT 68.58 2.5 68.75 2.95 ;
      RECT 68.34 1.76 68.51 2.11 ;
      RECT 68.1 2.5 68.27 2.83 ;
      RECT 67.79 5.02 67.96 8.31 ;
      RECT 67.36 5.02 67.53 7.23 ;
      RECT 67.36 7.8 67.53 8.31 ;
      RECT 67.35 3.49 67.52 3.82 ;
      RECT 66.66 2.5 66.83 2.95 ;
      RECT 66.18 2.5 66.35 2.83 ;
      RECT 65.99 5.95 66.16 7.225 ;
      RECT 65.7 2.5 65.87 2.83 ;
      RECT 65.22 2.5 65.39 2.95 ;
      RECT 64.98 3.49 65.15 3.82 ;
      RECT 64.74 2.5 64.91 3.23 ;
      RECT 64.26 2.5 64.43 2.83 ;
      RECT 64.02 1.76 64.19 2.11 ;
      RECT 63.54 3.06 63.71 3.48 ;
      RECT 63.3 2.5 63.47 2.83 ;
      RECT 63.06 3.15 63.23 3.51 ;
      RECT 62.82 2.5 62.99 2.95 ;
      RECT 62.34 2.5 62.51 2.95 ;
      RECT 62.13 1.76 62.3 2.11 ;
      RECT 62.13 3.15 62.3 3.51 ;
      RECT 60.5 0.58 60.67 1.09 ;
      RECT 60.5 2.4 60.67 3.87 ;
      RECT 60.5 5.02 60.67 6.49 ;
      RECT 60.5 7.8 60.67 8.31 ;
      RECT 59.51 0.58 59.68 1.09 ;
      RECT 59.51 2.4 59.68 3.87 ;
      RECT 59.51 5.02 59.68 6.49 ;
      RECT 59.51 7.8 59.68 8.31 ;
      RECT 58.145 0.58 58.315 3.87 ;
      RECT 58.145 5.02 58.315 8.31 ;
      RECT 57.715 0.58 57.885 1.09 ;
      RECT 57.715 1.66 57.885 3.87 ;
      RECT 57.715 5.02 57.885 7.23 ;
      RECT 57.715 7.8 57.885 8.31 ;
      RECT 56.345 1.665 56.515 2.94 ;
      RECT 56.345 5.95 56.515 7.225 ;
      RECT 54.04 1.76 54.21 2.11 ;
      RECT 53.8 2.5 53.97 2.83 ;
      RECT 53.32 2.5 53.49 2.95 ;
      RECT 53.08 1.76 53.25 2.11 ;
      RECT 52.84 2.5 53.01 2.83 ;
      RECT 52.53 5.02 52.7 8.31 ;
      RECT 52.1 5.02 52.27 7.23 ;
      RECT 52.1 7.8 52.27 8.31 ;
      RECT 52.09 3.49 52.26 3.82 ;
      RECT 51.4 2.5 51.57 2.95 ;
      RECT 50.92 2.5 51.09 2.83 ;
      RECT 50.73 5.95 50.9 7.225 ;
      RECT 50.44 2.5 50.61 2.83 ;
      RECT 49.96 2.5 50.13 2.95 ;
      RECT 49.72 3.49 49.89 3.82 ;
      RECT 49.48 2.5 49.65 3.23 ;
      RECT 49 2.5 49.17 2.83 ;
      RECT 48.76 1.76 48.93 2.11 ;
      RECT 48.28 3.06 48.45 3.48 ;
      RECT 48.04 2.5 48.21 2.83 ;
      RECT 47.8 3.15 47.97 3.51 ;
      RECT 47.56 2.5 47.73 2.95 ;
      RECT 47.08 2.5 47.25 2.95 ;
      RECT 46.87 1.76 47.04 2.11 ;
      RECT 46.87 3.15 47.04 3.51 ;
      RECT 45.24 0.58 45.41 1.09 ;
      RECT 45.24 2.4 45.41 3.87 ;
      RECT 45.24 5.02 45.41 6.49 ;
      RECT 45.24 7.8 45.41 8.31 ;
      RECT 44.25 0.58 44.42 1.09 ;
      RECT 44.25 2.4 44.42 3.87 ;
      RECT 44.25 5.02 44.42 6.49 ;
      RECT 44.25 7.8 44.42 8.31 ;
      RECT 42.885 0.58 43.055 3.87 ;
      RECT 42.885 5.02 43.055 8.31 ;
      RECT 42.455 0.58 42.625 1.09 ;
      RECT 42.455 1.66 42.625 3.87 ;
      RECT 42.455 5.02 42.625 7.23 ;
      RECT 42.455 7.8 42.625 8.31 ;
      RECT 41.085 1.665 41.255 2.94 ;
      RECT 41.085 5.95 41.255 7.225 ;
      RECT 38.78 1.76 38.95 2.11 ;
      RECT 38.54 2.5 38.71 2.83 ;
      RECT 38.06 2.5 38.23 2.95 ;
      RECT 37.82 1.76 37.99 2.11 ;
      RECT 37.58 2.5 37.75 2.83 ;
      RECT 37.27 5.02 37.44 8.31 ;
      RECT 36.84 5.02 37.01 7.23 ;
      RECT 36.84 7.8 37.01 8.31 ;
      RECT 36.83 3.49 37 3.82 ;
      RECT 36.14 2.5 36.31 2.95 ;
      RECT 35.66 2.5 35.83 2.83 ;
      RECT 35.47 5.95 35.64 7.225 ;
      RECT 35.18 2.5 35.35 2.83 ;
      RECT 34.7 2.5 34.87 2.95 ;
      RECT 34.46 3.49 34.63 3.82 ;
      RECT 34.22 2.5 34.39 3.23 ;
      RECT 33.74 2.5 33.91 2.83 ;
      RECT 33.5 1.76 33.67 2.11 ;
      RECT 33.02 3.06 33.19 3.48 ;
      RECT 32.78 2.5 32.95 2.83 ;
      RECT 32.54 3.15 32.71 3.51 ;
      RECT 32.3 2.5 32.47 2.95 ;
      RECT 31.82 2.5 31.99 2.95 ;
      RECT 31.61 1.76 31.78 2.11 ;
      RECT 31.61 3.15 31.78 3.51 ;
      RECT 29.98 0.58 30.15 1.09 ;
      RECT 29.98 2.4 30.15 3.87 ;
      RECT 29.98 5.02 30.15 6.49 ;
      RECT 29.98 7.8 30.15 8.31 ;
      RECT 28.99 0.58 29.16 1.09 ;
      RECT 28.99 2.4 29.16 3.87 ;
      RECT 28.99 5.02 29.16 6.49 ;
      RECT 28.99 7.8 29.16 8.31 ;
      RECT 27.625 0.58 27.795 3.87 ;
      RECT 27.625 5.02 27.795 8.31 ;
      RECT 27.195 0.58 27.365 1.09 ;
      RECT 27.195 1.66 27.365 3.87 ;
      RECT 27.195 5.02 27.365 7.23 ;
      RECT 27.195 7.8 27.365 8.31 ;
      RECT 25.825 1.665 25.995 2.94 ;
      RECT 25.825 5.95 25.995 7.225 ;
      RECT 23.52 1.76 23.69 2.11 ;
      RECT 23.28 2.5 23.45 2.83 ;
      RECT 22.8 2.5 22.97 2.95 ;
      RECT 22.56 1.76 22.73 2.11 ;
      RECT 22.32 2.5 22.49 2.83 ;
      RECT 22.01 5.02 22.18 8.31 ;
      RECT 21.58 5.02 21.75 7.23 ;
      RECT 21.58 7.8 21.75 8.31 ;
      RECT 21.57 3.49 21.74 3.82 ;
      RECT 20.88 2.5 21.05 2.95 ;
      RECT 20.4 2.5 20.57 2.83 ;
      RECT 20.21 5.95 20.38 7.225 ;
      RECT 19.92 2.5 20.09 2.83 ;
      RECT 19.44 2.5 19.61 2.95 ;
      RECT 19.2 3.49 19.37 3.82 ;
      RECT 18.96 2.5 19.13 3.23 ;
      RECT 18.48 2.5 18.65 2.83 ;
      RECT 18.24 1.76 18.41 2.11 ;
      RECT 17.76 3.06 17.93 3.48 ;
      RECT 17.52 2.5 17.69 2.83 ;
      RECT 17.28 3.15 17.45 3.51 ;
      RECT 17.04 2.5 17.21 2.95 ;
      RECT 16.56 2.5 16.73 2.95 ;
      RECT 16.35 1.76 16.52 2.11 ;
      RECT 16.35 3.15 16.52 3.51 ;
      RECT 14.72 0.58 14.89 1.09 ;
      RECT 14.72 2.4 14.89 3.87 ;
      RECT 14.72 5.02 14.89 6.49 ;
      RECT 14.72 7.8 14.89 8.31 ;
      RECT 13.73 0.58 13.9 1.09 ;
      RECT 13.73 2.4 13.9 3.87 ;
      RECT 13.73 5.02 13.9 6.49 ;
      RECT 13.73 7.8 13.9 8.31 ;
      RECT 12.365 0.58 12.535 3.87 ;
      RECT 12.365 5.02 12.535 8.31 ;
      RECT 11.935 0.58 12.105 1.09 ;
      RECT 11.935 1.66 12.105 3.87 ;
      RECT 11.935 5.02 12.105 7.23 ;
      RECT 11.935 7.8 12.105 8.31 ;
      RECT 10.565 1.665 10.735 2.94 ;
      RECT 10.565 5.95 10.735 7.225 ;
      RECT 8.26 1.76 8.43 2.11 ;
      RECT 8.02 2.5 8.19 2.83 ;
      RECT 7.54 2.5 7.71 2.95 ;
      RECT 7.3 1.76 7.47 2.11 ;
      RECT 7.06 2.5 7.23 2.83 ;
      RECT 6.75 5.02 6.92 8.31 ;
      RECT 6.32 5.02 6.49 7.23 ;
      RECT 6.32 7.8 6.49 8.31 ;
      RECT 6.31 3.49 6.48 3.82 ;
      RECT 5.62 2.5 5.79 2.95 ;
      RECT 5.14 2.5 5.31 2.83 ;
      RECT 4.95 5.95 5.12 7.225 ;
      RECT 4.66 2.5 4.83 2.83 ;
      RECT 4.18 2.5 4.35 2.95 ;
      RECT 3.94 3.49 4.11 3.82 ;
      RECT 3.7 2.5 3.87 3.23 ;
      RECT 3.22 2.5 3.39 2.83 ;
      RECT 2.98 1.76 3.15 2.11 ;
      RECT 2.5 3.06 2.67 3.48 ;
      RECT 2.26 2.5 2.43 2.83 ;
      RECT 2.02 3.15 2.19 3.51 ;
      RECT 1.78 2.5 1.95 2.95 ;
      RECT 1.3 2.5 1.47 2.95 ;
      RECT 1.09 1.76 1.26 2.11 ;
      RECT 1.09 3.15 1.26 3.51 ;
      RECT -1.195 5.02 -1.025 7.23 ;
      RECT -1.195 7.8 -1.025 8.31 ;
      RECT -2.565 5.95 -2.395 7.225 ;
  END
END sky130_osu_ring_oscillator_mpr2xa_8_b0r2

MACRO sky130_osu_ring_oscillator_mpr2ya_8_b0r1
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 2.795 0 ;
  SIZE 79.095 BY 8.88 ;
  SYMMETRY X Y R90 ;
  SITE CoreSite ;
  OBS
    LAYER met3 ;
      RECT 67.24 7.055 67.61 7.425 ;
      RECT 67.275 4.27 67.575 7.425 ;
      RECT 63.085 4.27 67.575 4.57 ;
      RECT 66.265 1.855 66.565 4.57 ;
      RECT 63.085 2.435 63.385 4.57 ;
      RECT 66.22 2.76 66.565 3.49 ;
      RECT 62.98 2.015 63.31 2.745 ;
      RECT 65.86 1.855 66.59 2.185 ;
      RECT 51.98 7.055 52.35 7.425 ;
      RECT 52.015 4.27 52.315 7.425 ;
      RECT 47.825 4.27 52.315 4.57 ;
      RECT 51.005 1.855 51.305 4.57 ;
      RECT 47.825 2.435 48.125 4.57 ;
      RECT 50.96 2.76 51.305 3.49 ;
      RECT 47.72 2.015 48.05 2.745 ;
      RECT 50.6 1.855 51.33 2.185 ;
      RECT 36.72 7.055 37.09 7.425 ;
      RECT 36.755 4.27 37.055 7.425 ;
      RECT 32.565 4.27 37.055 4.57 ;
      RECT 35.745 1.855 36.045 4.57 ;
      RECT 32.565 2.435 32.865 4.57 ;
      RECT 35.7 2.76 36.045 3.49 ;
      RECT 32.46 2.015 32.79 2.745 ;
      RECT 35.34 1.855 36.07 2.185 ;
      RECT 21.46 7.055 21.83 7.425 ;
      RECT 21.495 4.27 21.795 7.425 ;
      RECT 17.305 4.27 21.795 4.57 ;
      RECT 20.485 1.855 20.785 4.57 ;
      RECT 17.305 2.435 17.605 4.57 ;
      RECT 20.44 2.76 20.785 3.49 ;
      RECT 17.2 2.015 17.53 2.745 ;
      RECT 20.08 1.855 20.81 2.185 ;
      RECT 6.2 7.055 6.57 7.425 ;
      RECT 6.235 4.27 6.535 7.425 ;
      RECT 2.045 4.27 6.535 4.57 ;
      RECT 5.225 1.855 5.525 4.57 ;
      RECT 2.045 2.435 2.345 4.57 ;
      RECT 5.18 2.76 5.525 3.49 ;
      RECT 1.94 2.015 2.27 2.745 ;
      RECT 4.82 1.855 5.55 2.185 ;
      RECT 69.34 2.015 69.67 2.745 ;
      RECT 68.14 2.88 68.47 3.61 ;
      RECT 67.3 1.855 68.03 2.185 ;
      RECT 64.9 1.855 65.23 2.585 ;
      RECT 63.7 2.015 64.03 2.745 ;
      RECT 54.08 2.015 54.41 2.745 ;
      RECT 52.88 2.88 53.21 3.61 ;
      RECT 52.04 1.855 52.77 2.185 ;
      RECT 49.64 1.855 49.97 2.585 ;
      RECT 48.44 2.015 48.77 2.745 ;
      RECT 38.82 2.015 39.15 2.745 ;
      RECT 37.62 2.88 37.95 3.61 ;
      RECT 36.78 1.855 37.51 2.185 ;
      RECT 34.38 1.855 34.71 2.585 ;
      RECT 33.18 2.015 33.51 2.745 ;
      RECT 23.56 2.015 23.89 2.745 ;
      RECT 22.36 2.88 22.69 3.61 ;
      RECT 21.52 1.855 22.25 2.185 ;
      RECT 19.12 1.855 19.45 2.585 ;
      RECT 17.92 2.015 18.25 2.745 ;
      RECT 8.3 2.015 8.63 2.745 ;
      RECT 7.1 2.88 7.43 3.61 ;
      RECT 6.26 1.855 6.99 2.185 ;
      RECT 3.86 1.855 4.19 2.585 ;
      RECT 2.66 2.015 2.99 2.745 ;
    LAYER via2 ;
      RECT 69.405 2.48 69.605 2.68 ;
      RECT 68.205 3.04 68.405 3.24 ;
      RECT 67.365 1.92 67.565 2.12 ;
      RECT 67.325 7.14 67.525 7.34 ;
      RECT 66.285 2.825 66.485 3.025 ;
      RECT 65.925 1.92 66.125 2.12 ;
      RECT 64.965 1.92 65.165 2.12 ;
      RECT 63.765 2.48 63.965 2.68 ;
      RECT 63.045 2.48 63.245 2.68 ;
      RECT 54.145 2.48 54.345 2.68 ;
      RECT 52.945 3.04 53.145 3.24 ;
      RECT 52.105 1.92 52.305 2.12 ;
      RECT 52.065 7.14 52.265 7.34 ;
      RECT 51.025 2.825 51.225 3.025 ;
      RECT 50.665 1.92 50.865 2.12 ;
      RECT 49.705 1.92 49.905 2.12 ;
      RECT 48.505 2.48 48.705 2.68 ;
      RECT 47.785 2.48 47.985 2.68 ;
      RECT 38.885 2.48 39.085 2.68 ;
      RECT 37.685 3.04 37.885 3.24 ;
      RECT 36.845 1.92 37.045 2.12 ;
      RECT 36.805 7.14 37.005 7.34 ;
      RECT 35.765 2.825 35.965 3.025 ;
      RECT 35.405 1.92 35.605 2.12 ;
      RECT 34.445 1.92 34.645 2.12 ;
      RECT 33.245 2.48 33.445 2.68 ;
      RECT 32.525 2.48 32.725 2.68 ;
      RECT 23.625 2.48 23.825 2.68 ;
      RECT 22.425 3.04 22.625 3.24 ;
      RECT 21.585 1.92 21.785 2.12 ;
      RECT 21.545 7.14 21.745 7.34 ;
      RECT 20.505 2.825 20.705 3.025 ;
      RECT 20.145 1.92 20.345 2.12 ;
      RECT 19.185 1.92 19.385 2.12 ;
      RECT 17.985 2.48 18.185 2.68 ;
      RECT 17.265 2.48 17.465 2.68 ;
      RECT 8.365 2.48 8.565 2.68 ;
      RECT 7.165 3.04 7.365 3.24 ;
      RECT 6.325 1.92 6.525 2.12 ;
      RECT 6.285 7.14 6.485 7.34 ;
      RECT 5.245 2.825 5.445 3.025 ;
      RECT 4.885 1.92 5.085 2.12 ;
      RECT 3.925 1.92 4.125 2.12 ;
      RECT 2.725 2.48 2.925 2.68 ;
      RECT 2.005 2.48 2.205 2.68 ;
    LAYER met2 ;
      RECT -1.565 8.4 75.93 8.57 ;
      RECT 75.76 7.275 75.93 8.57 ;
      RECT -1.565 6.255 -1.395 8.57 ;
      RECT 75.73 7.275 76.08 7.625 ;
      RECT -1.63 6.255 -1.34 6.605 ;
      RECT 72.57 6.22 72.89 6.545 ;
      RECT 72.6 5.695 72.77 6.545 ;
      RECT 72.6 5.695 72.775 6.045 ;
      RECT 72.6 5.695 73.575 5.87 ;
      RECT 73.4 1.965 73.575 5.87 ;
      RECT 73.345 1.965 73.695 2.315 ;
      RECT 73.37 6.655 73.695 6.98 ;
      RECT 72.255 6.745 73.695 6.915 ;
      RECT 72.255 2.395 72.415 6.915 ;
      RECT 72.57 2.365 72.89 2.685 ;
      RECT 72.255 2.395 72.89 2.565 ;
      RECT 71.52 5.86 71.86 6.21 ;
      RECT 71.6 2.705 71.775 6.21 ;
      RECT 71.525 2.705 71.865 3.055 ;
      RECT 70.965 2.705 71.305 3.055 ;
      RECT 70.36 2.77 71.305 2.97 ;
      RECT 70.36 2.765 70.575 2.97 ;
      RECT 70.375 2.34 70.575 2.97 ;
      RECT 69.365 2.34 69.645 2.72 ;
      RECT 71.055 2.7 71.225 3.055 ;
      RECT 69.36 2.34 69.645 2.673 ;
      RECT 69.34 2.34 69.645 2.65 ;
      RECT 69.33 2.34 69.645 2.63 ;
      RECT 69.32 2.34 69.645 2.615 ;
      RECT 69.295 2.34 69.645 2.588 ;
      RECT 69.285 2.34 69.645 2.563 ;
      RECT 69.24 2.295 69.52 2.555 ;
      RECT 69.24 2.34 70.575 2.54 ;
      RECT 69.24 2.335 69.565 2.555 ;
      RECT 69.24 2.327 69.56 2.555 ;
      RECT 69.24 2.317 69.555 2.555 ;
      RECT 69.24 2.305 69.55 2.555 ;
      RECT 68.165 3 68.445 3.28 ;
      RECT 68.165 3 68.48 3.26 ;
      RECT 60.445 6.655 60.795 7.005 ;
      RECT 67.91 6.61 68.26 6.96 ;
      RECT 60.445 6.685 68.26 6.885 ;
      RECT 68.2 2.42 68.25 2.68 ;
      RECT 67.99 2.42 67.995 2.68 ;
      RECT 67.185 1.975 67.215 2.235 ;
      RECT 66.955 1.975 67.03 2.235 ;
      RECT 68.175 2.37 68.2 2.68 ;
      RECT 68.17 2.327 68.175 2.68 ;
      RECT 68.165 2.31 68.17 2.68 ;
      RECT 68.16 2.297 68.165 2.68 ;
      RECT 68.085 2.18 68.16 2.68 ;
      RECT 68.04 1.997 68.085 2.68 ;
      RECT 68.035 1.925 68.04 2.68 ;
      RECT 68.02 1.9 68.035 2.68 ;
      RECT 67.995 1.862 68.02 2.68 ;
      RECT 67.985 1.842 67.995 2.402 ;
      RECT 67.97 1.834 67.985 2.357 ;
      RECT 67.965 1.826 67.97 2.328 ;
      RECT 67.96 1.823 67.965 2.308 ;
      RECT 67.955 1.82 67.96 2.288 ;
      RECT 67.95 1.817 67.955 2.268 ;
      RECT 67.92 1.806 67.95 2.205 ;
      RECT 67.9 1.791 67.92 2.12 ;
      RECT 67.895 1.783 67.9 2.083 ;
      RECT 67.885 1.777 67.895 2.05 ;
      RECT 67.87 1.769 67.885 2.01 ;
      RECT 67.865 1.762 67.87 1.97 ;
      RECT 67.86 1.759 67.865 1.948 ;
      RECT 67.855 1.756 67.86 1.935 ;
      RECT 67.85 1.755 67.855 1.925 ;
      RECT 67.835 1.749 67.85 1.915 ;
      RECT 67.81 1.736 67.835 1.9 ;
      RECT 67.76 1.711 67.81 1.871 ;
      RECT 67.745 1.69 67.76 1.846 ;
      RECT 67.735 1.683 67.745 1.835 ;
      RECT 67.68 1.664 67.735 1.808 ;
      RECT 67.655 1.642 67.68 1.781 ;
      RECT 67.65 1.635 67.655 1.776 ;
      RECT 67.635 1.635 67.65 1.774 ;
      RECT 67.61 1.627 67.635 1.77 ;
      RECT 67.595 1.625 67.61 1.766 ;
      RECT 67.565 1.625 67.595 1.763 ;
      RECT 67.555 1.625 67.565 1.758 ;
      RECT 67.51 1.625 67.555 1.756 ;
      RECT 67.481 1.625 67.51 1.757 ;
      RECT 67.395 1.625 67.481 1.759 ;
      RECT 67.381 1.626 67.395 1.761 ;
      RECT 67.295 1.627 67.381 1.763 ;
      RECT 67.28 1.628 67.295 1.773 ;
      RECT 67.275 1.629 67.28 1.782 ;
      RECT 67.255 1.632 67.275 1.792 ;
      RECT 67.24 1.64 67.255 1.807 ;
      RECT 67.22 1.658 67.24 1.822 ;
      RECT 67.21 1.67 67.22 1.845 ;
      RECT 67.2 1.679 67.21 1.875 ;
      RECT 67.185 1.691 67.2 1.92 ;
      RECT 67.13 1.724 67.185 2.235 ;
      RECT 67.125 1.752 67.13 2.235 ;
      RECT 67.105 1.767 67.125 2.235 ;
      RECT 67.07 1.827 67.105 2.235 ;
      RECT 67.068 1.877 67.07 2.235 ;
      RECT 67.065 1.885 67.068 2.235 ;
      RECT 67.055 1.9 67.065 2.235 ;
      RECT 67.05 1.912 67.055 2.235 ;
      RECT 67.04 1.937 67.05 2.235 ;
      RECT 67.03 1.965 67.04 2.235 ;
      RECT 64.935 3.47 64.985 3.73 ;
      RECT 67.845 3.02 67.905 3.28 ;
      RECT 67.83 3.02 67.845 3.29 ;
      RECT 67.811 3.02 67.83 3.323 ;
      RECT 67.725 3.02 67.811 3.448 ;
      RECT 67.645 3.02 67.725 3.63 ;
      RECT 67.64 3.257 67.645 3.715 ;
      RECT 67.615 3.327 67.64 3.743 ;
      RECT 67.61 3.397 67.615 3.77 ;
      RECT 67.59 3.469 67.61 3.792 ;
      RECT 67.585 3.536 67.59 3.815 ;
      RECT 67.575 3.565 67.585 3.83 ;
      RECT 67.565 3.587 67.575 3.847 ;
      RECT 67.56 3.597 67.565 3.858 ;
      RECT 67.555 3.605 67.56 3.866 ;
      RECT 67.545 3.613 67.555 3.878 ;
      RECT 67.54 3.625 67.545 3.888 ;
      RECT 67.535 3.633 67.54 3.893 ;
      RECT 67.515 3.651 67.535 3.903 ;
      RECT 67.51 3.668 67.515 3.91 ;
      RECT 67.505 3.676 67.51 3.911 ;
      RECT 67.5 3.687 67.505 3.913 ;
      RECT 67.46 3.725 67.5 3.923 ;
      RECT 67.455 3.76 67.46 3.934 ;
      RECT 67.45 3.765 67.455 3.937 ;
      RECT 67.425 3.775 67.45 3.944 ;
      RECT 67.415 3.789 67.425 3.953 ;
      RECT 67.395 3.801 67.415 3.956 ;
      RECT 67.345 3.82 67.395 3.96 ;
      RECT 67.3 3.835 67.345 3.965 ;
      RECT 67.235 3.838 67.3 3.971 ;
      RECT 67.22 3.836 67.235 3.978 ;
      RECT 67.19 3.835 67.22 3.978 ;
      RECT 67.151 3.834 67.19 3.974 ;
      RECT 67.065 3.831 67.151 3.97 ;
      RECT 67.048 3.829 67.065 3.967 ;
      RECT 66.962 3.827 67.048 3.964 ;
      RECT 66.876 3.824 66.962 3.958 ;
      RECT 66.79 3.82 66.876 3.953 ;
      RECT 66.712 3.817 66.79 3.949 ;
      RECT 66.626 3.814 66.712 3.947 ;
      RECT 66.54 3.811 66.626 3.944 ;
      RECT 66.482 3.809 66.54 3.941 ;
      RECT 66.396 3.806 66.482 3.939 ;
      RECT 66.31 3.802 66.396 3.937 ;
      RECT 66.224 3.799 66.31 3.934 ;
      RECT 66.138 3.795 66.224 3.932 ;
      RECT 66.052 3.791 66.138 3.929 ;
      RECT 65.966 3.788 66.052 3.927 ;
      RECT 65.88 3.784 65.966 3.924 ;
      RECT 65.794 3.781 65.88 3.922 ;
      RECT 65.708 3.777 65.794 3.919 ;
      RECT 65.622 3.774 65.708 3.917 ;
      RECT 65.536 3.77 65.622 3.914 ;
      RECT 65.45 3.767 65.536 3.912 ;
      RECT 65.44 3.765 65.45 3.908 ;
      RECT 65.435 3.765 65.44 3.906 ;
      RECT 65.395 3.76 65.435 3.9 ;
      RECT 65.381 3.751 65.395 3.893 ;
      RECT 65.295 3.721 65.381 3.878 ;
      RECT 65.275 3.687 65.295 3.863 ;
      RECT 65.205 3.656 65.275 3.85 ;
      RECT 65.2 3.631 65.205 3.839 ;
      RECT 65.195 3.625 65.2 3.837 ;
      RECT 65.126 3.47 65.195 3.825 ;
      RECT 65.04 3.47 65.126 3.799 ;
      RECT 65.015 3.47 65.04 3.778 ;
      RECT 65.01 3.47 65.015 3.768 ;
      RECT 65.005 3.47 65.01 3.76 ;
      RECT 64.985 3.47 65.005 3.743 ;
      RECT 67.405 2.04 67.665 2.3 ;
      RECT 67.39 2.04 67.665 2.203 ;
      RECT 67.36 2.04 67.665 2.178 ;
      RECT 67.325 1.88 67.605 2.16 ;
      RECT 67.295 3.37 67.355 3.63 ;
      RECT 66.32 2.06 66.375 2.32 ;
      RECT 67.255 3.327 67.295 3.63 ;
      RECT 67.226 3.248 67.255 3.63 ;
      RECT 67.14 3.12 67.226 3.63 ;
      RECT 67.12 3 67.14 3.63 ;
      RECT 67.095 2.951 67.12 3.63 ;
      RECT 67.09 2.916 67.095 3.48 ;
      RECT 67.06 2.876 67.09 3.418 ;
      RECT 67.035 2.813 67.06 3.333 ;
      RECT 67.025 2.775 67.035 3.27 ;
      RECT 67.01 2.75 67.025 3.231 ;
      RECT 66.967 2.708 67.01 3.137 ;
      RECT 66.965 2.681 66.967 3.064 ;
      RECT 66.96 2.676 66.965 3.055 ;
      RECT 66.955 2.669 66.96 3.03 ;
      RECT 66.95 2.663 66.955 3.015 ;
      RECT 66.945 2.657 66.95 3.003 ;
      RECT 66.935 2.648 66.945 2.985 ;
      RECT 66.93 2.639 66.935 2.963 ;
      RECT 66.905 2.62 66.93 2.913 ;
      RECT 66.9 2.601 66.905 2.863 ;
      RECT 66.885 2.587 66.9 2.823 ;
      RECT 66.88 2.573 66.885 2.79 ;
      RECT 66.875 2.566 66.88 2.783 ;
      RECT 66.86 2.553 66.875 2.775 ;
      RECT 66.815 2.515 66.86 2.748 ;
      RECT 66.785 2.468 66.815 2.713 ;
      RECT 66.765 2.437 66.785 2.69 ;
      RECT 66.685 2.37 66.765 2.643 ;
      RECT 66.655 2.3 66.685 2.59 ;
      RECT 66.65 2.277 66.655 2.573 ;
      RECT 66.62 2.255 66.65 2.558 ;
      RECT 66.59 2.214 66.62 2.53 ;
      RECT 66.585 2.189 66.59 2.515 ;
      RECT 66.58 2.183 66.585 2.508 ;
      RECT 66.57 2.06 66.58 2.5 ;
      RECT 66.56 2.06 66.57 2.493 ;
      RECT 66.555 2.06 66.56 2.485 ;
      RECT 66.535 2.06 66.555 2.473 ;
      RECT 66.485 2.06 66.535 2.443 ;
      RECT 66.43 2.06 66.485 2.393 ;
      RECT 66.4 2.06 66.43 2.353 ;
      RECT 66.375 2.06 66.4 2.33 ;
      RECT 66.245 2.785 66.525 3.065 ;
      RECT 66.21 2.7 66.47 2.96 ;
      RECT 66.21 2.782 66.48 2.96 ;
      RECT 64.41 2.155 64.415 2.64 ;
      RECT 64.3 2.34 64.305 2.64 ;
      RECT 64.21 2.38 64.275 2.64 ;
      RECT 65.885 1.88 65.975 2.51 ;
      RECT 65.85 1.93 65.855 2.51 ;
      RECT 65.795 1.955 65.805 2.51 ;
      RECT 65.75 1.955 65.76 2.51 ;
      RECT 66.12 1.88 66.165 2.16 ;
      RECT 64.97 1.61 65.17 1.75 ;
      RECT 66.086 1.88 66.12 2.172 ;
      RECT 66 1.88 66.086 2.212 ;
      RECT 65.985 1.88 66 2.253 ;
      RECT 65.98 1.88 65.985 2.273 ;
      RECT 65.975 1.88 65.98 2.293 ;
      RECT 65.855 1.922 65.885 2.51 ;
      RECT 65.805 1.942 65.85 2.51 ;
      RECT 65.79 1.957 65.795 2.51 ;
      RECT 65.76 1.957 65.79 2.51 ;
      RECT 65.715 1.942 65.75 2.51 ;
      RECT 65.71 1.93 65.715 2.29 ;
      RECT 65.705 1.927 65.71 2.27 ;
      RECT 65.69 1.917 65.705 2.223 ;
      RECT 65.685 1.91 65.69 2.186 ;
      RECT 65.68 1.907 65.685 2.169 ;
      RECT 65.665 1.897 65.68 2.125 ;
      RECT 65.66 1.888 65.665 2.085 ;
      RECT 65.655 1.884 65.66 2.07 ;
      RECT 65.645 1.878 65.655 2.053 ;
      RECT 65.605 1.859 65.645 2.028 ;
      RECT 65.6 1.841 65.605 2.008 ;
      RECT 65.59 1.835 65.6 2.003 ;
      RECT 65.56 1.819 65.59 1.99 ;
      RECT 65.545 1.801 65.56 1.973 ;
      RECT 65.53 1.789 65.545 1.96 ;
      RECT 65.525 1.781 65.53 1.953 ;
      RECT 65.495 1.767 65.525 1.94 ;
      RECT 65.49 1.752 65.495 1.928 ;
      RECT 65.48 1.746 65.49 1.92 ;
      RECT 65.46 1.734 65.48 1.908 ;
      RECT 65.45 1.722 65.46 1.895 ;
      RECT 65.42 1.706 65.45 1.88 ;
      RECT 65.4 1.686 65.42 1.863 ;
      RECT 65.395 1.676 65.4 1.853 ;
      RECT 65.37 1.664 65.395 1.84 ;
      RECT 65.365 1.652 65.37 1.828 ;
      RECT 65.36 1.647 65.365 1.824 ;
      RECT 65.345 1.64 65.36 1.816 ;
      RECT 65.335 1.627 65.345 1.806 ;
      RECT 65.33 1.625 65.335 1.8 ;
      RECT 65.305 1.618 65.33 1.789 ;
      RECT 65.3 1.611 65.305 1.778 ;
      RECT 65.275 1.61 65.3 1.765 ;
      RECT 65.256 1.61 65.275 1.755 ;
      RECT 65.17 1.61 65.256 1.752 ;
      RECT 64.94 1.61 64.97 1.755 ;
      RECT 64.9 1.617 64.94 1.768 ;
      RECT 64.875 1.627 64.9 1.781 ;
      RECT 64.86 1.636 64.875 1.791 ;
      RECT 64.83 1.641 64.86 1.81 ;
      RECT 64.825 1.647 64.83 1.828 ;
      RECT 64.805 1.657 64.825 1.843 ;
      RECT 64.795 1.67 64.805 1.863 ;
      RECT 64.78 1.682 64.795 1.88 ;
      RECT 64.775 1.692 64.78 1.89 ;
      RECT 64.77 1.697 64.775 1.895 ;
      RECT 64.76 1.705 64.77 1.908 ;
      RECT 64.71 1.737 64.76 1.945 ;
      RECT 64.695 1.772 64.71 1.986 ;
      RECT 64.69 1.782 64.695 2.001 ;
      RECT 64.685 1.787 64.69 2.008 ;
      RECT 64.66 1.803 64.685 2.028 ;
      RECT 64.645 1.824 64.66 2.053 ;
      RECT 64.62 1.845 64.645 2.078 ;
      RECT 64.61 1.864 64.62 2.101 ;
      RECT 64.585 1.882 64.61 2.124 ;
      RECT 64.57 1.902 64.585 2.148 ;
      RECT 64.565 1.912 64.57 2.16 ;
      RECT 64.55 1.924 64.565 2.18 ;
      RECT 64.54 1.939 64.55 2.22 ;
      RECT 64.535 1.947 64.54 2.248 ;
      RECT 64.525 1.957 64.535 2.268 ;
      RECT 64.52 1.97 64.525 2.293 ;
      RECT 64.515 1.983 64.52 2.313 ;
      RECT 64.51 1.989 64.515 2.335 ;
      RECT 64.5 1.998 64.51 2.355 ;
      RECT 64.495 2.018 64.5 2.378 ;
      RECT 64.49 2.024 64.495 2.398 ;
      RECT 64.485 2.031 64.49 2.42 ;
      RECT 64.48 2.042 64.485 2.433 ;
      RECT 64.47 2.052 64.48 2.458 ;
      RECT 64.45 2.077 64.47 2.64 ;
      RECT 64.42 2.117 64.45 2.64 ;
      RECT 64.415 2.147 64.42 2.64 ;
      RECT 64.39 2.175 64.41 2.64 ;
      RECT 64.36 2.22 64.39 2.64 ;
      RECT 64.355 2.247 64.36 2.64 ;
      RECT 64.335 2.265 64.355 2.64 ;
      RECT 64.325 2.29 64.335 2.64 ;
      RECT 64.32 2.302 64.325 2.64 ;
      RECT 64.305 2.325 64.32 2.64 ;
      RECT 64.285 2.352 64.3 2.64 ;
      RECT 64.275 2.375 64.285 2.64 ;
      RECT 66.065 3.26 66.145 3.52 ;
      RECT 65.3 2.48 65.37 2.74 ;
      RECT 66.031 3.227 66.065 3.52 ;
      RECT 65.945 3.13 66.031 3.52 ;
      RECT 65.925 3.042 65.945 3.52 ;
      RECT 65.915 3.012 65.925 3.52 ;
      RECT 65.905 2.992 65.915 3.52 ;
      RECT 65.885 2.979 65.905 3.52 ;
      RECT 65.87 2.969 65.885 3.348 ;
      RECT 65.865 2.962 65.87 3.303 ;
      RECT 65.855 2.956 65.865 3.293 ;
      RECT 65.845 2.948 65.855 3.275 ;
      RECT 65.84 2.942 65.845 3.263 ;
      RECT 65.83 2.937 65.84 3.25 ;
      RECT 65.81 2.927 65.83 3.223 ;
      RECT 65.77 2.906 65.81 3.175 ;
      RECT 65.755 2.887 65.77 3.133 ;
      RECT 65.73 2.873 65.755 3.103 ;
      RECT 65.72 2.861 65.73 3.07 ;
      RECT 65.715 2.856 65.72 3.06 ;
      RECT 65.685 2.842 65.715 3.04 ;
      RECT 65.675 2.826 65.685 3.013 ;
      RECT 65.67 2.821 65.675 3.003 ;
      RECT 65.645 2.812 65.67 2.983 ;
      RECT 65.635 2.8 65.645 2.963 ;
      RECT 65.565 2.768 65.635 2.938 ;
      RECT 65.56 2.737 65.565 2.915 ;
      RECT 65.511 2.48 65.56 2.898 ;
      RECT 65.425 2.48 65.511 2.857 ;
      RECT 65.37 2.48 65.425 2.785 ;
      RECT 65.46 3.265 65.62 3.525 ;
      RECT 64.985 1.88 65.035 2.565 ;
      RECT 64.775 2.305 64.81 2.565 ;
      RECT 65.09 1.88 65.095 2.34 ;
      RECT 65.18 1.88 65.205 2.16 ;
      RECT 65.455 3.262 65.46 3.525 ;
      RECT 65.42 3.25 65.455 3.525 ;
      RECT 65.36 3.223 65.42 3.525 ;
      RECT 65.355 3.206 65.36 3.379 ;
      RECT 65.35 3.203 65.355 3.366 ;
      RECT 65.33 3.196 65.35 3.353 ;
      RECT 65.295 3.179 65.33 3.335 ;
      RECT 65.255 3.158 65.295 3.315 ;
      RECT 65.25 3.146 65.255 3.303 ;
      RECT 65.21 3.132 65.25 3.289 ;
      RECT 65.19 3.115 65.21 3.271 ;
      RECT 65.18 3.107 65.19 3.263 ;
      RECT 65.165 1.88 65.18 2.178 ;
      RECT 65.15 3.097 65.18 3.25 ;
      RECT 65.135 1.88 65.165 2.223 ;
      RECT 65.14 3.087 65.15 3.237 ;
      RECT 65.11 3.072 65.14 3.224 ;
      RECT 65.095 1.88 65.135 2.29 ;
      RECT 65.095 3.04 65.11 3.21 ;
      RECT 65.09 3.012 65.095 3.204 ;
      RECT 65.085 1.88 65.09 2.345 ;
      RECT 65.075 2.982 65.09 3.198 ;
      RECT 65.08 1.88 65.085 2.358 ;
      RECT 65.07 1.88 65.08 2.378 ;
      RECT 65.035 2.895 65.075 3.183 ;
      RECT 65.035 1.88 65.07 2.418 ;
      RECT 65.03 2.827 65.035 3.171 ;
      RECT 65.015 2.782 65.03 3.166 ;
      RECT 65.01 2.72 65.015 3.161 ;
      RECT 64.985 2.627 65.01 3.154 ;
      RECT 64.98 1.88 64.985 3.146 ;
      RECT 64.965 1.88 64.98 3.133 ;
      RECT 64.945 1.88 64.965 3.09 ;
      RECT 64.935 1.88 64.945 3.04 ;
      RECT 64.93 1.88 64.935 3.013 ;
      RECT 64.925 1.88 64.93 2.991 ;
      RECT 64.92 2.106 64.925 2.974 ;
      RECT 64.915 2.128 64.92 2.952 ;
      RECT 64.91 2.17 64.915 2.935 ;
      RECT 64.88 2.22 64.91 2.879 ;
      RECT 64.875 2.247 64.88 2.821 ;
      RECT 64.86 2.265 64.875 2.785 ;
      RECT 64.855 2.283 64.86 2.749 ;
      RECT 64.849 2.29 64.855 2.73 ;
      RECT 64.845 2.297 64.849 2.713 ;
      RECT 64.84 2.302 64.845 2.682 ;
      RECT 64.83 2.305 64.84 2.657 ;
      RECT 64.82 2.305 64.83 2.623 ;
      RECT 64.815 2.305 64.82 2.6 ;
      RECT 64.81 2.305 64.815 2.58 ;
      RECT 63.725 2.44 64.005 2.72 ;
      RECT 63.725 2.44 64.025 2.615 ;
      RECT 63.815 2.33 64.075 2.59 ;
      RECT 63.78 2.425 64.075 2.59 ;
      RECT 63.905 0.945 64.07 2.59 ;
      RECT 63.805 0.945 64.175 1.315 ;
      RECT 63.43 3.47 63.69 3.73 ;
      RECT 63.45 3.397 63.63 3.73 ;
      RECT 63.45 3.14 63.625 3.73 ;
      RECT 63.45 2.932 63.615 3.73 ;
      RECT 63.455 2.85 63.615 3.73 ;
      RECT 63.455 2.615 63.605 3.73 ;
      RECT 63.455 2.462 63.6 3.73 ;
      RECT 63.46 2.447 63.6 3.73 ;
      RECT 63.51 2.162 63.6 3.73 ;
      RECT 63.465 2.397 63.6 3.73 ;
      RECT 63.495 2.215 63.6 3.73 ;
      RECT 63.48 2.327 63.6 3.73 ;
      RECT 63.485 2.285 63.6 3.73 ;
      RECT 63.48 2.327 63.615 2.39 ;
      RECT 63.515 1.915 63.62 2.335 ;
      RECT 63.515 1.915 63.635 2.318 ;
      RECT 63.515 1.915 63.67 2.28 ;
      RECT 63.51 2.162 63.72 2.213 ;
      RECT 63.515 1.915 63.775 2.175 ;
      RECT 62.775 2.62 63.035 2.88 ;
      RECT 62.775 2.62 63.045 2.838 ;
      RECT 62.775 2.62 63.131 2.809 ;
      RECT 62.775 2.62 63.2 2.761 ;
      RECT 62.775 2.62 63.235 2.73 ;
      RECT 63.005 2.44 63.285 2.72 ;
      RECT 62.84 2.605 63.285 2.72 ;
      RECT 62.93 2.482 63.035 2.88 ;
      RECT 62.86 2.545 63.285 2.72 ;
      RECT 57.31 6.22 57.63 6.545 ;
      RECT 57.34 5.695 57.51 6.545 ;
      RECT 57.34 5.695 57.515 6.045 ;
      RECT 57.34 5.695 58.315 5.87 ;
      RECT 58.14 1.965 58.315 5.87 ;
      RECT 58.085 1.965 58.435 2.315 ;
      RECT 58.11 6.655 58.435 6.98 ;
      RECT 56.995 6.745 58.435 6.915 ;
      RECT 56.995 2.395 57.155 6.915 ;
      RECT 57.31 2.365 57.63 2.685 ;
      RECT 56.995 2.395 57.63 2.565 ;
      RECT 56.26 5.86 56.6 6.21 ;
      RECT 56.34 2.705 56.515 6.21 ;
      RECT 56.265 2.705 56.605 3.055 ;
      RECT 55.705 2.705 56.045 3.055 ;
      RECT 55.1 2.77 56.045 2.97 ;
      RECT 55.1 2.765 55.315 2.97 ;
      RECT 55.115 2.34 55.315 2.97 ;
      RECT 54.105 2.34 54.385 2.72 ;
      RECT 55.795 2.7 55.965 3.055 ;
      RECT 54.1 2.34 54.385 2.673 ;
      RECT 54.08 2.34 54.385 2.65 ;
      RECT 54.07 2.34 54.385 2.63 ;
      RECT 54.06 2.34 54.385 2.615 ;
      RECT 54.035 2.34 54.385 2.588 ;
      RECT 54.025 2.34 54.385 2.563 ;
      RECT 53.98 2.295 54.26 2.555 ;
      RECT 53.98 2.34 55.315 2.54 ;
      RECT 53.98 2.335 54.305 2.555 ;
      RECT 53.98 2.327 54.3 2.555 ;
      RECT 53.98 2.317 54.295 2.555 ;
      RECT 53.98 2.305 54.29 2.555 ;
      RECT 52.905 3 53.185 3.28 ;
      RECT 52.905 3 53.22 3.26 ;
      RECT 45.185 6.655 45.535 7.005 ;
      RECT 52.65 6.61 53 6.96 ;
      RECT 45.185 6.685 53 6.885 ;
      RECT 52.94 2.42 52.99 2.68 ;
      RECT 52.73 2.42 52.735 2.68 ;
      RECT 51.925 1.975 51.955 2.235 ;
      RECT 51.695 1.975 51.77 2.235 ;
      RECT 52.915 2.37 52.94 2.68 ;
      RECT 52.91 2.327 52.915 2.68 ;
      RECT 52.905 2.31 52.91 2.68 ;
      RECT 52.9 2.297 52.905 2.68 ;
      RECT 52.825 2.18 52.9 2.68 ;
      RECT 52.78 1.997 52.825 2.68 ;
      RECT 52.775 1.925 52.78 2.68 ;
      RECT 52.76 1.9 52.775 2.68 ;
      RECT 52.735 1.862 52.76 2.68 ;
      RECT 52.725 1.842 52.735 2.402 ;
      RECT 52.71 1.834 52.725 2.357 ;
      RECT 52.705 1.826 52.71 2.328 ;
      RECT 52.7 1.823 52.705 2.308 ;
      RECT 52.695 1.82 52.7 2.288 ;
      RECT 52.69 1.817 52.695 2.268 ;
      RECT 52.66 1.806 52.69 2.205 ;
      RECT 52.64 1.791 52.66 2.12 ;
      RECT 52.635 1.783 52.64 2.083 ;
      RECT 52.625 1.777 52.635 2.05 ;
      RECT 52.61 1.769 52.625 2.01 ;
      RECT 52.605 1.762 52.61 1.97 ;
      RECT 52.6 1.759 52.605 1.948 ;
      RECT 52.595 1.756 52.6 1.935 ;
      RECT 52.59 1.755 52.595 1.925 ;
      RECT 52.575 1.749 52.59 1.915 ;
      RECT 52.55 1.736 52.575 1.9 ;
      RECT 52.5 1.711 52.55 1.871 ;
      RECT 52.485 1.69 52.5 1.846 ;
      RECT 52.475 1.683 52.485 1.835 ;
      RECT 52.42 1.664 52.475 1.808 ;
      RECT 52.395 1.642 52.42 1.781 ;
      RECT 52.39 1.635 52.395 1.776 ;
      RECT 52.375 1.635 52.39 1.774 ;
      RECT 52.35 1.627 52.375 1.77 ;
      RECT 52.335 1.625 52.35 1.766 ;
      RECT 52.305 1.625 52.335 1.763 ;
      RECT 52.295 1.625 52.305 1.758 ;
      RECT 52.25 1.625 52.295 1.756 ;
      RECT 52.221 1.625 52.25 1.757 ;
      RECT 52.135 1.625 52.221 1.759 ;
      RECT 52.121 1.626 52.135 1.761 ;
      RECT 52.035 1.627 52.121 1.763 ;
      RECT 52.02 1.628 52.035 1.773 ;
      RECT 52.015 1.629 52.02 1.782 ;
      RECT 51.995 1.632 52.015 1.792 ;
      RECT 51.98 1.64 51.995 1.807 ;
      RECT 51.96 1.658 51.98 1.822 ;
      RECT 51.95 1.67 51.96 1.845 ;
      RECT 51.94 1.679 51.95 1.875 ;
      RECT 51.925 1.691 51.94 1.92 ;
      RECT 51.87 1.724 51.925 2.235 ;
      RECT 51.865 1.752 51.87 2.235 ;
      RECT 51.845 1.767 51.865 2.235 ;
      RECT 51.81 1.827 51.845 2.235 ;
      RECT 51.808 1.877 51.81 2.235 ;
      RECT 51.805 1.885 51.808 2.235 ;
      RECT 51.795 1.9 51.805 2.235 ;
      RECT 51.79 1.912 51.795 2.235 ;
      RECT 51.78 1.937 51.79 2.235 ;
      RECT 51.77 1.965 51.78 2.235 ;
      RECT 49.675 3.47 49.725 3.73 ;
      RECT 52.585 3.02 52.645 3.28 ;
      RECT 52.57 3.02 52.585 3.29 ;
      RECT 52.551 3.02 52.57 3.323 ;
      RECT 52.465 3.02 52.551 3.448 ;
      RECT 52.385 3.02 52.465 3.63 ;
      RECT 52.38 3.257 52.385 3.715 ;
      RECT 52.355 3.327 52.38 3.743 ;
      RECT 52.35 3.397 52.355 3.77 ;
      RECT 52.33 3.469 52.35 3.792 ;
      RECT 52.325 3.536 52.33 3.815 ;
      RECT 52.315 3.565 52.325 3.83 ;
      RECT 52.305 3.587 52.315 3.847 ;
      RECT 52.3 3.597 52.305 3.858 ;
      RECT 52.295 3.605 52.3 3.866 ;
      RECT 52.285 3.613 52.295 3.878 ;
      RECT 52.28 3.625 52.285 3.888 ;
      RECT 52.275 3.633 52.28 3.893 ;
      RECT 52.255 3.651 52.275 3.903 ;
      RECT 52.25 3.668 52.255 3.91 ;
      RECT 52.245 3.676 52.25 3.911 ;
      RECT 52.24 3.687 52.245 3.913 ;
      RECT 52.2 3.725 52.24 3.923 ;
      RECT 52.195 3.76 52.2 3.934 ;
      RECT 52.19 3.765 52.195 3.937 ;
      RECT 52.165 3.775 52.19 3.944 ;
      RECT 52.155 3.789 52.165 3.953 ;
      RECT 52.135 3.801 52.155 3.956 ;
      RECT 52.085 3.82 52.135 3.96 ;
      RECT 52.04 3.835 52.085 3.965 ;
      RECT 51.975 3.838 52.04 3.971 ;
      RECT 51.96 3.836 51.975 3.978 ;
      RECT 51.93 3.835 51.96 3.978 ;
      RECT 51.891 3.834 51.93 3.974 ;
      RECT 51.805 3.831 51.891 3.97 ;
      RECT 51.788 3.829 51.805 3.967 ;
      RECT 51.702 3.827 51.788 3.964 ;
      RECT 51.616 3.824 51.702 3.958 ;
      RECT 51.53 3.82 51.616 3.953 ;
      RECT 51.452 3.817 51.53 3.949 ;
      RECT 51.366 3.814 51.452 3.947 ;
      RECT 51.28 3.811 51.366 3.944 ;
      RECT 51.222 3.809 51.28 3.941 ;
      RECT 51.136 3.806 51.222 3.939 ;
      RECT 51.05 3.802 51.136 3.937 ;
      RECT 50.964 3.799 51.05 3.934 ;
      RECT 50.878 3.795 50.964 3.932 ;
      RECT 50.792 3.791 50.878 3.929 ;
      RECT 50.706 3.788 50.792 3.927 ;
      RECT 50.62 3.784 50.706 3.924 ;
      RECT 50.534 3.781 50.62 3.922 ;
      RECT 50.448 3.777 50.534 3.919 ;
      RECT 50.362 3.774 50.448 3.917 ;
      RECT 50.276 3.77 50.362 3.914 ;
      RECT 50.19 3.767 50.276 3.912 ;
      RECT 50.18 3.765 50.19 3.908 ;
      RECT 50.175 3.765 50.18 3.906 ;
      RECT 50.135 3.76 50.175 3.9 ;
      RECT 50.121 3.751 50.135 3.893 ;
      RECT 50.035 3.721 50.121 3.878 ;
      RECT 50.015 3.687 50.035 3.863 ;
      RECT 49.945 3.656 50.015 3.85 ;
      RECT 49.94 3.631 49.945 3.839 ;
      RECT 49.935 3.625 49.94 3.837 ;
      RECT 49.866 3.47 49.935 3.825 ;
      RECT 49.78 3.47 49.866 3.799 ;
      RECT 49.755 3.47 49.78 3.778 ;
      RECT 49.75 3.47 49.755 3.768 ;
      RECT 49.745 3.47 49.75 3.76 ;
      RECT 49.725 3.47 49.745 3.743 ;
      RECT 52.145 2.04 52.405 2.3 ;
      RECT 52.13 2.04 52.405 2.203 ;
      RECT 52.1 2.04 52.405 2.178 ;
      RECT 52.065 1.88 52.345 2.16 ;
      RECT 52.035 3.37 52.095 3.63 ;
      RECT 51.06 2.06 51.115 2.32 ;
      RECT 51.995 3.327 52.035 3.63 ;
      RECT 51.966 3.248 51.995 3.63 ;
      RECT 51.88 3.12 51.966 3.63 ;
      RECT 51.86 3 51.88 3.63 ;
      RECT 51.835 2.951 51.86 3.63 ;
      RECT 51.83 2.916 51.835 3.48 ;
      RECT 51.8 2.876 51.83 3.418 ;
      RECT 51.775 2.813 51.8 3.333 ;
      RECT 51.765 2.775 51.775 3.27 ;
      RECT 51.75 2.75 51.765 3.231 ;
      RECT 51.707 2.708 51.75 3.137 ;
      RECT 51.705 2.681 51.707 3.064 ;
      RECT 51.7 2.676 51.705 3.055 ;
      RECT 51.695 2.669 51.7 3.03 ;
      RECT 51.69 2.663 51.695 3.015 ;
      RECT 51.685 2.657 51.69 3.003 ;
      RECT 51.675 2.648 51.685 2.985 ;
      RECT 51.67 2.639 51.675 2.963 ;
      RECT 51.645 2.62 51.67 2.913 ;
      RECT 51.64 2.601 51.645 2.863 ;
      RECT 51.625 2.587 51.64 2.823 ;
      RECT 51.62 2.573 51.625 2.79 ;
      RECT 51.615 2.566 51.62 2.783 ;
      RECT 51.6 2.553 51.615 2.775 ;
      RECT 51.555 2.515 51.6 2.748 ;
      RECT 51.525 2.468 51.555 2.713 ;
      RECT 51.505 2.437 51.525 2.69 ;
      RECT 51.425 2.37 51.505 2.643 ;
      RECT 51.395 2.3 51.425 2.59 ;
      RECT 51.39 2.277 51.395 2.573 ;
      RECT 51.36 2.255 51.39 2.558 ;
      RECT 51.33 2.214 51.36 2.53 ;
      RECT 51.325 2.189 51.33 2.515 ;
      RECT 51.32 2.183 51.325 2.508 ;
      RECT 51.31 2.06 51.32 2.5 ;
      RECT 51.3 2.06 51.31 2.493 ;
      RECT 51.295 2.06 51.3 2.485 ;
      RECT 51.275 2.06 51.295 2.473 ;
      RECT 51.225 2.06 51.275 2.443 ;
      RECT 51.17 2.06 51.225 2.393 ;
      RECT 51.14 2.06 51.17 2.353 ;
      RECT 51.115 2.06 51.14 2.33 ;
      RECT 50.985 2.785 51.265 3.065 ;
      RECT 50.95 2.7 51.21 2.96 ;
      RECT 50.95 2.782 51.22 2.96 ;
      RECT 49.15 2.155 49.155 2.64 ;
      RECT 49.04 2.34 49.045 2.64 ;
      RECT 48.95 2.38 49.015 2.64 ;
      RECT 50.625 1.88 50.715 2.51 ;
      RECT 50.59 1.93 50.595 2.51 ;
      RECT 50.535 1.955 50.545 2.51 ;
      RECT 50.49 1.955 50.5 2.51 ;
      RECT 50.86 1.88 50.905 2.16 ;
      RECT 49.71 1.61 49.91 1.75 ;
      RECT 50.826 1.88 50.86 2.172 ;
      RECT 50.74 1.88 50.826 2.212 ;
      RECT 50.725 1.88 50.74 2.253 ;
      RECT 50.72 1.88 50.725 2.273 ;
      RECT 50.715 1.88 50.72 2.293 ;
      RECT 50.595 1.922 50.625 2.51 ;
      RECT 50.545 1.942 50.59 2.51 ;
      RECT 50.53 1.957 50.535 2.51 ;
      RECT 50.5 1.957 50.53 2.51 ;
      RECT 50.455 1.942 50.49 2.51 ;
      RECT 50.45 1.93 50.455 2.29 ;
      RECT 50.445 1.927 50.45 2.27 ;
      RECT 50.43 1.917 50.445 2.223 ;
      RECT 50.425 1.91 50.43 2.186 ;
      RECT 50.42 1.907 50.425 2.169 ;
      RECT 50.405 1.897 50.42 2.125 ;
      RECT 50.4 1.888 50.405 2.085 ;
      RECT 50.395 1.884 50.4 2.07 ;
      RECT 50.385 1.878 50.395 2.053 ;
      RECT 50.345 1.859 50.385 2.028 ;
      RECT 50.34 1.841 50.345 2.008 ;
      RECT 50.33 1.835 50.34 2.003 ;
      RECT 50.3 1.819 50.33 1.99 ;
      RECT 50.285 1.801 50.3 1.973 ;
      RECT 50.27 1.789 50.285 1.96 ;
      RECT 50.265 1.781 50.27 1.953 ;
      RECT 50.235 1.767 50.265 1.94 ;
      RECT 50.23 1.752 50.235 1.928 ;
      RECT 50.22 1.746 50.23 1.92 ;
      RECT 50.2 1.734 50.22 1.908 ;
      RECT 50.19 1.722 50.2 1.895 ;
      RECT 50.16 1.706 50.19 1.88 ;
      RECT 50.14 1.686 50.16 1.863 ;
      RECT 50.135 1.676 50.14 1.853 ;
      RECT 50.11 1.664 50.135 1.84 ;
      RECT 50.105 1.652 50.11 1.828 ;
      RECT 50.1 1.647 50.105 1.824 ;
      RECT 50.085 1.64 50.1 1.816 ;
      RECT 50.075 1.627 50.085 1.806 ;
      RECT 50.07 1.625 50.075 1.8 ;
      RECT 50.045 1.618 50.07 1.789 ;
      RECT 50.04 1.611 50.045 1.778 ;
      RECT 50.015 1.61 50.04 1.765 ;
      RECT 49.996 1.61 50.015 1.755 ;
      RECT 49.91 1.61 49.996 1.752 ;
      RECT 49.68 1.61 49.71 1.755 ;
      RECT 49.64 1.617 49.68 1.768 ;
      RECT 49.615 1.627 49.64 1.781 ;
      RECT 49.6 1.636 49.615 1.791 ;
      RECT 49.57 1.641 49.6 1.81 ;
      RECT 49.565 1.647 49.57 1.828 ;
      RECT 49.545 1.657 49.565 1.843 ;
      RECT 49.535 1.67 49.545 1.863 ;
      RECT 49.52 1.682 49.535 1.88 ;
      RECT 49.515 1.692 49.52 1.89 ;
      RECT 49.51 1.697 49.515 1.895 ;
      RECT 49.5 1.705 49.51 1.908 ;
      RECT 49.45 1.737 49.5 1.945 ;
      RECT 49.435 1.772 49.45 1.986 ;
      RECT 49.43 1.782 49.435 2.001 ;
      RECT 49.425 1.787 49.43 2.008 ;
      RECT 49.4 1.803 49.425 2.028 ;
      RECT 49.385 1.824 49.4 2.053 ;
      RECT 49.36 1.845 49.385 2.078 ;
      RECT 49.35 1.864 49.36 2.101 ;
      RECT 49.325 1.882 49.35 2.124 ;
      RECT 49.31 1.902 49.325 2.148 ;
      RECT 49.305 1.912 49.31 2.16 ;
      RECT 49.29 1.924 49.305 2.18 ;
      RECT 49.28 1.939 49.29 2.22 ;
      RECT 49.275 1.947 49.28 2.248 ;
      RECT 49.265 1.957 49.275 2.268 ;
      RECT 49.26 1.97 49.265 2.293 ;
      RECT 49.255 1.983 49.26 2.313 ;
      RECT 49.25 1.989 49.255 2.335 ;
      RECT 49.24 1.998 49.25 2.355 ;
      RECT 49.235 2.018 49.24 2.378 ;
      RECT 49.23 2.024 49.235 2.398 ;
      RECT 49.225 2.031 49.23 2.42 ;
      RECT 49.22 2.042 49.225 2.433 ;
      RECT 49.21 2.052 49.22 2.458 ;
      RECT 49.19 2.077 49.21 2.64 ;
      RECT 49.16 2.117 49.19 2.64 ;
      RECT 49.155 2.147 49.16 2.64 ;
      RECT 49.13 2.175 49.15 2.64 ;
      RECT 49.1 2.22 49.13 2.64 ;
      RECT 49.095 2.247 49.1 2.64 ;
      RECT 49.075 2.265 49.095 2.64 ;
      RECT 49.065 2.29 49.075 2.64 ;
      RECT 49.06 2.302 49.065 2.64 ;
      RECT 49.045 2.325 49.06 2.64 ;
      RECT 49.025 2.352 49.04 2.64 ;
      RECT 49.015 2.375 49.025 2.64 ;
      RECT 50.805 3.26 50.885 3.52 ;
      RECT 50.04 2.48 50.11 2.74 ;
      RECT 50.771 3.227 50.805 3.52 ;
      RECT 50.685 3.13 50.771 3.52 ;
      RECT 50.665 3.042 50.685 3.52 ;
      RECT 50.655 3.012 50.665 3.52 ;
      RECT 50.645 2.992 50.655 3.52 ;
      RECT 50.625 2.979 50.645 3.52 ;
      RECT 50.61 2.969 50.625 3.348 ;
      RECT 50.605 2.962 50.61 3.303 ;
      RECT 50.595 2.956 50.605 3.293 ;
      RECT 50.585 2.948 50.595 3.275 ;
      RECT 50.58 2.942 50.585 3.263 ;
      RECT 50.57 2.937 50.58 3.25 ;
      RECT 50.55 2.927 50.57 3.223 ;
      RECT 50.51 2.906 50.55 3.175 ;
      RECT 50.495 2.887 50.51 3.133 ;
      RECT 50.47 2.873 50.495 3.103 ;
      RECT 50.46 2.861 50.47 3.07 ;
      RECT 50.455 2.856 50.46 3.06 ;
      RECT 50.425 2.842 50.455 3.04 ;
      RECT 50.415 2.826 50.425 3.013 ;
      RECT 50.41 2.821 50.415 3.003 ;
      RECT 50.385 2.812 50.41 2.983 ;
      RECT 50.375 2.8 50.385 2.963 ;
      RECT 50.305 2.768 50.375 2.938 ;
      RECT 50.3 2.737 50.305 2.915 ;
      RECT 50.251 2.48 50.3 2.898 ;
      RECT 50.165 2.48 50.251 2.857 ;
      RECT 50.11 2.48 50.165 2.785 ;
      RECT 50.2 3.265 50.36 3.525 ;
      RECT 49.725 1.88 49.775 2.565 ;
      RECT 49.515 2.305 49.55 2.565 ;
      RECT 49.83 1.88 49.835 2.34 ;
      RECT 49.92 1.88 49.945 2.16 ;
      RECT 50.195 3.262 50.2 3.525 ;
      RECT 50.16 3.25 50.195 3.525 ;
      RECT 50.1 3.223 50.16 3.525 ;
      RECT 50.095 3.206 50.1 3.379 ;
      RECT 50.09 3.203 50.095 3.366 ;
      RECT 50.07 3.196 50.09 3.353 ;
      RECT 50.035 3.179 50.07 3.335 ;
      RECT 49.995 3.158 50.035 3.315 ;
      RECT 49.99 3.146 49.995 3.303 ;
      RECT 49.95 3.132 49.99 3.289 ;
      RECT 49.93 3.115 49.95 3.271 ;
      RECT 49.92 3.107 49.93 3.263 ;
      RECT 49.905 1.88 49.92 2.178 ;
      RECT 49.89 3.097 49.92 3.25 ;
      RECT 49.875 1.88 49.905 2.223 ;
      RECT 49.88 3.087 49.89 3.237 ;
      RECT 49.85 3.072 49.88 3.224 ;
      RECT 49.835 1.88 49.875 2.29 ;
      RECT 49.835 3.04 49.85 3.21 ;
      RECT 49.83 3.012 49.835 3.204 ;
      RECT 49.825 1.88 49.83 2.345 ;
      RECT 49.815 2.982 49.83 3.198 ;
      RECT 49.82 1.88 49.825 2.358 ;
      RECT 49.81 1.88 49.82 2.378 ;
      RECT 49.775 2.895 49.815 3.183 ;
      RECT 49.775 1.88 49.81 2.418 ;
      RECT 49.77 2.827 49.775 3.171 ;
      RECT 49.755 2.782 49.77 3.166 ;
      RECT 49.75 2.72 49.755 3.161 ;
      RECT 49.725 2.627 49.75 3.154 ;
      RECT 49.72 1.88 49.725 3.146 ;
      RECT 49.705 1.88 49.72 3.133 ;
      RECT 49.685 1.88 49.705 3.09 ;
      RECT 49.675 1.88 49.685 3.04 ;
      RECT 49.67 1.88 49.675 3.013 ;
      RECT 49.665 1.88 49.67 2.991 ;
      RECT 49.66 2.106 49.665 2.974 ;
      RECT 49.655 2.128 49.66 2.952 ;
      RECT 49.65 2.17 49.655 2.935 ;
      RECT 49.62 2.22 49.65 2.879 ;
      RECT 49.615 2.247 49.62 2.821 ;
      RECT 49.6 2.265 49.615 2.785 ;
      RECT 49.595 2.283 49.6 2.749 ;
      RECT 49.589 2.29 49.595 2.73 ;
      RECT 49.585 2.297 49.589 2.713 ;
      RECT 49.58 2.302 49.585 2.682 ;
      RECT 49.57 2.305 49.58 2.657 ;
      RECT 49.56 2.305 49.57 2.623 ;
      RECT 49.555 2.305 49.56 2.6 ;
      RECT 49.55 2.305 49.555 2.58 ;
      RECT 48.465 2.44 48.745 2.72 ;
      RECT 48.465 2.44 48.765 2.615 ;
      RECT 48.555 2.33 48.815 2.59 ;
      RECT 48.52 2.425 48.815 2.59 ;
      RECT 48.645 0.945 48.81 2.59 ;
      RECT 48.545 0.945 48.915 1.315 ;
      RECT 48.17 3.47 48.43 3.73 ;
      RECT 48.19 3.397 48.37 3.73 ;
      RECT 48.19 3.14 48.365 3.73 ;
      RECT 48.19 2.932 48.355 3.73 ;
      RECT 48.195 2.85 48.355 3.73 ;
      RECT 48.195 2.615 48.345 3.73 ;
      RECT 48.195 2.462 48.34 3.73 ;
      RECT 48.2 2.447 48.34 3.73 ;
      RECT 48.25 2.162 48.34 3.73 ;
      RECT 48.205 2.397 48.34 3.73 ;
      RECT 48.235 2.215 48.34 3.73 ;
      RECT 48.22 2.327 48.34 3.73 ;
      RECT 48.225 2.285 48.34 3.73 ;
      RECT 48.22 2.327 48.355 2.39 ;
      RECT 48.255 1.915 48.36 2.335 ;
      RECT 48.255 1.915 48.375 2.318 ;
      RECT 48.255 1.915 48.41 2.28 ;
      RECT 48.25 2.162 48.46 2.213 ;
      RECT 48.255 1.915 48.515 2.175 ;
      RECT 47.515 2.62 47.775 2.88 ;
      RECT 47.515 2.62 47.785 2.838 ;
      RECT 47.515 2.62 47.871 2.809 ;
      RECT 47.515 2.62 47.94 2.761 ;
      RECT 47.515 2.62 47.975 2.73 ;
      RECT 47.745 2.44 48.025 2.72 ;
      RECT 47.58 2.605 48.025 2.72 ;
      RECT 47.67 2.482 47.775 2.88 ;
      RECT 47.6 2.545 48.025 2.72 ;
      RECT 42.05 6.22 42.37 6.545 ;
      RECT 42.08 5.695 42.25 6.545 ;
      RECT 42.08 5.695 42.255 6.045 ;
      RECT 42.08 5.695 43.055 5.87 ;
      RECT 42.88 1.965 43.055 5.87 ;
      RECT 42.825 1.965 43.175 2.315 ;
      RECT 42.85 6.655 43.175 6.98 ;
      RECT 41.735 6.745 43.175 6.915 ;
      RECT 41.735 2.395 41.895 6.915 ;
      RECT 42.05 2.365 42.37 2.685 ;
      RECT 41.735 2.395 42.37 2.565 ;
      RECT 41 5.86 41.34 6.21 ;
      RECT 41.08 2.705 41.255 6.21 ;
      RECT 41.005 2.705 41.345 3.055 ;
      RECT 40.445 2.705 40.785 3.055 ;
      RECT 39.84 2.77 40.785 2.97 ;
      RECT 39.84 2.765 40.055 2.97 ;
      RECT 39.855 2.34 40.055 2.97 ;
      RECT 38.845 2.34 39.125 2.72 ;
      RECT 40.535 2.7 40.705 3.055 ;
      RECT 38.84 2.34 39.125 2.673 ;
      RECT 38.82 2.34 39.125 2.65 ;
      RECT 38.81 2.34 39.125 2.63 ;
      RECT 38.8 2.34 39.125 2.615 ;
      RECT 38.775 2.34 39.125 2.588 ;
      RECT 38.765 2.34 39.125 2.563 ;
      RECT 38.72 2.295 39 2.555 ;
      RECT 38.72 2.34 40.055 2.54 ;
      RECT 38.72 2.335 39.045 2.555 ;
      RECT 38.72 2.327 39.04 2.555 ;
      RECT 38.72 2.317 39.035 2.555 ;
      RECT 38.72 2.305 39.03 2.555 ;
      RECT 37.645 3 37.925 3.28 ;
      RECT 37.645 3 37.96 3.26 ;
      RECT 29.97 6.66 30.32 7.01 ;
      RECT 37.39 6.615 37.74 6.965 ;
      RECT 29.97 6.69 37.74 6.89 ;
      RECT 37.68 2.42 37.73 2.68 ;
      RECT 37.47 2.42 37.475 2.68 ;
      RECT 36.665 1.975 36.695 2.235 ;
      RECT 36.435 1.975 36.51 2.235 ;
      RECT 37.655 2.37 37.68 2.68 ;
      RECT 37.65 2.327 37.655 2.68 ;
      RECT 37.645 2.31 37.65 2.68 ;
      RECT 37.64 2.297 37.645 2.68 ;
      RECT 37.565 2.18 37.64 2.68 ;
      RECT 37.52 1.997 37.565 2.68 ;
      RECT 37.515 1.925 37.52 2.68 ;
      RECT 37.5 1.9 37.515 2.68 ;
      RECT 37.475 1.862 37.5 2.68 ;
      RECT 37.465 1.842 37.475 2.402 ;
      RECT 37.45 1.834 37.465 2.357 ;
      RECT 37.445 1.826 37.45 2.328 ;
      RECT 37.44 1.823 37.445 2.308 ;
      RECT 37.435 1.82 37.44 2.288 ;
      RECT 37.43 1.817 37.435 2.268 ;
      RECT 37.4 1.806 37.43 2.205 ;
      RECT 37.38 1.791 37.4 2.12 ;
      RECT 37.375 1.783 37.38 2.083 ;
      RECT 37.365 1.777 37.375 2.05 ;
      RECT 37.35 1.769 37.365 2.01 ;
      RECT 37.345 1.762 37.35 1.97 ;
      RECT 37.34 1.759 37.345 1.948 ;
      RECT 37.335 1.756 37.34 1.935 ;
      RECT 37.33 1.755 37.335 1.925 ;
      RECT 37.315 1.749 37.33 1.915 ;
      RECT 37.29 1.736 37.315 1.9 ;
      RECT 37.24 1.711 37.29 1.871 ;
      RECT 37.225 1.69 37.24 1.846 ;
      RECT 37.215 1.683 37.225 1.835 ;
      RECT 37.16 1.664 37.215 1.808 ;
      RECT 37.135 1.642 37.16 1.781 ;
      RECT 37.13 1.635 37.135 1.776 ;
      RECT 37.115 1.635 37.13 1.774 ;
      RECT 37.09 1.627 37.115 1.77 ;
      RECT 37.075 1.625 37.09 1.766 ;
      RECT 37.045 1.625 37.075 1.763 ;
      RECT 37.035 1.625 37.045 1.758 ;
      RECT 36.99 1.625 37.035 1.756 ;
      RECT 36.961 1.625 36.99 1.757 ;
      RECT 36.875 1.625 36.961 1.759 ;
      RECT 36.861 1.626 36.875 1.761 ;
      RECT 36.775 1.627 36.861 1.763 ;
      RECT 36.76 1.628 36.775 1.773 ;
      RECT 36.755 1.629 36.76 1.782 ;
      RECT 36.735 1.632 36.755 1.792 ;
      RECT 36.72 1.64 36.735 1.807 ;
      RECT 36.7 1.658 36.72 1.822 ;
      RECT 36.69 1.67 36.7 1.845 ;
      RECT 36.68 1.679 36.69 1.875 ;
      RECT 36.665 1.691 36.68 1.92 ;
      RECT 36.61 1.724 36.665 2.235 ;
      RECT 36.605 1.752 36.61 2.235 ;
      RECT 36.585 1.767 36.605 2.235 ;
      RECT 36.55 1.827 36.585 2.235 ;
      RECT 36.548 1.877 36.55 2.235 ;
      RECT 36.545 1.885 36.548 2.235 ;
      RECT 36.535 1.9 36.545 2.235 ;
      RECT 36.53 1.912 36.535 2.235 ;
      RECT 36.52 1.937 36.53 2.235 ;
      RECT 36.51 1.965 36.52 2.235 ;
      RECT 34.415 3.47 34.465 3.73 ;
      RECT 37.325 3.02 37.385 3.28 ;
      RECT 37.31 3.02 37.325 3.29 ;
      RECT 37.291 3.02 37.31 3.323 ;
      RECT 37.205 3.02 37.291 3.448 ;
      RECT 37.125 3.02 37.205 3.63 ;
      RECT 37.12 3.257 37.125 3.715 ;
      RECT 37.095 3.327 37.12 3.743 ;
      RECT 37.09 3.397 37.095 3.77 ;
      RECT 37.07 3.469 37.09 3.792 ;
      RECT 37.065 3.536 37.07 3.815 ;
      RECT 37.055 3.565 37.065 3.83 ;
      RECT 37.045 3.587 37.055 3.847 ;
      RECT 37.04 3.597 37.045 3.858 ;
      RECT 37.035 3.605 37.04 3.866 ;
      RECT 37.025 3.613 37.035 3.878 ;
      RECT 37.02 3.625 37.025 3.888 ;
      RECT 37.015 3.633 37.02 3.893 ;
      RECT 36.995 3.651 37.015 3.903 ;
      RECT 36.99 3.668 36.995 3.91 ;
      RECT 36.985 3.676 36.99 3.911 ;
      RECT 36.98 3.687 36.985 3.913 ;
      RECT 36.94 3.725 36.98 3.923 ;
      RECT 36.935 3.76 36.94 3.934 ;
      RECT 36.93 3.765 36.935 3.937 ;
      RECT 36.905 3.775 36.93 3.944 ;
      RECT 36.895 3.789 36.905 3.953 ;
      RECT 36.875 3.801 36.895 3.956 ;
      RECT 36.825 3.82 36.875 3.96 ;
      RECT 36.78 3.835 36.825 3.965 ;
      RECT 36.715 3.838 36.78 3.971 ;
      RECT 36.7 3.836 36.715 3.978 ;
      RECT 36.67 3.835 36.7 3.978 ;
      RECT 36.631 3.834 36.67 3.974 ;
      RECT 36.545 3.831 36.631 3.97 ;
      RECT 36.528 3.829 36.545 3.967 ;
      RECT 36.442 3.827 36.528 3.964 ;
      RECT 36.356 3.824 36.442 3.958 ;
      RECT 36.27 3.82 36.356 3.953 ;
      RECT 36.192 3.817 36.27 3.949 ;
      RECT 36.106 3.814 36.192 3.947 ;
      RECT 36.02 3.811 36.106 3.944 ;
      RECT 35.962 3.809 36.02 3.941 ;
      RECT 35.876 3.806 35.962 3.939 ;
      RECT 35.79 3.802 35.876 3.937 ;
      RECT 35.704 3.799 35.79 3.934 ;
      RECT 35.618 3.795 35.704 3.932 ;
      RECT 35.532 3.791 35.618 3.929 ;
      RECT 35.446 3.788 35.532 3.927 ;
      RECT 35.36 3.784 35.446 3.924 ;
      RECT 35.274 3.781 35.36 3.922 ;
      RECT 35.188 3.777 35.274 3.919 ;
      RECT 35.102 3.774 35.188 3.917 ;
      RECT 35.016 3.77 35.102 3.914 ;
      RECT 34.93 3.767 35.016 3.912 ;
      RECT 34.92 3.765 34.93 3.908 ;
      RECT 34.915 3.765 34.92 3.906 ;
      RECT 34.875 3.76 34.915 3.9 ;
      RECT 34.861 3.751 34.875 3.893 ;
      RECT 34.775 3.721 34.861 3.878 ;
      RECT 34.755 3.687 34.775 3.863 ;
      RECT 34.685 3.656 34.755 3.85 ;
      RECT 34.68 3.631 34.685 3.839 ;
      RECT 34.675 3.625 34.68 3.837 ;
      RECT 34.606 3.47 34.675 3.825 ;
      RECT 34.52 3.47 34.606 3.799 ;
      RECT 34.495 3.47 34.52 3.778 ;
      RECT 34.49 3.47 34.495 3.768 ;
      RECT 34.485 3.47 34.49 3.76 ;
      RECT 34.465 3.47 34.485 3.743 ;
      RECT 36.885 2.04 37.145 2.3 ;
      RECT 36.87 2.04 37.145 2.203 ;
      RECT 36.84 2.04 37.145 2.178 ;
      RECT 36.805 1.88 37.085 2.16 ;
      RECT 36.775 3.37 36.835 3.63 ;
      RECT 35.8 2.06 35.855 2.32 ;
      RECT 36.735 3.327 36.775 3.63 ;
      RECT 36.706 3.248 36.735 3.63 ;
      RECT 36.62 3.12 36.706 3.63 ;
      RECT 36.6 3 36.62 3.63 ;
      RECT 36.575 2.951 36.6 3.63 ;
      RECT 36.57 2.916 36.575 3.48 ;
      RECT 36.54 2.876 36.57 3.418 ;
      RECT 36.515 2.813 36.54 3.333 ;
      RECT 36.505 2.775 36.515 3.27 ;
      RECT 36.49 2.75 36.505 3.231 ;
      RECT 36.447 2.708 36.49 3.137 ;
      RECT 36.445 2.681 36.447 3.064 ;
      RECT 36.44 2.676 36.445 3.055 ;
      RECT 36.435 2.669 36.44 3.03 ;
      RECT 36.43 2.663 36.435 3.015 ;
      RECT 36.425 2.657 36.43 3.003 ;
      RECT 36.415 2.648 36.425 2.985 ;
      RECT 36.41 2.639 36.415 2.963 ;
      RECT 36.385 2.62 36.41 2.913 ;
      RECT 36.38 2.601 36.385 2.863 ;
      RECT 36.365 2.587 36.38 2.823 ;
      RECT 36.36 2.573 36.365 2.79 ;
      RECT 36.355 2.566 36.36 2.783 ;
      RECT 36.34 2.553 36.355 2.775 ;
      RECT 36.295 2.515 36.34 2.748 ;
      RECT 36.265 2.468 36.295 2.713 ;
      RECT 36.245 2.437 36.265 2.69 ;
      RECT 36.165 2.37 36.245 2.643 ;
      RECT 36.135 2.3 36.165 2.59 ;
      RECT 36.13 2.277 36.135 2.573 ;
      RECT 36.1 2.255 36.13 2.558 ;
      RECT 36.07 2.214 36.1 2.53 ;
      RECT 36.065 2.189 36.07 2.515 ;
      RECT 36.06 2.183 36.065 2.508 ;
      RECT 36.05 2.06 36.06 2.5 ;
      RECT 36.04 2.06 36.05 2.493 ;
      RECT 36.035 2.06 36.04 2.485 ;
      RECT 36.015 2.06 36.035 2.473 ;
      RECT 35.965 2.06 36.015 2.443 ;
      RECT 35.91 2.06 35.965 2.393 ;
      RECT 35.88 2.06 35.91 2.353 ;
      RECT 35.855 2.06 35.88 2.33 ;
      RECT 35.725 2.785 36.005 3.065 ;
      RECT 35.69 2.7 35.95 2.96 ;
      RECT 35.69 2.782 35.96 2.96 ;
      RECT 33.89 2.155 33.895 2.64 ;
      RECT 33.78 2.34 33.785 2.64 ;
      RECT 33.69 2.38 33.755 2.64 ;
      RECT 35.365 1.88 35.455 2.51 ;
      RECT 35.33 1.93 35.335 2.51 ;
      RECT 35.275 1.955 35.285 2.51 ;
      RECT 35.23 1.955 35.24 2.51 ;
      RECT 35.6 1.88 35.645 2.16 ;
      RECT 34.45 1.61 34.65 1.75 ;
      RECT 35.566 1.88 35.6 2.172 ;
      RECT 35.48 1.88 35.566 2.212 ;
      RECT 35.465 1.88 35.48 2.253 ;
      RECT 35.46 1.88 35.465 2.273 ;
      RECT 35.455 1.88 35.46 2.293 ;
      RECT 35.335 1.922 35.365 2.51 ;
      RECT 35.285 1.942 35.33 2.51 ;
      RECT 35.27 1.957 35.275 2.51 ;
      RECT 35.24 1.957 35.27 2.51 ;
      RECT 35.195 1.942 35.23 2.51 ;
      RECT 35.19 1.93 35.195 2.29 ;
      RECT 35.185 1.927 35.19 2.27 ;
      RECT 35.17 1.917 35.185 2.223 ;
      RECT 35.165 1.91 35.17 2.186 ;
      RECT 35.16 1.907 35.165 2.169 ;
      RECT 35.145 1.897 35.16 2.125 ;
      RECT 35.14 1.888 35.145 2.085 ;
      RECT 35.135 1.884 35.14 2.07 ;
      RECT 35.125 1.878 35.135 2.053 ;
      RECT 35.085 1.859 35.125 2.028 ;
      RECT 35.08 1.841 35.085 2.008 ;
      RECT 35.07 1.835 35.08 2.003 ;
      RECT 35.04 1.819 35.07 1.99 ;
      RECT 35.025 1.801 35.04 1.973 ;
      RECT 35.01 1.789 35.025 1.96 ;
      RECT 35.005 1.781 35.01 1.953 ;
      RECT 34.975 1.767 35.005 1.94 ;
      RECT 34.97 1.752 34.975 1.928 ;
      RECT 34.96 1.746 34.97 1.92 ;
      RECT 34.94 1.734 34.96 1.908 ;
      RECT 34.93 1.722 34.94 1.895 ;
      RECT 34.9 1.706 34.93 1.88 ;
      RECT 34.88 1.686 34.9 1.863 ;
      RECT 34.875 1.676 34.88 1.853 ;
      RECT 34.85 1.664 34.875 1.84 ;
      RECT 34.845 1.652 34.85 1.828 ;
      RECT 34.84 1.647 34.845 1.824 ;
      RECT 34.825 1.64 34.84 1.816 ;
      RECT 34.815 1.627 34.825 1.806 ;
      RECT 34.81 1.625 34.815 1.8 ;
      RECT 34.785 1.618 34.81 1.789 ;
      RECT 34.78 1.611 34.785 1.778 ;
      RECT 34.755 1.61 34.78 1.765 ;
      RECT 34.736 1.61 34.755 1.755 ;
      RECT 34.65 1.61 34.736 1.752 ;
      RECT 34.42 1.61 34.45 1.755 ;
      RECT 34.38 1.617 34.42 1.768 ;
      RECT 34.355 1.627 34.38 1.781 ;
      RECT 34.34 1.636 34.355 1.791 ;
      RECT 34.31 1.641 34.34 1.81 ;
      RECT 34.305 1.647 34.31 1.828 ;
      RECT 34.285 1.657 34.305 1.843 ;
      RECT 34.275 1.67 34.285 1.863 ;
      RECT 34.26 1.682 34.275 1.88 ;
      RECT 34.255 1.692 34.26 1.89 ;
      RECT 34.25 1.697 34.255 1.895 ;
      RECT 34.24 1.705 34.25 1.908 ;
      RECT 34.19 1.737 34.24 1.945 ;
      RECT 34.175 1.772 34.19 1.986 ;
      RECT 34.17 1.782 34.175 2.001 ;
      RECT 34.165 1.787 34.17 2.008 ;
      RECT 34.14 1.803 34.165 2.028 ;
      RECT 34.125 1.824 34.14 2.053 ;
      RECT 34.1 1.845 34.125 2.078 ;
      RECT 34.09 1.864 34.1 2.101 ;
      RECT 34.065 1.882 34.09 2.124 ;
      RECT 34.05 1.902 34.065 2.148 ;
      RECT 34.045 1.912 34.05 2.16 ;
      RECT 34.03 1.924 34.045 2.18 ;
      RECT 34.02 1.939 34.03 2.22 ;
      RECT 34.015 1.947 34.02 2.248 ;
      RECT 34.005 1.957 34.015 2.268 ;
      RECT 34 1.97 34.005 2.293 ;
      RECT 33.995 1.983 34 2.313 ;
      RECT 33.99 1.989 33.995 2.335 ;
      RECT 33.98 1.998 33.99 2.355 ;
      RECT 33.975 2.018 33.98 2.378 ;
      RECT 33.97 2.024 33.975 2.398 ;
      RECT 33.965 2.031 33.97 2.42 ;
      RECT 33.96 2.042 33.965 2.433 ;
      RECT 33.95 2.052 33.96 2.458 ;
      RECT 33.93 2.077 33.95 2.64 ;
      RECT 33.9 2.117 33.93 2.64 ;
      RECT 33.895 2.147 33.9 2.64 ;
      RECT 33.87 2.175 33.89 2.64 ;
      RECT 33.84 2.22 33.87 2.64 ;
      RECT 33.835 2.247 33.84 2.64 ;
      RECT 33.815 2.265 33.835 2.64 ;
      RECT 33.805 2.29 33.815 2.64 ;
      RECT 33.8 2.302 33.805 2.64 ;
      RECT 33.785 2.325 33.8 2.64 ;
      RECT 33.765 2.352 33.78 2.64 ;
      RECT 33.755 2.375 33.765 2.64 ;
      RECT 35.545 3.26 35.625 3.52 ;
      RECT 34.78 2.48 34.85 2.74 ;
      RECT 35.511 3.227 35.545 3.52 ;
      RECT 35.425 3.13 35.511 3.52 ;
      RECT 35.405 3.042 35.425 3.52 ;
      RECT 35.395 3.012 35.405 3.52 ;
      RECT 35.385 2.992 35.395 3.52 ;
      RECT 35.365 2.979 35.385 3.52 ;
      RECT 35.35 2.969 35.365 3.348 ;
      RECT 35.345 2.962 35.35 3.303 ;
      RECT 35.335 2.956 35.345 3.293 ;
      RECT 35.325 2.948 35.335 3.275 ;
      RECT 35.32 2.942 35.325 3.263 ;
      RECT 35.31 2.937 35.32 3.25 ;
      RECT 35.29 2.927 35.31 3.223 ;
      RECT 35.25 2.906 35.29 3.175 ;
      RECT 35.235 2.887 35.25 3.133 ;
      RECT 35.21 2.873 35.235 3.103 ;
      RECT 35.2 2.861 35.21 3.07 ;
      RECT 35.195 2.856 35.2 3.06 ;
      RECT 35.165 2.842 35.195 3.04 ;
      RECT 35.155 2.826 35.165 3.013 ;
      RECT 35.15 2.821 35.155 3.003 ;
      RECT 35.125 2.812 35.15 2.983 ;
      RECT 35.115 2.8 35.125 2.963 ;
      RECT 35.045 2.768 35.115 2.938 ;
      RECT 35.04 2.737 35.045 2.915 ;
      RECT 34.991 2.48 35.04 2.898 ;
      RECT 34.905 2.48 34.991 2.857 ;
      RECT 34.85 2.48 34.905 2.785 ;
      RECT 34.94 3.265 35.1 3.525 ;
      RECT 34.465 1.88 34.515 2.565 ;
      RECT 34.255 2.305 34.29 2.565 ;
      RECT 34.57 1.88 34.575 2.34 ;
      RECT 34.66 1.88 34.685 2.16 ;
      RECT 34.935 3.262 34.94 3.525 ;
      RECT 34.9 3.25 34.935 3.525 ;
      RECT 34.84 3.223 34.9 3.525 ;
      RECT 34.835 3.206 34.84 3.379 ;
      RECT 34.83 3.203 34.835 3.366 ;
      RECT 34.81 3.196 34.83 3.353 ;
      RECT 34.775 3.179 34.81 3.335 ;
      RECT 34.735 3.158 34.775 3.315 ;
      RECT 34.73 3.146 34.735 3.303 ;
      RECT 34.69 3.132 34.73 3.289 ;
      RECT 34.67 3.115 34.69 3.271 ;
      RECT 34.66 3.107 34.67 3.263 ;
      RECT 34.645 1.88 34.66 2.178 ;
      RECT 34.63 3.097 34.66 3.25 ;
      RECT 34.615 1.88 34.645 2.223 ;
      RECT 34.62 3.087 34.63 3.237 ;
      RECT 34.59 3.072 34.62 3.224 ;
      RECT 34.575 1.88 34.615 2.29 ;
      RECT 34.575 3.04 34.59 3.21 ;
      RECT 34.57 3.012 34.575 3.204 ;
      RECT 34.565 1.88 34.57 2.345 ;
      RECT 34.555 2.982 34.57 3.198 ;
      RECT 34.56 1.88 34.565 2.358 ;
      RECT 34.55 1.88 34.56 2.378 ;
      RECT 34.515 2.895 34.555 3.183 ;
      RECT 34.515 1.88 34.55 2.418 ;
      RECT 34.51 2.827 34.515 3.171 ;
      RECT 34.495 2.782 34.51 3.166 ;
      RECT 34.49 2.72 34.495 3.161 ;
      RECT 34.465 2.627 34.49 3.154 ;
      RECT 34.46 1.88 34.465 3.146 ;
      RECT 34.445 1.88 34.46 3.133 ;
      RECT 34.425 1.88 34.445 3.09 ;
      RECT 34.415 1.88 34.425 3.04 ;
      RECT 34.41 1.88 34.415 3.013 ;
      RECT 34.405 1.88 34.41 2.991 ;
      RECT 34.4 2.106 34.405 2.974 ;
      RECT 34.395 2.128 34.4 2.952 ;
      RECT 34.39 2.17 34.395 2.935 ;
      RECT 34.36 2.22 34.39 2.879 ;
      RECT 34.355 2.247 34.36 2.821 ;
      RECT 34.34 2.265 34.355 2.785 ;
      RECT 34.335 2.283 34.34 2.749 ;
      RECT 34.329 2.29 34.335 2.73 ;
      RECT 34.325 2.297 34.329 2.713 ;
      RECT 34.32 2.302 34.325 2.682 ;
      RECT 34.31 2.305 34.32 2.657 ;
      RECT 34.3 2.305 34.31 2.623 ;
      RECT 34.295 2.305 34.3 2.6 ;
      RECT 34.29 2.305 34.295 2.58 ;
      RECT 33.205 2.44 33.485 2.72 ;
      RECT 33.205 2.44 33.505 2.615 ;
      RECT 33.295 2.33 33.555 2.59 ;
      RECT 33.26 2.425 33.555 2.59 ;
      RECT 33.385 0.945 33.55 2.59 ;
      RECT 33.285 0.945 33.655 1.315 ;
      RECT 32.91 3.47 33.17 3.73 ;
      RECT 32.93 3.397 33.11 3.73 ;
      RECT 32.93 3.14 33.105 3.73 ;
      RECT 32.93 2.932 33.095 3.73 ;
      RECT 32.935 2.85 33.095 3.73 ;
      RECT 32.935 2.615 33.085 3.73 ;
      RECT 32.935 2.462 33.08 3.73 ;
      RECT 32.94 2.447 33.08 3.73 ;
      RECT 32.99 2.162 33.08 3.73 ;
      RECT 32.945 2.397 33.08 3.73 ;
      RECT 32.975 2.215 33.08 3.73 ;
      RECT 32.96 2.327 33.08 3.73 ;
      RECT 32.965 2.285 33.08 3.73 ;
      RECT 32.96 2.327 33.095 2.39 ;
      RECT 32.995 1.915 33.1 2.335 ;
      RECT 32.995 1.915 33.115 2.318 ;
      RECT 32.995 1.915 33.15 2.28 ;
      RECT 32.99 2.162 33.2 2.213 ;
      RECT 32.995 1.915 33.255 2.175 ;
      RECT 32.255 2.62 32.515 2.88 ;
      RECT 32.255 2.62 32.525 2.838 ;
      RECT 32.255 2.62 32.611 2.809 ;
      RECT 32.255 2.62 32.68 2.761 ;
      RECT 32.255 2.62 32.715 2.73 ;
      RECT 32.485 2.44 32.765 2.72 ;
      RECT 32.32 2.605 32.765 2.72 ;
      RECT 32.41 2.482 32.515 2.88 ;
      RECT 32.34 2.545 32.765 2.72 ;
      RECT 26.79 6.22 27.11 6.545 ;
      RECT 26.82 5.695 26.99 6.545 ;
      RECT 26.82 5.695 26.995 6.045 ;
      RECT 26.82 5.695 27.795 5.87 ;
      RECT 27.62 1.965 27.795 5.87 ;
      RECT 27.565 1.965 27.915 2.315 ;
      RECT 27.59 6.655 27.915 6.98 ;
      RECT 26.475 6.745 27.915 6.915 ;
      RECT 26.475 2.395 26.635 6.915 ;
      RECT 26.79 2.365 27.11 2.685 ;
      RECT 26.475 2.395 27.11 2.565 ;
      RECT 25.74 5.86 26.08 6.21 ;
      RECT 25.82 2.705 25.995 6.21 ;
      RECT 25.745 2.705 26.085 3.055 ;
      RECT 25.185 2.705 25.525 3.055 ;
      RECT 24.58 2.77 25.525 2.97 ;
      RECT 24.58 2.765 24.795 2.97 ;
      RECT 24.595 2.34 24.795 2.97 ;
      RECT 23.585 2.34 23.865 2.72 ;
      RECT 25.275 2.7 25.445 3.055 ;
      RECT 23.58 2.34 23.865 2.673 ;
      RECT 23.56 2.34 23.865 2.65 ;
      RECT 23.55 2.34 23.865 2.63 ;
      RECT 23.54 2.34 23.865 2.615 ;
      RECT 23.515 2.34 23.865 2.588 ;
      RECT 23.505 2.34 23.865 2.563 ;
      RECT 23.46 2.295 23.74 2.555 ;
      RECT 23.46 2.34 24.795 2.54 ;
      RECT 23.46 2.335 23.785 2.555 ;
      RECT 23.46 2.327 23.78 2.555 ;
      RECT 23.46 2.317 23.775 2.555 ;
      RECT 23.46 2.305 23.77 2.555 ;
      RECT 22.385 3 22.665 3.28 ;
      RECT 22.385 3 22.7 3.26 ;
      RECT 14.71 6.655 15.06 7.005 ;
      RECT 22.13 6.61 22.48 6.96 ;
      RECT 14.71 6.685 22.48 6.885 ;
      RECT 22.42 2.42 22.47 2.68 ;
      RECT 22.21 2.42 22.215 2.68 ;
      RECT 21.405 1.975 21.435 2.235 ;
      RECT 21.175 1.975 21.25 2.235 ;
      RECT 22.395 2.37 22.42 2.68 ;
      RECT 22.39 2.327 22.395 2.68 ;
      RECT 22.385 2.31 22.39 2.68 ;
      RECT 22.38 2.297 22.385 2.68 ;
      RECT 22.305 2.18 22.38 2.68 ;
      RECT 22.26 1.997 22.305 2.68 ;
      RECT 22.255 1.925 22.26 2.68 ;
      RECT 22.24 1.9 22.255 2.68 ;
      RECT 22.215 1.862 22.24 2.68 ;
      RECT 22.205 1.842 22.215 2.402 ;
      RECT 22.19 1.834 22.205 2.357 ;
      RECT 22.185 1.826 22.19 2.328 ;
      RECT 22.18 1.823 22.185 2.308 ;
      RECT 22.175 1.82 22.18 2.288 ;
      RECT 22.17 1.817 22.175 2.268 ;
      RECT 22.14 1.806 22.17 2.205 ;
      RECT 22.12 1.791 22.14 2.12 ;
      RECT 22.115 1.783 22.12 2.083 ;
      RECT 22.105 1.777 22.115 2.05 ;
      RECT 22.09 1.769 22.105 2.01 ;
      RECT 22.085 1.762 22.09 1.97 ;
      RECT 22.08 1.759 22.085 1.948 ;
      RECT 22.075 1.756 22.08 1.935 ;
      RECT 22.07 1.755 22.075 1.925 ;
      RECT 22.055 1.749 22.07 1.915 ;
      RECT 22.03 1.736 22.055 1.9 ;
      RECT 21.98 1.711 22.03 1.871 ;
      RECT 21.965 1.69 21.98 1.846 ;
      RECT 21.955 1.683 21.965 1.835 ;
      RECT 21.9 1.664 21.955 1.808 ;
      RECT 21.875 1.642 21.9 1.781 ;
      RECT 21.87 1.635 21.875 1.776 ;
      RECT 21.855 1.635 21.87 1.774 ;
      RECT 21.83 1.627 21.855 1.77 ;
      RECT 21.815 1.625 21.83 1.766 ;
      RECT 21.785 1.625 21.815 1.763 ;
      RECT 21.775 1.625 21.785 1.758 ;
      RECT 21.73 1.625 21.775 1.756 ;
      RECT 21.701 1.625 21.73 1.757 ;
      RECT 21.615 1.625 21.701 1.759 ;
      RECT 21.601 1.626 21.615 1.761 ;
      RECT 21.515 1.627 21.601 1.763 ;
      RECT 21.5 1.628 21.515 1.773 ;
      RECT 21.495 1.629 21.5 1.782 ;
      RECT 21.475 1.632 21.495 1.792 ;
      RECT 21.46 1.64 21.475 1.807 ;
      RECT 21.44 1.658 21.46 1.822 ;
      RECT 21.43 1.67 21.44 1.845 ;
      RECT 21.42 1.679 21.43 1.875 ;
      RECT 21.405 1.691 21.42 1.92 ;
      RECT 21.35 1.724 21.405 2.235 ;
      RECT 21.345 1.752 21.35 2.235 ;
      RECT 21.325 1.767 21.345 2.235 ;
      RECT 21.29 1.827 21.325 2.235 ;
      RECT 21.288 1.877 21.29 2.235 ;
      RECT 21.285 1.885 21.288 2.235 ;
      RECT 21.275 1.9 21.285 2.235 ;
      RECT 21.27 1.912 21.275 2.235 ;
      RECT 21.26 1.937 21.27 2.235 ;
      RECT 21.25 1.965 21.26 2.235 ;
      RECT 19.155 3.47 19.205 3.73 ;
      RECT 22.065 3.02 22.125 3.28 ;
      RECT 22.05 3.02 22.065 3.29 ;
      RECT 22.031 3.02 22.05 3.323 ;
      RECT 21.945 3.02 22.031 3.448 ;
      RECT 21.865 3.02 21.945 3.63 ;
      RECT 21.86 3.257 21.865 3.715 ;
      RECT 21.835 3.327 21.86 3.743 ;
      RECT 21.83 3.397 21.835 3.77 ;
      RECT 21.81 3.469 21.83 3.792 ;
      RECT 21.805 3.536 21.81 3.815 ;
      RECT 21.795 3.565 21.805 3.83 ;
      RECT 21.785 3.587 21.795 3.847 ;
      RECT 21.78 3.597 21.785 3.858 ;
      RECT 21.775 3.605 21.78 3.866 ;
      RECT 21.765 3.613 21.775 3.878 ;
      RECT 21.76 3.625 21.765 3.888 ;
      RECT 21.755 3.633 21.76 3.893 ;
      RECT 21.735 3.651 21.755 3.903 ;
      RECT 21.73 3.668 21.735 3.91 ;
      RECT 21.725 3.676 21.73 3.911 ;
      RECT 21.72 3.687 21.725 3.913 ;
      RECT 21.68 3.725 21.72 3.923 ;
      RECT 21.675 3.76 21.68 3.934 ;
      RECT 21.67 3.765 21.675 3.937 ;
      RECT 21.645 3.775 21.67 3.944 ;
      RECT 21.635 3.789 21.645 3.953 ;
      RECT 21.615 3.801 21.635 3.956 ;
      RECT 21.565 3.82 21.615 3.96 ;
      RECT 21.52 3.835 21.565 3.965 ;
      RECT 21.455 3.838 21.52 3.971 ;
      RECT 21.44 3.836 21.455 3.978 ;
      RECT 21.41 3.835 21.44 3.978 ;
      RECT 21.371 3.834 21.41 3.974 ;
      RECT 21.285 3.831 21.371 3.97 ;
      RECT 21.268 3.829 21.285 3.967 ;
      RECT 21.182 3.827 21.268 3.964 ;
      RECT 21.096 3.824 21.182 3.958 ;
      RECT 21.01 3.82 21.096 3.953 ;
      RECT 20.932 3.817 21.01 3.949 ;
      RECT 20.846 3.814 20.932 3.947 ;
      RECT 20.76 3.811 20.846 3.944 ;
      RECT 20.702 3.809 20.76 3.941 ;
      RECT 20.616 3.806 20.702 3.939 ;
      RECT 20.53 3.802 20.616 3.937 ;
      RECT 20.444 3.799 20.53 3.934 ;
      RECT 20.358 3.795 20.444 3.932 ;
      RECT 20.272 3.791 20.358 3.929 ;
      RECT 20.186 3.788 20.272 3.927 ;
      RECT 20.1 3.784 20.186 3.924 ;
      RECT 20.014 3.781 20.1 3.922 ;
      RECT 19.928 3.777 20.014 3.919 ;
      RECT 19.842 3.774 19.928 3.917 ;
      RECT 19.756 3.77 19.842 3.914 ;
      RECT 19.67 3.767 19.756 3.912 ;
      RECT 19.66 3.765 19.67 3.908 ;
      RECT 19.655 3.765 19.66 3.906 ;
      RECT 19.615 3.76 19.655 3.9 ;
      RECT 19.601 3.751 19.615 3.893 ;
      RECT 19.515 3.721 19.601 3.878 ;
      RECT 19.495 3.687 19.515 3.863 ;
      RECT 19.425 3.656 19.495 3.85 ;
      RECT 19.42 3.631 19.425 3.839 ;
      RECT 19.415 3.625 19.42 3.837 ;
      RECT 19.346 3.47 19.415 3.825 ;
      RECT 19.26 3.47 19.346 3.799 ;
      RECT 19.235 3.47 19.26 3.778 ;
      RECT 19.23 3.47 19.235 3.768 ;
      RECT 19.225 3.47 19.23 3.76 ;
      RECT 19.205 3.47 19.225 3.743 ;
      RECT 21.625 2.04 21.885 2.3 ;
      RECT 21.61 2.04 21.885 2.203 ;
      RECT 21.58 2.04 21.885 2.178 ;
      RECT 21.545 1.88 21.825 2.16 ;
      RECT 21.515 3.37 21.575 3.63 ;
      RECT 20.54 2.06 20.595 2.32 ;
      RECT 21.475 3.327 21.515 3.63 ;
      RECT 21.446 3.248 21.475 3.63 ;
      RECT 21.36 3.12 21.446 3.63 ;
      RECT 21.34 3 21.36 3.63 ;
      RECT 21.315 2.951 21.34 3.63 ;
      RECT 21.31 2.916 21.315 3.48 ;
      RECT 21.28 2.876 21.31 3.418 ;
      RECT 21.255 2.813 21.28 3.333 ;
      RECT 21.245 2.775 21.255 3.27 ;
      RECT 21.23 2.75 21.245 3.231 ;
      RECT 21.187 2.708 21.23 3.137 ;
      RECT 21.185 2.681 21.187 3.064 ;
      RECT 21.18 2.676 21.185 3.055 ;
      RECT 21.175 2.669 21.18 3.03 ;
      RECT 21.17 2.663 21.175 3.015 ;
      RECT 21.165 2.657 21.17 3.003 ;
      RECT 21.155 2.648 21.165 2.985 ;
      RECT 21.15 2.639 21.155 2.963 ;
      RECT 21.125 2.62 21.15 2.913 ;
      RECT 21.12 2.601 21.125 2.863 ;
      RECT 21.105 2.587 21.12 2.823 ;
      RECT 21.1 2.573 21.105 2.79 ;
      RECT 21.095 2.566 21.1 2.783 ;
      RECT 21.08 2.553 21.095 2.775 ;
      RECT 21.035 2.515 21.08 2.748 ;
      RECT 21.005 2.468 21.035 2.713 ;
      RECT 20.985 2.437 21.005 2.69 ;
      RECT 20.905 2.37 20.985 2.643 ;
      RECT 20.875 2.3 20.905 2.59 ;
      RECT 20.87 2.277 20.875 2.573 ;
      RECT 20.84 2.255 20.87 2.558 ;
      RECT 20.81 2.214 20.84 2.53 ;
      RECT 20.805 2.189 20.81 2.515 ;
      RECT 20.8 2.183 20.805 2.508 ;
      RECT 20.79 2.06 20.8 2.5 ;
      RECT 20.78 2.06 20.79 2.493 ;
      RECT 20.775 2.06 20.78 2.485 ;
      RECT 20.755 2.06 20.775 2.473 ;
      RECT 20.705 2.06 20.755 2.443 ;
      RECT 20.65 2.06 20.705 2.393 ;
      RECT 20.62 2.06 20.65 2.353 ;
      RECT 20.595 2.06 20.62 2.33 ;
      RECT 20.465 2.785 20.745 3.065 ;
      RECT 20.43 2.7 20.69 2.96 ;
      RECT 20.43 2.782 20.7 2.96 ;
      RECT 18.63 2.155 18.635 2.64 ;
      RECT 18.52 2.34 18.525 2.64 ;
      RECT 18.43 2.38 18.495 2.64 ;
      RECT 20.105 1.88 20.195 2.51 ;
      RECT 20.07 1.93 20.075 2.51 ;
      RECT 20.015 1.955 20.025 2.51 ;
      RECT 19.97 1.955 19.98 2.51 ;
      RECT 20.34 1.88 20.385 2.16 ;
      RECT 19.19 1.61 19.39 1.75 ;
      RECT 20.306 1.88 20.34 2.172 ;
      RECT 20.22 1.88 20.306 2.212 ;
      RECT 20.205 1.88 20.22 2.253 ;
      RECT 20.2 1.88 20.205 2.273 ;
      RECT 20.195 1.88 20.2 2.293 ;
      RECT 20.075 1.922 20.105 2.51 ;
      RECT 20.025 1.942 20.07 2.51 ;
      RECT 20.01 1.957 20.015 2.51 ;
      RECT 19.98 1.957 20.01 2.51 ;
      RECT 19.935 1.942 19.97 2.51 ;
      RECT 19.93 1.93 19.935 2.29 ;
      RECT 19.925 1.927 19.93 2.27 ;
      RECT 19.91 1.917 19.925 2.223 ;
      RECT 19.905 1.91 19.91 2.186 ;
      RECT 19.9 1.907 19.905 2.169 ;
      RECT 19.885 1.897 19.9 2.125 ;
      RECT 19.88 1.888 19.885 2.085 ;
      RECT 19.875 1.884 19.88 2.07 ;
      RECT 19.865 1.878 19.875 2.053 ;
      RECT 19.825 1.859 19.865 2.028 ;
      RECT 19.82 1.841 19.825 2.008 ;
      RECT 19.81 1.835 19.82 2.003 ;
      RECT 19.78 1.819 19.81 1.99 ;
      RECT 19.765 1.801 19.78 1.973 ;
      RECT 19.75 1.789 19.765 1.96 ;
      RECT 19.745 1.781 19.75 1.953 ;
      RECT 19.715 1.767 19.745 1.94 ;
      RECT 19.71 1.752 19.715 1.928 ;
      RECT 19.7 1.746 19.71 1.92 ;
      RECT 19.68 1.734 19.7 1.908 ;
      RECT 19.67 1.722 19.68 1.895 ;
      RECT 19.64 1.706 19.67 1.88 ;
      RECT 19.62 1.686 19.64 1.863 ;
      RECT 19.615 1.676 19.62 1.853 ;
      RECT 19.59 1.664 19.615 1.84 ;
      RECT 19.585 1.652 19.59 1.828 ;
      RECT 19.58 1.647 19.585 1.824 ;
      RECT 19.565 1.64 19.58 1.816 ;
      RECT 19.555 1.627 19.565 1.806 ;
      RECT 19.55 1.625 19.555 1.8 ;
      RECT 19.525 1.618 19.55 1.789 ;
      RECT 19.52 1.611 19.525 1.778 ;
      RECT 19.495 1.61 19.52 1.765 ;
      RECT 19.476 1.61 19.495 1.755 ;
      RECT 19.39 1.61 19.476 1.752 ;
      RECT 19.16 1.61 19.19 1.755 ;
      RECT 19.12 1.617 19.16 1.768 ;
      RECT 19.095 1.627 19.12 1.781 ;
      RECT 19.08 1.636 19.095 1.791 ;
      RECT 19.05 1.641 19.08 1.81 ;
      RECT 19.045 1.647 19.05 1.828 ;
      RECT 19.025 1.657 19.045 1.843 ;
      RECT 19.015 1.67 19.025 1.863 ;
      RECT 19 1.682 19.015 1.88 ;
      RECT 18.995 1.692 19 1.89 ;
      RECT 18.99 1.697 18.995 1.895 ;
      RECT 18.98 1.705 18.99 1.908 ;
      RECT 18.93 1.737 18.98 1.945 ;
      RECT 18.915 1.772 18.93 1.986 ;
      RECT 18.91 1.782 18.915 2.001 ;
      RECT 18.905 1.787 18.91 2.008 ;
      RECT 18.88 1.803 18.905 2.028 ;
      RECT 18.865 1.824 18.88 2.053 ;
      RECT 18.84 1.845 18.865 2.078 ;
      RECT 18.83 1.864 18.84 2.101 ;
      RECT 18.805 1.882 18.83 2.124 ;
      RECT 18.79 1.902 18.805 2.148 ;
      RECT 18.785 1.912 18.79 2.16 ;
      RECT 18.77 1.924 18.785 2.18 ;
      RECT 18.76 1.939 18.77 2.22 ;
      RECT 18.755 1.947 18.76 2.248 ;
      RECT 18.745 1.957 18.755 2.268 ;
      RECT 18.74 1.97 18.745 2.293 ;
      RECT 18.735 1.983 18.74 2.313 ;
      RECT 18.73 1.989 18.735 2.335 ;
      RECT 18.72 1.998 18.73 2.355 ;
      RECT 18.715 2.018 18.72 2.378 ;
      RECT 18.71 2.024 18.715 2.398 ;
      RECT 18.705 2.031 18.71 2.42 ;
      RECT 18.7 2.042 18.705 2.433 ;
      RECT 18.69 2.052 18.7 2.458 ;
      RECT 18.67 2.077 18.69 2.64 ;
      RECT 18.64 2.117 18.67 2.64 ;
      RECT 18.635 2.147 18.64 2.64 ;
      RECT 18.61 2.175 18.63 2.64 ;
      RECT 18.58 2.22 18.61 2.64 ;
      RECT 18.575 2.247 18.58 2.64 ;
      RECT 18.555 2.265 18.575 2.64 ;
      RECT 18.545 2.29 18.555 2.64 ;
      RECT 18.54 2.302 18.545 2.64 ;
      RECT 18.525 2.325 18.54 2.64 ;
      RECT 18.505 2.352 18.52 2.64 ;
      RECT 18.495 2.375 18.505 2.64 ;
      RECT 20.285 3.26 20.365 3.52 ;
      RECT 19.52 2.48 19.59 2.74 ;
      RECT 20.251 3.227 20.285 3.52 ;
      RECT 20.165 3.13 20.251 3.52 ;
      RECT 20.145 3.042 20.165 3.52 ;
      RECT 20.135 3.012 20.145 3.52 ;
      RECT 20.125 2.992 20.135 3.52 ;
      RECT 20.105 2.979 20.125 3.52 ;
      RECT 20.09 2.969 20.105 3.348 ;
      RECT 20.085 2.962 20.09 3.303 ;
      RECT 20.075 2.956 20.085 3.293 ;
      RECT 20.065 2.948 20.075 3.275 ;
      RECT 20.06 2.942 20.065 3.263 ;
      RECT 20.05 2.937 20.06 3.25 ;
      RECT 20.03 2.927 20.05 3.223 ;
      RECT 19.99 2.906 20.03 3.175 ;
      RECT 19.975 2.887 19.99 3.133 ;
      RECT 19.95 2.873 19.975 3.103 ;
      RECT 19.94 2.861 19.95 3.07 ;
      RECT 19.935 2.856 19.94 3.06 ;
      RECT 19.905 2.842 19.935 3.04 ;
      RECT 19.895 2.826 19.905 3.013 ;
      RECT 19.89 2.821 19.895 3.003 ;
      RECT 19.865 2.812 19.89 2.983 ;
      RECT 19.855 2.8 19.865 2.963 ;
      RECT 19.785 2.768 19.855 2.938 ;
      RECT 19.78 2.737 19.785 2.915 ;
      RECT 19.731 2.48 19.78 2.898 ;
      RECT 19.645 2.48 19.731 2.857 ;
      RECT 19.59 2.48 19.645 2.785 ;
      RECT 19.68 3.265 19.84 3.525 ;
      RECT 19.205 1.88 19.255 2.565 ;
      RECT 18.995 2.305 19.03 2.565 ;
      RECT 19.31 1.88 19.315 2.34 ;
      RECT 19.4 1.88 19.425 2.16 ;
      RECT 19.675 3.262 19.68 3.525 ;
      RECT 19.64 3.25 19.675 3.525 ;
      RECT 19.58 3.223 19.64 3.525 ;
      RECT 19.575 3.206 19.58 3.379 ;
      RECT 19.57 3.203 19.575 3.366 ;
      RECT 19.55 3.196 19.57 3.353 ;
      RECT 19.515 3.179 19.55 3.335 ;
      RECT 19.475 3.158 19.515 3.315 ;
      RECT 19.47 3.146 19.475 3.303 ;
      RECT 19.43 3.132 19.47 3.289 ;
      RECT 19.41 3.115 19.43 3.271 ;
      RECT 19.4 3.107 19.41 3.263 ;
      RECT 19.385 1.88 19.4 2.178 ;
      RECT 19.37 3.097 19.4 3.25 ;
      RECT 19.355 1.88 19.385 2.223 ;
      RECT 19.36 3.087 19.37 3.237 ;
      RECT 19.33 3.072 19.36 3.224 ;
      RECT 19.315 1.88 19.355 2.29 ;
      RECT 19.315 3.04 19.33 3.21 ;
      RECT 19.31 3.012 19.315 3.204 ;
      RECT 19.305 1.88 19.31 2.345 ;
      RECT 19.295 2.982 19.31 3.198 ;
      RECT 19.3 1.88 19.305 2.358 ;
      RECT 19.29 1.88 19.3 2.378 ;
      RECT 19.255 2.895 19.295 3.183 ;
      RECT 19.255 1.88 19.29 2.418 ;
      RECT 19.25 2.827 19.255 3.171 ;
      RECT 19.235 2.782 19.25 3.166 ;
      RECT 19.23 2.72 19.235 3.161 ;
      RECT 19.205 2.627 19.23 3.154 ;
      RECT 19.2 1.88 19.205 3.146 ;
      RECT 19.185 1.88 19.2 3.133 ;
      RECT 19.165 1.88 19.185 3.09 ;
      RECT 19.155 1.88 19.165 3.04 ;
      RECT 19.15 1.88 19.155 3.013 ;
      RECT 19.145 1.88 19.15 2.991 ;
      RECT 19.14 2.106 19.145 2.974 ;
      RECT 19.135 2.128 19.14 2.952 ;
      RECT 19.13 2.17 19.135 2.935 ;
      RECT 19.1 2.22 19.13 2.879 ;
      RECT 19.095 2.247 19.1 2.821 ;
      RECT 19.08 2.265 19.095 2.785 ;
      RECT 19.075 2.283 19.08 2.749 ;
      RECT 19.069 2.29 19.075 2.73 ;
      RECT 19.065 2.297 19.069 2.713 ;
      RECT 19.06 2.302 19.065 2.682 ;
      RECT 19.05 2.305 19.06 2.657 ;
      RECT 19.04 2.305 19.05 2.623 ;
      RECT 19.035 2.305 19.04 2.6 ;
      RECT 19.03 2.305 19.035 2.58 ;
      RECT 17.945 2.44 18.225 2.72 ;
      RECT 17.945 2.44 18.245 2.615 ;
      RECT 18.035 2.33 18.295 2.59 ;
      RECT 18 2.425 18.295 2.59 ;
      RECT 18.125 0.945 18.29 2.59 ;
      RECT 18.025 0.945 18.395 1.315 ;
      RECT 17.65 3.47 17.91 3.73 ;
      RECT 17.67 3.397 17.85 3.73 ;
      RECT 17.67 3.14 17.845 3.73 ;
      RECT 17.67 2.932 17.835 3.73 ;
      RECT 17.675 2.85 17.835 3.73 ;
      RECT 17.675 2.615 17.825 3.73 ;
      RECT 17.675 2.462 17.82 3.73 ;
      RECT 17.68 2.447 17.82 3.73 ;
      RECT 17.73 2.162 17.82 3.73 ;
      RECT 17.685 2.397 17.82 3.73 ;
      RECT 17.715 2.215 17.82 3.73 ;
      RECT 17.7 2.327 17.82 3.73 ;
      RECT 17.705 2.285 17.82 3.73 ;
      RECT 17.7 2.327 17.835 2.39 ;
      RECT 17.735 1.915 17.84 2.335 ;
      RECT 17.735 1.915 17.855 2.318 ;
      RECT 17.735 1.915 17.89 2.28 ;
      RECT 17.73 2.162 17.94 2.213 ;
      RECT 17.735 1.915 17.995 2.175 ;
      RECT 16.995 2.62 17.255 2.88 ;
      RECT 16.995 2.62 17.265 2.838 ;
      RECT 16.995 2.62 17.351 2.809 ;
      RECT 16.995 2.62 17.42 2.761 ;
      RECT 16.995 2.62 17.455 2.73 ;
      RECT 17.225 2.44 17.505 2.72 ;
      RECT 17.06 2.605 17.505 2.72 ;
      RECT 17.15 2.482 17.255 2.88 ;
      RECT 17.08 2.545 17.505 2.72 ;
      RECT 11.53 6.22 11.85 6.545 ;
      RECT 11.56 5.695 11.73 6.545 ;
      RECT 11.56 5.695 11.735 6.045 ;
      RECT 11.56 5.695 12.535 5.87 ;
      RECT 12.36 1.965 12.535 5.87 ;
      RECT 12.305 1.965 12.655 2.315 ;
      RECT 12.33 6.655 12.655 6.98 ;
      RECT 11.215 6.745 12.655 6.915 ;
      RECT 11.215 2.395 11.375 6.915 ;
      RECT 11.53 2.365 11.85 2.685 ;
      RECT 11.215 2.395 11.85 2.565 ;
      RECT 10.48 5.86 10.82 6.21 ;
      RECT 10.56 2.705 10.735 6.21 ;
      RECT 10.485 2.705 10.825 3.055 ;
      RECT 9.925 2.705 10.265 3.055 ;
      RECT 9.32 2.77 10.265 2.97 ;
      RECT 9.32 2.765 9.535 2.97 ;
      RECT 9.335 2.34 9.535 2.97 ;
      RECT 8.325 2.34 8.605 2.72 ;
      RECT 10.015 2.7 10.185 3.055 ;
      RECT 8.32 2.34 8.605 2.673 ;
      RECT 8.3 2.34 8.605 2.65 ;
      RECT 8.29 2.34 8.605 2.63 ;
      RECT 8.28 2.34 8.605 2.615 ;
      RECT 8.255 2.34 8.605 2.588 ;
      RECT 8.245 2.34 8.605 2.563 ;
      RECT 8.2 2.295 8.48 2.555 ;
      RECT 8.2 2.34 9.535 2.54 ;
      RECT 8.2 2.335 8.525 2.555 ;
      RECT 8.2 2.327 8.52 2.555 ;
      RECT 8.2 2.317 8.515 2.555 ;
      RECT 8.2 2.305 8.51 2.555 ;
      RECT 7.125 3 7.405 3.28 ;
      RECT 7.125 3 7.44 3.26 ;
      RECT -1.255 6.995 -0.965 7.345 ;
      RECT -1.255 7.055 0.075 7.225 ;
      RECT -0.095 6.685 0.075 7.225 ;
      RECT 6.87 6.605 7.22 6.955 ;
      RECT -0.095 6.685 7.22 6.855 ;
      RECT 7.16 2.42 7.21 2.68 ;
      RECT 6.95 2.42 6.955 2.68 ;
      RECT 6.145 1.975 6.175 2.235 ;
      RECT 5.915 1.975 5.99 2.235 ;
      RECT 7.135 2.37 7.16 2.68 ;
      RECT 7.13 2.327 7.135 2.68 ;
      RECT 7.125 2.31 7.13 2.68 ;
      RECT 7.12 2.297 7.125 2.68 ;
      RECT 7.045 2.18 7.12 2.68 ;
      RECT 7 1.997 7.045 2.68 ;
      RECT 6.995 1.925 7 2.68 ;
      RECT 6.98 1.9 6.995 2.68 ;
      RECT 6.955 1.862 6.98 2.68 ;
      RECT 6.945 1.842 6.955 2.402 ;
      RECT 6.93 1.834 6.945 2.357 ;
      RECT 6.925 1.826 6.93 2.328 ;
      RECT 6.92 1.823 6.925 2.308 ;
      RECT 6.915 1.82 6.92 2.288 ;
      RECT 6.91 1.817 6.915 2.268 ;
      RECT 6.88 1.806 6.91 2.205 ;
      RECT 6.86 1.791 6.88 2.12 ;
      RECT 6.855 1.783 6.86 2.083 ;
      RECT 6.845 1.777 6.855 2.05 ;
      RECT 6.83 1.769 6.845 2.01 ;
      RECT 6.825 1.762 6.83 1.97 ;
      RECT 6.82 1.759 6.825 1.948 ;
      RECT 6.815 1.756 6.82 1.935 ;
      RECT 6.81 1.755 6.815 1.925 ;
      RECT 6.795 1.749 6.81 1.915 ;
      RECT 6.77 1.736 6.795 1.9 ;
      RECT 6.72 1.711 6.77 1.871 ;
      RECT 6.705 1.69 6.72 1.846 ;
      RECT 6.695 1.683 6.705 1.835 ;
      RECT 6.64 1.664 6.695 1.808 ;
      RECT 6.615 1.642 6.64 1.781 ;
      RECT 6.61 1.635 6.615 1.776 ;
      RECT 6.595 1.635 6.61 1.774 ;
      RECT 6.57 1.627 6.595 1.77 ;
      RECT 6.555 1.625 6.57 1.766 ;
      RECT 6.525 1.625 6.555 1.763 ;
      RECT 6.515 1.625 6.525 1.758 ;
      RECT 6.47 1.625 6.515 1.756 ;
      RECT 6.441 1.625 6.47 1.757 ;
      RECT 6.355 1.625 6.441 1.759 ;
      RECT 6.341 1.626 6.355 1.761 ;
      RECT 6.255 1.627 6.341 1.763 ;
      RECT 6.24 1.628 6.255 1.773 ;
      RECT 6.235 1.629 6.24 1.782 ;
      RECT 6.215 1.632 6.235 1.792 ;
      RECT 6.2 1.64 6.215 1.807 ;
      RECT 6.18 1.658 6.2 1.822 ;
      RECT 6.17 1.67 6.18 1.845 ;
      RECT 6.16 1.679 6.17 1.875 ;
      RECT 6.145 1.691 6.16 1.92 ;
      RECT 6.09 1.724 6.145 2.235 ;
      RECT 6.085 1.752 6.09 2.235 ;
      RECT 6.065 1.767 6.085 2.235 ;
      RECT 6.03 1.827 6.065 2.235 ;
      RECT 6.028 1.877 6.03 2.235 ;
      RECT 6.025 1.885 6.028 2.235 ;
      RECT 6.015 1.9 6.025 2.235 ;
      RECT 6.01 1.912 6.015 2.235 ;
      RECT 6 1.937 6.01 2.235 ;
      RECT 5.99 1.965 6 2.235 ;
      RECT 3.895 3.47 3.945 3.73 ;
      RECT 6.805 3.02 6.865 3.28 ;
      RECT 6.79 3.02 6.805 3.29 ;
      RECT 6.771 3.02 6.79 3.323 ;
      RECT 6.685 3.02 6.771 3.448 ;
      RECT 6.605 3.02 6.685 3.63 ;
      RECT 6.6 3.257 6.605 3.715 ;
      RECT 6.575 3.327 6.6 3.743 ;
      RECT 6.57 3.397 6.575 3.77 ;
      RECT 6.55 3.469 6.57 3.792 ;
      RECT 6.545 3.536 6.55 3.815 ;
      RECT 6.535 3.565 6.545 3.83 ;
      RECT 6.525 3.587 6.535 3.847 ;
      RECT 6.52 3.597 6.525 3.858 ;
      RECT 6.515 3.605 6.52 3.866 ;
      RECT 6.505 3.613 6.515 3.878 ;
      RECT 6.5 3.625 6.505 3.888 ;
      RECT 6.495 3.633 6.5 3.893 ;
      RECT 6.475 3.651 6.495 3.903 ;
      RECT 6.47 3.668 6.475 3.91 ;
      RECT 6.465 3.676 6.47 3.911 ;
      RECT 6.46 3.687 6.465 3.913 ;
      RECT 6.42 3.725 6.46 3.923 ;
      RECT 6.415 3.76 6.42 3.934 ;
      RECT 6.41 3.765 6.415 3.937 ;
      RECT 6.385 3.775 6.41 3.944 ;
      RECT 6.375 3.789 6.385 3.953 ;
      RECT 6.355 3.801 6.375 3.956 ;
      RECT 6.305 3.82 6.355 3.96 ;
      RECT 6.26 3.835 6.305 3.965 ;
      RECT 6.195 3.838 6.26 3.971 ;
      RECT 6.18 3.836 6.195 3.978 ;
      RECT 6.15 3.835 6.18 3.978 ;
      RECT 6.111 3.834 6.15 3.974 ;
      RECT 6.025 3.831 6.111 3.97 ;
      RECT 6.008 3.829 6.025 3.967 ;
      RECT 5.922 3.827 6.008 3.964 ;
      RECT 5.836 3.824 5.922 3.958 ;
      RECT 5.75 3.82 5.836 3.953 ;
      RECT 5.672 3.817 5.75 3.949 ;
      RECT 5.586 3.814 5.672 3.947 ;
      RECT 5.5 3.811 5.586 3.944 ;
      RECT 5.442 3.809 5.5 3.941 ;
      RECT 5.356 3.806 5.442 3.939 ;
      RECT 5.27 3.802 5.356 3.937 ;
      RECT 5.184 3.799 5.27 3.934 ;
      RECT 5.098 3.795 5.184 3.932 ;
      RECT 5.012 3.791 5.098 3.929 ;
      RECT 4.926 3.788 5.012 3.927 ;
      RECT 4.84 3.784 4.926 3.924 ;
      RECT 4.754 3.781 4.84 3.922 ;
      RECT 4.668 3.777 4.754 3.919 ;
      RECT 4.582 3.774 4.668 3.917 ;
      RECT 4.496 3.77 4.582 3.914 ;
      RECT 4.41 3.767 4.496 3.912 ;
      RECT 4.4 3.765 4.41 3.908 ;
      RECT 4.395 3.765 4.4 3.906 ;
      RECT 4.355 3.76 4.395 3.9 ;
      RECT 4.341 3.751 4.355 3.893 ;
      RECT 4.255 3.721 4.341 3.878 ;
      RECT 4.235 3.687 4.255 3.863 ;
      RECT 4.165 3.656 4.235 3.85 ;
      RECT 4.16 3.631 4.165 3.839 ;
      RECT 4.155 3.625 4.16 3.837 ;
      RECT 4.086 3.47 4.155 3.825 ;
      RECT 4 3.47 4.086 3.799 ;
      RECT 3.975 3.47 4 3.778 ;
      RECT 3.97 3.47 3.975 3.768 ;
      RECT 3.965 3.47 3.97 3.76 ;
      RECT 3.945 3.47 3.965 3.743 ;
      RECT 6.365 2.04 6.625 2.3 ;
      RECT 6.35 2.04 6.625 2.203 ;
      RECT 6.32 2.04 6.625 2.178 ;
      RECT 6.285 1.88 6.565 2.16 ;
      RECT 6.255 3.37 6.315 3.63 ;
      RECT 5.28 2.06 5.335 2.32 ;
      RECT 6.215 3.327 6.255 3.63 ;
      RECT 6.186 3.248 6.215 3.63 ;
      RECT 6.1 3.12 6.186 3.63 ;
      RECT 6.08 3 6.1 3.63 ;
      RECT 6.055 2.951 6.08 3.63 ;
      RECT 6.05 2.916 6.055 3.48 ;
      RECT 6.02 2.876 6.05 3.418 ;
      RECT 5.995 2.813 6.02 3.333 ;
      RECT 5.985 2.775 5.995 3.27 ;
      RECT 5.97 2.75 5.985 3.231 ;
      RECT 5.927 2.708 5.97 3.137 ;
      RECT 5.925 2.681 5.927 3.064 ;
      RECT 5.92 2.676 5.925 3.055 ;
      RECT 5.915 2.669 5.92 3.03 ;
      RECT 5.91 2.663 5.915 3.015 ;
      RECT 5.905 2.657 5.91 3.003 ;
      RECT 5.895 2.648 5.905 2.985 ;
      RECT 5.89 2.639 5.895 2.963 ;
      RECT 5.865 2.62 5.89 2.913 ;
      RECT 5.86 2.601 5.865 2.863 ;
      RECT 5.845 2.587 5.86 2.823 ;
      RECT 5.84 2.573 5.845 2.79 ;
      RECT 5.835 2.566 5.84 2.783 ;
      RECT 5.82 2.553 5.835 2.775 ;
      RECT 5.775 2.515 5.82 2.748 ;
      RECT 5.745 2.468 5.775 2.713 ;
      RECT 5.725 2.437 5.745 2.69 ;
      RECT 5.645 2.37 5.725 2.643 ;
      RECT 5.615 2.3 5.645 2.59 ;
      RECT 5.61 2.277 5.615 2.573 ;
      RECT 5.58 2.255 5.61 2.558 ;
      RECT 5.55 2.214 5.58 2.53 ;
      RECT 5.545 2.189 5.55 2.515 ;
      RECT 5.54 2.183 5.545 2.508 ;
      RECT 5.53 2.06 5.54 2.5 ;
      RECT 5.52 2.06 5.53 2.493 ;
      RECT 5.515 2.06 5.52 2.485 ;
      RECT 5.495 2.06 5.515 2.473 ;
      RECT 5.445 2.06 5.495 2.443 ;
      RECT 5.39 2.06 5.445 2.393 ;
      RECT 5.36 2.06 5.39 2.353 ;
      RECT 5.335 2.06 5.36 2.33 ;
      RECT 5.205 2.785 5.485 3.065 ;
      RECT 5.17 2.7 5.43 2.96 ;
      RECT 5.17 2.782 5.44 2.96 ;
      RECT 3.37 2.155 3.375 2.64 ;
      RECT 3.26 2.34 3.265 2.64 ;
      RECT 3.17 2.38 3.235 2.64 ;
      RECT 4.845 1.88 4.935 2.51 ;
      RECT 4.81 1.93 4.815 2.51 ;
      RECT 4.755 1.955 4.765 2.51 ;
      RECT 4.71 1.955 4.72 2.51 ;
      RECT 5.08 1.88 5.125 2.16 ;
      RECT 3.93 1.61 4.13 1.75 ;
      RECT 5.046 1.88 5.08 2.172 ;
      RECT 4.96 1.88 5.046 2.212 ;
      RECT 4.945 1.88 4.96 2.253 ;
      RECT 4.94 1.88 4.945 2.273 ;
      RECT 4.935 1.88 4.94 2.293 ;
      RECT 4.815 1.922 4.845 2.51 ;
      RECT 4.765 1.942 4.81 2.51 ;
      RECT 4.75 1.957 4.755 2.51 ;
      RECT 4.72 1.957 4.75 2.51 ;
      RECT 4.675 1.942 4.71 2.51 ;
      RECT 4.67 1.93 4.675 2.29 ;
      RECT 4.665 1.927 4.67 2.27 ;
      RECT 4.65 1.917 4.665 2.223 ;
      RECT 4.645 1.91 4.65 2.186 ;
      RECT 4.64 1.907 4.645 2.169 ;
      RECT 4.625 1.897 4.64 2.125 ;
      RECT 4.62 1.888 4.625 2.085 ;
      RECT 4.615 1.884 4.62 2.07 ;
      RECT 4.605 1.878 4.615 2.053 ;
      RECT 4.565 1.859 4.605 2.028 ;
      RECT 4.56 1.841 4.565 2.008 ;
      RECT 4.55 1.835 4.56 2.003 ;
      RECT 4.52 1.819 4.55 1.99 ;
      RECT 4.505 1.801 4.52 1.973 ;
      RECT 4.49 1.789 4.505 1.96 ;
      RECT 4.485 1.781 4.49 1.953 ;
      RECT 4.455 1.767 4.485 1.94 ;
      RECT 4.45 1.752 4.455 1.928 ;
      RECT 4.44 1.746 4.45 1.92 ;
      RECT 4.42 1.734 4.44 1.908 ;
      RECT 4.41 1.722 4.42 1.895 ;
      RECT 4.38 1.706 4.41 1.88 ;
      RECT 4.36 1.686 4.38 1.863 ;
      RECT 4.355 1.676 4.36 1.853 ;
      RECT 4.33 1.664 4.355 1.84 ;
      RECT 4.325 1.652 4.33 1.828 ;
      RECT 4.32 1.647 4.325 1.824 ;
      RECT 4.305 1.64 4.32 1.816 ;
      RECT 4.295 1.627 4.305 1.806 ;
      RECT 4.29 1.625 4.295 1.8 ;
      RECT 4.265 1.618 4.29 1.789 ;
      RECT 4.26 1.611 4.265 1.778 ;
      RECT 4.235 1.61 4.26 1.765 ;
      RECT 4.216 1.61 4.235 1.755 ;
      RECT 4.13 1.61 4.216 1.752 ;
      RECT 3.9 1.61 3.93 1.755 ;
      RECT 3.86 1.617 3.9 1.768 ;
      RECT 3.835 1.627 3.86 1.781 ;
      RECT 3.82 1.636 3.835 1.791 ;
      RECT 3.79 1.641 3.82 1.81 ;
      RECT 3.785 1.647 3.79 1.828 ;
      RECT 3.765 1.657 3.785 1.843 ;
      RECT 3.755 1.67 3.765 1.863 ;
      RECT 3.74 1.682 3.755 1.88 ;
      RECT 3.735 1.692 3.74 1.89 ;
      RECT 3.73 1.697 3.735 1.895 ;
      RECT 3.72 1.705 3.73 1.908 ;
      RECT 3.67 1.737 3.72 1.945 ;
      RECT 3.655 1.772 3.67 1.986 ;
      RECT 3.65 1.782 3.655 2.001 ;
      RECT 3.645 1.787 3.65 2.008 ;
      RECT 3.62 1.803 3.645 2.028 ;
      RECT 3.605 1.824 3.62 2.053 ;
      RECT 3.58 1.845 3.605 2.078 ;
      RECT 3.57 1.864 3.58 2.101 ;
      RECT 3.545 1.882 3.57 2.124 ;
      RECT 3.53 1.902 3.545 2.148 ;
      RECT 3.525 1.912 3.53 2.16 ;
      RECT 3.51 1.924 3.525 2.18 ;
      RECT 3.5 1.939 3.51 2.22 ;
      RECT 3.495 1.947 3.5 2.248 ;
      RECT 3.485 1.957 3.495 2.268 ;
      RECT 3.48 1.97 3.485 2.293 ;
      RECT 3.475 1.983 3.48 2.313 ;
      RECT 3.47 1.989 3.475 2.335 ;
      RECT 3.46 1.998 3.47 2.355 ;
      RECT 3.455 2.018 3.46 2.378 ;
      RECT 3.45 2.024 3.455 2.398 ;
      RECT 3.445 2.031 3.45 2.42 ;
      RECT 3.44 2.042 3.445 2.433 ;
      RECT 3.43 2.052 3.44 2.458 ;
      RECT 3.41 2.077 3.43 2.64 ;
      RECT 3.38 2.117 3.41 2.64 ;
      RECT 3.375 2.147 3.38 2.64 ;
      RECT 3.35 2.175 3.37 2.64 ;
      RECT 3.32 2.22 3.35 2.64 ;
      RECT 3.315 2.247 3.32 2.64 ;
      RECT 3.295 2.265 3.315 2.64 ;
      RECT 3.285 2.29 3.295 2.64 ;
      RECT 3.28 2.302 3.285 2.64 ;
      RECT 3.265 2.325 3.28 2.64 ;
      RECT 3.245 2.352 3.26 2.64 ;
      RECT 3.235 2.375 3.245 2.64 ;
      RECT 5.025 3.26 5.105 3.52 ;
      RECT 4.26 2.48 4.33 2.74 ;
      RECT 4.991 3.227 5.025 3.52 ;
      RECT 4.905 3.13 4.991 3.52 ;
      RECT 4.885 3.042 4.905 3.52 ;
      RECT 4.875 3.012 4.885 3.52 ;
      RECT 4.865 2.992 4.875 3.52 ;
      RECT 4.845 2.979 4.865 3.52 ;
      RECT 4.83 2.969 4.845 3.348 ;
      RECT 4.825 2.962 4.83 3.303 ;
      RECT 4.815 2.956 4.825 3.293 ;
      RECT 4.805 2.948 4.815 3.275 ;
      RECT 4.8 2.942 4.805 3.263 ;
      RECT 4.79 2.937 4.8 3.25 ;
      RECT 4.77 2.927 4.79 3.223 ;
      RECT 4.73 2.906 4.77 3.175 ;
      RECT 4.715 2.887 4.73 3.133 ;
      RECT 4.69 2.873 4.715 3.103 ;
      RECT 4.68 2.861 4.69 3.07 ;
      RECT 4.675 2.856 4.68 3.06 ;
      RECT 4.645 2.842 4.675 3.04 ;
      RECT 4.635 2.826 4.645 3.013 ;
      RECT 4.63 2.821 4.635 3.003 ;
      RECT 4.605 2.812 4.63 2.983 ;
      RECT 4.595 2.8 4.605 2.963 ;
      RECT 4.525 2.768 4.595 2.938 ;
      RECT 4.52 2.737 4.525 2.915 ;
      RECT 4.471 2.48 4.52 2.898 ;
      RECT 4.385 2.48 4.471 2.857 ;
      RECT 4.33 2.48 4.385 2.785 ;
      RECT 4.42 3.265 4.58 3.525 ;
      RECT 3.945 1.88 3.995 2.565 ;
      RECT 3.735 2.305 3.77 2.565 ;
      RECT 4.05 1.88 4.055 2.34 ;
      RECT 4.14 1.88 4.165 2.16 ;
      RECT 4.415 3.262 4.42 3.525 ;
      RECT 4.38 3.25 4.415 3.525 ;
      RECT 4.32 3.223 4.38 3.525 ;
      RECT 4.315 3.206 4.32 3.379 ;
      RECT 4.31 3.203 4.315 3.366 ;
      RECT 4.29 3.196 4.31 3.353 ;
      RECT 4.255 3.179 4.29 3.335 ;
      RECT 4.215 3.158 4.255 3.315 ;
      RECT 4.21 3.146 4.215 3.303 ;
      RECT 4.17 3.132 4.21 3.289 ;
      RECT 4.15 3.115 4.17 3.271 ;
      RECT 4.14 3.107 4.15 3.263 ;
      RECT 4.125 1.88 4.14 2.178 ;
      RECT 4.11 3.097 4.14 3.25 ;
      RECT 4.095 1.88 4.125 2.223 ;
      RECT 4.1 3.087 4.11 3.237 ;
      RECT 4.07 3.072 4.1 3.224 ;
      RECT 4.055 1.88 4.095 2.29 ;
      RECT 4.055 3.04 4.07 3.21 ;
      RECT 4.05 3.012 4.055 3.204 ;
      RECT 4.045 1.88 4.05 2.345 ;
      RECT 4.035 2.982 4.05 3.198 ;
      RECT 4.04 1.88 4.045 2.358 ;
      RECT 4.03 1.88 4.04 2.378 ;
      RECT 3.995 2.895 4.035 3.183 ;
      RECT 3.995 1.88 4.03 2.418 ;
      RECT 3.99 2.827 3.995 3.171 ;
      RECT 3.975 2.782 3.99 3.166 ;
      RECT 3.97 2.72 3.975 3.161 ;
      RECT 3.945 2.627 3.97 3.154 ;
      RECT 3.94 1.88 3.945 3.146 ;
      RECT 3.925 1.88 3.94 3.133 ;
      RECT 3.905 1.88 3.925 3.09 ;
      RECT 3.895 1.88 3.905 3.04 ;
      RECT 3.89 1.88 3.895 3.013 ;
      RECT 3.885 1.88 3.89 2.991 ;
      RECT 3.88 2.106 3.885 2.974 ;
      RECT 3.875 2.128 3.88 2.952 ;
      RECT 3.87 2.17 3.875 2.935 ;
      RECT 3.84 2.22 3.87 2.879 ;
      RECT 3.835 2.247 3.84 2.821 ;
      RECT 3.82 2.265 3.835 2.785 ;
      RECT 3.815 2.283 3.82 2.749 ;
      RECT 3.809 2.29 3.815 2.73 ;
      RECT 3.805 2.297 3.809 2.713 ;
      RECT 3.8 2.302 3.805 2.682 ;
      RECT 3.79 2.305 3.8 2.657 ;
      RECT 3.78 2.305 3.79 2.623 ;
      RECT 3.775 2.305 3.78 2.6 ;
      RECT 3.77 2.305 3.775 2.58 ;
      RECT 2.685 2.44 2.965 2.72 ;
      RECT 2.685 2.44 2.985 2.615 ;
      RECT 2.775 2.33 3.035 2.59 ;
      RECT 2.74 2.425 3.035 2.59 ;
      RECT 2.865 0.945 3.03 2.59 ;
      RECT 2.765 0.945 3.135 1.315 ;
      RECT 2.39 3.47 2.65 3.73 ;
      RECT 2.41 3.397 2.59 3.73 ;
      RECT 2.41 3.14 2.585 3.73 ;
      RECT 2.41 2.932 2.575 3.73 ;
      RECT 2.415 2.85 2.575 3.73 ;
      RECT 2.415 2.615 2.565 3.73 ;
      RECT 2.415 2.462 2.56 3.73 ;
      RECT 2.42 2.447 2.56 3.73 ;
      RECT 2.47 2.162 2.56 3.73 ;
      RECT 2.425 2.397 2.56 3.73 ;
      RECT 2.455 2.215 2.56 3.73 ;
      RECT 2.44 2.327 2.56 3.73 ;
      RECT 2.445 2.285 2.56 3.73 ;
      RECT 2.44 2.327 2.575 2.39 ;
      RECT 2.475 1.915 2.58 2.335 ;
      RECT 2.475 1.915 2.595 2.318 ;
      RECT 2.475 1.915 2.63 2.28 ;
      RECT 2.47 2.162 2.68 2.213 ;
      RECT 2.475 1.915 2.735 2.175 ;
      RECT 1.735 2.62 1.995 2.88 ;
      RECT 1.735 2.62 2.005 2.838 ;
      RECT 1.735 2.62 2.091 2.809 ;
      RECT 1.735 2.62 2.16 2.761 ;
      RECT 1.735 2.62 2.195 2.73 ;
      RECT 1.965 2.44 2.245 2.72 ;
      RECT 1.8 2.605 2.245 2.72 ;
      RECT 1.89 2.482 1.995 2.88 ;
      RECT 1.82 2.545 2.245 2.72 ;
      RECT 67.24 7.055 67.61 7.425 ;
      RECT 51.98 7.055 52.35 7.425 ;
      RECT 36.72 7.055 37.09 7.425 ;
      RECT 21.46 7.055 21.83 7.425 ;
      RECT 6.2 7.055 6.57 7.425 ;
    LAYER via1 ;
      RECT 75.83 7.375 75.98 7.525 ;
      RECT 73.46 6.74 73.61 6.89 ;
      RECT 73.445 2.065 73.595 2.215 ;
      RECT 72.655 2.45 72.805 2.6 ;
      RECT 72.655 6.325 72.805 6.475 ;
      RECT 71.625 2.805 71.775 2.955 ;
      RECT 71.62 5.96 71.77 6.11 ;
      RECT 71.065 2.805 71.215 2.955 ;
      RECT 69.295 2.35 69.445 2.5 ;
      RECT 68.275 3.055 68.425 3.205 ;
      RECT 68.045 2.475 68.195 2.625 ;
      RECT 68.01 6.71 68.16 6.86 ;
      RECT 67.7 3.075 67.85 3.225 ;
      RECT 67.46 2.095 67.61 2.245 ;
      RECT 67.35 7.165 67.5 7.315 ;
      RECT 67.15 3.425 67.3 3.575 ;
      RECT 67.01 2.03 67.16 2.18 ;
      RECT 66.375 2.115 66.525 2.265 ;
      RECT 66.265 2.755 66.415 2.905 ;
      RECT 65.94 3.315 66.09 3.465 ;
      RECT 65.77 2.305 65.92 2.455 ;
      RECT 65.415 3.32 65.565 3.47 ;
      RECT 65.355 2.535 65.505 2.685 ;
      RECT 64.99 3.525 65.14 3.675 ;
      RECT 64.83 2.36 64.98 2.51 ;
      RECT 64.265 2.435 64.415 2.585 ;
      RECT 63.915 1.055 64.065 1.205 ;
      RECT 63.87 2.385 64.02 2.535 ;
      RECT 63.57 1.97 63.72 2.12 ;
      RECT 63.485 3.525 63.635 3.675 ;
      RECT 62.83 2.675 62.98 2.825 ;
      RECT 60.545 6.755 60.695 6.905 ;
      RECT 58.2 6.74 58.35 6.89 ;
      RECT 58.185 2.065 58.335 2.215 ;
      RECT 57.395 2.45 57.545 2.6 ;
      RECT 57.395 6.325 57.545 6.475 ;
      RECT 56.365 2.805 56.515 2.955 ;
      RECT 56.36 5.96 56.51 6.11 ;
      RECT 55.805 2.805 55.955 2.955 ;
      RECT 54.035 2.35 54.185 2.5 ;
      RECT 53.015 3.055 53.165 3.205 ;
      RECT 52.785 2.475 52.935 2.625 ;
      RECT 52.75 6.71 52.9 6.86 ;
      RECT 52.44 3.075 52.59 3.225 ;
      RECT 52.2 2.095 52.35 2.245 ;
      RECT 52.09 7.165 52.24 7.315 ;
      RECT 51.89 3.425 52.04 3.575 ;
      RECT 51.75 2.03 51.9 2.18 ;
      RECT 51.115 2.115 51.265 2.265 ;
      RECT 51.005 2.755 51.155 2.905 ;
      RECT 50.68 3.315 50.83 3.465 ;
      RECT 50.51 2.305 50.66 2.455 ;
      RECT 50.155 3.32 50.305 3.47 ;
      RECT 50.095 2.535 50.245 2.685 ;
      RECT 49.73 3.525 49.88 3.675 ;
      RECT 49.57 2.36 49.72 2.51 ;
      RECT 49.005 2.435 49.155 2.585 ;
      RECT 48.655 1.055 48.805 1.205 ;
      RECT 48.61 2.385 48.76 2.535 ;
      RECT 48.31 1.97 48.46 2.12 ;
      RECT 48.225 3.525 48.375 3.675 ;
      RECT 47.57 2.675 47.72 2.825 ;
      RECT 45.285 6.755 45.435 6.905 ;
      RECT 42.94 6.74 43.09 6.89 ;
      RECT 42.925 2.065 43.075 2.215 ;
      RECT 42.135 2.45 42.285 2.6 ;
      RECT 42.135 6.325 42.285 6.475 ;
      RECT 41.105 2.805 41.255 2.955 ;
      RECT 41.1 5.96 41.25 6.11 ;
      RECT 40.545 2.805 40.695 2.955 ;
      RECT 38.775 2.35 38.925 2.5 ;
      RECT 37.755 3.055 37.905 3.205 ;
      RECT 37.525 2.475 37.675 2.625 ;
      RECT 37.49 6.715 37.64 6.865 ;
      RECT 37.18 3.075 37.33 3.225 ;
      RECT 36.94 2.095 37.09 2.245 ;
      RECT 36.83 7.165 36.98 7.315 ;
      RECT 36.63 3.425 36.78 3.575 ;
      RECT 36.49 2.03 36.64 2.18 ;
      RECT 35.855 2.115 36.005 2.265 ;
      RECT 35.745 2.755 35.895 2.905 ;
      RECT 35.42 3.315 35.57 3.465 ;
      RECT 35.25 2.305 35.4 2.455 ;
      RECT 34.895 3.32 35.045 3.47 ;
      RECT 34.835 2.535 34.985 2.685 ;
      RECT 34.47 3.525 34.62 3.675 ;
      RECT 34.31 2.36 34.46 2.51 ;
      RECT 33.745 2.435 33.895 2.585 ;
      RECT 33.395 1.055 33.545 1.205 ;
      RECT 33.35 2.385 33.5 2.535 ;
      RECT 33.05 1.97 33.2 2.12 ;
      RECT 32.965 3.525 33.115 3.675 ;
      RECT 32.31 2.675 32.46 2.825 ;
      RECT 30.07 6.76 30.22 6.91 ;
      RECT 27.68 6.74 27.83 6.89 ;
      RECT 27.665 2.065 27.815 2.215 ;
      RECT 26.875 2.45 27.025 2.6 ;
      RECT 26.875 6.325 27.025 6.475 ;
      RECT 25.845 2.805 25.995 2.955 ;
      RECT 25.84 5.96 25.99 6.11 ;
      RECT 25.285 2.805 25.435 2.955 ;
      RECT 23.515 2.35 23.665 2.5 ;
      RECT 22.495 3.055 22.645 3.205 ;
      RECT 22.265 2.475 22.415 2.625 ;
      RECT 22.23 6.71 22.38 6.86 ;
      RECT 21.92 3.075 22.07 3.225 ;
      RECT 21.68 2.095 21.83 2.245 ;
      RECT 21.57 7.165 21.72 7.315 ;
      RECT 21.37 3.425 21.52 3.575 ;
      RECT 21.23 2.03 21.38 2.18 ;
      RECT 20.595 2.115 20.745 2.265 ;
      RECT 20.485 2.755 20.635 2.905 ;
      RECT 20.16 3.315 20.31 3.465 ;
      RECT 19.99 2.305 20.14 2.455 ;
      RECT 19.635 3.32 19.785 3.47 ;
      RECT 19.575 2.535 19.725 2.685 ;
      RECT 19.21 3.525 19.36 3.675 ;
      RECT 19.05 2.36 19.2 2.51 ;
      RECT 18.485 2.435 18.635 2.585 ;
      RECT 18.135 1.055 18.285 1.205 ;
      RECT 18.09 2.385 18.24 2.535 ;
      RECT 17.79 1.97 17.94 2.12 ;
      RECT 17.705 3.525 17.855 3.675 ;
      RECT 17.05 2.675 17.2 2.825 ;
      RECT 14.81 6.755 14.96 6.905 ;
      RECT 12.42 6.74 12.57 6.89 ;
      RECT 12.405 2.065 12.555 2.215 ;
      RECT 11.615 2.45 11.765 2.6 ;
      RECT 11.615 6.325 11.765 6.475 ;
      RECT 10.585 2.805 10.735 2.955 ;
      RECT 10.58 5.96 10.73 6.11 ;
      RECT 10.025 2.805 10.175 2.955 ;
      RECT 8.255 2.35 8.405 2.5 ;
      RECT 7.235 3.055 7.385 3.205 ;
      RECT 7.005 2.475 7.155 2.625 ;
      RECT 6.97 6.705 7.12 6.855 ;
      RECT 6.66 3.075 6.81 3.225 ;
      RECT 6.42 2.095 6.57 2.245 ;
      RECT 6.31 7.165 6.46 7.315 ;
      RECT 6.11 3.425 6.26 3.575 ;
      RECT 5.97 2.03 6.12 2.18 ;
      RECT 5.335 2.115 5.485 2.265 ;
      RECT 5.225 2.755 5.375 2.905 ;
      RECT 4.9 3.315 5.05 3.465 ;
      RECT 4.73 2.305 4.88 2.455 ;
      RECT 4.375 3.32 4.525 3.47 ;
      RECT 4.315 2.535 4.465 2.685 ;
      RECT 3.95 3.525 4.1 3.675 ;
      RECT 3.79 2.36 3.94 2.51 ;
      RECT 3.225 2.435 3.375 2.585 ;
      RECT 2.875 1.055 3.025 1.205 ;
      RECT 2.83 2.385 2.98 2.535 ;
      RECT 2.53 1.97 2.68 2.12 ;
      RECT 2.445 3.525 2.595 3.675 ;
      RECT 1.79 2.675 1.94 2.825 ;
      RECT -1.185 7.095 -1.035 7.245 ;
      RECT -1.56 6.355 -1.41 6.505 ;
    LAYER met1 ;
      RECT 61.79 0 70.53 1.74 ;
      RECT 46.53 0 55.27 1.74 ;
      RECT 31.27 0 40.01 1.74 ;
      RECT 16.01 0 24.75 1.74 ;
      RECT 0.75 0 9.49 1.74 ;
      RECT -2.75 0 76.3 0.305 ;
      RECT -2.75 4.14 76.3 4.745 ;
      RECT 61.79 4.135 76.3 4.745 ;
      RECT 46.53 4.135 61.04 4.745 ;
      RECT 31.27 4.135 45.78 4.745 ;
      RECT 16.01 4.135 30.52 4.745 ;
      RECT 0.75 4.135 15.26 4.745 ;
      RECT 61.79 3.98 70.53 4.745 ;
      RECT 46.53 3.98 55.27 4.745 ;
      RECT 31.27 3.98 40.01 4.745 ;
      RECT 16.01 3.98 24.75 4.745 ;
      RECT 0.75 3.98 9.49 4.745 ;
      RECT -2.75 8.575 76.3 8.88 ;
      RECT 66.735 6.315 66.905 8.88 ;
      RECT 51.475 6.315 51.645 8.88 ;
      RECT 36.215 6.315 36.385 8.88 ;
      RECT 20.955 6.315 21.125 8.88 ;
      RECT 5.695 6.315 5.865 8.88 ;
      RECT 66.905 6.285 67.195 6.515 ;
      RECT 51.645 6.285 51.935 6.515 ;
      RECT 36.385 6.285 36.675 6.515 ;
      RECT 21.125 6.285 21.415 6.515 ;
      RECT 5.865 6.285 6.155 6.515 ;
      RECT 75.7 7.765 75.99 7.995 ;
      RECT 75.76 6.285 75.93 7.995 ;
      RECT 75.73 7.275 76.08 7.625 ;
      RECT 75.7 6.285 75.99 6.515 ;
      RECT 75.7 2.365 75.99 2.595 ;
      RECT 75.76 0.885 75.93 2.595 ;
      RECT 75.7 0.885 75.99 1.115 ;
      RECT 75.29 2.735 75.62 2.965 ;
      RECT 75.29 2.765 75.79 2.935 ;
      RECT 75.29 2.395 75.48 2.965 ;
      RECT 74.71 2.365 75 2.595 ;
      RECT 74.71 2.395 75.48 2.565 ;
      RECT 74.77 0.885 74.94 2.595 ;
      RECT 74.71 0.885 75 1.115 ;
      RECT 74.71 7.765 75 7.995 ;
      RECT 74.77 6.285 74.94 7.995 ;
      RECT 74.71 6.285 75 6.515 ;
      RECT 74.71 6.325 75.56 6.485 ;
      RECT 75.39 5.915 75.56 6.485 ;
      RECT 74.71 6.32 75.1 6.485 ;
      RECT 75.33 5.915 75.62 6.145 ;
      RECT 75.33 5.945 75.79 6.115 ;
      RECT 74.34 2.735 74.63 2.965 ;
      RECT 74.34 2.765 74.8 2.935 ;
      RECT 74.4 1.655 74.565 2.965 ;
      RECT 72.915 1.625 73.205 1.855 ;
      RECT 72.915 1.655 74.565 1.825 ;
      RECT 72.975 0.885 73.145 1.855 ;
      RECT 72.915 0.885 73.205 1.115 ;
      RECT 72.915 7.765 73.205 7.995 ;
      RECT 72.975 7.025 73.145 7.995 ;
      RECT 72.975 7.12 74.565 7.29 ;
      RECT 74.395 5.915 74.565 7.29 ;
      RECT 72.915 7.025 73.205 7.255 ;
      RECT 74.34 5.915 74.63 6.145 ;
      RECT 74.34 5.945 74.8 6.115 ;
      RECT 70.965 2.705 71.305 3.055 ;
      RECT 71.055 2.025 71.225 3.055 ;
      RECT 73.345 1.965 73.695 2.315 ;
      RECT 71.055 2.025 73.695 2.195 ;
      RECT 73.37 6.655 73.695 6.98 ;
      RECT 67.91 6.61 68.26 6.96 ;
      RECT 73.345 6.655 73.695 6.885 ;
      RECT 67.71 6.655 68.26 6.885 ;
      RECT 67.54 6.685 73.695 6.855 ;
      RECT 72.57 2.365 72.89 2.685 ;
      RECT 72.54 2.365 72.89 2.595 ;
      RECT 72.37 2.395 72.89 2.565 ;
      RECT 72.57 6.255 72.89 6.545 ;
      RECT 72.54 6.285 72.89 6.515 ;
      RECT 72.37 6.315 72.89 6.485 ;
      RECT 71.525 2.705 71.865 3.055 ;
      RECT 71.525 2.765 72.005 2.935 ;
      RECT 71.52 5.86 71.86 6.21 ;
      RECT 65.91 5.915 66.2 6.145 ;
      RECT 65.91 5.945 72.005 6.115 ;
      RECT 68.26 2.985 68.41 3.26 ;
      RECT 68.8 2.065 68.805 2.285 ;
      RECT 69.95 2.265 69.965 2.463 ;
      RECT 69.915 2.257 69.95 2.47 ;
      RECT 69.885 2.25 69.915 2.47 ;
      RECT 69.83 2.215 69.885 2.47 ;
      RECT 69.765 2.152 69.83 2.47 ;
      RECT 69.76 2.117 69.765 2.468 ;
      RECT 69.755 2.112 69.76 2.46 ;
      RECT 69.75 2.107 69.755 2.446 ;
      RECT 69.745 2.104 69.75 2.439 ;
      RECT 69.7 2.094 69.745 2.39 ;
      RECT 69.68 2.081 69.7 2.325 ;
      RECT 69.675 2.076 69.68 2.298 ;
      RECT 69.67 2.075 69.675 2.291 ;
      RECT 69.665 2.074 69.67 2.284 ;
      RECT 69.58 2.059 69.665 2.23 ;
      RECT 69.55 2.04 69.58 2.18 ;
      RECT 69.47 2.023 69.55 2.165 ;
      RECT 69.435 2.01 69.47 2.15 ;
      RECT 69.427 2.01 69.435 2.145 ;
      RECT 69.341 2.011 69.427 2.145 ;
      RECT 69.255 2.013 69.341 2.145 ;
      RECT 69.23 2.014 69.255 2.149 ;
      RECT 69.155 2.02 69.23 2.164 ;
      RECT 69.072 2.032 69.155 2.188 ;
      RECT 68.986 2.045 69.072 2.214 ;
      RECT 68.9 2.058 68.986 2.24 ;
      RECT 68.865 2.067 68.9 2.259 ;
      RECT 68.815 2.067 68.865 2.272 ;
      RECT 68.805 2.065 68.815 2.283 ;
      RECT 68.79 2.062 68.8 2.285 ;
      RECT 68.775 2.054 68.79 2.293 ;
      RECT 68.76 2.046 68.775 2.313 ;
      RECT 68.755 2.041 68.76 2.37 ;
      RECT 68.74 2.036 68.755 2.443 ;
      RECT 68.735 2.031 68.74 2.485 ;
      RECT 68.73 2.029 68.735 2.513 ;
      RECT 68.725 2.027 68.73 2.535 ;
      RECT 68.715 2.023 68.725 2.578 ;
      RECT 68.71 2.02 68.715 2.603 ;
      RECT 68.705 2.018 68.71 2.623 ;
      RECT 68.7 2.016 68.705 2.647 ;
      RECT 68.695 2.012 68.7 2.67 ;
      RECT 68.69 2.008 68.695 2.693 ;
      RECT 68.655 1.998 68.69 2.8 ;
      RECT 68.65 1.988 68.655 2.898 ;
      RECT 68.645 1.986 68.65 2.925 ;
      RECT 68.64 1.985 68.645 2.945 ;
      RECT 68.635 1.977 68.64 2.965 ;
      RECT 68.63 1.972 68.635 3 ;
      RECT 68.625 1.97 68.63 3.018 ;
      RECT 68.62 1.97 68.625 3.043 ;
      RECT 68.615 1.97 68.62 3.065 ;
      RECT 68.58 1.97 68.615 3.108 ;
      RECT 68.555 1.97 68.58 3.137 ;
      RECT 68.545 1.97 68.555 2.323 ;
      RECT 68.548 2.38 68.555 3.147 ;
      RECT 68.545 2.437 68.548 3.15 ;
      RECT 68.54 1.97 68.545 2.295 ;
      RECT 68.54 2.487 68.545 3.153 ;
      RECT 68.53 1.97 68.54 2.285 ;
      RECT 68.535 2.54 68.54 3.156 ;
      RECT 68.53 2.625 68.535 3.16 ;
      RECT 68.52 1.97 68.53 2.273 ;
      RECT 68.525 2.672 68.53 3.164 ;
      RECT 68.52 2.747 68.525 3.168 ;
      RECT 68.485 1.97 68.52 2.248 ;
      RECT 68.51 2.83 68.52 3.173 ;
      RECT 68.5 2.897 68.51 3.18 ;
      RECT 68.495 2.925 68.5 3.185 ;
      RECT 68.485 2.938 68.495 3.191 ;
      RECT 68.44 1.97 68.485 2.205 ;
      RECT 68.48 2.943 68.485 3.198 ;
      RECT 68.44 2.96 68.48 3.26 ;
      RECT 68.435 1.972 68.44 2.178 ;
      RECT 68.41 2.98 68.44 3.26 ;
      RECT 68.43 1.977 68.435 2.15 ;
      RECT 68.22 2.989 68.26 3.26 ;
      RECT 68.195 2.997 68.22 3.23 ;
      RECT 68.15 3.005 68.195 3.23 ;
      RECT 68.135 3.01 68.15 3.225 ;
      RECT 68.125 3.01 68.135 3.219 ;
      RECT 68.115 3.017 68.125 3.216 ;
      RECT 68.11 3.055 68.115 3.205 ;
      RECT 68.105 3.117 68.11 3.183 ;
      RECT 69.375 2.992 69.56 3.215 ;
      RECT 69.375 3.007 69.565 3.211 ;
      RECT 69.365 2.28 69.45 3.21 ;
      RECT 69.365 3.007 69.57 3.204 ;
      RECT 69.36 3.015 69.57 3.203 ;
      RECT 69.565 2.735 69.885 3.055 ;
      RECT 69.36 2.907 69.53 2.998 ;
      RECT 69.355 2.907 69.53 2.98 ;
      RECT 69.345 2.715 69.48 2.955 ;
      RECT 69.34 2.715 69.48 2.9 ;
      RECT 69.3 2.295 69.47 2.8 ;
      RECT 69.285 2.295 69.47 2.67 ;
      RECT 69.28 2.295 69.47 2.623 ;
      RECT 69.275 2.295 69.47 2.603 ;
      RECT 69.27 2.295 69.47 2.578 ;
      RECT 69.24 2.295 69.5 2.555 ;
      RECT 69.25 2.292 69.46 2.555 ;
      RECT 69.375 2.287 69.46 3.215 ;
      RECT 69.26 2.28 69.45 2.555 ;
      RECT 69.255 2.285 69.45 2.555 ;
      RECT 68.085 2.497 68.27 2.71 ;
      RECT 68.085 2.505 68.28 2.703 ;
      RECT 68.065 2.505 68.28 2.7 ;
      RECT 68.06 2.505 68.28 2.685 ;
      RECT 67.99 2.42 68.25 2.68 ;
      RECT 67.99 2.565 68.285 2.593 ;
      RECT 67.645 3.02 67.905 3.28 ;
      RECT 67.67 2.965 67.865 3.28 ;
      RECT 67.665 2.714 67.845 3.008 ;
      RECT 67.665 2.72 67.855 3.008 ;
      RECT 67.645 2.722 67.855 2.953 ;
      RECT 67.64 2.732 67.855 2.82 ;
      RECT 67.67 2.712 67.845 3.28 ;
      RECT 67.756 2.71 67.845 3.28 ;
      RECT 67.615 1.93 67.65 2.3 ;
      RECT 67.405 2.04 67.41 2.3 ;
      RECT 67.65 1.937 67.665 2.3 ;
      RECT 67.54 1.93 67.615 2.378 ;
      RECT 67.53 1.93 67.54 2.463 ;
      RECT 67.505 1.93 67.53 2.498 ;
      RECT 67.465 1.93 67.505 2.566 ;
      RECT 67.455 1.937 67.465 2.618 ;
      RECT 67.425 2.04 67.455 2.659 ;
      RECT 67.42 2.04 67.425 2.698 ;
      RECT 67.41 2.04 67.42 2.718 ;
      RECT 67.405 2.335 67.41 2.755 ;
      RECT 67.4 2.352 67.405 2.775 ;
      RECT 67.385 2.415 67.4 2.815 ;
      RECT 67.38 2.458 67.385 2.85 ;
      RECT 67.375 2.466 67.38 2.863 ;
      RECT 67.365 2.48 67.375 2.885 ;
      RECT 67.34 2.515 67.365 2.95 ;
      RECT 67.33 2.55 67.34 3.013 ;
      RECT 67.31 2.58 67.33 3.074 ;
      RECT 67.295 2.616 67.31 3.141 ;
      RECT 67.285 2.644 67.295 3.18 ;
      RECT 67.275 2.666 67.285 3.2 ;
      RECT 67.27 2.676 67.275 3.211 ;
      RECT 67.265 2.685 67.27 3.214 ;
      RECT 67.255 2.703 67.265 3.218 ;
      RECT 67.245 2.721 67.255 3.219 ;
      RECT 67.22 2.76 67.245 3.216 ;
      RECT 67.2 2.802 67.22 3.213 ;
      RECT 67.185 2.84 67.2 3.212 ;
      RECT 67.15 2.875 67.185 3.209 ;
      RECT 67.145 2.897 67.15 3.207 ;
      RECT 67.08 2.937 67.145 3.204 ;
      RECT 67.075 2.977 67.08 3.2 ;
      RECT 67.06 2.987 67.075 3.191 ;
      RECT 67.05 3.107 67.06 3.176 ;
      RECT 67.53 3.52 67.54 3.78 ;
      RECT 67.53 3.523 67.55 3.779 ;
      RECT 67.52 3.513 67.53 3.778 ;
      RECT 67.51 3.528 67.59 3.774 ;
      RECT 67.495 3.507 67.51 3.772 ;
      RECT 67.47 3.532 67.595 3.768 ;
      RECT 67.455 3.492 67.47 3.763 ;
      RECT 67.455 3.534 67.605 3.762 ;
      RECT 67.455 3.542 67.62 3.755 ;
      RECT 67.395 3.479 67.455 3.745 ;
      RECT 67.385 3.466 67.395 3.727 ;
      RECT 67.36 3.456 67.385 3.717 ;
      RECT 67.355 3.446 67.36 3.709 ;
      RECT 67.29 3.542 67.62 3.691 ;
      RECT 67.205 3.542 67.62 3.653 ;
      RECT 67.095 3.37 67.355 3.63 ;
      RECT 67.47 3.5 67.495 3.768 ;
      RECT 67.51 3.51 67.52 3.774 ;
      RECT 67.095 3.518 67.535 3.63 ;
      RECT 67.28 7.765 67.57 7.995 ;
      RECT 67.34 7.025 67.51 7.995 ;
      RECT 67.24 7.055 67.61 7.425 ;
      RECT 67.28 7.025 67.57 7.425 ;
      RECT 66.31 3.275 66.34 3.575 ;
      RECT 66.085 3.26 66.09 3.535 ;
      RECT 65.885 3.26 66.04 3.52 ;
      RECT 67.185 1.975 67.215 2.235 ;
      RECT 67.175 1.975 67.185 2.343 ;
      RECT 67.155 1.975 67.175 2.353 ;
      RECT 67.14 1.975 67.155 2.365 ;
      RECT 67.085 1.975 67.14 2.415 ;
      RECT 67.07 1.975 67.085 2.463 ;
      RECT 67.04 1.975 67.07 2.498 ;
      RECT 66.985 1.975 67.04 2.56 ;
      RECT 66.965 1.975 66.985 2.628 ;
      RECT 66.96 1.975 66.965 2.658 ;
      RECT 66.955 1.975 66.96 2.67 ;
      RECT 66.95 2.092 66.955 2.688 ;
      RECT 66.93 2.11 66.95 2.713 ;
      RECT 66.91 2.137 66.93 2.763 ;
      RECT 66.905 2.157 66.91 2.794 ;
      RECT 66.9 2.165 66.905 2.811 ;
      RECT 66.885 2.191 66.9 2.84 ;
      RECT 66.87 2.233 66.885 2.875 ;
      RECT 66.865 2.262 66.87 2.898 ;
      RECT 66.86 2.277 66.865 2.911 ;
      RECT 66.855 2.3 66.86 2.922 ;
      RECT 66.845 2.32 66.855 2.94 ;
      RECT 66.835 2.35 66.845 2.963 ;
      RECT 66.83 2.372 66.835 2.983 ;
      RECT 66.825 2.387 66.83 2.998 ;
      RECT 66.81 2.417 66.825 3.025 ;
      RECT 66.805 2.447 66.81 3.051 ;
      RECT 66.8 2.465 66.805 3.063 ;
      RECT 66.79 2.495 66.8 3.082 ;
      RECT 66.78 2.52 66.79 3.107 ;
      RECT 66.775 2.54 66.78 3.126 ;
      RECT 66.77 2.557 66.775 3.139 ;
      RECT 66.76 2.583 66.77 3.158 ;
      RECT 66.75 2.621 66.76 3.185 ;
      RECT 66.745 2.647 66.75 3.205 ;
      RECT 66.74 2.657 66.745 3.215 ;
      RECT 66.735 2.67 66.74 3.23 ;
      RECT 66.73 2.685 66.735 3.24 ;
      RECT 66.725 2.707 66.73 3.255 ;
      RECT 66.72 2.725 66.725 3.266 ;
      RECT 66.715 2.735 66.72 3.277 ;
      RECT 66.71 2.743 66.715 3.289 ;
      RECT 66.705 2.751 66.71 3.3 ;
      RECT 66.7 2.777 66.705 3.313 ;
      RECT 66.69 2.805 66.7 3.326 ;
      RECT 66.685 2.835 66.69 3.335 ;
      RECT 66.68 2.85 66.685 3.342 ;
      RECT 66.665 2.875 66.68 3.349 ;
      RECT 66.66 2.897 66.665 3.355 ;
      RECT 66.655 2.922 66.66 3.358 ;
      RECT 66.646 2.95 66.655 3.362 ;
      RECT 66.64 2.967 66.646 3.367 ;
      RECT 66.635 2.985 66.64 3.371 ;
      RECT 66.63 2.997 66.635 3.374 ;
      RECT 66.625 3.018 66.63 3.378 ;
      RECT 66.62 3.036 66.625 3.381 ;
      RECT 66.615 3.05 66.62 3.384 ;
      RECT 66.61 3.067 66.615 3.387 ;
      RECT 66.605 3.08 66.61 3.39 ;
      RECT 66.58 3.117 66.605 3.398 ;
      RECT 66.575 3.162 66.58 3.407 ;
      RECT 66.57 3.19 66.575 3.41 ;
      RECT 66.56 3.21 66.57 3.414 ;
      RECT 66.555 3.23 66.56 3.419 ;
      RECT 66.55 3.245 66.555 3.422 ;
      RECT 66.53 3.255 66.55 3.429 ;
      RECT 66.465 3.262 66.53 3.455 ;
      RECT 66.43 3.265 66.465 3.483 ;
      RECT 66.415 3.268 66.43 3.498 ;
      RECT 66.405 3.269 66.415 3.513 ;
      RECT 66.395 3.27 66.405 3.53 ;
      RECT 66.39 3.27 66.395 3.545 ;
      RECT 66.385 3.27 66.39 3.553 ;
      RECT 66.37 3.271 66.385 3.568 ;
      RECT 66.34 3.273 66.37 3.575 ;
      RECT 66.23 3.28 66.31 3.575 ;
      RECT 66.185 3.285 66.23 3.575 ;
      RECT 66.175 3.286 66.185 3.565 ;
      RECT 66.165 3.287 66.175 3.558 ;
      RECT 66.145 3.289 66.165 3.553 ;
      RECT 66.135 3.26 66.145 3.548 ;
      RECT 66.09 3.26 66.135 3.54 ;
      RECT 66.06 3.26 66.085 3.53 ;
      RECT 66.04 3.26 66.06 3.523 ;
      RECT 66.32 2.06 66.58 2.32 ;
      RECT 66.2 2.075 66.21 2.24 ;
      RECT 66.185 2.075 66.19 2.235 ;
      RECT 63.55 1.915 63.735 2.205 ;
      RECT 65.365 2.04 65.38 2.195 ;
      RECT 63.515 1.915 63.54 2.175 ;
      RECT 65.93 1.965 65.935 2.107 ;
      RECT 65.845 1.96 65.87 2.1 ;
      RECT 66.245 2.077 66.32 2.27 ;
      RECT 66.23 2.075 66.245 2.253 ;
      RECT 66.21 2.075 66.23 2.245 ;
      RECT 66.19 2.075 66.2 2.238 ;
      RECT 66.145 2.07 66.185 2.228 ;
      RECT 66.105 2.045 66.145 2.213 ;
      RECT 66.09 2.02 66.105 2.203 ;
      RECT 66.085 2.014 66.09 2.201 ;
      RECT 66.05 2.006 66.085 2.184 ;
      RECT 66.045 1.999 66.05 2.172 ;
      RECT 66.025 1.994 66.045 2.16 ;
      RECT 66.015 1.988 66.025 2.145 ;
      RECT 65.995 1.983 66.015 2.13 ;
      RECT 65.985 1.978 65.995 2.123 ;
      RECT 65.98 1.976 65.985 2.118 ;
      RECT 65.975 1.975 65.98 2.115 ;
      RECT 65.935 1.97 65.975 2.111 ;
      RECT 65.915 1.964 65.93 2.106 ;
      RECT 65.88 1.961 65.915 2.103 ;
      RECT 65.87 1.96 65.88 2.101 ;
      RECT 65.81 1.96 65.845 2.098 ;
      RECT 65.765 1.96 65.81 2.098 ;
      RECT 65.715 1.96 65.765 2.101 ;
      RECT 65.7 1.962 65.715 2.103 ;
      RECT 65.685 1.965 65.7 2.104 ;
      RECT 65.675 1.97 65.685 2.105 ;
      RECT 65.645 1.975 65.675 2.11 ;
      RECT 65.635 1.981 65.645 2.118 ;
      RECT 65.625 1.983 65.635 2.122 ;
      RECT 65.615 1.987 65.625 2.126 ;
      RECT 65.59 1.993 65.615 2.134 ;
      RECT 65.58 1.998 65.59 2.142 ;
      RECT 65.565 2.002 65.58 2.146 ;
      RECT 65.53 2.008 65.565 2.154 ;
      RECT 65.51 2.013 65.53 2.164 ;
      RECT 65.48 2.02 65.51 2.173 ;
      RECT 65.435 2.029 65.48 2.187 ;
      RECT 65.43 2.034 65.435 2.198 ;
      RECT 65.41 2.037 65.43 2.199 ;
      RECT 65.38 2.04 65.41 2.197 ;
      RECT 65.345 2.04 65.365 2.193 ;
      RECT 65.275 2.04 65.345 2.184 ;
      RECT 65.26 2.037 65.275 2.176 ;
      RECT 65.22 2.03 65.26 2.171 ;
      RECT 65.195 2.02 65.22 2.164 ;
      RECT 65.19 2.014 65.195 2.161 ;
      RECT 65.15 2.008 65.19 2.158 ;
      RECT 65.135 2.001 65.15 2.153 ;
      RECT 65.115 1.997 65.135 2.148 ;
      RECT 65.1 1.992 65.115 2.144 ;
      RECT 65.085 1.987 65.1 2.142 ;
      RECT 65.07 1.983 65.085 2.141 ;
      RECT 65.055 1.981 65.07 2.137 ;
      RECT 65.045 1.979 65.055 2.132 ;
      RECT 65.03 1.976 65.045 2.128 ;
      RECT 65.02 1.974 65.03 2.123 ;
      RECT 65 1.971 65.02 2.119 ;
      RECT 64.955 1.97 65 2.117 ;
      RECT 64.895 1.972 64.955 2.118 ;
      RECT 64.875 1.974 64.895 2.12 ;
      RECT 64.845 1.977 64.875 2.121 ;
      RECT 64.795 1.982 64.845 2.123 ;
      RECT 64.79 1.985 64.795 2.125 ;
      RECT 64.78 1.987 64.79 2.128 ;
      RECT 64.775 1.989 64.78 2.131 ;
      RECT 64.725 1.992 64.775 2.138 ;
      RECT 64.705 1.996 64.725 2.15 ;
      RECT 64.695 1.999 64.705 2.156 ;
      RECT 64.685 2 64.695 2.159 ;
      RECT 64.646 2.003 64.685 2.161 ;
      RECT 64.56 2.01 64.646 2.164 ;
      RECT 64.486 2.02 64.56 2.168 ;
      RECT 64.4 2.031 64.486 2.173 ;
      RECT 64.385 2.038 64.4 2.175 ;
      RECT 64.33 2.042 64.385 2.176 ;
      RECT 64.316 2.045 64.33 2.178 ;
      RECT 64.23 2.045 64.316 2.18 ;
      RECT 64.19 2.042 64.23 2.183 ;
      RECT 64.166 2.038 64.19 2.185 ;
      RECT 64.08 2.028 64.166 2.188 ;
      RECT 64.05 2.017 64.08 2.189 ;
      RECT 64.031 2.013 64.05 2.188 ;
      RECT 63.945 2.006 64.031 2.185 ;
      RECT 63.885 1.995 63.945 2.182 ;
      RECT 63.865 1.987 63.885 2.18 ;
      RECT 63.83 1.982 63.865 2.179 ;
      RECT 63.805 1.977 63.83 2.178 ;
      RECT 63.775 1.972 63.805 2.177 ;
      RECT 63.75 1.915 63.775 2.176 ;
      RECT 63.735 1.915 63.75 2.2 ;
      RECT 63.54 1.915 63.55 2.2 ;
      RECT 65.315 2.935 65.32 3.075 ;
      RECT 64.975 2.935 65.01 3.073 ;
      RECT 64.55 2.92 64.565 3.065 ;
      RECT 66.38 2.7 66.47 2.96 ;
      RECT 66.21 2.565 66.31 2.96 ;
      RECT 63.245 2.54 63.325 2.75 ;
      RECT 66.335 2.677 66.38 2.96 ;
      RECT 66.325 2.647 66.335 2.96 ;
      RECT 66.31 2.57 66.325 2.96 ;
      RECT 66.125 2.565 66.21 2.925 ;
      RECT 66.12 2.567 66.125 2.92 ;
      RECT 66.115 2.572 66.12 2.92 ;
      RECT 66.08 2.672 66.115 2.92 ;
      RECT 66.07 2.7 66.08 2.92 ;
      RECT 66.06 2.715 66.07 2.92 ;
      RECT 66.05 2.727 66.06 2.92 ;
      RECT 66.045 2.737 66.05 2.92 ;
      RECT 66.03 2.747 66.045 2.922 ;
      RECT 66.025 2.762 66.03 2.924 ;
      RECT 66.01 2.775 66.025 2.926 ;
      RECT 66.005 2.79 66.01 2.929 ;
      RECT 65.985 2.8 66.005 2.933 ;
      RECT 65.97 2.81 65.985 2.936 ;
      RECT 65.935 2.817 65.97 2.941 ;
      RECT 65.891 2.824 65.935 2.949 ;
      RECT 65.805 2.836 65.891 2.962 ;
      RECT 65.78 2.847 65.805 2.973 ;
      RECT 65.75 2.852 65.78 2.978 ;
      RECT 65.715 2.857 65.75 2.986 ;
      RECT 65.685 2.862 65.715 2.993 ;
      RECT 65.66 2.867 65.685 2.998 ;
      RECT 65.595 2.874 65.66 3.007 ;
      RECT 65.525 2.887 65.595 3.023 ;
      RECT 65.495 2.897 65.525 3.035 ;
      RECT 65.47 2.902 65.495 3.042 ;
      RECT 65.415 2.909 65.47 3.05 ;
      RECT 65.41 2.916 65.415 3.055 ;
      RECT 65.405 2.918 65.41 3.056 ;
      RECT 65.39 2.92 65.405 3.058 ;
      RECT 65.385 2.92 65.39 3.061 ;
      RECT 65.32 2.927 65.385 3.068 ;
      RECT 65.285 2.937 65.315 3.078 ;
      RECT 65.268 2.94 65.285 3.08 ;
      RECT 65.182 2.939 65.268 3.079 ;
      RECT 65.096 2.937 65.182 3.076 ;
      RECT 65.01 2.936 65.096 3.074 ;
      RECT 64.909 2.934 64.975 3.073 ;
      RECT 64.823 2.931 64.909 3.071 ;
      RECT 64.737 2.927 64.823 3.069 ;
      RECT 64.651 2.924 64.737 3.068 ;
      RECT 64.565 2.921 64.651 3.066 ;
      RECT 64.465 2.92 64.55 3.063 ;
      RECT 64.415 2.918 64.465 3.061 ;
      RECT 64.395 2.915 64.415 3.059 ;
      RECT 64.375 2.913 64.395 3.056 ;
      RECT 64.35 2.909 64.375 3.053 ;
      RECT 64.305 2.903 64.35 3.048 ;
      RECT 64.265 2.897 64.305 3.04 ;
      RECT 64.24 2.892 64.265 3.033 ;
      RECT 64.185 2.885 64.24 3.025 ;
      RECT 64.161 2.878 64.185 3.018 ;
      RECT 64.075 2.869 64.161 3.008 ;
      RECT 64.045 2.861 64.075 2.998 ;
      RECT 64.015 2.857 64.045 2.993 ;
      RECT 64.01 2.854 64.015 2.99 ;
      RECT 64.005 2.853 64.01 2.99 ;
      RECT 63.93 2.846 64.005 2.983 ;
      RECT 63.891 2.837 63.93 2.972 ;
      RECT 63.805 2.827 63.891 2.96 ;
      RECT 63.765 2.817 63.805 2.948 ;
      RECT 63.726 2.812 63.765 2.941 ;
      RECT 63.64 2.802 63.726 2.93 ;
      RECT 63.6 2.79 63.64 2.919 ;
      RECT 63.565 2.775 63.6 2.912 ;
      RECT 63.555 2.765 63.565 2.909 ;
      RECT 63.535 2.75 63.555 2.907 ;
      RECT 63.505 2.72 63.535 2.903 ;
      RECT 63.495 2.7 63.505 2.898 ;
      RECT 63.49 2.692 63.495 2.895 ;
      RECT 63.485 2.685 63.49 2.893 ;
      RECT 63.47 2.672 63.485 2.886 ;
      RECT 63.465 2.662 63.47 2.878 ;
      RECT 63.46 2.655 63.465 2.873 ;
      RECT 63.455 2.65 63.46 2.869 ;
      RECT 63.44 2.637 63.455 2.861 ;
      RECT 63.435 2.547 63.44 2.85 ;
      RECT 63.43 2.542 63.435 2.843 ;
      RECT 63.355 2.54 63.43 2.803 ;
      RECT 63.325 2.54 63.355 2.758 ;
      RECT 63.23 2.545 63.245 2.745 ;
      RECT 65.715 2.25 65.975 2.51 ;
      RECT 65.7 2.238 65.88 2.475 ;
      RECT 65.695 2.239 65.88 2.473 ;
      RECT 65.68 2.243 65.89 2.463 ;
      RECT 65.675 2.248 65.895 2.433 ;
      RECT 65.68 2.245 65.895 2.463 ;
      RECT 65.695 2.24 65.89 2.473 ;
      RECT 65.715 2.237 65.88 2.51 ;
      RECT 65.715 2.236 65.87 2.51 ;
      RECT 65.74 2.235 65.87 2.51 ;
      RECT 65.3 2.48 65.56 2.74 ;
      RECT 65.175 2.525 65.56 2.735 ;
      RECT 65.165 2.53 65.56 2.73 ;
      RECT 65.18 3.47 65.195 3.78 ;
      RECT 63.775 3.24 63.785 3.37 ;
      RECT 63.555 3.235 63.66 3.37 ;
      RECT 63.47 3.24 63.52 3.37 ;
      RECT 62.02 1.975 62.025 3.08 ;
      RECT 65.275 3.562 65.28 3.698 ;
      RECT 65.27 3.557 65.275 3.758 ;
      RECT 65.265 3.555 65.27 3.771 ;
      RECT 65.25 3.552 65.265 3.773 ;
      RECT 65.245 3.547 65.25 3.775 ;
      RECT 65.24 3.543 65.245 3.778 ;
      RECT 65.225 3.538 65.24 3.78 ;
      RECT 65.195 3.53 65.225 3.78 ;
      RECT 65.156 3.47 65.18 3.78 ;
      RECT 65.07 3.47 65.156 3.777 ;
      RECT 65.04 3.47 65.07 3.77 ;
      RECT 65.015 3.47 65.04 3.763 ;
      RECT 64.99 3.47 65.015 3.755 ;
      RECT 64.975 3.47 64.99 3.748 ;
      RECT 64.95 3.47 64.975 3.74 ;
      RECT 64.935 3.47 64.95 3.733 ;
      RECT 64.895 3.48 64.935 3.722 ;
      RECT 64.885 3.475 64.895 3.712 ;
      RECT 64.881 3.474 64.885 3.709 ;
      RECT 64.795 3.466 64.881 3.692 ;
      RECT 64.762 3.455 64.795 3.669 ;
      RECT 64.676 3.444 64.762 3.647 ;
      RECT 64.59 3.428 64.676 3.616 ;
      RECT 64.52 3.413 64.59 3.588 ;
      RECT 64.51 3.406 64.52 3.575 ;
      RECT 64.48 3.403 64.51 3.565 ;
      RECT 64.455 3.399 64.48 3.558 ;
      RECT 64.44 3.396 64.455 3.553 ;
      RECT 64.435 3.395 64.44 3.548 ;
      RECT 64.405 3.39 64.435 3.541 ;
      RECT 64.4 3.385 64.405 3.536 ;
      RECT 64.385 3.382 64.4 3.531 ;
      RECT 64.38 3.377 64.385 3.526 ;
      RECT 64.36 3.372 64.38 3.523 ;
      RECT 64.345 3.367 64.36 3.515 ;
      RECT 64.33 3.361 64.345 3.51 ;
      RECT 64.3 3.352 64.33 3.503 ;
      RECT 64.295 3.345 64.3 3.495 ;
      RECT 64.29 3.343 64.295 3.493 ;
      RECT 64.285 3.342 64.29 3.49 ;
      RECT 64.245 3.335 64.285 3.483 ;
      RECT 64.231 3.325 64.245 3.473 ;
      RECT 64.18 3.314 64.231 3.461 ;
      RECT 64.155 3.3 64.18 3.447 ;
      RECT 64.13 3.289 64.155 3.439 ;
      RECT 64.11 3.278 64.13 3.433 ;
      RECT 64.1 3.272 64.11 3.428 ;
      RECT 64.095 3.27 64.1 3.424 ;
      RECT 64.075 3.265 64.095 3.419 ;
      RECT 64.045 3.255 64.075 3.409 ;
      RECT 64.04 3.247 64.045 3.402 ;
      RECT 64.025 3.245 64.04 3.398 ;
      RECT 64.005 3.245 64.025 3.393 ;
      RECT 64 3.244 64.005 3.391 ;
      RECT 63.995 3.244 64 3.388 ;
      RECT 63.955 3.243 63.995 3.383 ;
      RECT 63.93 3.242 63.955 3.378 ;
      RECT 63.87 3.241 63.93 3.375 ;
      RECT 63.785 3.24 63.87 3.373 ;
      RECT 63.746 3.239 63.775 3.37 ;
      RECT 63.66 3.237 63.746 3.37 ;
      RECT 63.52 3.237 63.555 3.37 ;
      RECT 63.43 3.241 63.47 3.373 ;
      RECT 63.415 3.244 63.43 3.38 ;
      RECT 63.405 3.245 63.415 3.387 ;
      RECT 63.38 3.248 63.405 3.392 ;
      RECT 63.375 3.25 63.38 3.395 ;
      RECT 63.325 3.252 63.375 3.396 ;
      RECT 63.286 3.256 63.325 3.398 ;
      RECT 63.2 3.258 63.286 3.401 ;
      RECT 63.182 3.26 63.2 3.403 ;
      RECT 63.096 3.263 63.182 3.405 ;
      RECT 63.01 3.267 63.096 3.408 ;
      RECT 62.973 3.271 63.01 3.411 ;
      RECT 62.887 3.274 62.973 3.414 ;
      RECT 62.801 3.278 62.887 3.417 ;
      RECT 62.715 3.283 62.801 3.421 ;
      RECT 62.695 3.285 62.715 3.424 ;
      RECT 62.675 3.284 62.695 3.425 ;
      RECT 62.626 3.281 62.675 3.426 ;
      RECT 62.54 3.276 62.626 3.429 ;
      RECT 62.49 3.271 62.54 3.431 ;
      RECT 62.466 3.269 62.49 3.432 ;
      RECT 62.38 3.264 62.466 3.434 ;
      RECT 62.355 3.26 62.38 3.433 ;
      RECT 62.345 3.257 62.355 3.431 ;
      RECT 62.335 3.25 62.345 3.428 ;
      RECT 62.33 3.23 62.335 3.423 ;
      RECT 62.32 3.2 62.33 3.418 ;
      RECT 62.305 3.07 62.32 3.409 ;
      RECT 62.3 3.062 62.305 3.402 ;
      RECT 62.28 3.055 62.3 3.394 ;
      RECT 62.275 3.037 62.28 3.386 ;
      RECT 62.265 3.017 62.275 3.381 ;
      RECT 62.26 2.99 62.265 3.377 ;
      RECT 62.255 2.967 62.26 3.374 ;
      RECT 62.235 2.925 62.255 3.366 ;
      RECT 62.2 2.84 62.235 3.35 ;
      RECT 62.195 2.772 62.2 3.338 ;
      RECT 62.18 2.742 62.195 3.332 ;
      RECT 62.175 1.987 62.18 2.233 ;
      RECT 62.165 2.712 62.18 3.323 ;
      RECT 62.17 1.982 62.175 2.265 ;
      RECT 62.165 1.977 62.17 2.308 ;
      RECT 62.16 1.975 62.165 2.343 ;
      RECT 62.145 2.675 62.165 3.313 ;
      RECT 62.155 1.975 62.16 2.38 ;
      RECT 62.14 1.975 62.155 2.478 ;
      RECT 62.14 2.648 62.145 3.306 ;
      RECT 62.135 1.975 62.14 2.553 ;
      RECT 62.135 2.636 62.14 3.303 ;
      RECT 62.13 1.975 62.135 2.585 ;
      RECT 62.13 2.615 62.135 3.3 ;
      RECT 62.125 1.975 62.13 3.297 ;
      RECT 62.09 1.975 62.125 3.283 ;
      RECT 62.075 1.975 62.09 3.265 ;
      RECT 62.055 1.975 62.075 3.255 ;
      RECT 62.03 1.975 62.055 3.238 ;
      RECT 62.025 1.975 62.03 3.188 ;
      RECT 62.015 1.975 62.02 3.018 ;
      RECT 62.01 1.975 62.015 2.925 ;
      RECT 62.005 1.975 62.01 2.838 ;
      RECT 62 1.975 62.005 2.77 ;
      RECT 61.995 1.975 62 2.713 ;
      RECT 61.985 1.975 61.995 2.608 ;
      RECT 61.98 1.975 61.985 2.48 ;
      RECT 61.975 1.975 61.98 2.398 ;
      RECT 61.97 1.977 61.975 2.315 ;
      RECT 61.965 1.982 61.97 2.248 ;
      RECT 61.96 1.987 61.965 2.175 ;
      RECT 64.775 2.305 65.035 2.565 ;
      RECT 64.795 2.272 65.005 2.565 ;
      RECT 64.795 2.27 64.995 2.565 ;
      RECT 64.805 2.257 64.995 2.565 ;
      RECT 64.805 2.255 64.92 2.565 ;
      RECT 64.28 2.38 64.455 2.66 ;
      RECT 64.275 2.38 64.455 2.658 ;
      RECT 64.275 2.38 64.47 2.655 ;
      RECT 64.265 2.38 64.47 2.653 ;
      RECT 64.21 2.38 64.47 2.64 ;
      RECT 64.21 2.455 64.475 2.618 ;
      RECT 63.755 2.392 63.775 2.635 ;
      RECT 63.755 2.392 63.815 2.634 ;
      RECT 63.75 2.394 63.815 2.633 ;
      RECT 63.75 2.394 63.901 2.632 ;
      RECT 63.75 2.394 63.97 2.631 ;
      RECT 63.75 2.394 63.99 2.623 ;
      RECT 63.73 2.397 63.99 2.621 ;
      RECT 63.715 2.407 63.99 2.606 ;
      RECT 63.715 2.407 64.005 2.605 ;
      RECT 63.71 2.416 64.005 2.597 ;
      RECT 63.71 2.416 64.01 2.593 ;
      RECT 63.815 2.33 64.075 2.59 ;
      RECT 63.705 2.418 64.075 2.475 ;
      RECT 63.775 2.385 64.075 2.59 ;
      RECT 63.74 3.578 63.745 3.785 ;
      RECT 63.69 3.572 63.74 3.784 ;
      RECT 63.657 3.586 63.75 3.783 ;
      RECT 63.571 3.586 63.75 3.782 ;
      RECT 63.485 3.586 63.75 3.781 ;
      RECT 63.485 3.685 63.755 3.778 ;
      RECT 63.48 3.685 63.755 3.773 ;
      RECT 63.475 3.685 63.755 3.755 ;
      RECT 63.47 3.685 63.755 3.738 ;
      RECT 63.43 3.47 63.69 3.73 ;
      RECT 62.89 2.62 62.976 3.034 ;
      RECT 62.89 2.62 63.015 3.031 ;
      RECT 62.89 2.62 63.035 3.021 ;
      RECT 62.845 2.62 63.035 3.018 ;
      RECT 62.845 2.772 63.045 3.008 ;
      RECT 62.845 2.793 63.05 3.002 ;
      RECT 62.845 2.811 63.055 2.998 ;
      RECT 62.845 2.831 63.065 2.993 ;
      RECT 62.82 2.831 63.065 2.99 ;
      RECT 62.81 2.831 63.065 2.968 ;
      RECT 62.81 2.847 63.07 2.938 ;
      RECT 62.775 2.62 63.035 2.925 ;
      RECT 62.775 2.859 63.075 2.88 ;
      RECT 60.44 7.765 60.73 7.995 ;
      RECT 60.5 6.285 60.67 7.995 ;
      RECT 60.445 6.655 60.795 7.005 ;
      RECT 60.44 6.285 60.73 6.515 ;
      RECT 60.44 2.365 60.73 2.595 ;
      RECT 60.5 0.885 60.67 2.595 ;
      RECT 60.44 0.885 60.73 1.115 ;
      RECT 60.03 2.735 60.36 2.965 ;
      RECT 60.03 2.765 60.53 2.935 ;
      RECT 60.03 2.395 60.22 2.965 ;
      RECT 59.45 2.365 59.74 2.595 ;
      RECT 59.45 2.395 60.22 2.565 ;
      RECT 59.51 0.885 59.68 2.595 ;
      RECT 59.45 0.885 59.74 1.115 ;
      RECT 59.45 7.765 59.74 7.995 ;
      RECT 59.51 6.285 59.68 7.995 ;
      RECT 59.45 6.285 59.74 6.515 ;
      RECT 59.45 6.325 60.3 6.485 ;
      RECT 60.13 5.915 60.3 6.485 ;
      RECT 59.45 6.32 59.84 6.485 ;
      RECT 60.07 5.915 60.36 6.145 ;
      RECT 60.07 5.945 60.53 6.115 ;
      RECT 59.08 2.735 59.37 2.965 ;
      RECT 59.08 2.765 59.54 2.935 ;
      RECT 59.14 1.655 59.305 2.965 ;
      RECT 57.655 1.625 57.945 1.855 ;
      RECT 57.655 1.655 59.305 1.825 ;
      RECT 57.715 0.885 57.885 1.855 ;
      RECT 57.655 0.885 57.945 1.115 ;
      RECT 57.655 7.765 57.945 7.995 ;
      RECT 57.715 7.025 57.885 7.995 ;
      RECT 57.715 7.12 59.305 7.29 ;
      RECT 59.135 5.915 59.305 7.29 ;
      RECT 57.655 7.025 57.945 7.255 ;
      RECT 59.08 5.915 59.37 6.145 ;
      RECT 59.08 5.945 59.54 6.115 ;
      RECT 55.705 2.705 56.045 3.055 ;
      RECT 55.795 2.025 55.965 3.055 ;
      RECT 58.085 1.965 58.435 2.315 ;
      RECT 55.795 2.025 58.435 2.195 ;
      RECT 58.11 6.655 58.435 6.98 ;
      RECT 52.65 6.61 53 6.96 ;
      RECT 58.085 6.655 58.435 6.885 ;
      RECT 52.45 6.655 53 6.885 ;
      RECT 52.28 6.685 58.435 6.855 ;
      RECT 57.31 2.365 57.63 2.685 ;
      RECT 57.28 2.365 57.63 2.595 ;
      RECT 57.11 2.395 57.63 2.565 ;
      RECT 57.31 6.255 57.63 6.545 ;
      RECT 57.28 6.285 57.63 6.515 ;
      RECT 57.11 6.315 57.63 6.485 ;
      RECT 56.265 2.705 56.605 3.055 ;
      RECT 56.265 2.765 56.745 2.935 ;
      RECT 56.26 5.86 56.6 6.21 ;
      RECT 50.65 5.915 50.94 6.145 ;
      RECT 50.65 5.945 56.745 6.115 ;
      RECT 53 2.985 53.15 3.26 ;
      RECT 53.54 2.065 53.545 2.285 ;
      RECT 54.69 2.265 54.705 2.463 ;
      RECT 54.655 2.257 54.69 2.47 ;
      RECT 54.625 2.25 54.655 2.47 ;
      RECT 54.57 2.215 54.625 2.47 ;
      RECT 54.505 2.152 54.57 2.47 ;
      RECT 54.5 2.117 54.505 2.468 ;
      RECT 54.495 2.112 54.5 2.46 ;
      RECT 54.49 2.107 54.495 2.446 ;
      RECT 54.485 2.104 54.49 2.439 ;
      RECT 54.44 2.094 54.485 2.39 ;
      RECT 54.42 2.081 54.44 2.325 ;
      RECT 54.415 2.076 54.42 2.298 ;
      RECT 54.41 2.075 54.415 2.291 ;
      RECT 54.405 2.074 54.41 2.284 ;
      RECT 54.32 2.059 54.405 2.23 ;
      RECT 54.29 2.04 54.32 2.18 ;
      RECT 54.21 2.023 54.29 2.165 ;
      RECT 54.175 2.01 54.21 2.15 ;
      RECT 54.167 2.01 54.175 2.145 ;
      RECT 54.081 2.011 54.167 2.145 ;
      RECT 53.995 2.013 54.081 2.145 ;
      RECT 53.97 2.014 53.995 2.149 ;
      RECT 53.895 2.02 53.97 2.164 ;
      RECT 53.812 2.032 53.895 2.188 ;
      RECT 53.726 2.045 53.812 2.214 ;
      RECT 53.64 2.058 53.726 2.24 ;
      RECT 53.605 2.067 53.64 2.259 ;
      RECT 53.555 2.067 53.605 2.272 ;
      RECT 53.545 2.065 53.555 2.283 ;
      RECT 53.53 2.062 53.54 2.285 ;
      RECT 53.515 2.054 53.53 2.293 ;
      RECT 53.5 2.046 53.515 2.313 ;
      RECT 53.495 2.041 53.5 2.37 ;
      RECT 53.48 2.036 53.495 2.443 ;
      RECT 53.475 2.031 53.48 2.485 ;
      RECT 53.47 2.029 53.475 2.513 ;
      RECT 53.465 2.027 53.47 2.535 ;
      RECT 53.455 2.023 53.465 2.578 ;
      RECT 53.45 2.02 53.455 2.603 ;
      RECT 53.445 2.018 53.45 2.623 ;
      RECT 53.44 2.016 53.445 2.647 ;
      RECT 53.435 2.012 53.44 2.67 ;
      RECT 53.43 2.008 53.435 2.693 ;
      RECT 53.395 1.998 53.43 2.8 ;
      RECT 53.39 1.988 53.395 2.898 ;
      RECT 53.385 1.986 53.39 2.925 ;
      RECT 53.38 1.985 53.385 2.945 ;
      RECT 53.375 1.977 53.38 2.965 ;
      RECT 53.37 1.972 53.375 3 ;
      RECT 53.365 1.97 53.37 3.018 ;
      RECT 53.36 1.97 53.365 3.043 ;
      RECT 53.355 1.97 53.36 3.065 ;
      RECT 53.32 1.97 53.355 3.108 ;
      RECT 53.295 1.97 53.32 3.137 ;
      RECT 53.285 1.97 53.295 2.323 ;
      RECT 53.288 2.38 53.295 3.147 ;
      RECT 53.285 2.437 53.288 3.15 ;
      RECT 53.28 1.97 53.285 2.295 ;
      RECT 53.28 2.487 53.285 3.153 ;
      RECT 53.27 1.97 53.28 2.285 ;
      RECT 53.275 2.54 53.28 3.156 ;
      RECT 53.27 2.625 53.275 3.16 ;
      RECT 53.26 1.97 53.27 2.273 ;
      RECT 53.265 2.672 53.27 3.164 ;
      RECT 53.26 2.747 53.265 3.168 ;
      RECT 53.225 1.97 53.26 2.248 ;
      RECT 53.25 2.83 53.26 3.173 ;
      RECT 53.24 2.897 53.25 3.18 ;
      RECT 53.235 2.925 53.24 3.185 ;
      RECT 53.225 2.938 53.235 3.191 ;
      RECT 53.18 1.97 53.225 2.205 ;
      RECT 53.22 2.943 53.225 3.198 ;
      RECT 53.18 2.96 53.22 3.26 ;
      RECT 53.175 1.972 53.18 2.178 ;
      RECT 53.15 2.98 53.18 3.26 ;
      RECT 53.17 1.977 53.175 2.15 ;
      RECT 52.96 2.989 53 3.26 ;
      RECT 52.935 2.997 52.96 3.23 ;
      RECT 52.89 3.005 52.935 3.23 ;
      RECT 52.875 3.01 52.89 3.225 ;
      RECT 52.865 3.01 52.875 3.219 ;
      RECT 52.855 3.017 52.865 3.216 ;
      RECT 52.85 3.055 52.855 3.205 ;
      RECT 52.845 3.117 52.85 3.183 ;
      RECT 54.115 2.992 54.3 3.215 ;
      RECT 54.115 3.007 54.305 3.211 ;
      RECT 54.105 2.28 54.19 3.21 ;
      RECT 54.105 3.007 54.31 3.204 ;
      RECT 54.1 3.015 54.31 3.203 ;
      RECT 54.305 2.735 54.625 3.055 ;
      RECT 54.1 2.907 54.27 2.998 ;
      RECT 54.095 2.907 54.27 2.98 ;
      RECT 54.085 2.715 54.22 2.955 ;
      RECT 54.08 2.715 54.22 2.9 ;
      RECT 54.04 2.295 54.21 2.8 ;
      RECT 54.025 2.295 54.21 2.67 ;
      RECT 54.02 2.295 54.21 2.623 ;
      RECT 54.015 2.295 54.21 2.603 ;
      RECT 54.01 2.295 54.21 2.578 ;
      RECT 53.98 2.295 54.24 2.555 ;
      RECT 53.99 2.292 54.2 2.555 ;
      RECT 54.115 2.287 54.2 3.215 ;
      RECT 54 2.28 54.19 2.555 ;
      RECT 53.995 2.285 54.19 2.555 ;
      RECT 52.825 2.497 53.01 2.71 ;
      RECT 52.825 2.505 53.02 2.703 ;
      RECT 52.805 2.505 53.02 2.7 ;
      RECT 52.8 2.505 53.02 2.685 ;
      RECT 52.73 2.42 52.99 2.68 ;
      RECT 52.73 2.565 53.025 2.593 ;
      RECT 52.385 3.02 52.645 3.28 ;
      RECT 52.41 2.965 52.605 3.28 ;
      RECT 52.405 2.714 52.585 3.008 ;
      RECT 52.405 2.72 52.595 3.008 ;
      RECT 52.385 2.722 52.595 2.953 ;
      RECT 52.38 2.732 52.595 2.82 ;
      RECT 52.41 2.712 52.585 3.28 ;
      RECT 52.496 2.71 52.585 3.28 ;
      RECT 52.355 1.93 52.39 2.3 ;
      RECT 52.145 2.04 52.15 2.3 ;
      RECT 52.39 1.937 52.405 2.3 ;
      RECT 52.28 1.93 52.355 2.378 ;
      RECT 52.27 1.93 52.28 2.463 ;
      RECT 52.245 1.93 52.27 2.498 ;
      RECT 52.205 1.93 52.245 2.566 ;
      RECT 52.195 1.937 52.205 2.618 ;
      RECT 52.165 2.04 52.195 2.659 ;
      RECT 52.16 2.04 52.165 2.698 ;
      RECT 52.15 2.04 52.16 2.718 ;
      RECT 52.145 2.335 52.15 2.755 ;
      RECT 52.14 2.352 52.145 2.775 ;
      RECT 52.125 2.415 52.14 2.815 ;
      RECT 52.12 2.458 52.125 2.85 ;
      RECT 52.115 2.466 52.12 2.863 ;
      RECT 52.105 2.48 52.115 2.885 ;
      RECT 52.08 2.515 52.105 2.95 ;
      RECT 52.07 2.55 52.08 3.013 ;
      RECT 52.05 2.58 52.07 3.074 ;
      RECT 52.035 2.616 52.05 3.141 ;
      RECT 52.025 2.644 52.035 3.18 ;
      RECT 52.015 2.666 52.025 3.2 ;
      RECT 52.01 2.676 52.015 3.211 ;
      RECT 52.005 2.685 52.01 3.214 ;
      RECT 51.995 2.703 52.005 3.218 ;
      RECT 51.985 2.721 51.995 3.219 ;
      RECT 51.96 2.76 51.985 3.216 ;
      RECT 51.94 2.802 51.96 3.213 ;
      RECT 51.925 2.84 51.94 3.212 ;
      RECT 51.89 2.875 51.925 3.209 ;
      RECT 51.885 2.897 51.89 3.207 ;
      RECT 51.82 2.937 51.885 3.204 ;
      RECT 51.815 2.977 51.82 3.2 ;
      RECT 51.8 2.987 51.815 3.191 ;
      RECT 51.79 3.107 51.8 3.176 ;
      RECT 52.27 3.52 52.28 3.78 ;
      RECT 52.27 3.523 52.29 3.779 ;
      RECT 52.26 3.513 52.27 3.778 ;
      RECT 52.25 3.528 52.33 3.774 ;
      RECT 52.235 3.507 52.25 3.772 ;
      RECT 52.21 3.532 52.335 3.768 ;
      RECT 52.195 3.492 52.21 3.763 ;
      RECT 52.195 3.534 52.345 3.762 ;
      RECT 52.195 3.542 52.36 3.755 ;
      RECT 52.135 3.479 52.195 3.745 ;
      RECT 52.125 3.466 52.135 3.727 ;
      RECT 52.1 3.456 52.125 3.717 ;
      RECT 52.095 3.446 52.1 3.709 ;
      RECT 52.03 3.542 52.36 3.691 ;
      RECT 51.945 3.542 52.36 3.653 ;
      RECT 51.835 3.37 52.095 3.63 ;
      RECT 52.21 3.5 52.235 3.768 ;
      RECT 52.25 3.51 52.26 3.774 ;
      RECT 51.835 3.518 52.275 3.63 ;
      RECT 52.02 7.765 52.31 7.995 ;
      RECT 52.08 7.025 52.25 7.995 ;
      RECT 51.98 7.055 52.35 7.425 ;
      RECT 52.02 7.025 52.31 7.425 ;
      RECT 51.05 3.275 51.08 3.575 ;
      RECT 50.825 3.26 50.83 3.535 ;
      RECT 50.625 3.26 50.78 3.52 ;
      RECT 51.925 1.975 51.955 2.235 ;
      RECT 51.915 1.975 51.925 2.343 ;
      RECT 51.895 1.975 51.915 2.353 ;
      RECT 51.88 1.975 51.895 2.365 ;
      RECT 51.825 1.975 51.88 2.415 ;
      RECT 51.81 1.975 51.825 2.463 ;
      RECT 51.78 1.975 51.81 2.498 ;
      RECT 51.725 1.975 51.78 2.56 ;
      RECT 51.705 1.975 51.725 2.628 ;
      RECT 51.7 1.975 51.705 2.658 ;
      RECT 51.695 1.975 51.7 2.67 ;
      RECT 51.69 2.092 51.695 2.688 ;
      RECT 51.67 2.11 51.69 2.713 ;
      RECT 51.65 2.137 51.67 2.763 ;
      RECT 51.645 2.157 51.65 2.794 ;
      RECT 51.64 2.165 51.645 2.811 ;
      RECT 51.625 2.191 51.64 2.84 ;
      RECT 51.61 2.233 51.625 2.875 ;
      RECT 51.605 2.262 51.61 2.898 ;
      RECT 51.6 2.277 51.605 2.911 ;
      RECT 51.595 2.3 51.6 2.922 ;
      RECT 51.585 2.32 51.595 2.94 ;
      RECT 51.575 2.35 51.585 2.963 ;
      RECT 51.57 2.372 51.575 2.983 ;
      RECT 51.565 2.387 51.57 2.998 ;
      RECT 51.55 2.417 51.565 3.025 ;
      RECT 51.545 2.447 51.55 3.051 ;
      RECT 51.54 2.465 51.545 3.063 ;
      RECT 51.53 2.495 51.54 3.082 ;
      RECT 51.52 2.52 51.53 3.107 ;
      RECT 51.515 2.54 51.52 3.126 ;
      RECT 51.51 2.557 51.515 3.139 ;
      RECT 51.5 2.583 51.51 3.158 ;
      RECT 51.49 2.621 51.5 3.185 ;
      RECT 51.485 2.647 51.49 3.205 ;
      RECT 51.48 2.657 51.485 3.215 ;
      RECT 51.475 2.67 51.48 3.23 ;
      RECT 51.47 2.685 51.475 3.24 ;
      RECT 51.465 2.707 51.47 3.255 ;
      RECT 51.46 2.725 51.465 3.266 ;
      RECT 51.455 2.735 51.46 3.277 ;
      RECT 51.45 2.743 51.455 3.289 ;
      RECT 51.445 2.751 51.45 3.3 ;
      RECT 51.44 2.777 51.445 3.313 ;
      RECT 51.43 2.805 51.44 3.326 ;
      RECT 51.425 2.835 51.43 3.335 ;
      RECT 51.42 2.85 51.425 3.342 ;
      RECT 51.405 2.875 51.42 3.349 ;
      RECT 51.4 2.897 51.405 3.355 ;
      RECT 51.395 2.922 51.4 3.358 ;
      RECT 51.386 2.95 51.395 3.362 ;
      RECT 51.38 2.967 51.386 3.367 ;
      RECT 51.375 2.985 51.38 3.371 ;
      RECT 51.37 2.997 51.375 3.374 ;
      RECT 51.365 3.018 51.37 3.378 ;
      RECT 51.36 3.036 51.365 3.381 ;
      RECT 51.355 3.05 51.36 3.384 ;
      RECT 51.35 3.067 51.355 3.387 ;
      RECT 51.345 3.08 51.35 3.39 ;
      RECT 51.32 3.117 51.345 3.398 ;
      RECT 51.315 3.162 51.32 3.407 ;
      RECT 51.31 3.19 51.315 3.41 ;
      RECT 51.3 3.21 51.31 3.414 ;
      RECT 51.295 3.23 51.3 3.419 ;
      RECT 51.29 3.245 51.295 3.422 ;
      RECT 51.27 3.255 51.29 3.429 ;
      RECT 51.205 3.262 51.27 3.455 ;
      RECT 51.17 3.265 51.205 3.483 ;
      RECT 51.155 3.268 51.17 3.498 ;
      RECT 51.145 3.269 51.155 3.513 ;
      RECT 51.135 3.27 51.145 3.53 ;
      RECT 51.13 3.27 51.135 3.545 ;
      RECT 51.125 3.27 51.13 3.553 ;
      RECT 51.11 3.271 51.125 3.568 ;
      RECT 51.08 3.273 51.11 3.575 ;
      RECT 50.97 3.28 51.05 3.575 ;
      RECT 50.925 3.285 50.97 3.575 ;
      RECT 50.915 3.286 50.925 3.565 ;
      RECT 50.905 3.287 50.915 3.558 ;
      RECT 50.885 3.289 50.905 3.553 ;
      RECT 50.875 3.26 50.885 3.548 ;
      RECT 50.83 3.26 50.875 3.54 ;
      RECT 50.8 3.26 50.825 3.53 ;
      RECT 50.78 3.26 50.8 3.523 ;
      RECT 51.06 2.06 51.32 2.32 ;
      RECT 50.94 2.075 50.95 2.24 ;
      RECT 50.925 2.075 50.93 2.235 ;
      RECT 48.29 1.915 48.475 2.205 ;
      RECT 50.105 2.04 50.12 2.195 ;
      RECT 48.255 1.915 48.28 2.175 ;
      RECT 50.67 1.965 50.675 2.107 ;
      RECT 50.585 1.96 50.61 2.1 ;
      RECT 50.985 2.077 51.06 2.27 ;
      RECT 50.97 2.075 50.985 2.253 ;
      RECT 50.95 2.075 50.97 2.245 ;
      RECT 50.93 2.075 50.94 2.238 ;
      RECT 50.885 2.07 50.925 2.228 ;
      RECT 50.845 2.045 50.885 2.213 ;
      RECT 50.83 2.02 50.845 2.203 ;
      RECT 50.825 2.014 50.83 2.201 ;
      RECT 50.79 2.006 50.825 2.184 ;
      RECT 50.785 1.999 50.79 2.172 ;
      RECT 50.765 1.994 50.785 2.16 ;
      RECT 50.755 1.988 50.765 2.145 ;
      RECT 50.735 1.983 50.755 2.13 ;
      RECT 50.725 1.978 50.735 2.123 ;
      RECT 50.72 1.976 50.725 2.118 ;
      RECT 50.715 1.975 50.72 2.115 ;
      RECT 50.675 1.97 50.715 2.111 ;
      RECT 50.655 1.964 50.67 2.106 ;
      RECT 50.62 1.961 50.655 2.103 ;
      RECT 50.61 1.96 50.62 2.101 ;
      RECT 50.55 1.96 50.585 2.098 ;
      RECT 50.505 1.96 50.55 2.098 ;
      RECT 50.455 1.96 50.505 2.101 ;
      RECT 50.44 1.962 50.455 2.103 ;
      RECT 50.425 1.965 50.44 2.104 ;
      RECT 50.415 1.97 50.425 2.105 ;
      RECT 50.385 1.975 50.415 2.11 ;
      RECT 50.375 1.981 50.385 2.118 ;
      RECT 50.365 1.983 50.375 2.122 ;
      RECT 50.355 1.987 50.365 2.126 ;
      RECT 50.33 1.993 50.355 2.134 ;
      RECT 50.32 1.998 50.33 2.142 ;
      RECT 50.305 2.002 50.32 2.146 ;
      RECT 50.27 2.008 50.305 2.154 ;
      RECT 50.25 2.013 50.27 2.164 ;
      RECT 50.22 2.02 50.25 2.173 ;
      RECT 50.175 2.029 50.22 2.187 ;
      RECT 50.17 2.034 50.175 2.198 ;
      RECT 50.15 2.037 50.17 2.199 ;
      RECT 50.12 2.04 50.15 2.197 ;
      RECT 50.085 2.04 50.105 2.193 ;
      RECT 50.015 2.04 50.085 2.184 ;
      RECT 50 2.037 50.015 2.176 ;
      RECT 49.96 2.03 50 2.171 ;
      RECT 49.935 2.02 49.96 2.164 ;
      RECT 49.93 2.014 49.935 2.161 ;
      RECT 49.89 2.008 49.93 2.158 ;
      RECT 49.875 2.001 49.89 2.153 ;
      RECT 49.855 1.997 49.875 2.148 ;
      RECT 49.84 1.992 49.855 2.144 ;
      RECT 49.825 1.987 49.84 2.142 ;
      RECT 49.81 1.983 49.825 2.141 ;
      RECT 49.795 1.981 49.81 2.137 ;
      RECT 49.785 1.979 49.795 2.132 ;
      RECT 49.77 1.976 49.785 2.128 ;
      RECT 49.76 1.974 49.77 2.123 ;
      RECT 49.74 1.971 49.76 2.119 ;
      RECT 49.695 1.97 49.74 2.117 ;
      RECT 49.635 1.972 49.695 2.118 ;
      RECT 49.615 1.974 49.635 2.12 ;
      RECT 49.585 1.977 49.615 2.121 ;
      RECT 49.535 1.982 49.585 2.123 ;
      RECT 49.53 1.985 49.535 2.125 ;
      RECT 49.52 1.987 49.53 2.128 ;
      RECT 49.515 1.989 49.52 2.131 ;
      RECT 49.465 1.992 49.515 2.138 ;
      RECT 49.445 1.996 49.465 2.15 ;
      RECT 49.435 1.999 49.445 2.156 ;
      RECT 49.425 2 49.435 2.159 ;
      RECT 49.386 2.003 49.425 2.161 ;
      RECT 49.3 2.01 49.386 2.164 ;
      RECT 49.226 2.02 49.3 2.168 ;
      RECT 49.14 2.031 49.226 2.173 ;
      RECT 49.125 2.038 49.14 2.175 ;
      RECT 49.07 2.042 49.125 2.176 ;
      RECT 49.056 2.045 49.07 2.178 ;
      RECT 48.97 2.045 49.056 2.18 ;
      RECT 48.93 2.042 48.97 2.183 ;
      RECT 48.906 2.038 48.93 2.185 ;
      RECT 48.82 2.028 48.906 2.188 ;
      RECT 48.79 2.017 48.82 2.189 ;
      RECT 48.771 2.013 48.79 2.188 ;
      RECT 48.685 2.006 48.771 2.185 ;
      RECT 48.625 1.995 48.685 2.182 ;
      RECT 48.605 1.987 48.625 2.18 ;
      RECT 48.57 1.982 48.605 2.179 ;
      RECT 48.545 1.977 48.57 2.178 ;
      RECT 48.515 1.972 48.545 2.177 ;
      RECT 48.49 1.915 48.515 2.176 ;
      RECT 48.475 1.915 48.49 2.2 ;
      RECT 48.28 1.915 48.29 2.2 ;
      RECT 50.055 2.935 50.06 3.075 ;
      RECT 49.715 2.935 49.75 3.073 ;
      RECT 49.29 2.92 49.305 3.065 ;
      RECT 51.12 2.7 51.21 2.96 ;
      RECT 50.95 2.565 51.05 2.96 ;
      RECT 47.985 2.54 48.065 2.75 ;
      RECT 51.075 2.677 51.12 2.96 ;
      RECT 51.065 2.647 51.075 2.96 ;
      RECT 51.05 2.57 51.065 2.96 ;
      RECT 50.865 2.565 50.95 2.925 ;
      RECT 50.86 2.567 50.865 2.92 ;
      RECT 50.855 2.572 50.86 2.92 ;
      RECT 50.82 2.672 50.855 2.92 ;
      RECT 50.81 2.7 50.82 2.92 ;
      RECT 50.8 2.715 50.81 2.92 ;
      RECT 50.79 2.727 50.8 2.92 ;
      RECT 50.785 2.737 50.79 2.92 ;
      RECT 50.77 2.747 50.785 2.922 ;
      RECT 50.765 2.762 50.77 2.924 ;
      RECT 50.75 2.775 50.765 2.926 ;
      RECT 50.745 2.79 50.75 2.929 ;
      RECT 50.725 2.8 50.745 2.933 ;
      RECT 50.71 2.81 50.725 2.936 ;
      RECT 50.675 2.817 50.71 2.941 ;
      RECT 50.631 2.824 50.675 2.949 ;
      RECT 50.545 2.836 50.631 2.962 ;
      RECT 50.52 2.847 50.545 2.973 ;
      RECT 50.49 2.852 50.52 2.978 ;
      RECT 50.455 2.857 50.49 2.986 ;
      RECT 50.425 2.862 50.455 2.993 ;
      RECT 50.4 2.867 50.425 2.998 ;
      RECT 50.335 2.874 50.4 3.007 ;
      RECT 50.265 2.887 50.335 3.023 ;
      RECT 50.235 2.897 50.265 3.035 ;
      RECT 50.21 2.902 50.235 3.042 ;
      RECT 50.155 2.909 50.21 3.05 ;
      RECT 50.15 2.916 50.155 3.055 ;
      RECT 50.145 2.918 50.15 3.056 ;
      RECT 50.13 2.92 50.145 3.058 ;
      RECT 50.125 2.92 50.13 3.061 ;
      RECT 50.06 2.927 50.125 3.068 ;
      RECT 50.025 2.937 50.055 3.078 ;
      RECT 50.008 2.94 50.025 3.08 ;
      RECT 49.922 2.939 50.008 3.079 ;
      RECT 49.836 2.937 49.922 3.076 ;
      RECT 49.75 2.936 49.836 3.074 ;
      RECT 49.649 2.934 49.715 3.073 ;
      RECT 49.563 2.931 49.649 3.071 ;
      RECT 49.477 2.927 49.563 3.069 ;
      RECT 49.391 2.924 49.477 3.068 ;
      RECT 49.305 2.921 49.391 3.066 ;
      RECT 49.205 2.92 49.29 3.063 ;
      RECT 49.155 2.918 49.205 3.061 ;
      RECT 49.135 2.915 49.155 3.059 ;
      RECT 49.115 2.913 49.135 3.056 ;
      RECT 49.09 2.909 49.115 3.053 ;
      RECT 49.045 2.903 49.09 3.048 ;
      RECT 49.005 2.897 49.045 3.04 ;
      RECT 48.98 2.892 49.005 3.033 ;
      RECT 48.925 2.885 48.98 3.025 ;
      RECT 48.901 2.878 48.925 3.018 ;
      RECT 48.815 2.869 48.901 3.008 ;
      RECT 48.785 2.861 48.815 2.998 ;
      RECT 48.755 2.857 48.785 2.993 ;
      RECT 48.75 2.854 48.755 2.99 ;
      RECT 48.745 2.853 48.75 2.99 ;
      RECT 48.67 2.846 48.745 2.983 ;
      RECT 48.631 2.837 48.67 2.972 ;
      RECT 48.545 2.827 48.631 2.96 ;
      RECT 48.505 2.817 48.545 2.948 ;
      RECT 48.466 2.812 48.505 2.941 ;
      RECT 48.38 2.802 48.466 2.93 ;
      RECT 48.34 2.79 48.38 2.919 ;
      RECT 48.305 2.775 48.34 2.912 ;
      RECT 48.295 2.765 48.305 2.909 ;
      RECT 48.275 2.75 48.295 2.907 ;
      RECT 48.245 2.72 48.275 2.903 ;
      RECT 48.235 2.7 48.245 2.898 ;
      RECT 48.23 2.692 48.235 2.895 ;
      RECT 48.225 2.685 48.23 2.893 ;
      RECT 48.21 2.672 48.225 2.886 ;
      RECT 48.205 2.662 48.21 2.878 ;
      RECT 48.2 2.655 48.205 2.873 ;
      RECT 48.195 2.65 48.2 2.869 ;
      RECT 48.18 2.637 48.195 2.861 ;
      RECT 48.175 2.547 48.18 2.85 ;
      RECT 48.17 2.542 48.175 2.843 ;
      RECT 48.095 2.54 48.17 2.803 ;
      RECT 48.065 2.54 48.095 2.758 ;
      RECT 47.97 2.545 47.985 2.745 ;
      RECT 50.455 2.25 50.715 2.51 ;
      RECT 50.44 2.238 50.62 2.475 ;
      RECT 50.435 2.239 50.62 2.473 ;
      RECT 50.42 2.243 50.63 2.463 ;
      RECT 50.415 2.248 50.635 2.433 ;
      RECT 50.42 2.245 50.635 2.463 ;
      RECT 50.435 2.24 50.63 2.473 ;
      RECT 50.455 2.237 50.62 2.51 ;
      RECT 50.455 2.236 50.61 2.51 ;
      RECT 50.48 2.235 50.61 2.51 ;
      RECT 50.04 2.48 50.3 2.74 ;
      RECT 49.915 2.525 50.3 2.735 ;
      RECT 49.905 2.53 50.3 2.73 ;
      RECT 49.92 3.47 49.935 3.78 ;
      RECT 48.515 3.24 48.525 3.37 ;
      RECT 48.295 3.235 48.4 3.37 ;
      RECT 48.21 3.24 48.26 3.37 ;
      RECT 46.76 1.975 46.765 3.08 ;
      RECT 50.015 3.562 50.02 3.698 ;
      RECT 50.01 3.557 50.015 3.758 ;
      RECT 50.005 3.555 50.01 3.771 ;
      RECT 49.99 3.552 50.005 3.773 ;
      RECT 49.985 3.547 49.99 3.775 ;
      RECT 49.98 3.543 49.985 3.778 ;
      RECT 49.965 3.538 49.98 3.78 ;
      RECT 49.935 3.53 49.965 3.78 ;
      RECT 49.896 3.47 49.92 3.78 ;
      RECT 49.81 3.47 49.896 3.777 ;
      RECT 49.78 3.47 49.81 3.77 ;
      RECT 49.755 3.47 49.78 3.763 ;
      RECT 49.73 3.47 49.755 3.755 ;
      RECT 49.715 3.47 49.73 3.748 ;
      RECT 49.69 3.47 49.715 3.74 ;
      RECT 49.675 3.47 49.69 3.733 ;
      RECT 49.635 3.48 49.675 3.722 ;
      RECT 49.625 3.475 49.635 3.712 ;
      RECT 49.621 3.474 49.625 3.709 ;
      RECT 49.535 3.466 49.621 3.692 ;
      RECT 49.502 3.455 49.535 3.669 ;
      RECT 49.416 3.444 49.502 3.647 ;
      RECT 49.33 3.428 49.416 3.616 ;
      RECT 49.26 3.413 49.33 3.588 ;
      RECT 49.25 3.406 49.26 3.575 ;
      RECT 49.22 3.403 49.25 3.565 ;
      RECT 49.195 3.399 49.22 3.558 ;
      RECT 49.18 3.396 49.195 3.553 ;
      RECT 49.175 3.395 49.18 3.548 ;
      RECT 49.145 3.39 49.175 3.541 ;
      RECT 49.14 3.385 49.145 3.536 ;
      RECT 49.125 3.382 49.14 3.531 ;
      RECT 49.12 3.377 49.125 3.526 ;
      RECT 49.1 3.372 49.12 3.523 ;
      RECT 49.085 3.367 49.1 3.515 ;
      RECT 49.07 3.361 49.085 3.51 ;
      RECT 49.04 3.352 49.07 3.503 ;
      RECT 49.035 3.345 49.04 3.495 ;
      RECT 49.03 3.343 49.035 3.493 ;
      RECT 49.025 3.342 49.03 3.49 ;
      RECT 48.985 3.335 49.025 3.483 ;
      RECT 48.971 3.325 48.985 3.473 ;
      RECT 48.92 3.314 48.971 3.461 ;
      RECT 48.895 3.3 48.92 3.447 ;
      RECT 48.87 3.289 48.895 3.439 ;
      RECT 48.85 3.278 48.87 3.433 ;
      RECT 48.84 3.272 48.85 3.428 ;
      RECT 48.835 3.27 48.84 3.424 ;
      RECT 48.815 3.265 48.835 3.419 ;
      RECT 48.785 3.255 48.815 3.409 ;
      RECT 48.78 3.247 48.785 3.402 ;
      RECT 48.765 3.245 48.78 3.398 ;
      RECT 48.745 3.245 48.765 3.393 ;
      RECT 48.74 3.244 48.745 3.391 ;
      RECT 48.735 3.244 48.74 3.388 ;
      RECT 48.695 3.243 48.735 3.383 ;
      RECT 48.67 3.242 48.695 3.378 ;
      RECT 48.61 3.241 48.67 3.375 ;
      RECT 48.525 3.24 48.61 3.373 ;
      RECT 48.486 3.239 48.515 3.37 ;
      RECT 48.4 3.237 48.486 3.37 ;
      RECT 48.26 3.237 48.295 3.37 ;
      RECT 48.17 3.241 48.21 3.373 ;
      RECT 48.155 3.244 48.17 3.38 ;
      RECT 48.145 3.245 48.155 3.387 ;
      RECT 48.12 3.248 48.145 3.392 ;
      RECT 48.115 3.25 48.12 3.395 ;
      RECT 48.065 3.252 48.115 3.396 ;
      RECT 48.026 3.256 48.065 3.398 ;
      RECT 47.94 3.258 48.026 3.401 ;
      RECT 47.922 3.26 47.94 3.403 ;
      RECT 47.836 3.263 47.922 3.405 ;
      RECT 47.75 3.267 47.836 3.408 ;
      RECT 47.713 3.271 47.75 3.411 ;
      RECT 47.627 3.274 47.713 3.414 ;
      RECT 47.541 3.278 47.627 3.417 ;
      RECT 47.455 3.283 47.541 3.421 ;
      RECT 47.435 3.285 47.455 3.424 ;
      RECT 47.415 3.284 47.435 3.425 ;
      RECT 47.366 3.281 47.415 3.426 ;
      RECT 47.28 3.276 47.366 3.429 ;
      RECT 47.23 3.271 47.28 3.431 ;
      RECT 47.206 3.269 47.23 3.432 ;
      RECT 47.12 3.264 47.206 3.434 ;
      RECT 47.095 3.26 47.12 3.433 ;
      RECT 47.085 3.257 47.095 3.431 ;
      RECT 47.075 3.25 47.085 3.428 ;
      RECT 47.07 3.23 47.075 3.423 ;
      RECT 47.06 3.2 47.07 3.418 ;
      RECT 47.045 3.07 47.06 3.409 ;
      RECT 47.04 3.062 47.045 3.402 ;
      RECT 47.02 3.055 47.04 3.394 ;
      RECT 47.015 3.037 47.02 3.386 ;
      RECT 47.005 3.017 47.015 3.381 ;
      RECT 47 2.99 47.005 3.377 ;
      RECT 46.995 2.967 47 3.374 ;
      RECT 46.975 2.925 46.995 3.366 ;
      RECT 46.94 2.84 46.975 3.35 ;
      RECT 46.935 2.772 46.94 3.338 ;
      RECT 46.92 2.742 46.935 3.332 ;
      RECT 46.915 1.987 46.92 2.233 ;
      RECT 46.905 2.712 46.92 3.323 ;
      RECT 46.91 1.982 46.915 2.265 ;
      RECT 46.905 1.977 46.91 2.308 ;
      RECT 46.9 1.975 46.905 2.343 ;
      RECT 46.885 2.675 46.905 3.313 ;
      RECT 46.895 1.975 46.9 2.38 ;
      RECT 46.88 1.975 46.895 2.478 ;
      RECT 46.88 2.648 46.885 3.306 ;
      RECT 46.875 1.975 46.88 2.553 ;
      RECT 46.875 2.636 46.88 3.303 ;
      RECT 46.87 1.975 46.875 2.585 ;
      RECT 46.87 2.615 46.875 3.3 ;
      RECT 46.865 1.975 46.87 3.297 ;
      RECT 46.83 1.975 46.865 3.283 ;
      RECT 46.815 1.975 46.83 3.265 ;
      RECT 46.795 1.975 46.815 3.255 ;
      RECT 46.77 1.975 46.795 3.238 ;
      RECT 46.765 1.975 46.77 3.188 ;
      RECT 46.755 1.975 46.76 3.018 ;
      RECT 46.75 1.975 46.755 2.925 ;
      RECT 46.745 1.975 46.75 2.838 ;
      RECT 46.74 1.975 46.745 2.77 ;
      RECT 46.735 1.975 46.74 2.713 ;
      RECT 46.725 1.975 46.735 2.608 ;
      RECT 46.72 1.975 46.725 2.48 ;
      RECT 46.715 1.975 46.72 2.398 ;
      RECT 46.71 1.977 46.715 2.315 ;
      RECT 46.705 1.982 46.71 2.248 ;
      RECT 46.7 1.987 46.705 2.175 ;
      RECT 49.515 2.305 49.775 2.565 ;
      RECT 49.535 2.272 49.745 2.565 ;
      RECT 49.535 2.27 49.735 2.565 ;
      RECT 49.545 2.257 49.735 2.565 ;
      RECT 49.545 2.255 49.66 2.565 ;
      RECT 49.02 2.38 49.195 2.66 ;
      RECT 49.015 2.38 49.195 2.658 ;
      RECT 49.015 2.38 49.21 2.655 ;
      RECT 49.005 2.38 49.21 2.653 ;
      RECT 48.95 2.38 49.21 2.64 ;
      RECT 48.95 2.455 49.215 2.618 ;
      RECT 48.495 2.392 48.515 2.635 ;
      RECT 48.495 2.392 48.555 2.634 ;
      RECT 48.49 2.394 48.555 2.633 ;
      RECT 48.49 2.394 48.641 2.632 ;
      RECT 48.49 2.394 48.71 2.631 ;
      RECT 48.49 2.394 48.73 2.623 ;
      RECT 48.47 2.397 48.73 2.621 ;
      RECT 48.455 2.407 48.73 2.606 ;
      RECT 48.455 2.407 48.745 2.605 ;
      RECT 48.45 2.416 48.745 2.597 ;
      RECT 48.45 2.416 48.75 2.593 ;
      RECT 48.555 2.33 48.815 2.59 ;
      RECT 48.445 2.418 48.815 2.475 ;
      RECT 48.515 2.385 48.815 2.59 ;
      RECT 48.48 3.578 48.485 3.785 ;
      RECT 48.43 3.572 48.48 3.784 ;
      RECT 48.397 3.586 48.49 3.783 ;
      RECT 48.311 3.586 48.49 3.782 ;
      RECT 48.225 3.586 48.49 3.781 ;
      RECT 48.225 3.685 48.495 3.778 ;
      RECT 48.22 3.685 48.495 3.773 ;
      RECT 48.215 3.685 48.495 3.755 ;
      RECT 48.21 3.685 48.495 3.738 ;
      RECT 48.17 3.47 48.43 3.73 ;
      RECT 47.63 2.62 47.716 3.034 ;
      RECT 47.63 2.62 47.755 3.031 ;
      RECT 47.63 2.62 47.775 3.021 ;
      RECT 47.585 2.62 47.775 3.018 ;
      RECT 47.585 2.772 47.785 3.008 ;
      RECT 47.585 2.793 47.79 3.002 ;
      RECT 47.585 2.811 47.795 2.998 ;
      RECT 47.585 2.831 47.805 2.993 ;
      RECT 47.56 2.831 47.805 2.99 ;
      RECT 47.55 2.831 47.805 2.968 ;
      RECT 47.55 2.847 47.81 2.938 ;
      RECT 47.515 2.62 47.775 2.925 ;
      RECT 47.515 2.859 47.815 2.88 ;
      RECT 45.18 7.765 45.47 7.995 ;
      RECT 45.24 6.285 45.41 7.995 ;
      RECT 45.185 6.655 45.535 7.005 ;
      RECT 45.18 6.285 45.47 6.515 ;
      RECT 45.18 2.365 45.47 2.595 ;
      RECT 45.24 0.885 45.41 2.595 ;
      RECT 45.18 0.885 45.47 1.115 ;
      RECT 44.77 2.735 45.1 2.965 ;
      RECT 44.77 2.765 45.27 2.935 ;
      RECT 44.77 2.395 44.96 2.965 ;
      RECT 44.19 2.365 44.48 2.595 ;
      RECT 44.19 2.395 44.96 2.565 ;
      RECT 44.25 0.885 44.42 2.595 ;
      RECT 44.19 0.885 44.48 1.115 ;
      RECT 44.19 7.765 44.48 7.995 ;
      RECT 44.25 6.285 44.42 7.995 ;
      RECT 44.19 6.285 44.48 6.515 ;
      RECT 44.19 6.325 45.04 6.485 ;
      RECT 44.87 5.915 45.04 6.485 ;
      RECT 44.19 6.32 44.58 6.485 ;
      RECT 44.81 5.915 45.1 6.145 ;
      RECT 44.81 5.945 45.27 6.115 ;
      RECT 43.82 2.735 44.11 2.965 ;
      RECT 43.82 2.765 44.28 2.935 ;
      RECT 43.88 1.655 44.045 2.965 ;
      RECT 42.395 1.625 42.685 1.855 ;
      RECT 42.395 1.655 44.045 1.825 ;
      RECT 42.455 0.885 42.625 1.855 ;
      RECT 42.395 0.885 42.685 1.115 ;
      RECT 42.395 7.765 42.685 7.995 ;
      RECT 42.455 7.025 42.625 7.995 ;
      RECT 42.455 7.12 44.045 7.29 ;
      RECT 43.875 5.915 44.045 7.29 ;
      RECT 42.395 7.025 42.685 7.255 ;
      RECT 43.82 5.915 44.11 6.145 ;
      RECT 43.82 5.945 44.28 6.115 ;
      RECT 40.445 2.705 40.785 3.055 ;
      RECT 40.535 2.025 40.705 3.055 ;
      RECT 42.825 1.965 43.175 2.315 ;
      RECT 40.535 2.025 43.175 2.195 ;
      RECT 42.85 6.655 43.175 6.98 ;
      RECT 37.39 6.615 37.74 6.965 ;
      RECT 42.825 6.655 43.175 6.885 ;
      RECT 37.19 6.655 37.74 6.885 ;
      RECT 37.02 6.685 43.175 6.855 ;
      RECT 42.05 2.365 42.37 2.685 ;
      RECT 42.02 2.365 42.37 2.595 ;
      RECT 41.85 2.395 42.37 2.565 ;
      RECT 42.05 6.255 42.37 6.545 ;
      RECT 42.02 6.285 42.37 6.515 ;
      RECT 41.85 6.315 42.37 6.485 ;
      RECT 41.005 2.705 41.345 3.055 ;
      RECT 41.005 2.765 41.485 2.935 ;
      RECT 41 5.86 41.34 6.21 ;
      RECT 35.39 5.915 35.68 6.145 ;
      RECT 35.39 5.945 41.485 6.115 ;
      RECT 37.74 2.985 37.89 3.26 ;
      RECT 38.28 2.065 38.285 2.285 ;
      RECT 39.43 2.265 39.445 2.463 ;
      RECT 39.395 2.257 39.43 2.47 ;
      RECT 39.365 2.25 39.395 2.47 ;
      RECT 39.31 2.215 39.365 2.47 ;
      RECT 39.245 2.152 39.31 2.47 ;
      RECT 39.24 2.117 39.245 2.468 ;
      RECT 39.235 2.112 39.24 2.46 ;
      RECT 39.23 2.107 39.235 2.446 ;
      RECT 39.225 2.104 39.23 2.439 ;
      RECT 39.18 2.094 39.225 2.39 ;
      RECT 39.16 2.081 39.18 2.325 ;
      RECT 39.155 2.076 39.16 2.298 ;
      RECT 39.15 2.075 39.155 2.291 ;
      RECT 39.145 2.074 39.15 2.284 ;
      RECT 39.06 2.059 39.145 2.23 ;
      RECT 39.03 2.04 39.06 2.18 ;
      RECT 38.95 2.023 39.03 2.165 ;
      RECT 38.915 2.01 38.95 2.15 ;
      RECT 38.907 2.01 38.915 2.145 ;
      RECT 38.821 2.011 38.907 2.145 ;
      RECT 38.735 2.013 38.821 2.145 ;
      RECT 38.71 2.014 38.735 2.149 ;
      RECT 38.635 2.02 38.71 2.164 ;
      RECT 38.552 2.032 38.635 2.188 ;
      RECT 38.466 2.045 38.552 2.214 ;
      RECT 38.38 2.058 38.466 2.24 ;
      RECT 38.345 2.067 38.38 2.259 ;
      RECT 38.295 2.067 38.345 2.272 ;
      RECT 38.285 2.065 38.295 2.283 ;
      RECT 38.27 2.062 38.28 2.285 ;
      RECT 38.255 2.054 38.27 2.293 ;
      RECT 38.24 2.046 38.255 2.313 ;
      RECT 38.235 2.041 38.24 2.37 ;
      RECT 38.22 2.036 38.235 2.443 ;
      RECT 38.215 2.031 38.22 2.485 ;
      RECT 38.21 2.029 38.215 2.513 ;
      RECT 38.205 2.027 38.21 2.535 ;
      RECT 38.195 2.023 38.205 2.578 ;
      RECT 38.19 2.02 38.195 2.603 ;
      RECT 38.185 2.018 38.19 2.623 ;
      RECT 38.18 2.016 38.185 2.647 ;
      RECT 38.175 2.012 38.18 2.67 ;
      RECT 38.17 2.008 38.175 2.693 ;
      RECT 38.135 1.998 38.17 2.8 ;
      RECT 38.13 1.988 38.135 2.898 ;
      RECT 38.125 1.986 38.13 2.925 ;
      RECT 38.12 1.985 38.125 2.945 ;
      RECT 38.115 1.977 38.12 2.965 ;
      RECT 38.11 1.972 38.115 3 ;
      RECT 38.105 1.97 38.11 3.018 ;
      RECT 38.1 1.97 38.105 3.043 ;
      RECT 38.095 1.97 38.1 3.065 ;
      RECT 38.06 1.97 38.095 3.108 ;
      RECT 38.035 1.97 38.06 3.137 ;
      RECT 38.025 1.97 38.035 2.323 ;
      RECT 38.028 2.38 38.035 3.147 ;
      RECT 38.025 2.437 38.028 3.15 ;
      RECT 38.02 1.97 38.025 2.295 ;
      RECT 38.02 2.487 38.025 3.153 ;
      RECT 38.01 1.97 38.02 2.285 ;
      RECT 38.015 2.54 38.02 3.156 ;
      RECT 38.01 2.625 38.015 3.16 ;
      RECT 38 1.97 38.01 2.273 ;
      RECT 38.005 2.672 38.01 3.164 ;
      RECT 38 2.747 38.005 3.168 ;
      RECT 37.965 1.97 38 2.248 ;
      RECT 37.99 2.83 38 3.173 ;
      RECT 37.98 2.897 37.99 3.18 ;
      RECT 37.975 2.925 37.98 3.185 ;
      RECT 37.965 2.938 37.975 3.191 ;
      RECT 37.92 1.97 37.965 2.205 ;
      RECT 37.96 2.943 37.965 3.198 ;
      RECT 37.92 2.96 37.96 3.26 ;
      RECT 37.915 1.972 37.92 2.178 ;
      RECT 37.89 2.98 37.92 3.26 ;
      RECT 37.91 1.977 37.915 2.15 ;
      RECT 37.7 2.989 37.74 3.26 ;
      RECT 37.675 2.997 37.7 3.23 ;
      RECT 37.63 3.005 37.675 3.23 ;
      RECT 37.615 3.01 37.63 3.225 ;
      RECT 37.605 3.01 37.615 3.219 ;
      RECT 37.595 3.017 37.605 3.216 ;
      RECT 37.59 3.055 37.595 3.205 ;
      RECT 37.585 3.117 37.59 3.183 ;
      RECT 38.855 2.992 39.04 3.215 ;
      RECT 38.855 3.007 39.045 3.211 ;
      RECT 38.845 2.28 38.93 3.21 ;
      RECT 38.845 3.007 39.05 3.204 ;
      RECT 38.84 3.015 39.05 3.203 ;
      RECT 39.045 2.735 39.365 3.055 ;
      RECT 38.84 2.907 39.01 2.998 ;
      RECT 38.835 2.907 39.01 2.98 ;
      RECT 38.825 2.715 38.96 2.955 ;
      RECT 38.82 2.715 38.96 2.9 ;
      RECT 38.78 2.295 38.95 2.8 ;
      RECT 38.765 2.295 38.95 2.67 ;
      RECT 38.76 2.295 38.95 2.623 ;
      RECT 38.755 2.295 38.95 2.603 ;
      RECT 38.75 2.295 38.95 2.578 ;
      RECT 38.72 2.295 38.98 2.555 ;
      RECT 38.73 2.292 38.94 2.555 ;
      RECT 38.855 2.287 38.94 3.215 ;
      RECT 38.74 2.28 38.93 2.555 ;
      RECT 38.735 2.285 38.93 2.555 ;
      RECT 37.565 2.497 37.75 2.71 ;
      RECT 37.565 2.505 37.76 2.703 ;
      RECT 37.545 2.505 37.76 2.7 ;
      RECT 37.54 2.505 37.76 2.685 ;
      RECT 37.47 2.42 37.73 2.68 ;
      RECT 37.47 2.565 37.765 2.593 ;
      RECT 37.125 3.02 37.385 3.28 ;
      RECT 37.15 2.965 37.345 3.28 ;
      RECT 37.145 2.714 37.325 3.008 ;
      RECT 37.145 2.72 37.335 3.008 ;
      RECT 37.125 2.722 37.335 2.953 ;
      RECT 37.12 2.732 37.335 2.82 ;
      RECT 37.15 2.712 37.325 3.28 ;
      RECT 37.236 2.71 37.325 3.28 ;
      RECT 37.095 1.93 37.13 2.3 ;
      RECT 36.885 2.04 36.89 2.3 ;
      RECT 37.13 1.937 37.145 2.3 ;
      RECT 37.02 1.93 37.095 2.378 ;
      RECT 37.01 1.93 37.02 2.463 ;
      RECT 36.985 1.93 37.01 2.498 ;
      RECT 36.945 1.93 36.985 2.566 ;
      RECT 36.935 1.937 36.945 2.618 ;
      RECT 36.905 2.04 36.935 2.659 ;
      RECT 36.9 2.04 36.905 2.698 ;
      RECT 36.89 2.04 36.9 2.718 ;
      RECT 36.885 2.335 36.89 2.755 ;
      RECT 36.88 2.352 36.885 2.775 ;
      RECT 36.865 2.415 36.88 2.815 ;
      RECT 36.86 2.458 36.865 2.85 ;
      RECT 36.855 2.466 36.86 2.863 ;
      RECT 36.845 2.48 36.855 2.885 ;
      RECT 36.82 2.515 36.845 2.95 ;
      RECT 36.81 2.55 36.82 3.013 ;
      RECT 36.79 2.58 36.81 3.074 ;
      RECT 36.775 2.616 36.79 3.141 ;
      RECT 36.765 2.644 36.775 3.18 ;
      RECT 36.755 2.666 36.765 3.2 ;
      RECT 36.75 2.676 36.755 3.211 ;
      RECT 36.745 2.685 36.75 3.214 ;
      RECT 36.735 2.703 36.745 3.218 ;
      RECT 36.725 2.721 36.735 3.219 ;
      RECT 36.7 2.76 36.725 3.216 ;
      RECT 36.68 2.802 36.7 3.213 ;
      RECT 36.665 2.84 36.68 3.212 ;
      RECT 36.63 2.875 36.665 3.209 ;
      RECT 36.625 2.897 36.63 3.207 ;
      RECT 36.56 2.937 36.625 3.204 ;
      RECT 36.555 2.977 36.56 3.2 ;
      RECT 36.54 2.987 36.555 3.191 ;
      RECT 36.53 3.107 36.54 3.176 ;
      RECT 37.01 3.52 37.02 3.78 ;
      RECT 37.01 3.523 37.03 3.779 ;
      RECT 37 3.513 37.01 3.778 ;
      RECT 36.99 3.528 37.07 3.774 ;
      RECT 36.975 3.507 36.99 3.772 ;
      RECT 36.95 3.532 37.075 3.768 ;
      RECT 36.935 3.492 36.95 3.763 ;
      RECT 36.935 3.534 37.085 3.762 ;
      RECT 36.935 3.542 37.1 3.755 ;
      RECT 36.875 3.479 36.935 3.745 ;
      RECT 36.865 3.466 36.875 3.727 ;
      RECT 36.84 3.456 36.865 3.717 ;
      RECT 36.835 3.446 36.84 3.709 ;
      RECT 36.77 3.542 37.1 3.691 ;
      RECT 36.685 3.542 37.1 3.653 ;
      RECT 36.575 3.37 36.835 3.63 ;
      RECT 36.95 3.5 36.975 3.768 ;
      RECT 36.99 3.51 37 3.774 ;
      RECT 36.575 3.518 37.015 3.63 ;
      RECT 36.76 7.765 37.05 7.995 ;
      RECT 36.82 7.025 36.99 7.995 ;
      RECT 36.72 7.055 37.09 7.425 ;
      RECT 36.76 7.025 37.05 7.425 ;
      RECT 35.79 3.275 35.82 3.575 ;
      RECT 35.565 3.26 35.57 3.535 ;
      RECT 35.365 3.26 35.52 3.52 ;
      RECT 36.665 1.975 36.695 2.235 ;
      RECT 36.655 1.975 36.665 2.343 ;
      RECT 36.635 1.975 36.655 2.353 ;
      RECT 36.62 1.975 36.635 2.365 ;
      RECT 36.565 1.975 36.62 2.415 ;
      RECT 36.55 1.975 36.565 2.463 ;
      RECT 36.52 1.975 36.55 2.498 ;
      RECT 36.465 1.975 36.52 2.56 ;
      RECT 36.445 1.975 36.465 2.628 ;
      RECT 36.44 1.975 36.445 2.658 ;
      RECT 36.435 1.975 36.44 2.67 ;
      RECT 36.43 2.092 36.435 2.688 ;
      RECT 36.41 2.11 36.43 2.713 ;
      RECT 36.39 2.137 36.41 2.763 ;
      RECT 36.385 2.157 36.39 2.794 ;
      RECT 36.38 2.165 36.385 2.811 ;
      RECT 36.365 2.191 36.38 2.84 ;
      RECT 36.35 2.233 36.365 2.875 ;
      RECT 36.345 2.262 36.35 2.898 ;
      RECT 36.34 2.277 36.345 2.911 ;
      RECT 36.335 2.3 36.34 2.922 ;
      RECT 36.325 2.32 36.335 2.94 ;
      RECT 36.315 2.35 36.325 2.963 ;
      RECT 36.31 2.372 36.315 2.983 ;
      RECT 36.305 2.387 36.31 2.998 ;
      RECT 36.29 2.417 36.305 3.025 ;
      RECT 36.285 2.447 36.29 3.051 ;
      RECT 36.28 2.465 36.285 3.063 ;
      RECT 36.27 2.495 36.28 3.082 ;
      RECT 36.26 2.52 36.27 3.107 ;
      RECT 36.255 2.54 36.26 3.126 ;
      RECT 36.25 2.557 36.255 3.139 ;
      RECT 36.24 2.583 36.25 3.158 ;
      RECT 36.23 2.621 36.24 3.185 ;
      RECT 36.225 2.647 36.23 3.205 ;
      RECT 36.22 2.657 36.225 3.215 ;
      RECT 36.215 2.67 36.22 3.23 ;
      RECT 36.21 2.685 36.215 3.24 ;
      RECT 36.205 2.707 36.21 3.255 ;
      RECT 36.2 2.725 36.205 3.266 ;
      RECT 36.195 2.735 36.2 3.277 ;
      RECT 36.19 2.743 36.195 3.289 ;
      RECT 36.185 2.751 36.19 3.3 ;
      RECT 36.18 2.777 36.185 3.313 ;
      RECT 36.17 2.805 36.18 3.326 ;
      RECT 36.165 2.835 36.17 3.335 ;
      RECT 36.16 2.85 36.165 3.342 ;
      RECT 36.145 2.875 36.16 3.349 ;
      RECT 36.14 2.897 36.145 3.355 ;
      RECT 36.135 2.922 36.14 3.358 ;
      RECT 36.126 2.95 36.135 3.362 ;
      RECT 36.12 2.967 36.126 3.367 ;
      RECT 36.115 2.985 36.12 3.371 ;
      RECT 36.11 2.997 36.115 3.374 ;
      RECT 36.105 3.018 36.11 3.378 ;
      RECT 36.1 3.036 36.105 3.381 ;
      RECT 36.095 3.05 36.1 3.384 ;
      RECT 36.09 3.067 36.095 3.387 ;
      RECT 36.085 3.08 36.09 3.39 ;
      RECT 36.06 3.117 36.085 3.398 ;
      RECT 36.055 3.162 36.06 3.407 ;
      RECT 36.05 3.19 36.055 3.41 ;
      RECT 36.04 3.21 36.05 3.414 ;
      RECT 36.035 3.23 36.04 3.419 ;
      RECT 36.03 3.245 36.035 3.422 ;
      RECT 36.01 3.255 36.03 3.429 ;
      RECT 35.945 3.262 36.01 3.455 ;
      RECT 35.91 3.265 35.945 3.483 ;
      RECT 35.895 3.268 35.91 3.498 ;
      RECT 35.885 3.269 35.895 3.513 ;
      RECT 35.875 3.27 35.885 3.53 ;
      RECT 35.87 3.27 35.875 3.545 ;
      RECT 35.865 3.27 35.87 3.553 ;
      RECT 35.85 3.271 35.865 3.568 ;
      RECT 35.82 3.273 35.85 3.575 ;
      RECT 35.71 3.28 35.79 3.575 ;
      RECT 35.665 3.285 35.71 3.575 ;
      RECT 35.655 3.286 35.665 3.565 ;
      RECT 35.645 3.287 35.655 3.558 ;
      RECT 35.625 3.289 35.645 3.553 ;
      RECT 35.615 3.26 35.625 3.548 ;
      RECT 35.57 3.26 35.615 3.54 ;
      RECT 35.54 3.26 35.565 3.53 ;
      RECT 35.52 3.26 35.54 3.523 ;
      RECT 35.8 2.06 36.06 2.32 ;
      RECT 35.68 2.075 35.69 2.24 ;
      RECT 35.665 2.075 35.67 2.235 ;
      RECT 33.03 1.915 33.215 2.205 ;
      RECT 34.845 2.04 34.86 2.195 ;
      RECT 32.995 1.915 33.02 2.175 ;
      RECT 35.41 1.965 35.415 2.107 ;
      RECT 35.325 1.96 35.35 2.1 ;
      RECT 35.725 2.077 35.8 2.27 ;
      RECT 35.71 2.075 35.725 2.253 ;
      RECT 35.69 2.075 35.71 2.245 ;
      RECT 35.67 2.075 35.68 2.238 ;
      RECT 35.625 2.07 35.665 2.228 ;
      RECT 35.585 2.045 35.625 2.213 ;
      RECT 35.57 2.02 35.585 2.203 ;
      RECT 35.565 2.014 35.57 2.201 ;
      RECT 35.53 2.006 35.565 2.184 ;
      RECT 35.525 1.999 35.53 2.172 ;
      RECT 35.505 1.994 35.525 2.16 ;
      RECT 35.495 1.988 35.505 2.145 ;
      RECT 35.475 1.983 35.495 2.13 ;
      RECT 35.465 1.978 35.475 2.123 ;
      RECT 35.46 1.976 35.465 2.118 ;
      RECT 35.455 1.975 35.46 2.115 ;
      RECT 35.415 1.97 35.455 2.111 ;
      RECT 35.395 1.964 35.41 2.106 ;
      RECT 35.36 1.961 35.395 2.103 ;
      RECT 35.35 1.96 35.36 2.101 ;
      RECT 35.29 1.96 35.325 2.098 ;
      RECT 35.245 1.96 35.29 2.098 ;
      RECT 35.195 1.96 35.245 2.101 ;
      RECT 35.18 1.962 35.195 2.103 ;
      RECT 35.165 1.965 35.18 2.104 ;
      RECT 35.155 1.97 35.165 2.105 ;
      RECT 35.125 1.975 35.155 2.11 ;
      RECT 35.115 1.981 35.125 2.118 ;
      RECT 35.105 1.983 35.115 2.122 ;
      RECT 35.095 1.987 35.105 2.126 ;
      RECT 35.07 1.993 35.095 2.134 ;
      RECT 35.06 1.998 35.07 2.142 ;
      RECT 35.045 2.002 35.06 2.146 ;
      RECT 35.01 2.008 35.045 2.154 ;
      RECT 34.99 2.013 35.01 2.164 ;
      RECT 34.96 2.02 34.99 2.173 ;
      RECT 34.915 2.029 34.96 2.187 ;
      RECT 34.91 2.034 34.915 2.198 ;
      RECT 34.89 2.037 34.91 2.199 ;
      RECT 34.86 2.04 34.89 2.197 ;
      RECT 34.825 2.04 34.845 2.193 ;
      RECT 34.755 2.04 34.825 2.184 ;
      RECT 34.74 2.037 34.755 2.176 ;
      RECT 34.7 2.03 34.74 2.171 ;
      RECT 34.675 2.02 34.7 2.164 ;
      RECT 34.67 2.014 34.675 2.161 ;
      RECT 34.63 2.008 34.67 2.158 ;
      RECT 34.615 2.001 34.63 2.153 ;
      RECT 34.595 1.997 34.615 2.148 ;
      RECT 34.58 1.992 34.595 2.144 ;
      RECT 34.565 1.987 34.58 2.142 ;
      RECT 34.55 1.983 34.565 2.141 ;
      RECT 34.535 1.981 34.55 2.137 ;
      RECT 34.525 1.979 34.535 2.132 ;
      RECT 34.51 1.976 34.525 2.128 ;
      RECT 34.5 1.974 34.51 2.123 ;
      RECT 34.48 1.971 34.5 2.119 ;
      RECT 34.435 1.97 34.48 2.117 ;
      RECT 34.375 1.972 34.435 2.118 ;
      RECT 34.355 1.974 34.375 2.12 ;
      RECT 34.325 1.977 34.355 2.121 ;
      RECT 34.275 1.982 34.325 2.123 ;
      RECT 34.27 1.985 34.275 2.125 ;
      RECT 34.26 1.987 34.27 2.128 ;
      RECT 34.255 1.989 34.26 2.131 ;
      RECT 34.205 1.992 34.255 2.138 ;
      RECT 34.185 1.996 34.205 2.15 ;
      RECT 34.175 1.999 34.185 2.156 ;
      RECT 34.165 2 34.175 2.159 ;
      RECT 34.126 2.003 34.165 2.161 ;
      RECT 34.04 2.01 34.126 2.164 ;
      RECT 33.966 2.02 34.04 2.168 ;
      RECT 33.88 2.031 33.966 2.173 ;
      RECT 33.865 2.038 33.88 2.175 ;
      RECT 33.81 2.042 33.865 2.176 ;
      RECT 33.796 2.045 33.81 2.178 ;
      RECT 33.71 2.045 33.796 2.18 ;
      RECT 33.67 2.042 33.71 2.183 ;
      RECT 33.646 2.038 33.67 2.185 ;
      RECT 33.56 2.028 33.646 2.188 ;
      RECT 33.53 2.017 33.56 2.189 ;
      RECT 33.511 2.013 33.53 2.188 ;
      RECT 33.425 2.006 33.511 2.185 ;
      RECT 33.365 1.995 33.425 2.182 ;
      RECT 33.345 1.987 33.365 2.18 ;
      RECT 33.31 1.982 33.345 2.179 ;
      RECT 33.285 1.977 33.31 2.178 ;
      RECT 33.255 1.972 33.285 2.177 ;
      RECT 33.23 1.915 33.255 2.176 ;
      RECT 33.215 1.915 33.23 2.2 ;
      RECT 33.02 1.915 33.03 2.2 ;
      RECT 34.795 2.935 34.8 3.075 ;
      RECT 34.455 2.935 34.49 3.073 ;
      RECT 34.03 2.92 34.045 3.065 ;
      RECT 35.86 2.7 35.95 2.96 ;
      RECT 35.69 2.565 35.79 2.96 ;
      RECT 32.725 2.54 32.805 2.75 ;
      RECT 35.815 2.677 35.86 2.96 ;
      RECT 35.805 2.647 35.815 2.96 ;
      RECT 35.79 2.57 35.805 2.96 ;
      RECT 35.605 2.565 35.69 2.925 ;
      RECT 35.6 2.567 35.605 2.92 ;
      RECT 35.595 2.572 35.6 2.92 ;
      RECT 35.56 2.672 35.595 2.92 ;
      RECT 35.55 2.7 35.56 2.92 ;
      RECT 35.54 2.715 35.55 2.92 ;
      RECT 35.53 2.727 35.54 2.92 ;
      RECT 35.525 2.737 35.53 2.92 ;
      RECT 35.51 2.747 35.525 2.922 ;
      RECT 35.505 2.762 35.51 2.924 ;
      RECT 35.49 2.775 35.505 2.926 ;
      RECT 35.485 2.79 35.49 2.929 ;
      RECT 35.465 2.8 35.485 2.933 ;
      RECT 35.45 2.81 35.465 2.936 ;
      RECT 35.415 2.817 35.45 2.941 ;
      RECT 35.371 2.824 35.415 2.949 ;
      RECT 35.285 2.836 35.371 2.962 ;
      RECT 35.26 2.847 35.285 2.973 ;
      RECT 35.23 2.852 35.26 2.978 ;
      RECT 35.195 2.857 35.23 2.986 ;
      RECT 35.165 2.862 35.195 2.993 ;
      RECT 35.14 2.867 35.165 2.998 ;
      RECT 35.075 2.874 35.14 3.007 ;
      RECT 35.005 2.887 35.075 3.023 ;
      RECT 34.975 2.897 35.005 3.035 ;
      RECT 34.95 2.902 34.975 3.042 ;
      RECT 34.895 2.909 34.95 3.05 ;
      RECT 34.89 2.916 34.895 3.055 ;
      RECT 34.885 2.918 34.89 3.056 ;
      RECT 34.87 2.92 34.885 3.058 ;
      RECT 34.865 2.92 34.87 3.061 ;
      RECT 34.8 2.927 34.865 3.068 ;
      RECT 34.765 2.937 34.795 3.078 ;
      RECT 34.748 2.94 34.765 3.08 ;
      RECT 34.662 2.939 34.748 3.079 ;
      RECT 34.576 2.937 34.662 3.076 ;
      RECT 34.49 2.936 34.576 3.074 ;
      RECT 34.389 2.934 34.455 3.073 ;
      RECT 34.303 2.931 34.389 3.071 ;
      RECT 34.217 2.927 34.303 3.069 ;
      RECT 34.131 2.924 34.217 3.068 ;
      RECT 34.045 2.921 34.131 3.066 ;
      RECT 33.945 2.92 34.03 3.063 ;
      RECT 33.895 2.918 33.945 3.061 ;
      RECT 33.875 2.915 33.895 3.059 ;
      RECT 33.855 2.913 33.875 3.056 ;
      RECT 33.83 2.909 33.855 3.053 ;
      RECT 33.785 2.903 33.83 3.048 ;
      RECT 33.745 2.897 33.785 3.04 ;
      RECT 33.72 2.892 33.745 3.033 ;
      RECT 33.665 2.885 33.72 3.025 ;
      RECT 33.641 2.878 33.665 3.018 ;
      RECT 33.555 2.869 33.641 3.008 ;
      RECT 33.525 2.861 33.555 2.998 ;
      RECT 33.495 2.857 33.525 2.993 ;
      RECT 33.49 2.854 33.495 2.99 ;
      RECT 33.485 2.853 33.49 2.99 ;
      RECT 33.41 2.846 33.485 2.983 ;
      RECT 33.371 2.837 33.41 2.972 ;
      RECT 33.285 2.827 33.371 2.96 ;
      RECT 33.245 2.817 33.285 2.948 ;
      RECT 33.206 2.812 33.245 2.941 ;
      RECT 33.12 2.802 33.206 2.93 ;
      RECT 33.08 2.79 33.12 2.919 ;
      RECT 33.045 2.775 33.08 2.912 ;
      RECT 33.035 2.765 33.045 2.909 ;
      RECT 33.015 2.75 33.035 2.907 ;
      RECT 32.985 2.72 33.015 2.903 ;
      RECT 32.975 2.7 32.985 2.898 ;
      RECT 32.97 2.692 32.975 2.895 ;
      RECT 32.965 2.685 32.97 2.893 ;
      RECT 32.95 2.672 32.965 2.886 ;
      RECT 32.945 2.662 32.95 2.878 ;
      RECT 32.94 2.655 32.945 2.873 ;
      RECT 32.935 2.65 32.94 2.869 ;
      RECT 32.92 2.637 32.935 2.861 ;
      RECT 32.915 2.547 32.92 2.85 ;
      RECT 32.91 2.542 32.915 2.843 ;
      RECT 32.835 2.54 32.91 2.803 ;
      RECT 32.805 2.54 32.835 2.758 ;
      RECT 32.71 2.545 32.725 2.745 ;
      RECT 35.195 2.25 35.455 2.51 ;
      RECT 35.18 2.238 35.36 2.475 ;
      RECT 35.175 2.239 35.36 2.473 ;
      RECT 35.16 2.243 35.37 2.463 ;
      RECT 35.155 2.248 35.375 2.433 ;
      RECT 35.16 2.245 35.375 2.463 ;
      RECT 35.175 2.24 35.37 2.473 ;
      RECT 35.195 2.237 35.36 2.51 ;
      RECT 35.195 2.236 35.35 2.51 ;
      RECT 35.22 2.235 35.35 2.51 ;
      RECT 34.78 2.48 35.04 2.74 ;
      RECT 34.655 2.525 35.04 2.735 ;
      RECT 34.645 2.53 35.04 2.73 ;
      RECT 34.66 3.47 34.675 3.78 ;
      RECT 33.255 3.24 33.265 3.37 ;
      RECT 33.035 3.235 33.14 3.37 ;
      RECT 32.95 3.24 33 3.37 ;
      RECT 31.5 1.975 31.505 3.08 ;
      RECT 34.755 3.562 34.76 3.698 ;
      RECT 34.75 3.557 34.755 3.758 ;
      RECT 34.745 3.555 34.75 3.771 ;
      RECT 34.73 3.552 34.745 3.773 ;
      RECT 34.725 3.547 34.73 3.775 ;
      RECT 34.72 3.543 34.725 3.778 ;
      RECT 34.705 3.538 34.72 3.78 ;
      RECT 34.675 3.53 34.705 3.78 ;
      RECT 34.636 3.47 34.66 3.78 ;
      RECT 34.55 3.47 34.636 3.777 ;
      RECT 34.52 3.47 34.55 3.77 ;
      RECT 34.495 3.47 34.52 3.763 ;
      RECT 34.47 3.47 34.495 3.755 ;
      RECT 34.455 3.47 34.47 3.748 ;
      RECT 34.43 3.47 34.455 3.74 ;
      RECT 34.415 3.47 34.43 3.733 ;
      RECT 34.375 3.48 34.415 3.722 ;
      RECT 34.365 3.475 34.375 3.712 ;
      RECT 34.361 3.474 34.365 3.709 ;
      RECT 34.275 3.466 34.361 3.692 ;
      RECT 34.242 3.455 34.275 3.669 ;
      RECT 34.156 3.444 34.242 3.647 ;
      RECT 34.07 3.428 34.156 3.616 ;
      RECT 34 3.413 34.07 3.588 ;
      RECT 33.99 3.406 34 3.575 ;
      RECT 33.96 3.403 33.99 3.565 ;
      RECT 33.935 3.399 33.96 3.558 ;
      RECT 33.92 3.396 33.935 3.553 ;
      RECT 33.915 3.395 33.92 3.548 ;
      RECT 33.885 3.39 33.915 3.541 ;
      RECT 33.88 3.385 33.885 3.536 ;
      RECT 33.865 3.382 33.88 3.531 ;
      RECT 33.86 3.377 33.865 3.526 ;
      RECT 33.84 3.372 33.86 3.523 ;
      RECT 33.825 3.367 33.84 3.515 ;
      RECT 33.81 3.361 33.825 3.51 ;
      RECT 33.78 3.352 33.81 3.503 ;
      RECT 33.775 3.345 33.78 3.495 ;
      RECT 33.77 3.343 33.775 3.493 ;
      RECT 33.765 3.342 33.77 3.49 ;
      RECT 33.725 3.335 33.765 3.483 ;
      RECT 33.711 3.325 33.725 3.473 ;
      RECT 33.66 3.314 33.711 3.461 ;
      RECT 33.635 3.3 33.66 3.447 ;
      RECT 33.61 3.289 33.635 3.439 ;
      RECT 33.59 3.278 33.61 3.433 ;
      RECT 33.58 3.272 33.59 3.428 ;
      RECT 33.575 3.27 33.58 3.424 ;
      RECT 33.555 3.265 33.575 3.419 ;
      RECT 33.525 3.255 33.555 3.409 ;
      RECT 33.52 3.247 33.525 3.402 ;
      RECT 33.505 3.245 33.52 3.398 ;
      RECT 33.485 3.245 33.505 3.393 ;
      RECT 33.48 3.244 33.485 3.391 ;
      RECT 33.475 3.244 33.48 3.388 ;
      RECT 33.435 3.243 33.475 3.383 ;
      RECT 33.41 3.242 33.435 3.378 ;
      RECT 33.35 3.241 33.41 3.375 ;
      RECT 33.265 3.24 33.35 3.373 ;
      RECT 33.226 3.239 33.255 3.37 ;
      RECT 33.14 3.237 33.226 3.37 ;
      RECT 33 3.237 33.035 3.37 ;
      RECT 32.91 3.241 32.95 3.373 ;
      RECT 32.895 3.244 32.91 3.38 ;
      RECT 32.885 3.245 32.895 3.387 ;
      RECT 32.86 3.248 32.885 3.392 ;
      RECT 32.855 3.25 32.86 3.395 ;
      RECT 32.805 3.252 32.855 3.396 ;
      RECT 32.766 3.256 32.805 3.398 ;
      RECT 32.68 3.258 32.766 3.401 ;
      RECT 32.662 3.26 32.68 3.403 ;
      RECT 32.576 3.263 32.662 3.405 ;
      RECT 32.49 3.267 32.576 3.408 ;
      RECT 32.453 3.271 32.49 3.411 ;
      RECT 32.367 3.274 32.453 3.414 ;
      RECT 32.281 3.278 32.367 3.417 ;
      RECT 32.195 3.283 32.281 3.421 ;
      RECT 32.175 3.285 32.195 3.424 ;
      RECT 32.155 3.284 32.175 3.425 ;
      RECT 32.106 3.281 32.155 3.426 ;
      RECT 32.02 3.276 32.106 3.429 ;
      RECT 31.97 3.271 32.02 3.431 ;
      RECT 31.946 3.269 31.97 3.432 ;
      RECT 31.86 3.264 31.946 3.434 ;
      RECT 31.835 3.26 31.86 3.433 ;
      RECT 31.825 3.257 31.835 3.431 ;
      RECT 31.815 3.25 31.825 3.428 ;
      RECT 31.81 3.23 31.815 3.423 ;
      RECT 31.8 3.2 31.81 3.418 ;
      RECT 31.785 3.07 31.8 3.409 ;
      RECT 31.78 3.062 31.785 3.402 ;
      RECT 31.76 3.055 31.78 3.394 ;
      RECT 31.755 3.037 31.76 3.386 ;
      RECT 31.745 3.017 31.755 3.381 ;
      RECT 31.74 2.99 31.745 3.377 ;
      RECT 31.735 2.967 31.74 3.374 ;
      RECT 31.715 2.925 31.735 3.366 ;
      RECT 31.68 2.84 31.715 3.35 ;
      RECT 31.675 2.772 31.68 3.338 ;
      RECT 31.66 2.742 31.675 3.332 ;
      RECT 31.655 1.987 31.66 2.233 ;
      RECT 31.645 2.712 31.66 3.323 ;
      RECT 31.65 1.982 31.655 2.265 ;
      RECT 31.645 1.977 31.65 2.308 ;
      RECT 31.64 1.975 31.645 2.343 ;
      RECT 31.625 2.675 31.645 3.313 ;
      RECT 31.635 1.975 31.64 2.38 ;
      RECT 31.62 1.975 31.635 2.478 ;
      RECT 31.62 2.648 31.625 3.306 ;
      RECT 31.615 1.975 31.62 2.553 ;
      RECT 31.615 2.636 31.62 3.303 ;
      RECT 31.61 1.975 31.615 2.585 ;
      RECT 31.61 2.615 31.615 3.3 ;
      RECT 31.605 1.975 31.61 3.297 ;
      RECT 31.57 1.975 31.605 3.283 ;
      RECT 31.555 1.975 31.57 3.265 ;
      RECT 31.535 1.975 31.555 3.255 ;
      RECT 31.51 1.975 31.535 3.238 ;
      RECT 31.505 1.975 31.51 3.188 ;
      RECT 31.495 1.975 31.5 3.018 ;
      RECT 31.49 1.975 31.495 2.925 ;
      RECT 31.485 1.975 31.49 2.838 ;
      RECT 31.48 1.975 31.485 2.77 ;
      RECT 31.475 1.975 31.48 2.713 ;
      RECT 31.465 1.975 31.475 2.608 ;
      RECT 31.46 1.975 31.465 2.48 ;
      RECT 31.455 1.975 31.46 2.398 ;
      RECT 31.45 1.977 31.455 2.315 ;
      RECT 31.445 1.982 31.45 2.248 ;
      RECT 31.44 1.987 31.445 2.175 ;
      RECT 34.255 2.305 34.515 2.565 ;
      RECT 34.275 2.272 34.485 2.565 ;
      RECT 34.275 2.27 34.475 2.565 ;
      RECT 34.285 2.257 34.475 2.565 ;
      RECT 34.285 2.255 34.4 2.565 ;
      RECT 33.76 2.38 33.935 2.66 ;
      RECT 33.755 2.38 33.935 2.658 ;
      RECT 33.755 2.38 33.95 2.655 ;
      RECT 33.745 2.38 33.95 2.653 ;
      RECT 33.69 2.38 33.95 2.64 ;
      RECT 33.69 2.455 33.955 2.618 ;
      RECT 33.235 2.392 33.255 2.635 ;
      RECT 33.235 2.392 33.295 2.634 ;
      RECT 33.23 2.394 33.295 2.633 ;
      RECT 33.23 2.394 33.381 2.632 ;
      RECT 33.23 2.394 33.45 2.631 ;
      RECT 33.23 2.394 33.47 2.623 ;
      RECT 33.21 2.397 33.47 2.621 ;
      RECT 33.195 2.407 33.47 2.606 ;
      RECT 33.195 2.407 33.485 2.605 ;
      RECT 33.19 2.416 33.485 2.597 ;
      RECT 33.19 2.416 33.49 2.593 ;
      RECT 33.295 2.33 33.555 2.59 ;
      RECT 33.185 2.418 33.555 2.475 ;
      RECT 33.255 2.385 33.555 2.59 ;
      RECT 33.22 3.578 33.225 3.785 ;
      RECT 33.17 3.572 33.22 3.784 ;
      RECT 33.137 3.586 33.23 3.783 ;
      RECT 33.051 3.586 33.23 3.782 ;
      RECT 32.965 3.586 33.23 3.781 ;
      RECT 32.965 3.685 33.235 3.778 ;
      RECT 32.96 3.685 33.235 3.773 ;
      RECT 32.955 3.685 33.235 3.755 ;
      RECT 32.95 3.685 33.235 3.738 ;
      RECT 32.91 3.47 33.17 3.73 ;
      RECT 32.37 2.62 32.456 3.034 ;
      RECT 32.37 2.62 32.495 3.031 ;
      RECT 32.37 2.62 32.515 3.021 ;
      RECT 32.325 2.62 32.515 3.018 ;
      RECT 32.325 2.772 32.525 3.008 ;
      RECT 32.325 2.793 32.53 3.002 ;
      RECT 32.325 2.811 32.535 2.998 ;
      RECT 32.325 2.831 32.545 2.993 ;
      RECT 32.3 2.831 32.545 2.99 ;
      RECT 32.29 2.831 32.545 2.968 ;
      RECT 32.29 2.847 32.55 2.938 ;
      RECT 32.255 2.62 32.515 2.925 ;
      RECT 32.255 2.859 32.555 2.88 ;
      RECT 29.92 7.765 30.21 7.995 ;
      RECT 29.98 6.285 30.15 7.995 ;
      RECT 29.965 6.66 30.32 7.015 ;
      RECT 29.92 6.285 30.21 6.515 ;
      RECT 29.92 2.365 30.21 2.595 ;
      RECT 29.98 0.885 30.15 2.595 ;
      RECT 29.92 0.885 30.21 1.115 ;
      RECT 29.51 2.735 29.84 2.965 ;
      RECT 29.51 2.765 30.01 2.935 ;
      RECT 29.51 2.395 29.7 2.965 ;
      RECT 28.93 2.365 29.22 2.595 ;
      RECT 28.93 2.395 29.7 2.565 ;
      RECT 28.99 0.885 29.16 2.595 ;
      RECT 28.93 0.885 29.22 1.115 ;
      RECT 28.93 7.765 29.22 7.995 ;
      RECT 28.99 6.285 29.16 7.995 ;
      RECT 28.93 6.285 29.22 6.515 ;
      RECT 28.93 6.325 29.78 6.485 ;
      RECT 29.61 5.915 29.78 6.485 ;
      RECT 28.93 6.32 29.32 6.485 ;
      RECT 29.55 5.915 29.84 6.145 ;
      RECT 29.55 5.945 30.01 6.115 ;
      RECT 28.56 2.735 28.85 2.965 ;
      RECT 28.56 2.765 29.02 2.935 ;
      RECT 28.62 1.655 28.785 2.965 ;
      RECT 27.135 1.625 27.425 1.855 ;
      RECT 27.135 1.655 28.785 1.825 ;
      RECT 27.195 0.885 27.365 1.855 ;
      RECT 27.135 0.885 27.425 1.115 ;
      RECT 27.135 7.765 27.425 7.995 ;
      RECT 27.195 7.025 27.365 7.995 ;
      RECT 27.195 7.12 28.785 7.29 ;
      RECT 28.615 5.915 28.785 7.29 ;
      RECT 27.135 7.025 27.425 7.255 ;
      RECT 28.56 5.915 28.85 6.145 ;
      RECT 28.56 5.945 29.02 6.115 ;
      RECT 25.185 2.705 25.525 3.055 ;
      RECT 25.275 2.025 25.445 3.055 ;
      RECT 27.565 1.965 27.915 2.315 ;
      RECT 25.275 2.025 27.915 2.195 ;
      RECT 27.59 6.655 27.915 6.98 ;
      RECT 22.13 6.61 22.48 6.96 ;
      RECT 27.565 6.655 27.915 6.885 ;
      RECT 21.93 6.655 22.48 6.885 ;
      RECT 21.76 6.685 27.915 6.855 ;
      RECT 26.79 2.365 27.11 2.685 ;
      RECT 26.76 2.365 27.11 2.595 ;
      RECT 26.59 2.395 27.11 2.565 ;
      RECT 26.79 6.255 27.11 6.545 ;
      RECT 26.76 6.285 27.11 6.515 ;
      RECT 26.59 6.315 27.11 6.485 ;
      RECT 25.745 2.705 26.085 3.055 ;
      RECT 25.745 2.765 26.225 2.935 ;
      RECT 25.74 5.86 26.08 6.21 ;
      RECT 20.13 5.915 20.42 6.145 ;
      RECT 20.13 5.945 26.225 6.115 ;
      RECT 22.48 2.985 22.63 3.26 ;
      RECT 23.02 2.065 23.025 2.285 ;
      RECT 24.17 2.265 24.185 2.463 ;
      RECT 24.135 2.257 24.17 2.47 ;
      RECT 24.105 2.25 24.135 2.47 ;
      RECT 24.05 2.215 24.105 2.47 ;
      RECT 23.985 2.152 24.05 2.47 ;
      RECT 23.98 2.117 23.985 2.468 ;
      RECT 23.975 2.112 23.98 2.46 ;
      RECT 23.97 2.107 23.975 2.446 ;
      RECT 23.965 2.104 23.97 2.439 ;
      RECT 23.92 2.094 23.965 2.39 ;
      RECT 23.9 2.081 23.92 2.325 ;
      RECT 23.895 2.076 23.9 2.298 ;
      RECT 23.89 2.075 23.895 2.291 ;
      RECT 23.885 2.074 23.89 2.284 ;
      RECT 23.8 2.059 23.885 2.23 ;
      RECT 23.77 2.04 23.8 2.18 ;
      RECT 23.69 2.023 23.77 2.165 ;
      RECT 23.655 2.01 23.69 2.15 ;
      RECT 23.647 2.01 23.655 2.145 ;
      RECT 23.561 2.011 23.647 2.145 ;
      RECT 23.475 2.013 23.561 2.145 ;
      RECT 23.45 2.014 23.475 2.149 ;
      RECT 23.375 2.02 23.45 2.164 ;
      RECT 23.292 2.032 23.375 2.188 ;
      RECT 23.206 2.045 23.292 2.214 ;
      RECT 23.12 2.058 23.206 2.24 ;
      RECT 23.085 2.067 23.12 2.259 ;
      RECT 23.035 2.067 23.085 2.272 ;
      RECT 23.025 2.065 23.035 2.283 ;
      RECT 23.01 2.062 23.02 2.285 ;
      RECT 22.995 2.054 23.01 2.293 ;
      RECT 22.98 2.046 22.995 2.313 ;
      RECT 22.975 2.041 22.98 2.37 ;
      RECT 22.96 2.036 22.975 2.443 ;
      RECT 22.955 2.031 22.96 2.485 ;
      RECT 22.95 2.029 22.955 2.513 ;
      RECT 22.945 2.027 22.95 2.535 ;
      RECT 22.935 2.023 22.945 2.578 ;
      RECT 22.93 2.02 22.935 2.603 ;
      RECT 22.925 2.018 22.93 2.623 ;
      RECT 22.92 2.016 22.925 2.647 ;
      RECT 22.915 2.012 22.92 2.67 ;
      RECT 22.91 2.008 22.915 2.693 ;
      RECT 22.875 1.998 22.91 2.8 ;
      RECT 22.87 1.988 22.875 2.898 ;
      RECT 22.865 1.986 22.87 2.925 ;
      RECT 22.86 1.985 22.865 2.945 ;
      RECT 22.855 1.977 22.86 2.965 ;
      RECT 22.85 1.972 22.855 3 ;
      RECT 22.845 1.97 22.85 3.018 ;
      RECT 22.84 1.97 22.845 3.043 ;
      RECT 22.835 1.97 22.84 3.065 ;
      RECT 22.8 1.97 22.835 3.108 ;
      RECT 22.775 1.97 22.8 3.137 ;
      RECT 22.765 1.97 22.775 2.323 ;
      RECT 22.768 2.38 22.775 3.147 ;
      RECT 22.765 2.437 22.768 3.15 ;
      RECT 22.76 1.97 22.765 2.295 ;
      RECT 22.76 2.487 22.765 3.153 ;
      RECT 22.75 1.97 22.76 2.285 ;
      RECT 22.755 2.54 22.76 3.156 ;
      RECT 22.75 2.625 22.755 3.16 ;
      RECT 22.74 1.97 22.75 2.273 ;
      RECT 22.745 2.672 22.75 3.164 ;
      RECT 22.74 2.747 22.745 3.168 ;
      RECT 22.705 1.97 22.74 2.248 ;
      RECT 22.73 2.83 22.74 3.173 ;
      RECT 22.72 2.897 22.73 3.18 ;
      RECT 22.715 2.925 22.72 3.185 ;
      RECT 22.705 2.938 22.715 3.191 ;
      RECT 22.66 1.97 22.705 2.205 ;
      RECT 22.7 2.943 22.705 3.198 ;
      RECT 22.66 2.96 22.7 3.26 ;
      RECT 22.655 1.972 22.66 2.178 ;
      RECT 22.63 2.98 22.66 3.26 ;
      RECT 22.65 1.977 22.655 2.15 ;
      RECT 22.44 2.989 22.48 3.26 ;
      RECT 22.415 2.997 22.44 3.23 ;
      RECT 22.37 3.005 22.415 3.23 ;
      RECT 22.355 3.01 22.37 3.225 ;
      RECT 22.345 3.01 22.355 3.219 ;
      RECT 22.335 3.017 22.345 3.216 ;
      RECT 22.33 3.055 22.335 3.205 ;
      RECT 22.325 3.117 22.33 3.183 ;
      RECT 23.595 2.992 23.78 3.215 ;
      RECT 23.595 3.007 23.785 3.211 ;
      RECT 23.585 2.28 23.67 3.21 ;
      RECT 23.585 3.007 23.79 3.204 ;
      RECT 23.58 3.015 23.79 3.203 ;
      RECT 23.785 2.735 24.105 3.055 ;
      RECT 23.58 2.907 23.75 2.998 ;
      RECT 23.575 2.907 23.75 2.98 ;
      RECT 23.565 2.715 23.7 2.955 ;
      RECT 23.56 2.715 23.7 2.9 ;
      RECT 23.52 2.295 23.69 2.8 ;
      RECT 23.505 2.295 23.69 2.67 ;
      RECT 23.5 2.295 23.69 2.623 ;
      RECT 23.495 2.295 23.69 2.603 ;
      RECT 23.49 2.295 23.69 2.578 ;
      RECT 23.46 2.295 23.72 2.555 ;
      RECT 23.47 2.292 23.68 2.555 ;
      RECT 23.595 2.287 23.68 3.215 ;
      RECT 23.48 2.28 23.67 2.555 ;
      RECT 23.475 2.285 23.67 2.555 ;
      RECT 22.305 2.497 22.49 2.71 ;
      RECT 22.305 2.505 22.5 2.703 ;
      RECT 22.285 2.505 22.5 2.7 ;
      RECT 22.28 2.505 22.5 2.685 ;
      RECT 22.21 2.42 22.47 2.68 ;
      RECT 22.21 2.565 22.505 2.593 ;
      RECT 21.865 3.02 22.125 3.28 ;
      RECT 21.89 2.965 22.085 3.28 ;
      RECT 21.885 2.714 22.065 3.008 ;
      RECT 21.885 2.72 22.075 3.008 ;
      RECT 21.865 2.722 22.075 2.953 ;
      RECT 21.86 2.732 22.075 2.82 ;
      RECT 21.89 2.712 22.065 3.28 ;
      RECT 21.976 2.71 22.065 3.28 ;
      RECT 21.835 1.93 21.87 2.3 ;
      RECT 21.625 2.04 21.63 2.3 ;
      RECT 21.87 1.937 21.885 2.3 ;
      RECT 21.76 1.93 21.835 2.378 ;
      RECT 21.75 1.93 21.76 2.463 ;
      RECT 21.725 1.93 21.75 2.498 ;
      RECT 21.685 1.93 21.725 2.566 ;
      RECT 21.675 1.937 21.685 2.618 ;
      RECT 21.645 2.04 21.675 2.659 ;
      RECT 21.64 2.04 21.645 2.698 ;
      RECT 21.63 2.04 21.64 2.718 ;
      RECT 21.625 2.335 21.63 2.755 ;
      RECT 21.62 2.352 21.625 2.775 ;
      RECT 21.605 2.415 21.62 2.815 ;
      RECT 21.6 2.458 21.605 2.85 ;
      RECT 21.595 2.466 21.6 2.863 ;
      RECT 21.585 2.48 21.595 2.885 ;
      RECT 21.56 2.515 21.585 2.95 ;
      RECT 21.55 2.55 21.56 3.013 ;
      RECT 21.53 2.58 21.55 3.074 ;
      RECT 21.515 2.616 21.53 3.141 ;
      RECT 21.505 2.644 21.515 3.18 ;
      RECT 21.495 2.666 21.505 3.2 ;
      RECT 21.49 2.676 21.495 3.211 ;
      RECT 21.485 2.685 21.49 3.214 ;
      RECT 21.475 2.703 21.485 3.218 ;
      RECT 21.465 2.721 21.475 3.219 ;
      RECT 21.44 2.76 21.465 3.216 ;
      RECT 21.42 2.802 21.44 3.213 ;
      RECT 21.405 2.84 21.42 3.212 ;
      RECT 21.37 2.875 21.405 3.209 ;
      RECT 21.365 2.897 21.37 3.207 ;
      RECT 21.3 2.937 21.365 3.204 ;
      RECT 21.295 2.977 21.3 3.2 ;
      RECT 21.28 2.987 21.295 3.191 ;
      RECT 21.27 3.107 21.28 3.176 ;
      RECT 21.75 3.52 21.76 3.78 ;
      RECT 21.75 3.523 21.77 3.779 ;
      RECT 21.74 3.513 21.75 3.778 ;
      RECT 21.73 3.528 21.81 3.774 ;
      RECT 21.715 3.507 21.73 3.772 ;
      RECT 21.69 3.532 21.815 3.768 ;
      RECT 21.675 3.492 21.69 3.763 ;
      RECT 21.675 3.534 21.825 3.762 ;
      RECT 21.675 3.542 21.84 3.755 ;
      RECT 21.615 3.479 21.675 3.745 ;
      RECT 21.605 3.466 21.615 3.727 ;
      RECT 21.58 3.456 21.605 3.717 ;
      RECT 21.575 3.446 21.58 3.709 ;
      RECT 21.51 3.542 21.84 3.691 ;
      RECT 21.425 3.542 21.84 3.653 ;
      RECT 21.315 3.37 21.575 3.63 ;
      RECT 21.69 3.5 21.715 3.768 ;
      RECT 21.73 3.51 21.74 3.774 ;
      RECT 21.315 3.518 21.755 3.63 ;
      RECT 21.5 7.765 21.79 7.995 ;
      RECT 21.56 7.025 21.73 7.995 ;
      RECT 21.46 7.055 21.83 7.425 ;
      RECT 21.5 7.025 21.79 7.425 ;
      RECT 20.53 3.275 20.56 3.575 ;
      RECT 20.305 3.26 20.31 3.535 ;
      RECT 20.105 3.26 20.26 3.52 ;
      RECT 21.405 1.975 21.435 2.235 ;
      RECT 21.395 1.975 21.405 2.343 ;
      RECT 21.375 1.975 21.395 2.353 ;
      RECT 21.36 1.975 21.375 2.365 ;
      RECT 21.305 1.975 21.36 2.415 ;
      RECT 21.29 1.975 21.305 2.463 ;
      RECT 21.26 1.975 21.29 2.498 ;
      RECT 21.205 1.975 21.26 2.56 ;
      RECT 21.185 1.975 21.205 2.628 ;
      RECT 21.18 1.975 21.185 2.658 ;
      RECT 21.175 1.975 21.18 2.67 ;
      RECT 21.17 2.092 21.175 2.688 ;
      RECT 21.15 2.11 21.17 2.713 ;
      RECT 21.13 2.137 21.15 2.763 ;
      RECT 21.125 2.157 21.13 2.794 ;
      RECT 21.12 2.165 21.125 2.811 ;
      RECT 21.105 2.191 21.12 2.84 ;
      RECT 21.09 2.233 21.105 2.875 ;
      RECT 21.085 2.262 21.09 2.898 ;
      RECT 21.08 2.277 21.085 2.911 ;
      RECT 21.075 2.3 21.08 2.922 ;
      RECT 21.065 2.32 21.075 2.94 ;
      RECT 21.055 2.35 21.065 2.963 ;
      RECT 21.05 2.372 21.055 2.983 ;
      RECT 21.045 2.387 21.05 2.998 ;
      RECT 21.03 2.417 21.045 3.025 ;
      RECT 21.025 2.447 21.03 3.051 ;
      RECT 21.02 2.465 21.025 3.063 ;
      RECT 21.01 2.495 21.02 3.082 ;
      RECT 21 2.52 21.01 3.107 ;
      RECT 20.995 2.54 21 3.126 ;
      RECT 20.99 2.557 20.995 3.139 ;
      RECT 20.98 2.583 20.99 3.158 ;
      RECT 20.97 2.621 20.98 3.185 ;
      RECT 20.965 2.647 20.97 3.205 ;
      RECT 20.96 2.657 20.965 3.215 ;
      RECT 20.955 2.67 20.96 3.23 ;
      RECT 20.95 2.685 20.955 3.24 ;
      RECT 20.945 2.707 20.95 3.255 ;
      RECT 20.94 2.725 20.945 3.266 ;
      RECT 20.935 2.735 20.94 3.277 ;
      RECT 20.93 2.743 20.935 3.289 ;
      RECT 20.925 2.751 20.93 3.3 ;
      RECT 20.92 2.777 20.925 3.313 ;
      RECT 20.91 2.805 20.92 3.326 ;
      RECT 20.905 2.835 20.91 3.335 ;
      RECT 20.9 2.85 20.905 3.342 ;
      RECT 20.885 2.875 20.9 3.349 ;
      RECT 20.88 2.897 20.885 3.355 ;
      RECT 20.875 2.922 20.88 3.358 ;
      RECT 20.866 2.95 20.875 3.362 ;
      RECT 20.86 2.967 20.866 3.367 ;
      RECT 20.855 2.985 20.86 3.371 ;
      RECT 20.85 2.997 20.855 3.374 ;
      RECT 20.845 3.018 20.85 3.378 ;
      RECT 20.84 3.036 20.845 3.381 ;
      RECT 20.835 3.05 20.84 3.384 ;
      RECT 20.83 3.067 20.835 3.387 ;
      RECT 20.825 3.08 20.83 3.39 ;
      RECT 20.8 3.117 20.825 3.398 ;
      RECT 20.795 3.162 20.8 3.407 ;
      RECT 20.79 3.19 20.795 3.41 ;
      RECT 20.78 3.21 20.79 3.414 ;
      RECT 20.775 3.23 20.78 3.419 ;
      RECT 20.77 3.245 20.775 3.422 ;
      RECT 20.75 3.255 20.77 3.429 ;
      RECT 20.685 3.262 20.75 3.455 ;
      RECT 20.65 3.265 20.685 3.483 ;
      RECT 20.635 3.268 20.65 3.498 ;
      RECT 20.625 3.269 20.635 3.513 ;
      RECT 20.615 3.27 20.625 3.53 ;
      RECT 20.61 3.27 20.615 3.545 ;
      RECT 20.605 3.27 20.61 3.553 ;
      RECT 20.59 3.271 20.605 3.568 ;
      RECT 20.56 3.273 20.59 3.575 ;
      RECT 20.45 3.28 20.53 3.575 ;
      RECT 20.405 3.285 20.45 3.575 ;
      RECT 20.395 3.286 20.405 3.565 ;
      RECT 20.385 3.287 20.395 3.558 ;
      RECT 20.365 3.289 20.385 3.553 ;
      RECT 20.355 3.26 20.365 3.548 ;
      RECT 20.31 3.26 20.355 3.54 ;
      RECT 20.28 3.26 20.305 3.53 ;
      RECT 20.26 3.26 20.28 3.523 ;
      RECT 20.54 2.06 20.8 2.32 ;
      RECT 20.42 2.075 20.43 2.24 ;
      RECT 20.405 2.075 20.41 2.235 ;
      RECT 17.77 1.915 17.955 2.205 ;
      RECT 19.585 2.04 19.6 2.195 ;
      RECT 17.735 1.915 17.76 2.175 ;
      RECT 20.15 1.965 20.155 2.107 ;
      RECT 20.065 1.96 20.09 2.1 ;
      RECT 20.465 2.077 20.54 2.27 ;
      RECT 20.45 2.075 20.465 2.253 ;
      RECT 20.43 2.075 20.45 2.245 ;
      RECT 20.41 2.075 20.42 2.238 ;
      RECT 20.365 2.07 20.405 2.228 ;
      RECT 20.325 2.045 20.365 2.213 ;
      RECT 20.31 2.02 20.325 2.203 ;
      RECT 20.305 2.014 20.31 2.201 ;
      RECT 20.27 2.006 20.305 2.184 ;
      RECT 20.265 1.999 20.27 2.172 ;
      RECT 20.245 1.994 20.265 2.16 ;
      RECT 20.235 1.988 20.245 2.145 ;
      RECT 20.215 1.983 20.235 2.13 ;
      RECT 20.205 1.978 20.215 2.123 ;
      RECT 20.2 1.976 20.205 2.118 ;
      RECT 20.195 1.975 20.2 2.115 ;
      RECT 20.155 1.97 20.195 2.111 ;
      RECT 20.135 1.964 20.15 2.106 ;
      RECT 20.1 1.961 20.135 2.103 ;
      RECT 20.09 1.96 20.1 2.101 ;
      RECT 20.03 1.96 20.065 2.098 ;
      RECT 19.985 1.96 20.03 2.098 ;
      RECT 19.935 1.96 19.985 2.101 ;
      RECT 19.92 1.962 19.935 2.103 ;
      RECT 19.905 1.965 19.92 2.104 ;
      RECT 19.895 1.97 19.905 2.105 ;
      RECT 19.865 1.975 19.895 2.11 ;
      RECT 19.855 1.981 19.865 2.118 ;
      RECT 19.845 1.983 19.855 2.122 ;
      RECT 19.835 1.987 19.845 2.126 ;
      RECT 19.81 1.993 19.835 2.134 ;
      RECT 19.8 1.998 19.81 2.142 ;
      RECT 19.785 2.002 19.8 2.146 ;
      RECT 19.75 2.008 19.785 2.154 ;
      RECT 19.73 2.013 19.75 2.164 ;
      RECT 19.7 2.02 19.73 2.173 ;
      RECT 19.655 2.029 19.7 2.187 ;
      RECT 19.65 2.034 19.655 2.198 ;
      RECT 19.63 2.037 19.65 2.199 ;
      RECT 19.6 2.04 19.63 2.197 ;
      RECT 19.565 2.04 19.585 2.193 ;
      RECT 19.495 2.04 19.565 2.184 ;
      RECT 19.48 2.037 19.495 2.176 ;
      RECT 19.44 2.03 19.48 2.171 ;
      RECT 19.415 2.02 19.44 2.164 ;
      RECT 19.41 2.014 19.415 2.161 ;
      RECT 19.37 2.008 19.41 2.158 ;
      RECT 19.355 2.001 19.37 2.153 ;
      RECT 19.335 1.997 19.355 2.148 ;
      RECT 19.32 1.992 19.335 2.144 ;
      RECT 19.305 1.987 19.32 2.142 ;
      RECT 19.29 1.983 19.305 2.141 ;
      RECT 19.275 1.981 19.29 2.137 ;
      RECT 19.265 1.979 19.275 2.132 ;
      RECT 19.25 1.976 19.265 2.128 ;
      RECT 19.24 1.974 19.25 2.123 ;
      RECT 19.22 1.971 19.24 2.119 ;
      RECT 19.175 1.97 19.22 2.117 ;
      RECT 19.115 1.972 19.175 2.118 ;
      RECT 19.095 1.974 19.115 2.12 ;
      RECT 19.065 1.977 19.095 2.121 ;
      RECT 19.015 1.982 19.065 2.123 ;
      RECT 19.01 1.985 19.015 2.125 ;
      RECT 19 1.987 19.01 2.128 ;
      RECT 18.995 1.989 19 2.131 ;
      RECT 18.945 1.992 18.995 2.138 ;
      RECT 18.925 1.996 18.945 2.15 ;
      RECT 18.915 1.999 18.925 2.156 ;
      RECT 18.905 2 18.915 2.159 ;
      RECT 18.866 2.003 18.905 2.161 ;
      RECT 18.78 2.01 18.866 2.164 ;
      RECT 18.706 2.02 18.78 2.168 ;
      RECT 18.62 2.031 18.706 2.173 ;
      RECT 18.605 2.038 18.62 2.175 ;
      RECT 18.55 2.042 18.605 2.176 ;
      RECT 18.536 2.045 18.55 2.178 ;
      RECT 18.45 2.045 18.536 2.18 ;
      RECT 18.41 2.042 18.45 2.183 ;
      RECT 18.386 2.038 18.41 2.185 ;
      RECT 18.3 2.028 18.386 2.188 ;
      RECT 18.27 2.017 18.3 2.189 ;
      RECT 18.251 2.013 18.27 2.188 ;
      RECT 18.165 2.006 18.251 2.185 ;
      RECT 18.105 1.995 18.165 2.182 ;
      RECT 18.085 1.987 18.105 2.18 ;
      RECT 18.05 1.982 18.085 2.179 ;
      RECT 18.025 1.977 18.05 2.178 ;
      RECT 17.995 1.972 18.025 2.177 ;
      RECT 17.97 1.915 17.995 2.176 ;
      RECT 17.955 1.915 17.97 2.2 ;
      RECT 17.76 1.915 17.77 2.2 ;
      RECT 19.535 2.935 19.54 3.075 ;
      RECT 19.195 2.935 19.23 3.073 ;
      RECT 18.77 2.92 18.785 3.065 ;
      RECT 20.6 2.7 20.69 2.96 ;
      RECT 20.43 2.565 20.53 2.96 ;
      RECT 17.465 2.54 17.545 2.75 ;
      RECT 20.555 2.677 20.6 2.96 ;
      RECT 20.545 2.647 20.555 2.96 ;
      RECT 20.53 2.57 20.545 2.96 ;
      RECT 20.345 2.565 20.43 2.925 ;
      RECT 20.34 2.567 20.345 2.92 ;
      RECT 20.335 2.572 20.34 2.92 ;
      RECT 20.3 2.672 20.335 2.92 ;
      RECT 20.29 2.7 20.3 2.92 ;
      RECT 20.28 2.715 20.29 2.92 ;
      RECT 20.27 2.727 20.28 2.92 ;
      RECT 20.265 2.737 20.27 2.92 ;
      RECT 20.25 2.747 20.265 2.922 ;
      RECT 20.245 2.762 20.25 2.924 ;
      RECT 20.23 2.775 20.245 2.926 ;
      RECT 20.225 2.79 20.23 2.929 ;
      RECT 20.205 2.8 20.225 2.933 ;
      RECT 20.19 2.81 20.205 2.936 ;
      RECT 20.155 2.817 20.19 2.941 ;
      RECT 20.111 2.824 20.155 2.949 ;
      RECT 20.025 2.836 20.111 2.962 ;
      RECT 20 2.847 20.025 2.973 ;
      RECT 19.97 2.852 20 2.978 ;
      RECT 19.935 2.857 19.97 2.986 ;
      RECT 19.905 2.862 19.935 2.993 ;
      RECT 19.88 2.867 19.905 2.998 ;
      RECT 19.815 2.874 19.88 3.007 ;
      RECT 19.745 2.887 19.815 3.023 ;
      RECT 19.715 2.897 19.745 3.035 ;
      RECT 19.69 2.902 19.715 3.042 ;
      RECT 19.635 2.909 19.69 3.05 ;
      RECT 19.63 2.916 19.635 3.055 ;
      RECT 19.625 2.918 19.63 3.056 ;
      RECT 19.61 2.92 19.625 3.058 ;
      RECT 19.605 2.92 19.61 3.061 ;
      RECT 19.54 2.927 19.605 3.068 ;
      RECT 19.505 2.937 19.535 3.078 ;
      RECT 19.488 2.94 19.505 3.08 ;
      RECT 19.402 2.939 19.488 3.079 ;
      RECT 19.316 2.937 19.402 3.076 ;
      RECT 19.23 2.936 19.316 3.074 ;
      RECT 19.129 2.934 19.195 3.073 ;
      RECT 19.043 2.931 19.129 3.071 ;
      RECT 18.957 2.927 19.043 3.069 ;
      RECT 18.871 2.924 18.957 3.068 ;
      RECT 18.785 2.921 18.871 3.066 ;
      RECT 18.685 2.92 18.77 3.063 ;
      RECT 18.635 2.918 18.685 3.061 ;
      RECT 18.615 2.915 18.635 3.059 ;
      RECT 18.595 2.913 18.615 3.056 ;
      RECT 18.57 2.909 18.595 3.053 ;
      RECT 18.525 2.903 18.57 3.048 ;
      RECT 18.485 2.897 18.525 3.04 ;
      RECT 18.46 2.892 18.485 3.033 ;
      RECT 18.405 2.885 18.46 3.025 ;
      RECT 18.381 2.878 18.405 3.018 ;
      RECT 18.295 2.869 18.381 3.008 ;
      RECT 18.265 2.861 18.295 2.998 ;
      RECT 18.235 2.857 18.265 2.993 ;
      RECT 18.23 2.854 18.235 2.99 ;
      RECT 18.225 2.853 18.23 2.99 ;
      RECT 18.15 2.846 18.225 2.983 ;
      RECT 18.111 2.837 18.15 2.972 ;
      RECT 18.025 2.827 18.111 2.96 ;
      RECT 17.985 2.817 18.025 2.948 ;
      RECT 17.946 2.812 17.985 2.941 ;
      RECT 17.86 2.802 17.946 2.93 ;
      RECT 17.82 2.79 17.86 2.919 ;
      RECT 17.785 2.775 17.82 2.912 ;
      RECT 17.775 2.765 17.785 2.909 ;
      RECT 17.755 2.75 17.775 2.907 ;
      RECT 17.725 2.72 17.755 2.903 ;
      RECT 17.715 2.7 17.725 2.898 ;
      RECT 17.71 2.692 17.715 2.895 ;
      RECT 17.705 2.685 17.71 2.893 ;
      RECT 17.69 2.672 17.705 2.886 ;
      RECT 17.685 2.662 17.69 2.878 ;
      RECT 17.68 2.655 17.685 2.873 ;
      RECT 17.675 2.65 17.68 2.869 ;
      RECT 17.66 2.637 17.675 2.861 ;
      RECT 17.655 2.547 17.66 2.85 ;
      RECT 17.65 2.542 17.655 2.843 ;
      RECT 17.575 2.54 17.65 2.803 ;
      RECT 17.545 2.54 17.575 2.758 ;
      RECT 17.45 2.545 17.465 2.745 ;
      RECT 19.935 2.25 20.195 2.51 ;
      RECT 19.92 2.238 20.1 2.475 ;
      RECT 19.915 2.239 20.1 2.473 ;
      RECT 19.9 2.243 20.11 2.463 ;
      RECT 19.895 2.248 20.115 2.433 ;
      RECT 19.9 2.245 20.115 2.463 ;
      RECT 19.915 2.24 20.11 2.473 ;
      RECT 19.935 2.237 20.1 2.51 ;
      RECT 19.935 2.236 20.09 2.51 ;
      RECT 19.96 2.235 20.09 2.51 ;
      RECT 19.52 2.48 19.78 2.74 ;
      RECT 19.395 2.525 19.78 2.735 ;
      RECT 19.385 2.53 19.78 2.73 ;
      RECT 19.4 3.47 19.415 3.78 ;
      RECT 17.995 3.24 18.005 3.37 ;
      RECT 17.775 3.235 17.88 3.37 ;
      RECT 17.69 3.24 17.74 3.37 ;
      RECT 16.24 1.975 16.245 3.08 ;
      RECT 19.495 3.562 19.5 3.698 ;
      RECT 19.49 3.557 19.495 3.758 ;
      RECT 19.485 3.555 19.49 3.771 ;
      RECT 19.47 3.552 19.485 3.773 ;
      RECT 19.465 3.547 19.47 3.775 ;
      RECT 19.46 3.543 19.465 3.778 ;
      RECT 19.445 3.538 19.46 3.78 ;
      RECT 19.415 3.53 19.445 3.78 ;
      RECT 19.376 3.47 19.4 3.78 ;
      RECT 19.29 3.47 19.376 3.777 ;
      RECT 19.26 3.47 19.29 3.77 ;
      RECT 19.235 3.47 19.26 3.763 ;
      RECT 19.21 3.47 19.235 3.755 ;
      RECT 19.195 3.47 19.21 3.748 ;
      RECT 19.17 3.47 19.195 3.74 ;
      RECT 19.155 3.47 19.17 3.733 ;
      RECT 19.115 3.48 19.155 3.722 ;
      RECT 19.105 3.475 19.115 3.712 ;
      RECT 19.101 3.474 19.105 3.709 ;
      RECT 19.015 3.466 19.101 3.692 ;
      RECT 18.982 3.455 19.015 3.669 ;
      RECT 18.896 3.444 18.982 3.647 ;
      RECT 18.81 3.428 18.896 3.616 ;
      RECT 18.74 3.413 18.81 3.588 ;
      RECT 18.73 3.406 18.74 3.575 ;
      RECT 18.7 3.403 18.73 3.565 ;
      RECT 18.675 3.399 18.7 3.558 ;
      RECT 18.66 3.396 18.675 3.553 ;
      RECT 18.655 3.395 18.66 3.548 ;
      RECT 18.625 3.39 18.655 3.541 ;
      RECT 18.62 3.385 18.625 3.536 ;
      RECT 18.605 3.382 18.62 3.531 ;
      RECT 18.6 3.377 18.605 3.526 ;
      RECT 18.58 3.372 18.6 3.523 ;
      RECT 18.565 3.367 18.58 3.515 ;
      RECT 18.55 3.361 18.565 3.51 ;
      RECT 18.52 3.352 18.55 3.503 ;
      RECT 18.515 3.345 18.52 3.495 ;
      RECT 18.51 3.343 18.515 3.493 ;
      RECT 18.505 3.342 18.51 3.49 ;
      RECT 18.465 3.335 18.505 3.483 ;
      RECT 18.451 3.325 18.465 3.473 ;
      RECT 18.4 3.314 18.451 3.461 ;
      RECT 18.375 3.3 18.4 3.447 ;
      RECT 18.35 3.289 18.375 3.439 ;
      RECT 18.33 3.278 18.35 3.433 ;
      RECT 18.32 3.272 18.33 3.428 ;
      RECT 18.315 3.27 18.32 3.424 ;
      RECT 18.295 3.265 18.315 3.419 ;
      RECT 18.265 3.255 18.295 3.409 ;
      RECT 18.26 3.247 18.265 3.402 ;
      RECT 18.245 3.245 18.26 3.398 ;
      RECT 18.225 3.245 18.245 3.393 ;
      RECT 18.22 3.244 18.225 3.391 ;
      RECT 18.215 3.244 18.22 3.388 ;
      RECT 18.175 3.243 18.215 3.383 ;
      RECT 18.15 3.242 18.175 3.378 ;
      RECT 18.09 3.241 18.15 3.375 ;
      RECT 18.005 3.24 18.09 3.373 ;
      RECT 17.966 3.239 17.995 3.37 ;
      RECT 17.88 3.237 17.966 3.37 ;
      RECT 17.74 3.237 17.775 3.37 ;
      RECT 17.65 3.241 17.69 3.373 ;
      RECT 17.635 3.244 17.65 3.38 ;
      RECT 17.625 3.245 17.635 3.387 ;
      RECT 17.6 3.248 17.625 3.392 ;
      RECT 17.595 3.25 17.6 3.395 ;
      RECT 17.545 3.252 17.595 3.396 ;
      RECT 17.506 3.256 17.545 3.398 ;
      RECT 17.42 3.258 17.506 3.401 ;
      RECT 17.402 3.26 17.42 3.403 ;
      RECT 17.316 3.263 17.402 3.405 ;
      RECT 17.23 3.267 17.316 3.408 ;
      RECT 17.193 3.271 17.23 3.411 ;
      RECT 17.107 3.274 17.193 3.414 ;
      RECT 17.021 3.278 17.107 3.417 ;
      RECT 16.935 3.283 17.021 3.421 ;
      RECT 16.915 3.285 16.935 3.424 ;
      RECT 16.895 3.284 16.915 3.425 ;
      RECT 16.846 3.281 16.895 3.426 ;
      RECT 16.76 3.276 16.846 3.429 ;
      RECT 16.71 3.271 16.76 3.431 ;
      RECT 16.686 3.269 16.71 3.432 ;
      RECT 16.6 3.264 16.686 3.434 ;
      RECT 16.575 3.26 16.6 3.433 ;
      RECT 16.565 3.257 16.575 3.431 ;
      RECT 16.555 3.25 16.565 3.428 ;
      RECT 16.55 3.23 16.555 3.423 ;
      RECT 16.54 3.2 16.55 3.418 ;
      RECT 16.525 3.07 16.54 3.409 ;
      RECT 16.52 3.062 16.525 3.402 ;
      RECT 16.5 3.055 16.52 3.394 ;
      RECT 16.495 3.037 16.5 3.386 ;
      RECT 16.485 3.017 16.495 3.381 ;
      RECT 16.48 2.99 16.485 3.377 ;
      RECT 16.475 2.967 16.48 3.374 ;
      RECT 16.455 2.925 16.475 3.366 ;
      RECT 16.42 2.84 16.455 3.35 ;
      RECT 16.415 2.772 16.42 3.338 ;
      RECT 16.4 2.742 16.415 3.332 ;
      RECT 16.395 1.987 16.4 2.233 ;
      RECT 16.385 2.712 16.4 3.323 ;
      RECT 16.39 1.982 16.395 2.265 ;
      RECT 16.385 1.977 16.39 2.308 ;
      RECT 16.38 1.975 16.385 2.343 ;
      RECT 16.365 2.675 16.385 3.313 ;
      RECT 16.375 1.975 16.38 2.38 ;
      RECT 16.36 1.975 16.375 2.478 ;
      RECT 16.36 2.648 16.365 3.306 ;
      RECT 16.355 1.975 16.36 2.553 ;
      RECT 16.355 2.636 16.36 3.303 ;
      RECT 16.35 1.975 16.355 2.585 ;
      RECT 16.35 2.615 16.355 3.3 ;
      RECT 16.345 1.975 16.35 3.297 ;
      RECT 16.31 1.975 16.345 3.283 ;
      RECT 16.295 1.975 16.31 3.265 ;
      RECT 16.275 1.975 16.295 3.255 ;
      RECT 16.25 1.975 16.275 3.238 ;
      RECT 16.245 1.975 16.25 3.188 ;
      RECT 16.235 1.975 16.24 3.018 ;
      RECT 16.23 1.975 16.235 2.925 ;
      RECT 16.225 1.975 16.23 2.838 ;
      RECT 16.22 1.975 16.225 2.77 ;
      RECT 16.215 1.975 16.22 2.713 ;
      RECT 16.205 1.975 16.215 2.608 ;
      RECT 16.2 1.975 16.205 2.48 ;
      RECT 16.195 1.975 16.2 2.398 ;
      RECT 16.19 1.977 16.195 2.315 ;
      RECT 16.185 1.982 16.19 2.248 ;
      RECT 16.18 1.987 16.185 2.175 ;
      RECT 18.995 2.305 19.255 2.565 ;
      RECT 19.015 2.272 19.225 2.565 ;
      RECT 19.015 2.27 19.215 2.565 ;
      RECT 19.025 2.257 19.215 2.565 ;
      RECT 19.025 2.255 19.14 2.565 ;
      RECT 18.5 2.38 18.675 2.66 ;
      RECT 18.495 2.38 18.675 2.658 ;
      RECT 18.495 2.38 18.69 2.655 ;
      RECT 18.485 2.38 18.69 2.653 ;
      RECT 18.43 2.38 18.69 2.64 ;
      RECT 18.43 2.455 18.695 2.618 ;
      RECT 17.975 2.392 17.995 2.635 ;
      RECT 17.975 2.392 18.035 2.634 ;
      RECT 17.97 2.394 18.035 2.633 ;
      RECT 17.97 2.394 18.121 2.632 ;
      RECT 17.97 2.394 18.19 2.631 ;
      RECT 17.97 2.394 18.21 2.623 ;
      RECT 17.95 2.397 18.21 2.621 ;
      RECT 17.935 2.407 18.21 2.606 ;
      RECT 17.935 2.407 18.225 2.605 ;
      RECT 17.93 2.416 18.225 2.597 ;
      RECT 17.93 2.416 18.23 2.593 ;
      RECT 18.035 2.33 18.295 2.59 ;
      RECT 17.925 2.418 18.295 2.475 ;
      RECT 17.995 2.385 18.295 2.59 ;
      RECT 17.96 3.578 17.965 3.785 ;
      RECT 17.91 3.572 17.96 3.784 ;
      RECT 17.877 3.586 17.97 3.783 ;
      RECT 17.791 3.586 17.97 3.782 ;
      RECT 17.705 3.586 17.97 3.781 ;
      RECT 17.705 3.685 17.975 3.778 ;
      RECT 17.7 3.685 17.975 3.773 ;
      RECT 17.695 3.685 17.975 3.755 ;
      RECT 17.69 3.685 17.975 3.738 ;
      RECT 17.65 3.47 17.91 3.73 ;
      RECT 17.11 2.62 17.196 3.034 ;
      RECT 17.11 2.62 17.235 3.031 ;
      RECT 17.11 2.62 17.255 3.021 ;
      RECT 17.065 2.62 17.255 3.018 ;
      RECT 17.065 2.772 17.265 3.008 ;
      RECT 17.065 2.793 17.27 3.002 ;
      RECT 17.065 2.811 17.275 2.998 ;
      RECT 17.065 2.831 17.285 2.993 ;
      RECT 17.04 2.831 17.285 2.99 ;
      RECT 17.03 2.831 17.285 2.968 ;
      RECT 17.03 2.847 17.29 2.938 ;
      RECT 16.995 2.62 17.255 2.925 ;
      RECT 16.995 2.859 17.295 2.88 ;
      RECT 14.66 7.765 14.95 7.995 ;
      RECT 14.72 6.285 14.89 7.995 ;
      RECT 14.71 6.655 15.06 7.005 ;
      RECT 14.66 6.285 14.95 6.515 ;
      RECT 14.66 2.365 14.95 2.595 ;
      RECT 14.72 0.885 14.89 2.595 ;
      RECT 14.66 0.885 14.95 1.115 ;
      RECT 14.25 2.735 14.58 2.965 ;
      RECT 14.25 2.765 14.75 2.935 ;
      RECT 14.25 2.395 14.44 2.965 ;
      RECT 13.67 2.365 13.96 2.595 ;
      RECT 13.67 2.395 14.44 2.565 ;
      RECT 13.73 0.885 13.9 2.595 ;
      RECT 13.67 0.885 13.96 1.115 ;
      RECT 13.67 7.765 13.96 7.995 ;
      RECT 13.73 6.285 13.9 7.995 ;
      RECT 13.67 6.285 13.96 6.515 ;
      RECT 13.67 6.325 14.52 6.485 ;
      RECT 14.35 5.915 14.52 6.485 ;
      RECT 13.67 6.32 14.06 6.485 ;
      RECT 14.29 5.915 14.58 6.145 ;
      RECT 14.29 5.945 14.75 6.115 ;
      RECT 13.3 2.735 13.59 2.965 ;
      RECT 13.3 2.765 13.76 2.935 ;
      RECT 13.36 1.655 13.525 2.965 ;
      RECT 11.875 1.625 12.165 1.855 ;
      RECT 11.875 1.655 13.525 1.825 ;
      RECT 11.935 0.885 12.105 1.855 ;
      RECT 11.875 0.885 12.165 1.115 ;
      RECT 11.875 7.765 12.165 7.995 ;
      RECT 11.935 7.025 12.105 7.995 ;
      RECT 11.935 7.12 13.525 7.29 ;
      RECT 13.355 5.915 13.525 7.29 ;
      RECT 11.875 7.025 12.165 7.255 ;
      RECT 13.3 5.915 13.59 6.145 ;
      RECT 13.3 5.945 13.76 6.115 ;
      RECT 9.925 2.705 10.265 3.055 ;
      RECT 10.015 2.025 10.185 3.055 ;
      RECT 12.305 1.965 12.655 2.315 ;
      RECT 10.015 2.025 12.655 2.195 ;
      RECT 12.33 6.655 12.655 6.98 ;
      RECT 6.87 6.605 7.22 6.955 ;
      RECT 12.305 6.655 12.655 6.885 ;
      RECT 6.67 6.655 7.22 6.885 ;
      RECT 6.5 6.685 12.655 6.855 ;
      RECT 11.53 2.365 11.85 2.685 ;
      RECT 11.5 2.365 11.85 2.595 ;
      RECT 11.33 2.395 11.85 2.565 ;
      RECT 11.53 6.255 11.85 6.545 ;
      RECT 11.5 6.285 11.85 6.515 ;
      RECT 11.33 6.315 11.85 6.485 ;
      RECT 10.485 2.705 10.825 3.055 ;
      RECT 10.485 2.765 10.965 2.935 ;
      RECT 10.48 5.86 10.82 6.21 ;
      RECT 4.87 5.915 5.16 6.145 ;
      RECT 4.87 5.945 10.965 6.115 ;
      RECT 7.22 2.985 7.37 3.26 ;
      RECT 7.76 2.065 7.765 2.285 ;
      RECT 8.91 2.265 8.925 2.463 ;
      RECT 8.875 2.257 8.91 2.47 ;
      RECT 8.845 2.25 8.875 2.47 ;
      RECT 8.79 2.215 8.845 2.47 ;
      RECT 8.725 2.152 8.79 2.47 ;
      RECT 8.72 2.117 8.725 2.468 ;
      RECT 8.715 2.112 8.72 2.46 ;
      RECT 8.71 2.107 8.715 2.446 ;
      RECT 8.705 2.104 8.71 2.439 ;
      RECT 8.66 2.094 8.705 2.39 ;
      RECT 8.64 2.081 8.66 2.325 ;
      RECT 8.635 2.076 8.64 2.298 ;
      RECT 8.63 2.075 8.635 2.291 ;
      RECT 8.625 2.074 8.63 2.284 ;
      RECT 8.54 2.059 8.625 2.23 ;
      RECT 8.51 2.04 8.54 2.18 ;
      RECT 8.43 2.023 8.51 2.165 ;
      RECT 8.395 2.01 8.43 2.15 ;
      RECT 8.387 2.01 8.395 2.145 ;
      RECT 8.301 2.011 8.387 2.145 ;
      RECT 8.215 2.013 8.301 2.145 ;
      RECT 8.19 2.014 8.215 2.149 ;
      RECT 8.115 2.02 8.19 2.164 ;
      RECT 8.032 2.032 8.115 2.188 ;
      RECT 7.946 2.045 8.032 2.214 ;
      RECT 7.86 2.058 7.946 2.24 ;
      RECT 7.825 2.067 7.86 2.259 ;
      RECT 7.775 2.067 7.825 2.272 ;
      RECT 7.765 2.065 7.775 2.283 ;
      RECT 7.75 2.062 7.76 2.285 ;
      RECT 7.735 2.054 7.75 2.293 ;
      RECT 7.72 2.046 7.735 2.313 ;
      RECT 7.715 2.041 7.72 2.37 ;
      RECT 7.7 2.036 7.715 2.443 ;
      RECT 7.695 2.031 7.7 2.485 ;
      RECT 7.69 2.029 7.695 2.513 ;
      RECT 7.685 2.027 7.69 2.535 ;
      RECT 7.675 2.023 7.685 2.578 ;
      RECT 7.67 2.02 7.675 2.603 ;
      RECT 7.665 2.018 7.67 2.623 ;
      RECT 7.66 2.016 7.665 2.647 ;
      RECT 7.655 2.012 7.66 2.67 ;
      RECT 7.65 2.008 7.655 2.693 ;
      RECT 7.615 1.998 7.65 2.8 ;
      RECT 7.61 1.988 7.615 2.898 ;
      RECT 7.605 1.986 7.61 2.925 ;
      RECT 7.6 1.985 7.605 2.945 ;
      RECT 7.595 1.977 7.6 2.965 ;
      RECT 7.59 1.972 7.595 3 ;
      RECT 7.585 1.97 7.59 3.018 ;
      RECT 7.58 1.97 7.585 3.043 ;
      RECT 7.575 1.97 7.58 3.065 ;
      RECT 7.54 1.97 7.575 3.108 ;
      RECT 7.515 1.97 7.54 3.137 ;
      RECT 7.505 1.97 7.515 2.323 ;
      RECT 7.508 2.38 7.515 3.147 ;
      RECT 7.505 2.437 7.508 3.15 ;
      RECT 7.5 1.97 7.505 2.295 ;
      RECT 7.5 2.487 7.505 3.153 ;
      RECT 7.49 1.97 7.5 2.285 ;
      RECT 7.495 2.54 7.5 3.156 ;
      RECT 7.49 2.625 7.495 3.16 ;
      RECT 7.48 1.97 7.49 2.273 ;
      RECT 7.485 2.672 7.49 3.164 ;
      RECT 7.48 2.747 7.485 3.168 ;
      RECT 7.445 1.97 7.48 2.248 ;
      RECT 7.47 2.83 7.48 3.173 ;
      RECT 7.46 2.897 7.47 3.18 ;
      RECT 7.455 2.925 7.46 3.185 ;
      RECT 7.445 2.938 7.455 3.191 ;
      RECT 7.4 1.97 7.445 2.205 ;
      RECT 7.44 2.943 7.445 3.198 ;
      RECT 7.4 2.96 7.44 3.26 ;
      RECT 7.395 1.972 7.4 2.178 ;
      RECT 7.37 2.98 7.4 3.26 ;
      RECT 7.39 1.977 7.395 2.15 ;
      RECT 7.18 2.989 7.22 3.26 ;
      RECT 7.155 2.997 7.18 3.23 ;
      RECT 7.11 3.005 7.155 3.23 ;
      RECT 7.095 3.01 7.11 3.225 ;
      RECT 7.085 3.01 7.095 3.219 ;
      RECT 7.075 3.017 7.085 3.216 ;
      RECT 7.07 3.055 7.075 3.205 ;
      RECT 7.065 3.117 7.07 3.183 ;
      RECT 8.335 2.992 8.52 3.215 ;
      RECT 8.335 3.007 8.525 3.211 ;
      RECT 8.325 2.28 8.41 3.21 ;
      RECT 8.325 3.007 8.53 3.204 ;
      RECT 8.32 3.015 8.53 3.203 ;
      RECT 8.525 2.735 8.845 3.055 ;
      RECT 8.32 2.907 8.49 2.998 ;
      RECT 8.315 2.907 8.49 2.98 ;
      RECT 8.305 2.715 8.44 2.955 ;
      RECT 8.3 2.715 8.44 2.9 ;
      RECT 8.26 2.295 8.43 2.8 ;
      RECT 8.245 2.295 8.43 2.67 ;
      RECT 8.24 2.295 8.43 2.623 ;
      RECT 8.235 2.295 8.43 2.603 ;
      RECT 8.23 2.295 8.43 2.578 ;
      RECT 8.2 2.295 8.46 2.555 ;
      RECT 8.21 2.292 8.42 2.555 ;
      RECT 8.335 2.287 8.42 3.215 ;
      RECT 8.22 2.28 8.41 2.555 ;
      RECT 8.215 2.285 8.41 2.555 ;
      RECT 7.045 2.497 7.23 2.71 ;
      RECT 7.045 2.505 7.24 2.703 ;
      RECT 7.025 2.505 7.24 2.7 ;
      RECT 7.02 2.505 7.24 2.685 ;
      RECT 6.95 2.42 7.21 2.68 ;
      RECT 6.95 2.565 7.245 2.593 ;
      RECT 6.605 3.02 6.865 3.28 ;
      RECT 6.63 2.965 6.825 3.28 ;
      RECT 6.625 2.714 6.805 3.008 ;
      RECT 6.625 2.72 6.815 3.008 ;
      RECT 6.605 2.722 6.815 2.953 ;
      RECT 6.6 2.732 6.815 2.82 ;
      RECT 6.63 2.712 6.805 3.28 ;
      RECT 6.716 2.71 6.805 3.28 ;
      RECT 6.575 1.93 6.61 2.3 ;
      RECT 6.365 2.04 6.37 2.3 ;
      RECT 6.61 1.937 6.625 2.3 ;
      RECT 6.5 1.93 6.575 2.378 ;
      RECT 6.49 1.93 6.5 2.463 ;
      RECT 6.465 1.93 6.49 2.498 ;
      RECT 6.425 1.93 6.465 2.566 ;
      RECT 6.415 1.937 6.425 2.618 ;
      RECT 6.385 2.04 6.415 2.659 ;
      RECT 6.38 2.04 6.385 2.698 ;
      RECT 6.37 2.04 6.38 2.718 ;
      RECT 6.365 2.335 6.37 2.755 ;
      RECT 6.36 2.352 6.365 2.775 ;
      RECT 6.345 2.415 6.36 2.815 ;
      RECT 6.34 2.458 6.345 2.85 ;
      RECT 6.335 2.466 6.34 2.863 ;
      RECT 6.325 2.48 6.335 2.885 ;
      RECT 6.3 2.515 6.325 2.95 ;
      RECT 6.29 2.55 6.3 3.013 ;
      RECT 6.27 2.58 6.29 3.074 ;
      RECT 6.255 2.616 6.27 3.141 ;
      RECT 6.245 2.644 6.255 3.18 ;
      RECT 6.235 2.666 6.245 3.2 ;
      RECT 6.23 2.676 6.235 3.211 ;
      RECT 6.225 2.685 6.23 3.214 ;
      RECT 6.215 2.703 6.225 3.218 ;
      RECT 6.205 2.721 6.215 3.219 ;
      RECT 6.18 2.76 6.205 3.216 ;
      RECT 6.16 2.802 6.18 3.213 ;
      RECT 6.145 2.84 6.16 3.212 ;
      RECT 6.11 2.875 6.145 3.209 ;
      RECT 6.105 2.897 6.11 3.207 ;
      RECT 6.04 2.937 6.105 3.204 ;
      RECT 6.035 2.977 6.04 3.2 ;
      RECT 6.02 2.987 6.035 3.191 ;
      RECT 6.01 3.107 6.02 3.176 ;
      RECT 6.49 3.52 6.5 3.78 ;
      RECT 6.49 3.523 6.51 3.779 ;
      RECT 6.48 3.513 6.49 3.778 ;
      RECT 6.47 3.528 6.55 3.774 ;
      RECT 6.455 3.507 6.47 3.772 ;
      RECT 6.43 3.532 6.555 3.768 ;
      RECT 6.415 3.492 6.43 3.763 ;
      RECT 6.415 3.534 6.565 3.762 ;
      RECT 6.415 3.542 6.58 3.755 ;
      RECT 6.355 3.479 6.415 3.745 ;
      RECT 6.345 3.466 6.355 3.727 ;
      RECT 6.32 3.456 6.345 3.717 ;
      RECT 6.315 3.446 6.32 3.709 ;
      RECT 6.25 3.542 6.58 3.691 ;
      RECT 6.165 3.542 6.58 3.653 ;
      RECT 6.055 3.37 6.315 3.63 ;
      RECT 6.43 3.5 6.455 3.768 ;
      RECT 6.47 3.51 6.48 3.774 ;
      RECT 6.055 3.518 6.495 3.63 ;
      RECT 6.24 7.765 6.53 7.995 ;
      RECT 6.3 7.025 6.47 7.995 ;
      RECT 6.2 7.055 6.57 7.425 ;
      RECT 6.24 7.025 6.53 7.425 ;
      RECT 5.27 3.275 5.3 3.575 ;
      RECT 5.045 3.26 5.05 3.535 ;
      RECT 4.845 3.26 5 3.52 ;
      RECT 6.145 1.975 6.175 2.235 ;
      RECT 6.135 1.975 6.145 2.343 ;
      RECT 6.115 1.975 6.135 2.353 ;
      RECT 6.1 1.975 6.115 2.365 ;
      RECT 6.045 1.975 6.1 2.415 ;
      RECT 6.03 1.975 6.045 2.463 ;
      RECT 6 1.975 6.03 2.498 ;
      RECT 5.945 1.975 6 2.56 ;
      RECT 5.925 1.975 5.945 2.628 ;
      RECT 5.92 1.975 5.925 2.658 ;
      RECT 5.915 1.975 5.92 2.67 ;
      RECT 5.91 2.092 5.915 2.688 ;
      RECT 5.89 2.11 5.91 2.713 ;
      RECT 5.87 2.137 5.89 2.763 ;
      RECT 5.865 2.157 5.87 2.794 ;
      RECT 5.86 2.165 5.865 2.811 ;
      RECT 5.845 2.191 5.86 2.84 ;
      RECT 5.83 2.233 5.845 2.875 ;
      RECT 5.825 2.262 5.83 2.898 ;
      RECT 5.82 2.277 5.825 2.911 ;
      RECT 5.815 2.3 5.82 2.922 ;
      RECT 5.805 2.32 5.815 2.94 ;
      RECT 5.795 2.35 5.805 2.963 ;
      RECT 5.79 2.372 5.795 2.983 ;
      RECT 5.785 2.387 5.79 2.998 ;
      RECT 5.77 2.417 5.785 3.025 ;
      RECT 5.765 2.447 5.77 3.051 ;
      RECT 5.76 2.465 5.765 3.063 ;
      RECT 5.75 2.495 5.76 3.082 ;
      RECT 5.74 2.52 5.75 3.107 ;
      RECT 5.735 2.54 5.74 3.126 ;
      RECT 5.73 2.557 5.735 3.139 ;
      RECT 5.72 2.583 5.73 3.158 ;
      RECT 5.71 2.621 5.72 3.185 ;
      RECT 5.705 2.647 5.71 3.205 ;
      RECT 5.7 2.657 5.705 3.215 ;
      RECT 5.695 2.67 5.7 3.23 ;
      RECT 5.69 2.685 5.695 3.24 ;
      RECT 5.685 2.707 5.69 3.255 ;
      RECT 5.68 2.725 5.685 3.266 ;
      RECT 5.675 2.735 5.68 3.277 ;
      RECT 5.67 2.743 5.675 3.289 ;
      RECT 5.665 2.751 5.67 3.3 ;
      RECT 5.66 2.777 5.665 3.313 ;
      RECT 5.65 2.805 5.66 3.326 ;
      RECT 5.645 2.835 5.65 3.335 ;
      RECT 5.64 2.85 5.645 3.342 ;
      RECT 5.625 2.875 5.64 3.349 ;
      RECT 5.62 2.897 5.625 3.355 ;
      RECT 5.615 2.922 5.62 3.358 ;
      RECT 5.606 2.95 5.615 3.362 ;
      RECT 5.6 2.967 5.606 3.367 ;
      RECT 5.595 2.985 5.6 3.371 ;
      RECT 5.59 2.997 5.595 3.374 ;
      RECT 5.585 3.018 5.59 3.378 ;
      RECT 5.58 3.036 5.585 3.381 ;
      RECT 5.575 3.05 5.58 3.384 ;
      RECT 5.57 3.067 5.575 3.387 ;
      RECT 5.565 3.08 5.57 3.39 ;
      RECT 5.54 3.117 5.565 3.398 ;
      RECT 5.535 3.162 5.54 3.407 ;
      RECT 5.53 3.19 5.535 3.41 ;
      RECT 5.52 3.21 5.53 3.414 ;
      RECT 5.515 3.23 5.52 3.419 ;
      RECT 5.51 3.245 5.515 3.422 ;
      RECT 5.49 3.255 5.51 3.429 ;
      RECT 5.425 3.262 5.49 3.455 ;
      RECT 5.39 3.265 5.425 3.483 ;
      RECT 5.375 3.268 5.39 3.498 ;
      RECT 5.365 3.269 5.375 3.513 ;
      RECT 5.355 3.27 5.365 3.53 ;
      RECT 5.35 3.27 5.355 3.545 ;
      RECT 5.345 3.27 5.35 3.553 ;
      RECT 5.33 3.271 5.345 3.568 ;
      RECT 5.3 3.273 5.33 3.575 ;
      RECT 5.19 3.28 5.27 3.575 ;
      RECT 5.145 3.285 5.19 3.575 ;
      RECT 5.135 3.286 5.145 3.565 ;
      RECT 5.125 3.287 5.135 3.558 ;
      RECT 5.105 3.289 5.125 3.553 ;
      RECT 5.095 3.26 5.105 3.548 ;
      RECT 5.05 3.26 5.095 3.54 ;
      RECT 5.02 3.26 5.045 3.53 ;
      RECT 5 3.26 5.02 3.523 ;
      RECT 5.28 2.06 5.54 2.32 ;
      RECT 5.16 2.075 5.17 2.24 ;
      RECT 5.145 2.075 5.15 2.235 ;
      RECT 2.51 1.915 2.695 2.205 ;
      RECT 4.325 2.04 4.34 2.195 ;
      RECT 2.475 1.915 2.5 2.175 ;
      RECT 4.89 1.965 4.895 2.107 ;
      RECT 4.805 1.96 4.83 2.1 ;
      RECT 5.205 2.077 5.28 2.27 ;
      RECT 5.19 2.075 5.205 2.253 ;
      RECT 5.17 2.075 5.19 2.245 ;
      RECT 5.15 2.075 5.16 2.238 ;
      RECT 5.105 2.07 5.145 2.228 ;
      RECT 5.065 2.045 5.105 2.213 ;
      RECT 5.05 2.02 5.065 2.203 ;
      RECT 5.045 2.014 5.05 2.201 ;
      RECT 5.01 2.006 5.045 2.184 ;
      RECT 5.005 1.999 5.01 2.172 ;
      RECT 4.985 1.994 5.005 2.16 ;
      RECT 4.975 1.988 4.985 2.145 ;
      RECT 4.955 1.983 4.975 2.13 ;
      RECT 4.945 1.978 4.955 2.123 ;
      RECT 4.94 1.976 4.945 2.118 ;
      RECT 4.935 1.975 4.94 2.115 ;
      RECT 4.895 1.97 4.935 2.111 ;
      RECT 4.875 1.964 4.89 2.106 ;
      RECT 4.84 1.961 4.875 2.103 ;
      RECT 4.83 1.96 4.84 2.101 ;
      RECT 4.77 1.96 4.805 2.098 ;
      RECT 4.725 1.96 4.77 2.098 ;
      RECT 4.675 1.96 4.725 2.101 ;
      RECT 4.66 1.962 4.675 2.103 ;
      RECT 4.645 1.965 4.66 2.104 ;
      RECT 4.635 1.97 4.645 2.105 ;
      RECT 4.605 1.975 4.635 2.11 ;
      RECT 4.595 1.981 4.605 2.118 ;
      RECT 4.585 1.983 4.595 2.122 ;
      RECT 4.575 1.987 4.585 2.126 ;
      RECT 4.55 1.993 4.575 2.134 ;
      RECT 4.54 1.998 4.55 2.142 ;
      RECT 4.525 2.002 4.54 2.146 ;
      RECT 4.49 2.008 4.525 2.154 ;
      RECT 4.47 2.013 4.49 2.164 ;
      RECT 4.44 2.02 4.47 2.173 ;
      RECT 4.395 2.029 4.44 2.187 ;
      RECT 4.39 2.034 4.395 2.198 ;
      RECT 4.37 2.037 4.39 2.199 ;
      RECT 4.34 2.04 4.37 2.197 ;
      RECT 4.305 2.04 4.325 2.193 ;
      RECT 4.235 2.04 4.305 2.184 ;
      RECT 4.22 2.037 4.235 2.176 ;
      RECT 4.18 2.03 4.22 2.171 ;
      RECT 4.155 2.02 4.18 2.164 ;
      RECT 4.15 2.014 4.155 2.161 ;
      RECT 4.11 2.008 4.15 2.158 ;
      RECT 4.095 2.001 4.11 2.153 ;
      RECT 4.075 1.997 4.095 2.148 ;
      RECT 4.06 1.992 4.075 2.144 ;
      RECT 4.045 1.987 4.06 2.142 ;
      RECT 4.03 1.983 4.045 2.141 ;
      RECT 4.015 1.981 4.03 2.137 ;
      RECT 4.005 1.979 4.015 2.132 ;
      RECT 3.99 1.976 4.005 2.128 ;
      RECT 3.98 1.974 3.99 2.123 ;
      RECT 3.96 1.971 3.98 2.119 ;
      RECT 3.915 1.97 3.96 2.117 ;
      RECT 3.855 1.972 3.915 2.118 ;
      RECT 3.835 1.974 3.855 2.12 ;
      RECT 3.805 1.977 3.835 2.121 ;
      RECT 3.755 1.982 3.805 2.123 ;
      RECT 3.75 1.985 3.755 2.125 ;
      RECT 3.74 1.987 3.75 2.128 ;
      RECT 3.735 1.989 3.74 2.131 ;
      RECT 3.685 1.992 3.735 2.138 ;
      RECT 3.665 1.996 3.685 2.15 ;
      RECT 3.655 1.999 3.665 2.156 ;
      RECT 3.645 2 3.655 2.159 ;
      RECT 3.606 2.003 3.645 2.161 ;
      RECT 3.52 2.01 3.606 2.164 ;
      RECT 3.446 2.02 3.52 2.168 ;
      RECT 3.36 2.031 3.446 2.173 ;
      RECT 3.345 2.038 3.36 2.175 ;
      RECT 3.29 2.042 3.345 2.176 ;
      RECT 3.276 2.045 3.29 2.178 ;
      RECT 3.19 2.045 3.276 2.18 ;
      RECT 3.15 2.042 3.19 2.183 ;
      RECT 3.126 2.038 3.15 2.185 ;
      RECT 3.04 2.028 3.126 2.188 ;
      RECT 3.01 2.017 3.04 2.189 ;
      RECT 2.991 2.013 3.01 2.188 ;
      RECT 2.905 2.006 2.991 2.185 ;
      RECT 2.845 1.995 2.905 2.182 ;
      RECT 2.825 1.987 2.845 2.18 ;
      RECT 2.79 1.982 2.825 2.179 ;
      RECT 2.765 1.977 2.79 2.178 ;
      RECT 2.735 1.972 2.765 2.177 ;
      RECT 2.71 1.915 2.735 2.176 ;
      RECT 2.695 1.915 2.71 2.2 ;
      RECT 2.5 1.915 2.51 2.2 ;
      RECT 4.275 2.935 4.28 3.075 ;
      RECT 3.935 2.935 3.97 3.073 ;
      RECT 3.51 2.92 3.525 3.065 ;
      RECT 5.34 2.7 5.43 2.96 ;
      RECT 5.17 2.565 5.27 2.96 ;
      RECT 2.205 2.54 2.285 2.75 ;
      RECT 5.295 2.677 5.34 2.96 ;
      RECT 5.285 2.647 5.295 2.96 ;
      RECT 5.27 2.57 5.285 2.96 ;
      RECT 5.085 2.565 5.17 2.925 ;
      RECT 5.08 2.567 5.085 2.92 ;
      RECT 5.075 2.572 5.08 2.92 ;
      RECT 5.04 2.672 5.075 2.92 ;
      RECT 5.03 2.7 5.04 2.92 ;
      RECT 5.02 2.715 5.03 2.92 ;
      RECT 5.01 2.727 5.02 2.92 ;
      RECT 5.005 2.737 5.01 2.92 ;
      RECT 4.99 2.747 5.005 2.922 ;
      RECT 4.985 2.762 4.99 2.924 ;
      RECT 4.97 2.775 4.985 2.926 ;
      RECT 4.965 2.79 4.97 2.929 ;
      RECT 4.945 2.8 4.965 2.933 ;
      RECT 4.93 2.81 4.945 2.936 ;
      RECT 4.895 2.817 4.93 2.941 ;
      RECT 4.851 2.824 4.895 2.949 ;
      RECT 4.765 2.836 4.851 2.962 ;
      RECT 4.74 2.847 4.765 2.973 ;
      RECT 4.71 2.852 4.74 2.978 ;
      RECT 4.675 2.857 4.71 2.986 ;
      RECT 4.645 2.862 4.675 2.993 ;
      RECT 4.62 2.867 4.645 2.998 ;
      RECT 4.555 2.874 4.62 3.007 ;
      RECT 4.485 2.887 4.555 3.023 ;
      RECT 4.455 2.897 4.485 3.035 ;
      RECT 4.43 2.902 4.455 3.042 ;
      RECT 4.375 2.909 4.43 3.05 ;
      RECT 4.37 2.916 4.375 3.055 ;
      RECT 4.365 2.918 4.37 3.056 ;
      RECT 4.35 2.92 4.365 3.058 ;
      RECT 4.345 2.92 4.35 3.061 ;
      RECT 4.28 2.927 4.345 3.068 ;
      RECT 4.245 2.937 4.275 3.078 ;
      RECT 4.228 2.94 4.245 3.08 ;
      RECT 4.142 2.939 4.228 3.079 ;
      RECT 4.056 2.937 4.142 3.076 ;
      RECT 3.97 2.936 4.056 3.074 ;
      RECT 3.869 2.934 3.935 3.073 ;
      RECT 3.783 2.931 3.869 3.071 ;
      RECT 3.697 2.927 3.783 3.069 ;
      RECT 3.611 2.924 3.697 3.068 ;
      RECT 3.525 2.921 3.611 3.066 ;
      RECT 3.425 2.92 3.51 3.063 ;
      RECT 3.375 2.918 3.425 3.061 ;
      RECT 3.355 2.915 3.375 3.059 ;
      RECT 3.335 2.913 3.355 3.056 ;
      RECT 3.31 2.909 3.335 3.053 ;
      RECT 3.265 2.903 3.31 3.048 ;
      RECT 3.225 2.897 3.265 3.04 ;
      RECT 3.2 2.892 3.225 3.033 ;
      RECT 3.145 2.885 3.2 3.025 ;
      RECT 3.121 2.878 3.145 3.018 ;
      RECT 3.035 2.869 3.121 3.008 ;
      RECT 3.005 2.861 3.035 2.998 ;
      RECT 2.975 2.857 3.005 2.993 ;
      RECT 2.97 2.854 2.975 2.99 ;
      RECT 2.965 2.853 2.97 2.99 ;
      RECT 2.89 2.846 2.965 2.983 ;
      RECT 2.851 2.837 2.89 2.972 ;
      RECT 2.765 2.827 2.851 2.96 ;
      RECT 2.725 2.817 2.765 2.948 ;
      RECT 2.686 2.812 2.725 2.941 ;
      RECT 2.6 2.802 2.686 2.93 ;
      RECT 2.56 2.79 2.6 2.919 ;
      RECT 2.525 2.775 2.56 2.912 ;
      RECT 2.515 2.765 2.525 2.909 ;
      RECT 2.495 2.75 2.515 2.907 ;
      RECT 2.465 2.72 2.495 2.903 ;
      RECT 2.455 2.7 2.465 2.898 ;
      RECT 2.45 2.692 2.455 2.895 ;
      RECT 2.445 2.685 2.45 2.893 ;
      RECT 2.43 2.672 2.445 2.886 ;
      RECT 2.425 2.662 2.43 2.878 ;
      RECT 2.42 2.655 2.425 2.873 ;
      RECT 2.415 2.65 2.42 2.869 ;
      RECT 2.4 2.637 2.415 2.861 ;
      RECT 2.395 2.547 2.4 2.85 ;
      RECT 2.39 2.542 2.395 2.843 ;
      RECT 2.315 2.54 2.39 2.803 ;
      RECT 2.285 2.54 2.315 2.758 ;
      RECT 2.19 2.545 2.205 2.745 ;
      RECT 4.675 2.25 4.935 2.51 ;
      RECT 4.66 2.238 4.84 2.475 ;
      RECT 4.655 2.239 4.84 2.473 ;
      RECT 4.64 2.243 4.85 2.463 ;
      RECT 4.635 2.248 4.855 2.433 ;
      RECT 4.64 2.245 4.855 2.463 ;
      RECT 4.655 2.24 4.85 2.473 ;
      RECT 4.675 2.237 4.84 2.51 ;
      RECT 4.675 2.236 4.83 2.51 ;
      RECT 4.7 2.235 4.83 2.51 ;
      RECT 4.26 2.48 4.52 2.74 ;
      RECT 4.135 2.525 4.52 2.735 ;
      RECT 4.125 2.53 4.52 2.73 ;
      RECT 4.14 3.47 4.155 3.78 ;
      RECT 2.735 3.24 2.745 3.37 ;
      RECT 2.515 3.235 2.62 3.37 ;
      RECT 2.43 3.24 2.48 3.37 ;
      RECT 0.98 1.975 0.985 3.08 ;
      RECT 4.235 3.562 4.24 3.698 ;
      RECT 4.23 3.557 4.235 3.758 ;
      RECT 4.225 3.555 4.23 3.771 ;
      RECT 4.21 3.552 4.225 3.773 ;
      RECT 4.205 3.547 4.21 3.775 ;
      RECT 4.2 3.543 4.205 3.778 ;
      RECT 4.185 3.538 4.2 3.78 ;
      RECT 4.155 3.53 4.185 3.78 ;
      RECT 4.116 3.47 4.14 3.78 ;
      RECT 4.03 3.47 4.116 3.777 ;
      RECT 4 3.47 4.03 3.77 ;
      RECT 3.975 3.47 4 3.763 ;
      RECT 3.95 3.47 3.975 3.755 ;
      RECT 3.935 3.47 3.95 3.748 ;
      RECT 3.91 3.47 3.935 3.74 ;
      RECT 3.895 3.47 3.91 3.733 ;
      RECT 3.855 3.48 3.895 3.722 ;
      RECT 3.845 3.475 3.855 3.712 ;
      RECT 3.841 3.474 3.845 3.709 ;
      RECT 3.755 3.466 3.841 3.692 ;
      RECT 3.722 3.455 3.755 3.669 ;
      RECT 3.636 3.444 3.722 3.647 ;
      RECT 3.55 3.428 3.636 3.616 ;
      RECT 3.48 3.413 3.55 3.588 ;
      RECT 3.47 3.406 3.48 3.575 ;
      RECT 3.44 3.403 3.47 3.565 ;
      RECT 3.415 3.399 3.44 3.558 ;
      RECT 3.4 3.396 3.415 3.553 ;
      RECT 3.395 3.395 3.4 3.548 ;
      RECT 3.365 3.39 3.395 3.541 ;
      RECT 3.36 3.385 3.365 3.536 ;
      RECT 3.345 3.382 3.36 3.531 ;
      RECT 3.34 3.377 3.345 3.526 ;
      RECT 3.32 3.372 3.34 3.523 ;
      RECT 3.305 3.367 3.32 3.515 ;
      RECT 3.29 3.361 3.305 3.51 ;
      RECT 3.26 3.352 3.29 3.503 ;
      RECT 3.255 3.345 3.26 3.495 ;
      RECT 3.25 3.343 3.255 3.493 ;
      RECT 3.245 3.342 3.25 3.49 ;
      RECT 3.205 3.335 3.245 3.483 ;
      RECT 3.191 3.325 3.205 3.473 ;
      RECT 3.14 3.314 3.191 3.461 ;
      RECT 3.115 3.3 3.14 3.447 ;
      RECT 3.09 3.289 3.115 3.439 ;
      RECT 3.07 3.278 3.09 3.433 ;
      RECT 3.06 3.272 3.07 3.428 ;
      RECT 3.055 3.27 3.06 3.424 ;
      RECT 3.035 3.265 3.055 3.419 ;
      RECT 3.005 3.255 3.035 3.409 ;
      RECT 3 3.247 3.005 3.402 ;
      RECT 2.985 3.245 3 3.398 ;
      RECT 2.965 3.245 2.985 3.393 ;
      RECT 2.96 3.244 2.965 3.391 ;
      RECT 2.955 3.244 2.96 3.388 ;
      RECT 2.915 3.243 2.955 3.383 ;
      RECT 2.89 3.242 2.915 3.378 ;
      RECT 2.83 3.241 2.89 3.375 ;
      RECT 2.745 3.24 2.83 3.373 ;
      RECT 2.706 3.239 2.735 3.37 ;
      RECT 2.62 3.237 2.706 3.37 ;
      RECT 2.48 3.237 2.515 3.37 ;
      RECT 2.39 3.241 2.43 3.373 ;
      RECT 2.375 3.244 2.39 3.38 ;
      RECT 2.365 3.245 2.375 3.387 ;
      RECT 2.34 3.248 2.365 3.392 ;
      RECT 2.335 3.25 2.34 3.395 ;
      RECT 2.285 3.252 2.335 3.396 ;
      RECT 2.246 3.256 2.285 3.398 ;
      RECT 2.16 3.258 2.246 3.401 ;
      RECT 2.142 3.26 2.16 3.403 ;
      RECT 2.056 3.263 2.142 3.405 ;
      RECT 1.97 3.267 2.056 3.408 ;
      RECT 1.933 3.271 1.97 3.411 ;
      RECT 1.847 3.274 1.933 3.414 ;
      RECT 1.761 3.278 1.847 3.417 ;
      RECT 1.675 3.283 1.761 3.421 ;
      RECT 1.655 3.285 1.675 3.424 ;
      RECT 1.635 3.284 1.655 3.425 ;
      RECT 1.586 3.281 1.635 3.426 ;
      RECT 1.5 3.276 1.586 3.429 ;
      RECT 1.45 3.271 1.5 3.431 ;
      RECT 1.426 3.269 1.45 3.432 ;
      RECT 1.34 3.264 1.426 3.434 ;
      RECT 1.315 3.26 1.34 3.433 ;
      RECT 1.305 3.257 1.315 3.431 ;
      RECT 1.295 3.25 1.305 3.428 ;
      RECT 1.29 3.23 1.295 3.423 ;
      RECT 1.28 3.2 1.29 3.418 ;
      RECT 1.265 3.07 1.28 3.409 ;
      RECT 1.26 3.062 1.265 3.402 ;
      RECT 1.24 3.055 1.26 3.394 ;
      RECT 1.235 3.037 1.24 3.386 ;
      RECT 1.225 3.017 1.235 3.381 ;
      RECT 1.22 2.99 1.225 3.377 ;
      RECT 1.215 2.967 1.22 3.374 ;
      RECT 1.195 2.925 1.215 3.366 ;
      RECT 1.16 2.84 1.195 3.35 ;
      RECT 1.155 2.772 1.16 3.338 ;
      RECT 1.14 2.742 1.155 3.332 ;
      RECT 1.135 1.987 1.14 2.233 ;
      RECT 1.125 2.712 1.14 3.323 ;
      RECT 1.13 1.982 1.135 2.265 ;
      RECT 1.125 1.977 1.13 2.308 ;
      RECT 1.12 1.975 1.125 2.343 ;
      RECT 1.105 2.675 1.125 3.313 ;
      RECT 1.115 1.975 1.12 2.38 ;
      RECT 1.1 1.975 1.115 2.478 ;
      RECT 1.1 2.648 1.105 3.306 ;
      RECT 1.095 1.975 1.1 2.553 ;
      RECT 1.095 2.636 1.1 3.303 ;
      RECT 1.09 1.975 1.095 2.585 ;
      RECT 1.09 2.615 1.095 3.3 ;
      RECT 1.085 1.975 1.09 3.297 ;
      RECT 1.05 1.975 1.085 3.283 ;
      RECT 1.035 1.975 1.05 3.265 ;
      RECT 1.015 1.975 1.035 3.255 ;
      RECT 0.99 1.975 1.015 3.238 ;
      RECT 0.985 1.975 0.99 3.188 ;
      RECT 0.975 1.975 0.98 3.018 ;
      RECT 0.97 1.975 0.975 2.925 ;
      RECT 0.965 1.975 0.97 2.838 ;
      RECT 0.96 1.975 0.965 2.77 ;
      RECT 0.955 1.975 0.96 2.713 ;
      RECT 0.945 1.975 0.955 2.608 ;
      RECT 0.94 1.975 0.945 2.48 ;
      RECT 0.935 1.975 0.94 2.398 ;
      RECT 0.93 1.977 0.935 2.315 ;
      RECT 0.925 1.982 0.93 2.248 ;
      RECT 0.92 1.987 0.925 2.175 ;
      RECT 3.735 2.305 3.995 2.565 ;
      RECT 3.755 2.272 3.965 2.565 ;
      RECT 3.755 2.27 3.955 2.565 ;
      RECT 3.765 2.257 3.955 2.565 ;
      RECT 3.765 2.255 3.88 2.565 ;
      RECT 3.24 2.38 3.415 2.66 ;
      RECT 3.235 2.38 3.415 2.658 ;
      RECT 3.235 2.38 3.43 2.655 ;
      RECT 3.225 2.38 3.43 2.653 ;
      RECT 3.17 2.38 3.43 2.64 ;
      RECT 3.17 2.455 3.435 2.618 ;
      RECT 2.715 2.392 2.735 2.635 ;
      RECT 2.715 2.392 2.775 2.634 ;
      RECT 2.71 2.394 2.775 2.633 ;
      RECT 2.71 2.394 2.861 2.632 ;
      RECT 2.71 2.394 2.93 2.631 ;
      RECT 2.71 2.394 2.95 2.623 ;
      RECT 2.69 2.397 2.95 2.621 ;
      RECT 2.675 2.407 2.95 2.606 ;
      RECT 2.675 2.407 2.965 2.605 ;
      RECT 2.67 2.416 2.965 2.597 ;
      RECT 2.67 2.416 2.97 2.593 ;
      RECT 2.775 2.33 3.035 2.59 ;
      RECT 2.665 2.418 3.035 2.475 ;
      RECT 2.735 2.385 3.035 2.59 ;
      RECT 2.7 3.578 2.705 3.785 ;
      RECT 2.65 3.572 2.7 3.784 ;
      RECT 2.617 3.586 2.71 3.783 ;
      RECT 2.531 3.586 2.71 3.782 ;
      RECT 2.445 3.586 2.71 3.781 ;
      RECT 2.445 3.685 2.715 3.778 ;
      RECT 2.44 3.685 2.715 3.773 ;
      RECT 2.435 3.685 2.715 3.755 ;
      RECT 2.43 3.685 2.715 3.738 ;
      RECT 2.39 3.47 2.65 3.73 ;
      RECT 1.85 2.62 1.936 3.034 ;
      RECT 1.85 2.62 1.975 3.031 ;
      RECT 1.85 2.62 1.995 3.021 ;
      RECT 1.805 2.62 1.995 3.018 ;
      RECT 1.805 2.772 2.005 3.008 ;
      RECT 1.805 2.793 2.01 3.002 ;
      RECT 1.805 2.811 2.015 2.998 ;
      RECT 1.805 2.831 2.025 2.993 ;
      RECT 1.78 2.831 2.025 2.99 ;
      RECT 1.77 2.831 2.025 2.968 ;
      RECT 1.77 2.847 2.03 2.938 ;
      RECT 1.735 2.62 1.995 2.925 ;
      RECT 1.735 2.859 2.035 2.88 ;
      RECT -0.825 6.655 -0.535 6.885 ;
      RECT -0.995 6.685 -0.535 6.855 ;
      RECT -1.255 7.765 -0.965 7.995 ;
      RECT -1.195 7.025 -1.025 7.995 ;
      RECT -1.285 7.025 -0.935 7.315 ;
      RECT -1.66 6.285 -1.31 6.575 ;
      RECT -1.8 6.315 -1.31 6.485 ;
      RECT -2.625 5.915 -2.335 6.145 ;
      RECT -2.625 5.945 -2.165 6.115 ;
      RECT 65.36 3.265 65.62 3.525 ;
      RECT 50.1 3.265 50.36 3.525 ;
      RECT 34.84 3.265 35.1 3.525 ;
      RECT 19.58 3.265 19.84 3.525 ;
      RECT 4.32 3.265 4.58 3.525 ;
    LAYER mcon ;
      RECT 75.76 0.915 75.93 1.085 ;
      RECT 75.76 2.395 75.93 2.565 ;
      RECT 75.76 6.315 75.93 6.485 ;
      RECT 75.76 7.795 75.93 7.965 ;
      RECT 75.41 0.105 75.58 0.275 ;
      RECT 75.41 4.165 75.58 4.335 ;
      RECT 75.41 4.545 75.58 4.715 ;
      RECT 75.41 8.605 75.58 8.775 ;
      RECT 75.39 2.765 75.56 2.935 ;
      RECT 75.39 5.945 75.56 6.115 ;
      RECT 74.77 0.915 74.94 1.085 ;
      RECT 74.77 2.395 74.94 2.565 ;
      RECT 74.77 6.315 74.94 6.485 ;
      RECT 74.77 7.795 74.94 7.965 ;
      RECT 74.42 0.105 74.59 0.275 ;
      RECT 74.42 4.165 74.59 4.335 ;
      RECT 74.42 4.545 74.59 4.715 ;
      RECT 74.42 8.605 74.59 8.775 ;
      RECT 74.4 2.765 74.57 2.935 ;
      RECT 74.4 5.945 74.57 6.115 ;
      RECT 73.715 0.105 73.885 0.275 ;
      RECT 73.715 4.165 73.885 4.335 ;
      RECT 73.715 4.545 73.885 4.715 ;
      RECT 73.715 8.605 73.885 8.775 ;
      RECT 73.405 2.025 73.575 2.195 ;
      RECT 73.405 6.685 73.575 6.855 ;
      RECT 73.035 0.105 73.205 0.275 ;
      RECT 73.035 8.605 73.205 8.775 ;
      RECT 72.975 0.915 73.145 1.085 ;
      RECT 72.975 1.655 73.145 1.825 ;
      RECT 72.975 7.055 73.145 7.225 ;
      RECT 72.975 7.795 73.145 7.965 ;
      RECT 72.6 2.395 72.77 2.565 ;
      RECT 72.6 6.315 72.77 6.485 ;
      RECT 72.355 0.105 72.525 0.275 ;
      RECT 72.355 8.605 72.525 8.775 ;
      RECT 71.675 0.105 71.845 0.275 ;
      RECT 71.675 8.605 71.845 8.775 ;
      RECT 71.605 2.765 71.775 2.935 ;
      RECT 71.605 5.945 71.775 6.115 ;
      RECT 70.215 1.415 70.385 1.585 ;
      RECT 70.215 4.135 70.385 4.305 ;
      RECT 69.775 2.28 69.945 2.45 ;
      RECT 69.755 1.415 69.925 1.585 ;
      RECT 69.755 4.135 69.925 4.305 ;
      RECT 69.38 3.025 69.55 3.195 ;
      RECT 69.295 1.415 69.465 1.585 ;
      RECT 69.295 4.135 69.465 4.305 ;
      RECT 69.27 2.3 69.44 2.47 ;
      RECT 68.835 1.415 69.005 1.585 ;
      RECT 68.835 4.135 69.005 4.305 ;
      RECT 68.45 1.99 68.62 2.16 ;
      RECT 68.375 1.415 68.545 1.585 ;
      RECT 68.375 4.135 68.545 4.305 ;
      RECT 68.135 3.03 68.305 3.2 ;
      RECT 68.09 2.52 68.26 2.69 ;
      RECT 68.08 4.545 68.25 4.715 ;
      RECT 68.08 8.605 68.25 8.775 ;
      RECT 67.915 1.415 68.085 1.585 ;
      RECT 67.915 4.135 68.085 4.305 ;
      RECT 67.77 6.685 67.94 6.855 ;
      RECT 67.665 2.73 67.835 2.9 ;
      RECT 67.475 1.95 67.645 2.12 ;
      RECT 67.455 1.415 67.625 1.585 ;
      RECT 67.455 4.135 67.625 4.305 ;
      RECT 67.425 3.56 67.595 3.73 ;
      RECT 67.4 8.605 67.57 8.775 ;
      RECT 67.34 7.055 67.51 7.225 ;
      RECT 67.34 7.795 67.51 7.965 ;
      RECT 67.09 3 67.26 3.17 ;
      RECT 66.995 1.415 67.165 1.585 ;
      RECT 66.995 2.16 67.165 2.33 ;
      RECT 66.995 4.135 67.165 4.305 ;
      RECT 66.965 6.315 67.135 6.485 ;
      RECT 66.72 8.605 66.89 8.775 ;
      RECT 66.535 1.415 66.705 1.585 ;
      RECT 66.535 4.135 66.705 4.305 ;
      RECT 66.195 3.385 66.365 3.555 ;
      RECT 66.135 2.585 66.305 2.755 ;
      RECT 66.075 1.415 66.245 1.585 ;
      RECT 66.075 4.135 66.245 4.305 ;
      RECT 66.04 8.605 66.21 8.775 ;
      RECT 65.97 5.945 66.14 6.115 ;
      RECT 65.695 2.255 65.865 2.425 ;
      RECT 65.615 1.415 65.785 1.585 ;
      RECT 65.615 4.135 65.785 4.305 ;
      RECT 65.43 3.305 65.6 3.475 ;
      RECT 65.185 2.545 65.355 2.715 ;
      RECT 65.155 1.415 65.325 1.585 ;
      RECT 65.155 4.135 65.325 4.305 ;
      RECT 65.09 3.575 65.26 3.745 ;
      RECT 64.815 2.27 64.985 2.44 ;
      RECT 64.695 1.415 64.865 1.585 ;
      RECT 64.695 4.135 64.865 4.305 ;
      RECT 64.285 2.47 64.455 2.64 ;
      RECT 64.235 1.415 64.405 1.585 ;
      RECT 64.235 4.135 64.405 4.305 ;
      RECT 63.775 1.415 63.945 1.585 ;
      RECT 63.775 4.135 63.945 4.305 ;
      RECT 63.765 2.415 63.935 2.585 ;
      RECT 63.56 2.015 63.73 2.185 ;
      RECT 63.56 3.595 63.73 3.765 ;
      RECT 63.315 1.415 63.485 1.585 ;
      RECT 63.315 4.135 63.485 4.305 ;
      RECT 63.25 2.56 63.42 2.73 ;
      RECT 62.855 1.415 63.025 1.585 ;
      RECT 62.855 4.135 63.025 4.305 ;
      RECT 62.84 2.785 63.01 2.955 ;
      RECT 62.395 1.415 62.565 1.585 ;
      RECT 62.395 4.135 62.565 4.305 ;
      RECT 62.13 3.085 62.3 3.255 ;
      RECT 61.985 1.995 62.155 2.165 ;
      RECT 61.935 1.415 62.105 1.585 ;
      RECT 61.935 4.135 62.105 4.305 ;
      RECT 60.5 0.915 60.67 1.085 ;
      RECT 60.5 2.395 60.67 2.565 ;
      RECT 60.5 6.315 60.67 6.485 ;
      RECT 60.5 7.795 60.67 7.965 ;
      RECT 60.15 0.105 60.32 0.275 ;
      RECT 60.15 4.165 60.32 4.335 ;
      RECT 60.15 4.545 60.32 4.715 ;
      RECT 60.15 8.605 60.32 8.775 ;
      RECT 60.13 2.765 60.3 2.935 ;
      RECT 60.13 5.945 60.3 6.115 ;
      RECT 59.51 0.915 59.68 1.085 ;
      RECT 59.51 2.395 59.68 2.565 ;
      RECT 59.51 6.315 59.68 6.485 ;
      RECT 59.51 7.795 59.68 7.965 ;
      RECT 59.16 0.105 59.33 0.275 ;
      RECT 59.16 4.165 59.33 4.335 ;
      RECT 59.16 4.545 59.33 4.715 ;
      RECT 59.16 8.605 59.33 8.775 ;
      RECT 59.14 2.765 59.31 2.935 ;
      RECT 59.14 5.945 59.31 6.115 ;
      RECT 58.455 0.105 58.625 0.275 ;
      RECT 58.455 4.165 58.625 4.335 ;
      RECT 58.455 4.545 58.625 4.715 ;
      RECT 58.455 8.605 58.625 8.775 ;
      RECT 58.145 2.025 58.315 2.195 ;
      RECT 58.145 6.685 58.315 6.855 ;
      RECT 57.775 0.105 57.945 0.275 ;
      RECT 57.775 8.605 57.945 8.775 ;
      RECT 57.715 0.915 57.885 1.085 ;
      RECT 57.715 1.655 57.885 1.825 ;
      RECT 57.715 7.055 57.885 7.225 ;
      RECT 57.715 7.795 57.885 7.965 ;
      RECT 57.34 2.395 57.51 2.565 ;
      RECT 57.34 6.315 57.51 6.485 ;
      RECT 57.095 0.105 57.265 0.275 ;
      RECT 57.095 8.605 57.265 8.775 ;
      RECT 56.415 0.105 56.585 0.275 ;
      RECT 56.415 8.605 56.585 8.775 ;
      RECT 56.345 2.765 56.515 2.935 ;
      RECT 56.345 5.945 56.515 6.115 ;
      RECT 54.955 1.415 55.125 1.585 ;
      RECT 54.955 4.135 55.125 4.305 ;
      RECT 54.515 2.28 54.685 2.45 ;
      RECT 54.495 1.415 54.665 1.585 ;
      RECT 54.495 4.135 54.665 4.305 ;
      RECT 54.12 3.025 54.29 3.195 ;
      RECT 54.035 1.415 54.205 1.585 ;
      RECT 54.035 4.135 54.205 4.305 ;
      RECT 54.01 2.3 54.18 2.47 ;
      RECT 53.575 1.415 53.745 1.585 ;
      RECT 53.575 4.135 53.745 4.305 ;
      RECT 53.19 1.99 53.36 2.16 ;
      RECT 53.115 1.415 53.285 1.585 ;
      RECT 53.115 4.135 53.285 4.305 ;
      RECT 52.875 3.03 53.045 3.2 ;
      RECT 52.83 2.52 53 2.69 ;
      RECT 52.82 4.545 52.99 4.715 ;
      RECT 52.82 8.605 52.99 8.775 ;
      RECT 52.655 1.415 52.825 1.585 ;
      RECT 52.655 4.135 52.825 4.305 ;
      RECT 52.51 6.685 52.68 6.855 ;
      RECT 52.405 2.73 52.575 2.9 ;
      RECT 52.215 1.95 52.385 2.12 ;
      RECT 52.195 1.415 52.365 1.585 ;
      RECT 52.195 4.135 52.365 4.305 ;
      RECT 52.165 3.56 52.335 3.73 ;
      RECT 52.14 8.605 52.31 8.775 ;
      RECT 52.08 7.055 52.25 7.225 ;
      RECT 52.08 7.795 52.25 7.965 ;
      RECT 51.83 3 52 3.17 ;
      RECT 51.735 1.415 51.905 1.585 ;
      RECT 51.735 2.16 51.905 2.33 ;
      RECT 51.735 4.135 51.905 4.305 ;
      RECT 51.705 6.315 51.875 6.485 ;
      RECT 51.46 8.605 51.63 8.775 ;
      RECT 51.275 1.415 51.445 1.585 ;
      RECT 51.275 4.135 51.445 4.305 ;
      RECT 50.935 3.385 51.105 3.555 ;
      RECT 50.875 2.585 51.045 2.755 ;
      RECT 50.815 1.415 50.985 1.585 ;
      RECT 50.815 4.135 50.985 4.305 ;
      RECT 50.78 8.605 50.95 8.775 ;
      RECT 50.71 5.945 50.88 6.115 ;
      RECT 50.435 2.255 50.605 2.425 ;
      RECT 50.355 1.415 50.525 1.585 ;
      RECT 50.355 4.135 50.525 4.305 ;
      RECT 50.17 3.305 50.34 3.475 ;
      RECT 49.925 2.545 50.095 2.715 ;
      RECT 49.895 1.415 50.065 1.585 ;
      RECT 49.895 4.135 50.065 4.305 ;
      RECT 49.83 3.575 50 3.745 ;
      RECT 49.555 2.27 49.725 2.44 ;
      RECT 49.435 1.415 49.605 1.585 ;
      RECT 49.435 4.135 49.605 4.305 ;
      RECT 49.025 2.47 49.195 2.64 ;
      RECT 48.975 1.415 49.145 1.585 ;
      RECT 48.975 4.135 49.145 4.305 ;
      RECT 48.515 1.415 48.685 1.585 ;
      RECT 48.515 4.135 48.685 4.305 ;
      RECT 48.505 2.415 48.675 2.585 ;
      RECT 48.3 2.015 48.47 2.185 ;
      RECT 48.3 3.595 48.47 3.765 ;
      RECT 48.055 1.415 48.225 1.585 ;
      RECT 48.055 4.135 48.225 4.305 ;
      RECT 47.99 2.56 48.16 2.73 ;
      RECT 47.595 1.415 47.765 1.585 ;
      RECT 47.595 4.135 47.765 4.305 ;
      RECT 47.58 2.785 47.75 2.955 ;
      RECT 47.135 1.415 47.305 1.585 ;
      RECT 47.135 4.135 47.305 4.305 ;
      RECT 46.87 3.085 47.04 3.255 ;
      RECT 46.725 1.995 46.895 2.165 ;
      RECT 46.675 1.415 46.845 1.585 ;
      RECT 46.675 4.135 46.845 4.305 ;
      RECT 45.24 0.915 45.41 1.085 ;
      RECT 45.24 2.395 45.41 2.565 ;
      RECT 45.24 6.315 45.41 6.485 ;
      RECT 45.24 7.795 45.41 7.965 ;
      RECT 44.89 0.105 45.06 0.275 ;
      RECT 44.89 4.165 45.06 4.335 ;
      RECT 44.89 4.545 45.06 4.715 ;
      RECT 44.89 8.605 45.06 8.775 ;
      RECT 44.87 2.765 45.04 2.935 ;
      RECT 44.87 5.945 45.04 6.115 ;
      RECT 44.25 0.915 44.42 1.085 ;
      RECT 44.25 2.395 44.42 2.565 ;
      RECT 44.25 6.315 44.42 6.485 ;
      RECT 44.25 7.795 44.42 7.965 ;
      RECT 43.9 0.105 44.07 0.275 ;
      RECT 43.9 4.165 44.07 4.335 ;
      RECT 43.9 4.545 44.07 4.715 ;
      RECT 43.9 8.605 44.07 8.775 ;
      RECT 43.88 2.765 44.05 2.935 ;
      RECT 43.88 5.945 44.05 6.115 ;
      RECT 43.195 0.105 43.365 0.275 ;
      RECT 43.195 4.165 43.365 4.335 ;
      RECT 43.195 4.545 43.365 4.715 ;
      RECT 43.195 8.605 43.365 8.775 ;
      RECT 42.885 2.025 43.055 2.195 ;
      RECT 42.885 6.685 43.055 6.855 ;
      RECT 42.515 0.105 42.685 0.275 ;
      RECT 42.515 8.605 42.685 8.775 ;
      RECT 42.455 0.915 42.625 1.085 ;
      RECT 42.455 1.655 42.625 1.825 ;
      RECT 42.455 7.055 42.625 7.225 ;
      RECT 42.455 7.795 42.625 7.965 ;
      RECT 42.08 2.395 42.25 2.565 ;
      RECT 42.08 6.315 42.25 6.485 ;
      RECT 41.835 0.105 42.005 0.275 ;
      RECT 41.835 8.605 42.005 8.775 ;
      RECT 41.155 0.105 41.325 0.275 ;
      RECT 41.155 8.605 41.325 8.775 ;
      RECT 41.085 2.765 41.255 2.935 ;
      RECT 41.085 5.945 41.255 6.115 ;
      RECT 39.695 1.415 39.865 1.585 ;
      RECT 39.695 4.135 39.865 4.305 ;
      RECT 39.255 2.28 39.425 2.45 ;
      RECT 39.235 1.415 39.405 1.585 ;
      RECT 39.235 4.135 39.405 4.305 ;
      RECT 38.86 3.025 39.03 3.195 ;
      RECT 38.775 1.415 38.945 1.585 ;
      RECT 38.775 4.135 38.945 4.305 ;
      RECT 38.75 2.3 38.92 2.47 ;
      RECT 38.315 1.415 38.485 1.585 ;
      RECT 38.315 4.135 38.485 4.305 ;
      RECT 37.93 1.99 38.1 2.16 ;
      RECT 37.855 1.415 38.025 1.585 ;
      RECT 37.855 4.135 38.025 4.305 ;
      RECT 37.615 3.03 37.785 3.2 ;
      RECT 37.57 2.52 37.74 2.69 ;
      RECT 37.56 4.545 37.73 4.715 ;
      RECT 37.56 8.605 37.73 8.775 ;
      RECT 37.395 1.415 37.565 1.585 ;
      RECT 37.395 4.135 37.565 4.305 ;
      RECT 37.25 6.685 37.42 6.855 ;
      RECT 37.145 2.73 37.315 2.9 ;
      RECT 36.955 1.95 37.125 2.12 ;
      RECT 36.935 1.415 37.105 1.585 ;
      RECT 36.935 4.135 37.105 4.305 ;
      RECT 36.905 3.56 37.075 3.73 ;
      RECT 36.88 8.605 37.05 8.775 ;
      RECT 36.82 7.055 36.99 7.225 ;
      RECT 36.82 7.795 36.99 7.965 ;
      RECT 36.57 3 36.74 3.17 ;
      RECT 36.475 1.415 36.645 1.585 ;
      RECT 36.475 2.16 36.645 2.33 ;
      RECT 36.475 4.135 36.645 4.305 ;
      RECT 36.445 6.315 36.615 6.485 ;
      RECT 36.2 8.605 36.37 8.775 ;
      RECT 36.015 1.415 36.185 1.585 ;
      RECT 36.015 4.135 36.185 4.305 ;
      RECT 35.675 3.385 35.845 3.555 ;
      RECT 35.615 2.585 35.785 2.755 ;
      RECT 35.555 1.415 35.725 1.585 ;
      RECT 35.555 4.135 35.725 4.305 ;
      RECT 35.52 8.605 35.69 8.775 ;
      RECT 35.45 5.945 35.62 6.115 ;
      RECT 35.175 2.255 35.345 2.425 ;
      RECT 35.095 1.415 35.265 1.585 ;
      RECT 35.095 4.135 35.265 4.305 ;
      RECT 34.91 3.305 35.08 3.475 ;
      RECT 34.665 2.545 34.835 2.715 ;
      RECT 34.635 1.415 34.805 1.585 ;
      RECT 34.635 4.135 34.805 4.305 ;
      RECT 34.57 3.575 34.74 3.745 ;
      RECT 34.295 2.27 34.465 2.44 ;
      RECT 34.175 1.415 34.345 1.585 ;
      RECT 34.175 4.135 34.345 4.305 ;
      RECT 33.765 2.47 33.935 2.64 ;
      RECT 33.715 1.415 33.885 1.585 ;
      RECT 33.715 4.135 33.885 4.305 ;
      RECT 33.255 1.415 33.425 1.585 ;
      RECT 33.255 4.135 33.425 4.305 ;
      RECT 33.245 2.415 33.415 2.585 ;
      RECT 33.04 2.015 33.21 2.185 ;
      RECT 33.04 3.595 33.21 3.765 ;
      RECT 32.795 1.415 32.965 1.585 ;
      RECT 32.795 4.135 32.965 4.305 ;
      RECT 32.73 2.56 32.9 2.73 ;
      RECT 32.335 1.415 32.505 1.585 ;
      RECT 32.335 4.135 32.505 4.305 ;
      RECT 32.32 2.785 32.49 2.955 ;
      RECT 31.875 1.415 32.045 1.585 ;
      RECT 31.875 4.135 32.045 4.305 ;
      RECT 31.61 3.085 31.78 3.255 ;
      RECT 31.465 1.995 31.635 2.165 ;
      RECT 31.415 1.415 31.585 1.585 ;
      RECT 31.415 4.135 31.585 4.305 ;
      RECT 29.98 0.915 30.15 1.085 ;
      RECT 29.98 2.395 30.15 2.565 ;
      RECT 29.98 6.315 30.15 6.485 ;
      RECT 29.98 7.795 30.15 7.965 ;
      RECT 29.63 0.105 29.8 0.275 ;
      RECT 29.63 4.165 29.8 4.335 ;
      RECT 29.63 4.545 29.8 4.715 ;
      RECT 29.63 8.605 29.8 8.775 ;
      RECT 29.61 2.765 29.78 2.935 ;
      RECT 29.61 5.945 29.78 6.115 ;
      RECT 28.99 0.915 29.16 1.085 ;
      RECT 28.99 2.395 29.16 2.565 ;
      RECT 28.99 6.315 29.16 6.485 ;
      RECT 28.99 7.795 29.16 7.965 ;
      RECT 28.64 0.105 28.81 0.275 ;
      RECT 28.64 4.165 28.81 4.335 ;
      RECT 28.64 4.545 28.81 4.715 ;
      RECT 28.64 8.605 28.81 8.775 ;
      RECT 28.62 2.765 28.79 2.935 ;
      RECT 28.62 5.945 28.79 6.115 ;
      RECT 27.935 0.105 28.105 0.275 ;
      RECT 27.935 4.165 28.105 4.335 ;
      RECT 27.935 4.545 28.105 4.715 ;
      RECT 27.935 8.605 28.105 8.775 ;
      RECT 27.625 2.025 27.795 2.195 ;
      RECT 27.625 6.685 27.795 6.855 ;
      RECT 27.255 0.105 27.425 0.275 ;
      RECT 27.255 8.605 27.425 8.775 ;
      RECT 27.195 0.915 27.365 1.085 ;
      RECT 27.195 1.655 27.365 1.825 ;
      RECT 27.195 7.055 27.365 7.225 ;
      RECT 27.195 7.795 27.365 7.965 ;
      RECT 26.82 2.395 26.99 2.565 ;
      RECT 26.82 6.315 26.99 6.485 ;
      RECT 26.575 0.105 26.745 0.275 ;
      RECT 26.575 8.605 26.745 8.775 ;
      RECT 25.895 0.105 26.065 0.275 ;
      RECT 25.895 8.605 26.065 8.775 ;
      RECT 25.825 2.765 25.995 2.935 ;
      RECT 25.825 5.945 25.995 6.115 ;
      RECT 24.435 1.415 24.605 1.585 ;
      RECT 24.435 4.135 24.605 4.305 ;
      RECT 23.995 2.28 24.165 2.45 ;
      RECT 23.975 1.415 24.145 1.585 ;
      RECT 23.975 4.135 24.145 4.305 ;
      RECT 23.6 3.025 23.77 3.195 ;
      RECT 23.515 1.415 23.685 1.585 ;
      RECT 23.515 4.135 23.685 4.305 ;
      RECT 23.49 2.3 23.66 2.47 ;
      RECT 23.055 1.415 23.225 1.585 ;
      RECT 23.055 4.135 23.225 4.305 ;
      RECT 22.67 1.99 22.84 2.16 ;
      RECT 22.595 1.415 22.765 1.585 ;
      RECT 22.595 4.135 22.765 4.305 ;
      RECT 22.355 3.03 22.525 3.2 ;
      RECT 22.31 2.52 22.48 2.69 ;
      RECT 22.3 4.545 22.47 4.715 ;
      RECT 22.3 8.605 22.47 8.775 ;
      RECT 22.135 1.415 22.305 1.585 ;
      RECT 22.135 4.135 22.305 4.305 ;
      RECT 21.99 6.685 22.16 6.855 ;
      RECT 21.885 2.73 22.055 2.9 ;
      RECT 21.695 1.95 21.865 2.12 ;
      RECT 21.675 1.415 21.845 1.585 ;
      RECT 21.675 4.135 21.845 4.305 ;
      RECT 21.645 3.56 21.815 3.73 ;
      RECT 21.62 8.605 21.79 8.775 ;
      RECT 21.56 7.055 21.73 7.225 ;
      RECT 21.56 7.795 21.73 7.965 ;
      RECT 21.31 3 21.48 3.17 ;
      RECT 21.215 1.415 21.385 1.585 ;
      RECT 21.215 2.16 21.385 2.33 ;
      RECT 21.215 4.135 21.385 4.305 ;
      RECT 21.185 6.315 21.355 6.485 ;
      RECT 20.94 8.605 21.11 8.775 ;
      RECT 20.755 1.415 20.925 1.585 ;
      RECT 20.755 4.135 20.925 4.305 ;
      RECT 20.415 3.385 20.585 3.555 ;
      RECT 20.355 2.585 20.525 2.755 ;
      RECT 20.295 1.415 20.465 1.585 ;
      RECT 20.295 4.135 20.465 4.305 ;
      RECT 20.26 8.605 20.43 8.775 ;
      RECT 20.19 5.945 20.36 6.115 ;
      RECT 19.915 2.255 20.085 2.425 ;
      RECT 19.835 1.415 20.005 1.585 ;
      RECT 19.835 4.135 20.005 4.305 ;
      RECT 19.65 3.305 19.82 3.475 ;
      RECT 19.405 2.545 19.575 2.715 ;
      RECT 19.375 1.415 19.545 1.585 ;
      RECT 19.375 4.135 19.545 4.305 ;
      RECT 19.31 3.575 19.48 3.745 ;
      RECT 19.035 2.27 19.205 2.44 ;
      RECT 18.915 1.415 19.085 1.585 ;
      RECT 18.915 4.135 19.085 4.305 ;
      RECT 18.505 2.47 18.675 2.64 ;
      RECT 18.455 1.415 18.625 1.585 ;
      RECT 18.455 4.135 18.625 4.305 ;
      RECT 17.995 1.415 18.165 1.585 ;
      RECT 17.995 4.135 18.165 4.305 ;
      RECT 17.985 2.415 18.155 2.585 ;
      RECT 17.78 2.015 17.95 2.185 ;
      RECT 17.78 3.595 17.95 3.765 ;
      RECT 17.535 1.415 17.705 1.585 ;
      RECT 17.535 4.135 17.705 4.305 ;
      RECT 17.47 2.56 17.64 2.73 ;
      RECT 17.075 1.415 17.245 1.585 ;
      RECT 17.075 4.135 17.245 4.305 ;
      RECT 17.06 2.785 17.23 2.955 ;
      RECT 16.615 1.415 16.785 1.585 ;
      RECT 16.615 4.135 16.785 4.305 ;
      RECT 16.35 3.085 16.52 3.255 ;
      RECT 16.205 1.995 16.375 2.165 ;
      RECT 16.155 1.415 16.325 1.585 ;
      RECT 16.155 4.135 16.325 4.305 ;
      RECT 14.72 0.915 14.89 1.085 ;
      RECT 14.72 2.395 14.89 2.565 ;
      RECT 14.72 6.315 14.89 6.485 ;
      RECT 14.72 7.795 14.89 7.965 ;
      RECT 14.37 0.105 14.54 0.275 ;
      RECT 14.37 4.165 14.54 4.335 ;
      RECT 14.37 4.545 14.54 4.715 ;
      RECT 14.37 8.605 14.54 8.775 ;
      RECT 14.35 2.765 14.52 2.935 ;
      RECT 14.35 5.945 14.52 6.115 ;
      RECT 13.73 0.915 13.9 1.085 ;
      RECT 13.73 2.395 13.9 2.565 ;
      RECT 13.73 6.315 13.9 6.485 ;
      RECT 13.73 7.795 13.9 7.965 ;
      RECT 13.38 0.105 13.55 0.275 ;
      RECT 13.38 4.165 13.55 4.335 ;
      RECT 13.38 4.545 13.55 4.715 ;
      RECT 13.38 8.605 13.55 8.775 ;
      RECT 13.36 2.765 13.53 2.935 ;
      RECT 13.36 5.945 13.53 6.115 ;
      RECT 12.675 0.105 12.845 0.275 ;
      RECT 12.675 4.165 12.845 4.335 ;
      RECT 12.675 4.545 12.845 4.715 ;
      RECT 12.675 8.605 12.845 8.775 ;
      RECT 12.365 2.025 12.535 2.195 ;
      RECT 12.365 6.685 12.535 6.855 ;
      RECT 11.995 0.105 12.165 0.275 ;
      RECT 11.995 8.605 12.165 8.775 ;
      RECT 11.935 0.915 12.105 1.085 ;
      RECT 11.935 1.655 12.105 1.825 ;
      RECT 11.935 7.055 12.105 7.225 ;
      RECT 11.935 7.795 12.105 7.965 ;
      RECT 11.56 2.395 11.73 2.565 ;
      RECT 11.56 6.315 11.73 6.485 ;
      RECT 11.315 0.105 11.485 0.275 ;
      RECT 11.315 8.605 11.485 8.775 ;
      RECT 10.635 0.105 10.805 0.275 ;
      RECT 10.635 8.605 10.805 8.775 ;
      RECT 10.565 2.765 10.735 2.935 ;
      RECT 10.565 5.945 10.735 6.115 ;
      RECT 9.175 1.415 9.345 1.585 ;
      RECT 9.175 4.135 9.345 4.305 ;
      RECT 8.735 2.28 8.905 2.45 ;
      RECT 8.715 1.415 8.885 1.585 ;
      RECT 8.715 4.135 8.885 4.305 ;
      RECT 8.34 3.025 8.51 3.195 ;
      RECT 8.255 1.415 8.425 1.585 ;
      RECT 8.255 4.135 8.425 4.305 ;
      RECT 8.23 2.3 8.4 2.47 ;
      RECT 7.795 1.415 7.965 1.585 ;
      RECT 7.795 4.135 7.965 4.305 ;
      RECT 7.41 1.99 7.58 2.16 ;
      RECT 7.335 1.415 7.505 1.585 ;
      RECT 7.335 4.135 7.505 4.305 ;
      RECT 7.095 3.03 7.265 3.2 ;
      RECT 7.05 2.52 7.22 2.69 ;
      RECT 7.04 4.545 7.21 4.715 ;
      RECT 7.04 8.605 7.21 8.775 ;
      RECT 6.875 1.415 7.045 1.585 ;
      RECT 6.875 4.135 7.045 4.305 ;
      RECT 6.73 6.685 6.9 6.855 ;
      RECT 6.625 2.73 6.795 2.9 ;
      RECT 6.435 1.95 6.605 2.12 ;
      RECT 6.415 1.415 6.585 1.585 ;
      RECT 6.415 4.135 6.585 4.305 ;
      RECT 6.385 3.56 6.555 3.73 ;
      RECT 6.36 8.605 6.53 8.775 ;
      RECT 6.3 7.055 6.47 7.225 ;
      RECT 6.3 7.795 6.47 7.965 ;
      RECT 6.05 3 6.22 3.17 ;
      RECT 5.955 1.415 6.125 1.585 ;
      RECT 5.955 2.16 6.125 2.33 ;
      RECT 5.955 4.135 6.125 4.305 ;
      RECT 5.925 6.315 6.095 6.485 ;
      RECT 5.68 8.605 5.85 8.775 ;
      RECT 5.495 1.415 5.665 1.585 ;
      RECT 5.495 4.135 5.665 4.305 ;
      RECT 5.155 3.385 5.325 3.555 ;
      RECT 5.095 2.585 5.265 2.755 ;
      RECT 5.035 1.415 5.205 1.585 ;
      RECT 5.035 4.135 5.205 4.305 ;
      RECT 5 8.605 5.17 8.775 ;
      RECT 4.93 5.945 5.1 6.115 ;
      RECT 4.655 2.255 4.825 2.425 ;
      RECT 4.575 1.415 4.745 1.585 ;
      RECT 4.575 4.135 4.745 4.305 ;
      RECT 4.39 3.305 4.56 3.475 ;
      RECT 4.145 2.545 4.315 2.715 ;
      RECT 4.115 1.415 4.285 1.585 ;
      RECT 4.115 4.135 4.285 4.305 ;
      RECT 4.05 3.575 4.22 3.745 ;
      RECT 3.775 2.27 3.945 2.44 ;
      RECT 3.655 1.415 3.825 1.585 ;
      RECT 3.655 4.135 3.825 4.305 ;
      RECT 3.245 2.47 3.415 2.64 ;
      RECT 3.195 1.415 3.365 1.585 ;
      RECT 3.195 4.135 3.365 4.305 ;
      RECT 2.735 1.415 2.905 1.585 ;
      RECT 2.735 4.135 2.905 4.305 ;
      RECT 2.725 2.415 2.895 2.585 ;
      RECT 2.52 2.015 2.69 2.185 ;
      RECT 2.52 3.595 2.69 3.765 ;
      RECT 2.275 1.415 2.445 1.585 ;
      RECT 2.275 4.135 2.445 4.305 ;
      RECT 2.21 2.56 2.38 2.73 ;
      RECT 1.815 1.415 1.985 1.585 ;
      RECT 1.815 4.135 1.985 4.305 ;
      RECT 1.8 2.785 1.97 2.955 ;
      RECT 1.355 1.415 1.525 1.585 ;
      RECT 1.355 4.135 1.525 4.305 ;
      RECT 1.09 3.085 1.26 3.255 ;
      RECT 0.945 1.995 1.115 2.165 ;
      RECT 0.895 1.415 1.065 1.585 ;
      RECT 0.895 4.135 1.065 4.305 ;
      RECT -0.455 4.545 -0.285 4.715 ;
      RECT -0.455 8.605 -0.285 8.775 ;
      RECT -0.765 6.685 -0.595 6.855 ;
      RECT -1.135 8.605 -0.965 8.775 ;
      RECT -1.195 7.055 -1.025 7.225 ;
      RECT -1.195 7.795 -1.025 7.965 ;
      RECT -1.57 6.315 -1.4 6.485 ;
      RECT -1.815 8.605 -1.645 8.775 ;
      RECT -2.495 8.605 -2.325 8.775 ;
      RECT -2.565 5.945 -2.395 6.115 ;
    LAYER li ;
      RECT 69.76 0 69.93 2.085 ;
      RECT 68.82 0 68.99 2.085 ;
      RECT 67.86 0 68.03 2.085 ;
      RECT 65.94 0 66.11 2.085 ;
      RECT 64.98 0 65.15 2.085 ;
      RECT 63.06 0 63.23 2.085 ;
      RECT 54.5 0 54.67 2.085 ;
      RECT 53.56 0 53.73 2.085 ;
      RECT 52.6 0 52.77 2.085 ;
      RECT 50.68 0 50.85 2.085 ;
      RECT 49.72 0 49.89 2.085 ;
      RECT 47.8 0 47.97 2.085 ;
      RECT 39.24 0 39.41 2.085 ;
      RECT 38.3 0 38.47 2.085 ;
      RECT 37.34 0 37.51 2.085 ;
      RECT 35.42 0 35.59 2.085 ;
      RECT 34.46 0 34.63 2.085 ;
      RECT 32.54 0 32.71 2.085 ;
      RECT 23.98 0 24.15 2.085 ;
      RECT 23.04 0 23.21 2.085 ;
      RECT 22.08 0 22.25 2.085 ;
      RECT 20.16 0 20.33 2.085 ;
      RECT 19.2 0 19.37 2.085 ;
      RECT 17.28 0 17.45 2.085 ;
      RECT 8.72 0 8.89 2.085 ;
      RECT 7.78 0 7.95 2.085 ;
      RECT 6.82 0 6.99 2.085 ;
      RECT 4.9 0 5.07 2.085 ;
      RECT 3.94 0 4.11 2.085 ;
      RECT 2.02 0 2.19 2.085 ;
      RECT 66.815 0 67.01 1.595 ;
      RECT 63.06 0 63.335 1.595 ;
      RECT 51.555 0 51.75 1.595 ;
      RECT 47.8 0 48.075 1.595 ;
      RECT 36.295 0 36.49 1.595 ;
      RECT 32.54 0 32.815 1.595 ;
      RECT 21.035 0 21.23 1.595 ;
      RECT 17.28 0 17.555 1.595 ;
      RECT 5.775 0 5.97 1.595 ;
      RECT 2.02 0 2.295 1.595 ;
      RECT 61.79 0 70.53 1.585 ;
      RECT 46.53 0 55.27 1.585 ;
      RECT 31.27 0 40.01 1.585 ;
      RECT 16.01 0 24.75 1.585 ;
      RECT 0.75 0 9.49 1.585 ;
      RECT 75.33 0 75.5 0.935 ;
      RECT 74.34 0 74.51 0.935 ;
      RECT 71.595 0 71.765 0.935 ;
      RECT 60.07 0 60.24 0.935 ;
      RECT 59.08 0 59.25 0.935 ;
      RECT 56.335 0 56.505 0.935 ;
      RECT 44.81 0 44.98 0.935 ;
      RECT 43.82 0 43.99 0.935 ;
      RECT 41.075 0 41.245 0.935 ;
      RECT 29.55 0 29.72 0.935 ;
      RECT 28.56 0 28.73 0.935 ;
      RECT 25.815 0 25.985 0.935 ;
      RECT 14.29 0 14.46 0.935 ;
      RECT 13.3 0 13.47 0.935 ;
      RECT 10.555 0 10.725 0.935 ;
      RECT -2.75 0 76.3 0.305 ;
      RECT -0.765 4.14 -0.595 8.305 ;
      RECT 75.33 3.405 75.5 5.475 ;
      RECT 74.34 3.405 74.51 5.475 ;
      RECT 71.595 3.405 71.765 5.475 ;
      RECT 65.96 3.635 66.13 5.475 ;
      RECT 60.07 3.405 60.24 5.475 ;
      RECT 59.08 3.405 59.25 5.475 ;
      RECT 56.335 3.405 56.505 5.475 ;
      RECT 50.7 3.635 50.87 5.475 ;
      RECT 44.81 3.405 44.98 5.475 ;
      RECT 43.82 3.405 43.99 5.475 ;
      RECT 41.075 3.405 41.245 5.475 ;
      RECT 35.44 3.635 35.61 5.475 ;
      RECT 29.55 3.405 29.72 5.475 ;
      RECT 28.56 3.405 28.73 5.475 ;
      RECT 25.815 3.405 25.985 5.475 ;
      RECT 20.18 3.635 20.35 5.475 ;
      RECT 14.29 3.405 14.46 5.475 ;
      RECT 13.3 3.405 13.47 5.475 ;
      RECT 10.555 3.405 10.725 5.475 ;
      RECT 4.92 3.635 5.09 5.475 ;
      RECT -2.575 4.14 -2.405 5.475 ;
      RECT -2.75 4.14 76.3 4.745 ;
      RECT 61.79 4.135 76.3 4.745 ;
      RECT 46.53 4.135 61.04 4.745 ;
      RECT 31.27 4.135 45.78 4.745 ;
      RECT 16.01 4.135 30.52 4.745 ;
      RECT 0.75 4.135 15.26 4.745 ;
      RECT 68.82 3.635 68.99 4.745 ;
      RECT 66.9 3.635 67.07 4.745 ;
      RECT 64.5 3.635 64.67 4.745 ;
      RECT 62.58 3.635 62.75 4.745 ;
      RECT 53.56 3.635 53.73 4.745 ;
      RECT 51.64 3.635 51.81 4.745 ;
      RECT 49.24 3.635 49.41 4.745 ;
      RECT 47.32 3.635 47.49 4.745 ;
      RECT 38.3 3.635 38.47 4.745 ;
      RECT 36.38 3.635 36.55 4.745 ;
      RECT 33.98 3.635 34.15 4.745 ;
      RECT 32.06 3.635 32.23 4.745 ;
      RECT 23.04 3.635 23.21 4.745 ;
      RECT 21.12 3.635 21.29 4.745 ;
      RECT 18.72 3.635 18.89 4.745 ;
      RECT 16.8 3.635 16.97 4.745 ;
      RECT 7.78 3.635 7.95 4.745 ;
      RECT 5.86 3.635 6.03 4.745 ;
      RECT 3.46 3.635 3.63 4.745 ;
      RECT 1.54 3.635 1.71 4.745 ;
      RECT -2.75 8.575 76.3 8.88 ;
      RECT 75.33 7.945 75.5 8.88 ;
      RECT 74.34 7.945 74.51 8.88 ;
      RECT 71.595 7.945 71.765 8.88 ;
      RECT 65.96 7.945 66.13 8.88 ;
      RECT 60.07 7.945 60.24 8.88 ;
      RECT 59.08 7.945 59.25 8.88 ;
      RECT 56.335 7.945 56.505 8.88 ;
      RECT 50.7 7.945 50.87 8.88 ;
      RECT 44.81 7.945 44.98 8.88 ;
      RECT 43.82 7.945 43.99 8.88 ;
      RECT 41.075 7.945 41.245 8.88 ;
      RECT 35.44 7.945 35.61 8.88 ;
      RECT 29.55 7.945 29.72 8.88 ;
      RECT 28.56 7.945 28.73 8.88 ;
      RECT 25.815 7.945 25.985 8.88 ;
      RECT 20.18 7.945 20.35 8.88 ;
      RECT 14.29 7.945 14.46 8.88 ;
      RECT 13.3 7.945 13.47 8.88 ;
      RECT 10.555 7.945 10.725 8.88 ;
      RECT 4.92 7.945 5.09 8.88 ;
      RECT -2.575 7.945 -2.405 8.88 ;
      RECT 75.39 1.74 75.56 2.935 ;
      RECT 75.39 1.74 75.855 1.91 ;
      RECT 75.39 6.97 75.855 7.14 ;
      RECT 75.39 5.945 75.56 7.14 ;
      RECT 74.4 1.74 74.57 2.935 ;
      RECT 74.4 1.74 74.865 1.91 ;
      RECT 74.4 6.97 74.865 7.14 ;
      RECT 74.4 5.945 74.57 7.14 ;
      RECT 72.545 2.635 72.715 3.865 ;
      RECT 72.6 0.855 72.77 2.805 ;
      RECT 72.545 0.575 72.715 1.025 ;
      RECT 72.545 7.855 72.715 8.305 ;
      RECT 72.6 6.075 72.77 8.025 ;
      RECT 72.545 5.015 72.715 6.245 ;
      RECT 72.025 0.575 72.195 3.865 ;
      RECT 72.025 2.075 72.43 2.405 ;
      RECT 72.025 1.235 72.43 1.565 ;
      RECT 72.025 5.015 72.195 8.305 ;
      RECT 72.025 7.315 72.43 7.645 ;
      RECT 72.025 6.475 72.43 6.805 ;
      RECT 69.95 3.126 69.955 3.298 ;
      RECT 69.945 3.119 69.95 3.388 ;
      RECT 69.94 3.113 69.945 3.407 ;
      RECT 69.92 3.107 69.94 3.417 ;
      RECT 69.905 3.102 69.92 3.425 ;
      RECT 69.868 3.096 69.905 3.423 ;
      RECT 69.782 3.082 69.868 3.419 ;
      RECT 69.696 3.064 69.782 3.414 ;
      RECT 69.61 3.045 69.696 3.408 ;
      RECT 69.58 3.033 69.61 3.404 ;
      RECT 69.56 3.027 69.58 3.403 ;
      RECT 69.495 3.025 69.56 3.401 ;
      RECT 69.48 3.025 69.495 3.393 ;
      RECT 69.465 3.025 69.48 3.38 ;
      RECT 69.46 3.025 69.465 3.37 ;
      RECT 69.445 3.025 69.46 3.348 ;
      RECT 69.43 3.025 69.445 3.315 ;
      RECT 69.425 3.025 69.43 3.293 ;
      RECT 69.415 3.025 69.425 3.275 ;
      RECT 69.4 3.025 69.415 3.253 ;
      RECT 69.38 3.025 69.4 3.215 ;
      RECT 69.73 2.31 69.765 2.749 ;
      RECT 69.73 2.31 69.77 2.748 ;
      RECT 69.675 2.37 69.77 2.747 ;
      RECT 69.54 2.542 69.77 2.746 ;
      RECT 69.65 2.42 69.77 2.746 ;
      RECT 69.54 2.542 69.795 2.736 ;
      RECT 69.595 2.487 69.875 2.653 ;
      RECT 69.77 2.281 69.775 2.744 ;
      RECT 69.625 2.457 69.915 2.53 ;
      RECT 69.64 2.44 69.77 2.746 ;
      RECT 69.775 2.28 69.945 2.468 ;
      RECT 69.765 2.283 69.945 2.468 ;
      RECT 69.27 2.16 69.44 2.47 ;
      RECT 69.27 2.16 69.445 2.443 ;
      RECT 69.27 2.16 69.45 2.42 ;
      RECT 69.27 2.16 69.46 2.37 ;
      RECT 69.265 2.265 69.46 2.34 ;
      RECT 69.3 1.835 69.47 2.313 ;
      RECT 69.3 1.835 69.485 2.234 ;
      RECT 69.29 2.045 69.485 2.234 ;
      RECT 69.3 1.845 69.495 2.149 ;
      RECT 69.23 2.587 69.235 2.79 ;
      RECT 69.22 2.575 69.23 2.9 ;
      RECT 69.195 2.575 69.22 2.94 ;
      RECT 69.115 2.575 69.195 3.025 ;
      RECT 69.105 2.575 69.115 3.095 ;
      RECT 69.08 2.575 69.105 3.118 ;
      RECT 69.06 2.575 69.08 3.153 ;
      RECT 69.015 2.585 69.06 3.196 ;
      RECT 69.005 2.597 69.015 3.233 ;
      RECT 68.985 2.611 69.005 3.253 ;
      RECT 68.975 2.629 68.985 3.269 ;
      RECT 68.96 2.655 68.975 3.279 ;
      RECT 68.945 2.696 68.96 3.293 ;
      RECT 68.935 2.731 68.945 3.303 ;
      RECT 68.93 2.747 68.935 3.308 ;
      RECT 68.92 2.762 68.93 3.313 ;
      RECT 68.9 2.805 68.92 3.323 ;
      RECT 68.88 2.842 68.9 3.336 ;
      RECT 68.845 2.865 68.88 3.354 ;
      RECT 68.835 2.879 68.845 3.37 ;
      RECT 68.815 2.889 68.835 3.38 ;
      RECT 68.81 2.898 68.815 3.388 ;
      RECT 68.8 2.905 68.81 3.395 ;
      RECT 68.79 2.912 68.8 3.403 ;
      RECT 68.775 2.922 68.79 3.411 ;
      RECT 68.765 2.936 68.775 3.421 ;
      RECT 68.755 2.948 68.765 3.433 ;
      RECT 68.74 2.97 68.755 3.446 ;
      RECT 68.73 2.992 68.74 3.457 ;
      RECT 68.72 3.012 68.73 3.466 ;
      RECT 68.715 3.027 68.72 3.473 ;
      RECT 68.685 3.06 68.715 3.487 ;
      RECT 68.675 3.095 68.685 3.502 ;
      RECT 68.67 3.102 68.675 3.508 ;
      RECT 68.65 3.117 68.67 3.515 ;
      RECT 68.645 3.132 68.65 3.523 ;
      RECT 68.64 3.141 68.645 3.528 ;
      RECT 68.625 3.147 68.64 3.535 ;
      RECT 68.62 3.153 68.625 3.543 ;
      RECT 68.615 3.157 68.62 3.55 ;
      RECT 68.61 3.161 68.615 3.56 ;
      RECT 68.6 3.166 68.61 3.57 ;
      RECT 68.58 3.177 68.6 3.598 ;
      RECT 68.565 3.189 68.58 3.625 ;
      RECT 68.545 3.202 68.565 3.65 ;
      RECT 68.525 3.217 68.545 3.674 ;
      RECT 68.51 3.232 68.525 3.689 ;
      RECT 68.505 3.243 68.51 3.698 ;
      RECT 68.44 3.288 68.505 3.708 ;
      RECT 68.405 3.347 68.44 3.721 ;
      RECT 68.4 3.37 68.405 3.727 ;
      RECT 68.395 3.377 68.4 3.729 ;
      RECT 68.38 3.387 68.395 3.732 ;
      RECT 68.35 3.412 68.38 3.736 ;
      RECT 68.345 3.43 68.35 3.74 ;
      RECT 68.34 3.437 68.345 3.741 ;
      RECT 68.32 3.445 68.34 3.745 ;
      RECT 68.31 3.452 68.32 3.749 ;
      RECT 68.266 3.463 68.31 3.756 ;
      RECT 68.18 3.491 68.266 3.772 ;
      RECT 68.12 3.515 68.18 3.79 ;
      RECT 68.075 3.525 68.12 3.804 ;
      RECT 68.016 3.533 68.075 3.818 ;
      RECT 67.93 3.54 68.016 3.837 ;
      RECT 67.905 3.545 67.93 3.852 ;
      RECT 67.825 3.548 67.905 3.855 ;
      RECT 67.745 3.552 67.825 3.842 ;
      RECT 67.736 3.555 67.745 3.827 ;
      RECT 67.65 3.555 67.736 3.812 ;
      RECT 67.59 3.557 67.65 3.789 ;
      RECT 67.586 3.56 67.59 3.779 ;
      RECT 67.5 3.56 67.586 3.764 ;
      RECT 67.425 3.56 67.5 3.74 ;
      RECT 68.74 2.569 68.75 2.745 ;
      RECT 68.695 2.536 68.74 2.745 ;
      RECT 68.65 2.487 68.695 2.745 ;
      RECT 68.62 2.457 68.65 2.746 ;
      RECT 68.615 2.44 68.62 2.747 ;
      RECT 68.59 2.42 68.615 2.748 ;
      RECT 68.575 2.395 68.59 2.749 ;
      RECT 68.57 2.382 68.575 2.75 ;
      RECT 68.565 2.376 68.57 2.748 ;
      RECT 68.56 2.368 68.565 2.742 ;
      RECT 68.535 2.36 68.56 2.722 ;
      RECT 68.515 2.349 68.535 2.693 ;
      RECT 68.485 2.334 68.515 2.664 ;
      RECT 68.465 2.32 68.485 2.636 ;
      RECT 68.455 2.314 68.465 2.615 ;
      RECT 68.45 2.311 68.455 2.598 ;
      RECT 68.445 2.308 68.45 2.583 ;
      RECT 68.43 2.303 68.445 2.548 ;
      RECT 68.425 2.299 68.43 2.515 ;
      RECT 68.405 2.294 68.425 2.491 ;
      RECT 68.375 2.286 68.405 2.456 ;
      RECT 68.36 2.28 68.375 2.433 ;
      RECT 68.32 2.273 68.36 2.418 ;
      RECT 68.295 2.265 68.32 2.398 ;
      RECT 68.275 2.26 68.295 2.388 ;
      RECT 68.24 2.254 68.275 2.383 ;
      RECT 68.195 2.245 68.24 2.382 ;
      RECT 68.165 2.241 68.195 2.384 ;
      RECT 68.08 2.249 68.165 2.388 ;
      RECT 68.01 2.26 68.08 2.41 ;
      RECT 67.997 2.266 68.01 2.433 ;
      RECT 67.911 2.273 67.997 2.455 ;
      RECT 67.825 2.285 67.911 2.492 ;
      RECT 67.825 2.662 67.835 2.9 ;
      RECT 67.82 2.291 67.825 2.515 ;
      RECT 67.815 2.547 67.825 2.9 ;
      RECT 67.815 2.292 67.82 2.52 ;
      RECT 67.81 2.293 67.815 2.9 ;
      RECT 67.786 2.295 67.81 2.901 ;
      RECT 67.7 2.303 67.786 2.903 ;
      RECT 67.68 2.317 67.7 2.906 ;
      RECT 67.675 2.345 67.68 2.907 ;
      RECT 67.67 2.357 67.675 2.908 ;
      RECT 67.665 2.372 67.67 2.909 ;
      RECT 67.655 2.402 67.665 2.91 ;
      RECT 67.65 2.44 67.655 2.908 ;
      RECT 67.645 2.46 67.65 2.903 ;
      RECT 67.63 2.495 67.645 2.888 ;
      RECT 67.62 2.547 67.63 2.868 ;
      RECT 67.615 2.577 67.62 2.856 ;
      RECT 67.6 2.59 67.615 2.839 ;
      RECT 67.575 2.594 67.6 2.806 ;
      RECT 67.56 2.592 67.575 2.783 ;
      RECT 67.545 2.591 67.56 2.78 ;
      RECT 67.485 2.589 67.545 2.778 ;
      RECT 67.475 2.587 67.485 2.773 ;
      RECT 67.435 2.586 67.475 2.77 ;
      RECT 67.365 2.583 67.435 2.768 ;
      RECT 67.31 2.581 67.365 2.763 ;
      RECT 67.24 2.575 67.31 2.758 ;
      RECT 67.231 2.575 67.24 2.755 ;
      RECT 67.145 2.575 67.231 2.75 ;
      RECT 67.14 2.575 67.145 2.745 ;
      RECT 68.445 1.81 68.62 2.16 ;
      RECT 68.445 1.825 68.63 2.158 ;
      RECT 68.42 1.775 68.565 2.155 ;
      RECT 68.4 1.776 68.565 2.148 ;
      RECT 68.39 1.777 68.575 2.143 ;
      RECT 68.36 1.778 68.575 2.13 ;
      RECT 68.31 1.779 68.575 2.106 ;
      RECT 68.305 1.781 68.575 2.091 ;
      RECT 68.305 1.847 68.635 2.085 ;
      RECT 68.285 1.788 68.59 2.065 ;
      RECT 68.275 1.797 68.6 1.92 ;
      RECT 68.285 1.792 68.6 2.065 ;
      RECT 68.305 1.782 68.59 2.091 ;
      RECT 67.89 3.107 68.06 3.395 ;
      RECT 67.885 3.125 68.07 3.39 ;
      RECT 67.85 3.133 68.135 3.31 ;
      RECT 67.85 3.133 68.221 3.3 ;
      RECT 67.85 3.133 68.275 3.246 ;
      RECT 68.135 3.03 68.305 3.214 ;
      RECT 67.85 3.185 68.31 3.202 ;
      RECT 67.835 3.155 68.305 3.198 ;
      RECT 68.095 3.037 68.135 3.349 ;
      RECT 67.975 3.074 68.305 3.214 ;
      RECT 68.07 3.049 68.095 3.375 ;
      RECT 68.06 3.056 68.305 3.214 ;
      RECT 68.191 2.52 68.26 2.779 ;
      RECT 68.191 2.575 68.265 2.778 ;
      RECT 68.105 2.575 68.265 2.777 ;
      RECT 68.1 2.575 68.27 2.77 ;
      RECT 68.09 2.52 68.26 2.765 ;
      RECT 67.47 1.819 67.645 2.12 ;
      RECT 67.455 1.807 67.47 2.105 ;
      RECT 67.425 1.806 67.455 2.058 ;
      RECT 67.425 1.824 67.65 2.053 ;
      RECT 67.41 1.808 67.47 2.018 ;
      RECT 67.405 1.83 67.66 1.918 ;
      RECT 67.405 1.813 67.556 1.918 ;
      RECT 67.405 1.815 67.56 1.918 ;
      RECT 67.41 1.811 67.556 2.018 ;
      RECT 67.515 3.047 67.52 3.395 ;
      RECT 67.505 3.037 67.515 3.401 ;
      RECT 67.47 3.027 67.505 3.403 ;
      RECT 67.432 3.022 67.47 3.407 ;
      RECT 67.346 3.015 67.432 3.414 ;
      RECT 67.26 3.005 67.346 3.424 ;
      RECT 67.215 3 67.26 3.432 ;
      RECT 67.211 3 67.215 3.436 ;
      RECT 67.125 3 67.211 3.443 ;
      RECT 67.11 3 67.125 3.443 ;
      RECT 67.1 2.998 67.11 3.415 ;
      RECT 67.09 2.994 67.1 3.358 ;
      RECT 67.07 2.988 67.09 3.29 ;
      RECT 67.065 2.984 67.07 3.238 ;
      RECT 67.055 2.983 67.065 3.205 ;
      RECT 67.005 2.981 67.055 3.19 ;
      RECT 66.98 2.979 67.005 3.185 ;
      RECT 66.937 2.977 66.98 3.181 ;
      RECT 66.851 2.973 66.937 3.169 ;
      RECT 66.765 2.968 66.851 3.153 ;
      RECT 66.735 2.965 66.765 3.14 ;
      RECT 66.71 2.964 66.735 3.128 ;
      RECT 66.705 2.964 66.71 3.118 ;
      RECT 66.665 2.963 66.705 3.11 ;
      RECT 66.65 2.962 66.665 3.103 ;
      RECT 66.6 2.961 66.65 3.095 ;
      RECT 66.598 2.96 66.6 3.09 ;
      RECT 66.512 2.958 66.598 3.09 ;
      RECT 66.426 2.953 66.512 3.09 ;
      RECT 66.34 2.949 66.426 3.09 ;
      RECT 66.291 2.945 66.34 3.088 ;
      RECT 66.205 2.942 66.291 3.083 ;
      RECT 66.182 2.939 66.205 3.079 ;
      RECT 66.096 2.936 66.182 3.074 ;
      RECT 66.01 2.932 66.096 3.065 ;
      RECT 65.985 2.925 66.01 3.06 ;
      RECT 65.925 2.89 65.985 3.057 ;
      RECT 65.905 2.815 65.925 3.054 ;
      RECT 65.9 2.757 65.905 3.053 ;
      RECT 65.875 2.697 65.9 3.052 ;
      RECT 65.8 2.575 65.875 3.048 ;
      RECT 65.79 2.575 65.8 3.04 ;
      RECT 65.775 2.575 65.79 3.03 ;
      RECT 65.76 2.575 65.775 3 ;
      RECT 65.745 2.575 65.76 2.945 ;
      RECT 65.73 2.575 65.745 2.883 ;
      RECT 65.705 2.575 65.73 2.808 ;
      RECT 65.7 2.575 65.705 2.758 ;
      RECT 67.045 2.12 67.065 2.429 ;
      RECT 67.031 2.122 67.08 2.426 ;
      RECT 67.031 2.127 67.1 2.417 ;
      RECT 66.945 2.125 67.08 2.411 ;
      RECT 66.945 2.133 67.135 2.394 ;
      RECT 66.91 2.135 67.135 2.393 ;
      RECT 66.88 2.143 67.135 2.384 ;
      RECT 66.87 2.148 67.155 2.37 ;
      RECT 66.91 2.138 67.155 2.37 ;
      RECT 66.91 2.141 67.165 2.358 ;
      RECT 66.88 2.143 67.175 2.345 ;
      RECT 66.88 2.147 67.185 2.288 ;
      RECT 66.87 2.152 67.19 2.203 ;
      RECT 67.031 2.12 67.065 2.426 ;
      RECT 66.91 7.855 67.08 8.305 ;
      RECT 66.965 6.075 67.135 8.025 ;
      RECT 66.91 5.015 67.08 6.245 ;
      RECT 66.47 2.223 66.475 2.435 ;
      RECT 66.345 2.22 66.36 2.435 ;
      RECT 65.81 2.25 65.88 2.435 ;
      RECT 65.695 2.25 65.73 2.43 ;
      RECT 66.816 2.552 66.835 2.746 ;
      RECT 66.73 2.507 66.816 2.747 ;
      RECT 66.72 2.46 66.73 2.749 ;
      RECT 66.715 2.44 66.72 2.75 ;
      RECT 66.695 2.405 66.715 2.751 ;
      RECT 66.68 2.355 66.695 2.752 ;
      RECT 66.66 2.292 66.68 2.753 ;
      RECT 66.65 2.255 66.66 2.754 ;
      RECT 66.635 2.244 66.65 2.755 ;
      RECT 66.63 2.236 66.635 2.753 ;
      RECT 66.62 2.235 66.63 2.745 ;
      RECT 66.59 2.232 66.62 2.724 ;
      RECT 66.515 2.227 66.59 2.669 ;
      RECT 66.5 2.223 66.515 2.615 ;
      RECT 66.49 2.223 66.5 2.51 ;
      RECT 66.475 2.223 66.49 2.443 ;
      RECT 66.46 2.223 66.47 2.433 ;
      RECT 66.405 2.222 66.46 2.43 ;
      RECT 66.36 2.22 66.405 2.433 ;
      RECT 66.332 2.22 66.345 2.436 ;
      RECT 66.246 2.224 66.332 2.438 ;
      RECT 66.16 2.23 66.246 2.443 ;
      RECT 66.14 2.234 66.16 2.445 ;
      RECT 66.138 2.235 66.14 2.444 ;
      RECT 66.052 2.237 66.138 2.443 ;
      RECT 65.966 2.242 66.052 2.44 ;
      RECT 65.88 2.247 65.966 2.437 ;
      RECT 65.73 2.25 65.81 2.433 ;
      RECT 66.39 5.015 66.56 8.305 ;
      RECT 66.39 7.315 66.795 7.645 ;
      RECT 66.39 6.475 66.795 6.805 ;
      RECT 66.506 3.225 66.555 3.559 ;
      RECT 66.506 3.225 66.56 3.558 ;
      RECT 66.42 3.225 66.56 3.557 ;
      RECT 66.195 3.333 66.565 3.555 ;
      RECT 66.42 3.225 66.59 3.548 ;
      RECT 66.39 3.237 66.595 3.539 ;
      RECT 66.375 3.255 66.6 3.536 ;
      RECT 66.19 3.339 66.6 3.463 ;
      RECT 66.185 3.346 66.6 3.423 ;
      RECT 66.2 3.312 66.6 3.536 ;
      RECT 66.361 3.258 66.565 3.555 ;
      RECT 66.275 3.278 66.6 3.536 ;
      RECT 66.375 3.252 66.595 3.539 ;
      RECT 66.145 2.576 66.335 2.77 ;
      RECT 66.14 2.578 66.335 2.769 ;
      RECT 66.135 2.582 66.35 2.766 ;
      RECT 66.15 2.575 66.35 2.766 ;
      RECT 66.135 2.685 66.355 2.761 ;
      RECT 65.43 3.185 65.521 3.483 ;
      RECT 65.425 3.187 65.6 3.478 ;
      RECT 65.43 3.185 65.6 3.478 ;
      RECT 65.425 3.191 65.62 3.476 ;
      RECT 65.425 3.246 65.66 3.475 ;
      RECT 65.425 3.281 65.675 3.469 ;
      RECT 65.425 3.315 65.685 3.459 ;
      RECT 65.415 3.195 65.62 3.31 ;
      RECT 65.415 3.215 65.635 3.31 ;
      RECT 65.415 3.198 65.625 3.31 ;
      RECT 65.64 1.966 65.645 2.028 ;
      RECT 65.635 1.888 65.64 2.051 ;
      RECT 65.63 1.845 65.635 2.062 ;
      RECT 65.625 1.835 65.63 2.074 ;
      RECT 65.62 1.835 65.625 2.083 ;
      RECT 65.595 1.835 65.62 2.115 ;
      RECT 65.59 1.835 65.595 2.148 ;
      RECT 65.575 1.835 65.59 2.173 ;
      RECT 65.565 1.835 65.575 2.2 ;
      RECT 65.56 1.835 65.565 2.213 ;
      RECT 65.555 1.835 65.56 2.228 ;
      RECT 65.545 1.835 65.555 2.243 ;
      RECT 65.54 1.835 65.545 2.263 ;
      RECT 65.515 1.835 65.54 2.298 ;
      RECT 65.47 1.835 65.515 2.343 ;
      RECT 65.46 1.835 65.47 2.356 ;
      RECT 65.375 1.92 65.46 2.363 ;
      RECT 65.34 2.042 65.375 2.372 ;
      RECT 65.335 2.082 65.34 2.376 ;
      RECT 65.315 2.105 65.335 2.378 ;
      RECT 65.31 2.135 65.315 2.381 ;
      RECT 65.3 2.147 65.31 2.382 ;
      RECT 65.255 2.17 65.3 2.387 ;
      RECT 65.215 2.2 65.255 2.395 ;
      RECT 65.18 2.212 65.215 2.401 ;
      RECT 65.175 2.217 65.18 2.405 ;
      RECT 65.105 2.227 65.175 2.412 ;
      RECT 65.065 2.237 65.105 2.422 ;
      RECT 65.045 2.242 65.065 2.428 ;
      RECT 65.035 2.246 65.045 2.433 ;
      RECT 65.03 2.249 65.035 2.436 ;
      RECT 65.02 2.25 65.03 2.437 ;
      RECT 64.995 2.252 65.02 2.441 ;
      RECT 64.985 2.257 64.995 2.444 ;
      RECT 64.94 2.265 64.985 2.445 ;
      RECT 64.815 2.27 64.94 2.445 ;
      RECT 65.37 2.567 65.39 2.749 ;
      RECT 65.321 2.552 65.37 2.748 ;
      RECT 65.235 2.567 65.39 2.746 ;
      RECT 65.22 2.567 65.39 2.745 ;
      RECT 65.185 2.545 65.355 2.73 ;
      RECT 65.255 3.565 65.27 3.774 ;
      RECT 65.255 3.573 65.275 3.773 ;
      RECT 65.2 3.573 65.275 3.772 ;
      RECT 65.18 3.577 65.28 3.77 ;
      RECT 65.16 3.527 65.2 3.769 ;
      RECT 65.105 3.585 65.285 3.767 ;
      RECT 65.07 3.542 65.2 3.765 ;
      RECT 65.066 3.545 65.255 3.764 ;
      RECT 64.98 3.553 65.255 3.762 ;
      RECT 64.98 3.597 65.29 3.755 ;
      RECT 64.97 3.69 65.29 3.753 ;
      RECT 64.98 3.609 65.295 3.738 ;
      RECT 64.98 3.63 65.31 3.708 ;
      RECT 64.98 3.657 65.315 3.678 ;
      RECT 65.105 3.535 65.2 3.767 ;
      RECT 64.735 2.58 64.74 3.118 ;
      RECT 64.54 2.91 64.545 3.105 ;
      RECT 62.84 2.575 62.855 2.955 ;
      RECT 64.905 2.575 64.91 2.745 ;
      RECT 64.9 2.575 64.905 2.755 ;
      RECT 64.895 2.575 64.9 2.768 ;
      RECT 64.87 2.575 64.895 2.81 ;
      RECT 64.845 2.575 64.87 2.883 ;
      RECT 64.83 2.575 64.845 2.935 ;
      RECT 64.825 2.575 64.83 2.965 ;
      RECT 64.8 2.575 64.825 3.005 ;
      RECT 64.785 2.575 64.8 3.06 ;
      RECT 64.78 2.575 64.785 3.093 ;
      RECT 64.755 2.575 64.78 3.113 ;
      RECT 64.74 2.575 64.755 3.119 ;
      RECT 64.67 2.61 64.735 3.115 ;
      RECT 64.62 2.665 64.67 3.11 ;
      RECT 64.61 2.697 64.62 3.108 ;
      RECT 64.605 2.722 64.61 3.108 ;
      RECT 64.585 2.795 64.605 3.108 ;
      RECT 64.575 2.875 64.585 3.107 ;
      RECT 64.56 2.905 64.575 3.107 ;
      RECT 64.545 2.91 64.56 3.106 ;
      RECT 64.485 2.912 64.54 3.103 ;
      RECT 64.455 2.917 64.485 3.099 ;
      RECT 64.453 2.92 64.455 3.098 ;
      RECT 64.367 2.922 64.453 3.095 ;
      RECT 64.281 2.928 64.367 3.089 ;
      RECT 64.195 2.933 64.281 3.083 ;
      RECT 64.122 2.938 64.195 3.084 ;
      RECT 64.036 2.944 64.122 3.092 ;
      RECT 63.95 2.95 64.036 3.101 ;
      RECT 63.93 2.954 63.95 3.106 ;
      RECT 63.883 2.956 63.93 3.109 ;
      RECT 63.797 2.961 63.883 3.115 ;
      RECT 63.711 2.966 63.797 3.124 ;
      RECT 63.625 2.972 63.711 3.132 ;
      RECT 63.54 2.97 63.625 3.141 ;
      RECT 63.536 2.965 63.54 3.145 ;
      RECT 63.45 2.96 63.536 3.137 ;
      RECT 63.386 2.951 63.45 3.125 ;
      RECT 63.3 2.942 63.386 3.112 ;
      RECT 63.276 2.935 63.3 3.103 ;
      RECT 63.19 2.929 63.276 3.09 ;
      RECT 63.15 2.922 63.19 3.076 ;
      RECT 63.145 2.912 63.15 3.072 ;
      RECT 63.135 2.9 63.145 3.071 ;
      RECT 63.115 2.87 63.135 3.068 ;
      RECT 63.06 2.79 63.115 3.062 ;
      RECT 63.04 2.709 63.06 3.057 ;
      RECT 63.02 2.667 63.04 3.053 ;
      RECT 62.995 2.62 63.02 3.047 ;
      RECT 62.99 2.595 62.995 3.044 ;
      RECT 62.955 2.575 62.99 3.039 ;
      RECT 62.946 2.575 62.955 3.032 ;
      RECT 62.86 2.575 62.946 3.002 ;
      RECT 62.855 2.575 62.86 2.965 ;
      RECT 62.82 2.575 62.84 2.887 ;
      RECT 62.815 2.617 62.82 2.852 ;
      RECT 62.81 2.692 62.815 2.808 ;
      RECT 64.26 2.497 64.435 2.745 ;
      RECT 64.26 2.497 64.44 2.743 ;
      RECT 64.255 2.529 64.44 2.703 ;
      RECT 64.285 2.47 64.455 2.69 ;
      RECT 64.25 2.547 64.455 2.623 ;
      RECT 63.56 2.01 63.73 2.185 ;
      RECT 63.56 2.01 63.902 2.177 ;
      RECT 63.56 2.01 63.985 2.171 ;
      RECT 63.56 2.01 64.02 2.167 ;
      RECT 63.56 2.01 64.04 2.166 ;
      RECT 63.56 2.01 64.126 2.162 ;
      RECT 64.02 1.835 64.19 2.157 ;
      RECT 63.595 1.942 64.22 2.155 ;
      RECT 63.585 1.997 64.225 2.153 ;
      RECT 63.56 2.033 64.235 2.148 ;
      RECT 63.56 2.06 64.24 2.078 ;
      RECT 63.625 1.885 64.2 2.155 ;
      RECT 63.816 1.87 64.2 2.155 ;
      RECT 63.65 1.873 64.2 2.155 ;
      RECT 63.73 1.871 63.816 2.182 ;
      RECT 63.816 1.868 64.195 2.155 ;
      RECT 64 1.845 64.195 2.155 ;
      RECT 63.902 1.866 64.195 2.155 ;
      RECT 63.985 1.86 64 2.168 ;
      RECT 64.135 3.225 64.14 3.425 ;
      RECT 63.6 3.29 63.645 3.425 ;
      RECT 64.17 3.225 64.19 3.398 ;
      RECT 64.14 3.225 64.17 3.413 ;
      RECT 64.075 3.225 64.135 3.45 ;
      RECT 64.06 3.225 64.075 3.48 ;
      RECT 64.045 3.225 64.06 3.493 ;
      RECT 64.025 3.225 64.045 3.508 ;
      RECT 64.02 3.225 64.025 3.517 ;
      RECT 64.01 3.229 64.02 3.522 ;
      RECT 63.995 3.239 64.01 3.533 ;
      RECT 63.97 3.255 63.995 3.543 ;
      RECT 63.96 3.269 63.97 3.545 ;
      RECT 63.94 3.281 63.96 3.542 ;
      RECT 63.91 3.302 63.94 3.536 ;
      RECT 63.9 3.314 63.91 3.531 ;
      RECT 63.89 3.312 63.9 3.528 ;
      RECT 63.875 3.311 63.89 3.523 ;
      RECT 63.87 3.31 63.875 3.518 ;
      RECT 63.835 3.308 63.87 3.508 ;
      RECT 63.815 3.305 63.835 3.49 ;
      RECT 63.805 3.303 63.815 3.485 ;
      RECT 63.795 3.302 63.805 3.48 ;
      RECT 63.76 3.3 63.795 3.468 ;
      RECT 63.705 3.296 63.76 3.448 ;
      RECT 63.695 3.294 63.705 3.433 ;
      RECT 63.69 3.294 63.695 3.428 ;
      RECT 63.645 3.292 63.69 3.425 ;
      RECT 63.55 3.29 63.6 3.429 ;
      RECT 63.54 3.291 63.55 3.434 ;
      RECT 63.48 3.298 63.54 3.448 ;
      RECT 63.455 3.306 63.48 3.468 ;
      RECT 63.445 3.31 63.455 3.48 ;
      RECT 63.44 3.311 63.445 3.485 ;
      RECT 63.425 3.313 63.44 3.488 ;
      RECT 63.41 3.315 63.425 3.493 ;
      RECT 63.405 3.315 63.41 3.496 ;
      RECT 63.36 3.32 63.405 3.507 ;
      RECT 63.355 3.324 63.36 3.519 ;
      RECT 63.33 3.32 63.355 3.523 ;
      RECT 63.32 3.316 63.33 3.527 ;
      RECT 63.31 3.315 63.32 3.531 ;
      RECT 63.295 3.305 63.31 3.537 ;
      RECT 63.29 3.293 63.295 3.541 ;
      RECT 63.285 3.29 63.29 3.542 ;
      RECT 63.28 3.287 63.285 3.544 ;
      RECT 63.265 3.275 63.28 3.543 ;
      RECT 63.25 3.257 63.265 3.54 ;
      RECT 63.23 3.236 63.25 3.533 ;
      RECT 63.165 3.225 63.23 3.505 ;
      RECT 63.161 3.225 63.165 3.484 ;
      RECT 63.075 3.225 63.161 3.454 ;
      RECT 63.06 3.225 63.075 3.41 ;
      RECT 63.635 2.325 63.64 2.56 ;
      RECT 62.765 2.241 62.77 2.445 ;
      RECT 63.345 2.27 63.35 2.425 ;
      RECT 63.265 2.25 63.27 2.425 ;
      RECT 63.935 2.392 63.95 2.745 ;
      RECT 63.861 2.377 63.935 2.745 ;
      RECT 63.775 2.36 63.861 2.745 ;
      RECT 63.765 2.35 63.775 2.743 ;
      RECT 63.76 2.348 63.765 2.738 ;
      RECT 63.745 2.346 63.76 2.724 ;
      RECT 63.675 2.338 63.745 2.664 ;
      RECT 63.655 2.329 63.675 2.598 ;
      RECT 63.65 2.326 63.655 2.578 ;
      RECT 63.64 2.325 63.65 2.568 ;
      RECT 63.63 2.325 63.635 2.552 ;
      RECT 63.62 2.324 63.63 2.542 ;
      RECT 63.61 2.322 63.62 2.53 ;
      RECT 63.595 2.319 63.61 2.51 ;
      RECT 63.585 2.317 63.595 2.495 ;
      RECT 63.565 2.314 63.585 2.483 ;
      RECT 63.56 2.312 63.565 2.473 ;
      RECT 63.535 2.31 63.56 2.46 ;
      RECT 63.505 2.305 63.535 2.445 ;
      RECT 63.425 2.296 63.505 2.436 ;
      RECT 63.38 2.285 63.425 2.429 ;
      RECT 63.36 2.276 63.38 2.426 ;
      RECT 63.35 2.271 63.36 2.425 ;
      RECT 63.305 2.265 63.345 2.425 ;
      RECT 63.29 2.257 63.305 2.425 ;
      RECT 63.27 2.252 63.29 2.425 ;
      RECT 63.25 2.249 63.265 2.425 ;
      RECT 63.167 2.248 63.25 2.424 ;
      RECT 63.081 2.247 63.167 2.42 ;
      RECT 62.995 2.245 63.081 2.417 ;
      RECT 62.942 2.244 62.995 2.419 ;
      RECT 62.856 2.243 62.942 2.428 ;
      RECT 62.77 2.242 62.856 2.44 ;
      RECT 62.75 2.241 62.765 2.448 ;
      RECT 62.67 2.24 62.75 2.46 ;
      RECT 62.645 2.24 62.67 2.473 ;
      RECT 62.62 2.24 62.645 2.488 ;
      RECT 62.615 2.24 62.62 2.51 ;
      RECT 62.61 2.24 62.615 2.528 ;
      RECT 62.605 2.24 62.61 2.545 ;
      RECT 62.6 2.24 62.605 2.558 ;
      RECT 62.595 2.24 62.6 2.568 ;
      RECT 62.555 2.24 62.595 2.653 ;
      RECT 62.54 2.24 62.555 2.738 ;
      RECT 62.53 2.241 62.54 2.75 ;
      RECT 62.495 2.246 62.53 2.755 ;
      RECT 62.455 2.255 62.495 2.755 ;
      RECT 62.44 2.265 62.455 2.755 ;
      RECT 62.435 2.275 62.44 2.755 ;
      RECT 62.415 2.302 62.435 2.755 ;
      RECT 62.365 2.385 62.415 2.755 ;
      RECT 62.36 2.447 62.365 2.755 ;
      RECT 62.35 2.46 62.36 2.755 ;
      RECT 62.34 2.482 62.35 2.755 ;
      RECT 62.33 2.507 62.34 2.75 ;
      RECT 62.325 2.545 62.33 2.743 ;
      RECT 62.315 2.655 62.325 2.738 ;
      RECT 63.71 3.576 63.725 3.835 ;
      RECT 63.71 3.591 63.73 3.834 ;
      RECT 63.626 3.591 63.73 3.832 ;
      RECT 63.626 3.605 63.735 3.831 ;
      RECT 63.54 3.647 63.74 3.828 ;
      RECT 63.535 3.59 63.725 3.823 ;
      RECT 63.535 3.661 63.745 3.82 ;
      RECT 63.53 3.692 63.745 3.818 ;
      RECT 63.535 3.689 63.76 3.808 ;
      RECT 63.53 3.735 63.775 3.793 ;
      RECT 63.53 3.763 63.78 3.778 ;
      RECT 63.54 3.565 63.71 3.828 ;
      RECT 63.3 2.575 63.47 2.745 ;
      RECT 63.265 2.575 63.47 2.74 ;
      RECT 63.255 2.575 63.47 2.733 ;
      RECT 63.25 2.56 63.42 2.73 ;
      RECT 62.08 3.097 62.345 3.54 ;
      RECT 62.075 3.068 62.29 3.538 ;
      RECT 62.07 3.222 62.35 3.533 ;
      RECT 62.075 3.117 62.35 3.533 ;
      RECT 62.075 3.128 62.36 3.52 ;
      RECT 62.075 3.075 62.32 3.538 ;
      RECT 62.08 3.062 62.29 3.54 ;
      RECT 62.08 3.06 62.24 3.54 ;
      RECT 62.181 3.052 62.24 3.54 ;
      RECT 62.095 3.053 62.24 3.54 ;
      RECT 62.181 3.051 62.23 3.54 ;
      RECT 61.985 1.866 62.16 2.165 ;
      RECT 62.035 1.828 62.16 2.165 ;
      RECT 62.02 1.83 62.246 2.157 ;
      RECT 62.02 1.833 62.285 2.144 ;
      RECT 62.02 1.834 62.295 2.13 ;
      RECT 61.975 1.885 62.295 2.12 ;
      RECT 62.02 1.835 62.3 2.115 ;
      RECT 61.975 2.045 62.305 2.105 ;
      RECT 61.96 1.905 62.3 2.045 ;
      RECT 61.955 1.921 62.3 1.985 ;
      RECT 62 1.845 62.3 2.115 ;
      RECT 62.035 1.826 62.121 2.165 ;
      RECT 60.13 1.74 60.3 2.935 ;
      RECT 60.13 1.74 60.595 1.91 ;
      RECT 60.13 6.97 60.595 7.14 ;
      RECT 60.13 5.945 60.3 7.14 ;
      RECT 59.14 1.74 59.31 2.935 ;
      RECT 59.14 1.74 59.605 1.91 ;
      RECT 59.14 6.97 59.605 7.14 ;
      RECT 59.14 5.945 59.31 7.14 ;
      RECT 57.285 2.635 57.455 3.865 ;
      RECT 57.34 0.855 57.51 2.805 ;
      RECT 57.285 0.575 57.455 1.025 ;
      RECT 57.285 7.855 57.455 8.305 ;
      RECT 57.34 6.075 57.51 8.025 ;
      RECT 57.285 5.015 57.455 6.245 ;
      RECT 56.765 0.575 56.935 3.865 ;
      RECT 56.765 2.075 57.17 2.405 ;
      RECT 56.765 1.235 57.17 1.565 ;
      RECT 56.765 5.015 56.935 8.305 ;
      RECT 56.765 7.315 57.17 7.645 ;
      RECT 56.765 6.475 57.17 6.805 ;
      RECT 54.69 3.126 54.695 3.298 ;
      RECT 54.685 3.119 54.69 3.388 ;
      RECT 54.68 3.113 54.685 3.407 ;
      RECT 54.66 3.107 54.68 3.417 ;
      RECT 54.645 3.102 54.66 3.425 ;
      RECT 54.608 3.096 54.645 3.423 ;
      RECT 54.522 3.082 54.608 3.419 ;
      RECT 54.436 3.064 54.522 3.414 ;
      RECT 54.35 3.045 54.436 3.408 ;
      RECT 54.32 3.033 54.35 3.404 ;
      RECT 54.3 3.027 54.32 3.403 ;
      RECT 54.235 3.025 54.3 3.401 ;
      RECT 54.22 3.025 54.235 3.393 ;
      RECT 54.205 3.025 54.22 3.38 ;
      RECT 54.2 3.025 54.205 3.37 ;
      RECT 54.185 3.025 54.2 3.348 ;
      RECT 54.17 3.025 54.185 3.315 ;
      RECT 54.165 3.025 54.17 3.293 ;
      RECT 54.155 3.025 54.165 3.275 ;
      RECT 54.14 3.025 54.155 3.253 ;
      RECT 54.12 3.025 54.14 3.215 ;
      RECT 54.47 2.31 54.505 2.749 ;
      RECT 54.47 2.31 54.51 2.748 ;
      RECT 54.415 2.37 54.51 2.747 ;
      RECT 54.28 2.542 54.51 2.746 ;
      RECT 54.39 2.42 54.51 2.746 ;
      RECT 54.28 2.542 54.535 2.736 ;
      RECT 54.335 2.487 54.615 2.653 ;
      RECT 54.51 2.281 54.515 2.744 ;
      RECT 54.365 2.457 54.655 2.53 ;
      RECT 54.38 2.44 54.51 2.746 ;
      RECT 54.515 2.28 54.685 2.468 ;
      RECT 54.505 2.283 54.685 2.468 ;
      RECT 54.01 2.16 54.18 2.47 ;
      RECT 54.01 2.16 54.185 2.443 ;
      RECT 54.01 2.16 54.19 2.42 ;
      RECT 54.01 2.16 54.2 2.37 ;
      RECT 54.005 2.265 54.2 2.34 ;
      RECT 54.04 1.835 54.21 2.313 ;
      RECT 54.04 1.835 54.225 2.234 ;
      RECT 54.03 2.045 54.225 2.234 ;
      RECT 54.04 1.845 54.235 2.149 ;
      RECT 53.97 2.587 53.975 2.79 ;
      RECT 53.96 2.575 53.97 2.9 ;
      RECT 53.935 2.575 53.96 2.94 ;
      RECT 53.855 2.575 53.935 3.025 ;
      RECT 53.845 2.575 53.855 3.095 ;
      RECT 53.82 2.575 53.845 3.118 ;
      RECT 53.8 2.575 53.82 3.153 ;
      RECT 53.755 2.585 53.8 3.196 ;
      RECT 53.745 2.597 53.755 3.233 ;
      RECT 53.725 2.611 53.745 3.253 ;
      RECT 53.715 2.629 53.725 3.269 ;
      RECT 53.7 2.655 53.715 3.279 ;
      RECT 53.685 2.696 53.7 3.293 ;
      RECT 53.675 2.731 53.685 3.303 ;
      RECT 53.67 2.747 53.675 3.308 ;
      RECT 53.66 2.762 53.67 3.313 ;
      RECT 53.64 2.805 53.66 3.323 ;
      RECT 53.62 2.842 53.64 3.336 ;
      RECT 53.585 2.865 53.62 3.354 ;
      RECT 53.575 2.879 53.585 3.37 ;
      RECT 53.555 2.889 53.575 3.38 ;
      RECT 53.55 2.898 53.555 3.388 ;
      RECT 53.54 2.905 53.55 3.395 ;
      RECT 53.53 2.912 53.54 3.403 ;
      RECT 53.515 2.922 53.53 3.411 ;
      RECT 53.505 2.936 53.515 3.421 ;
      RECT 53.495 2.948 53.505 3.433 ;
      RECT 53.48 2.97 53.495 3.446 ;
      RECT 53.47 2.992 53.48 3.457 ;
      RECT 53.46 3.012 53.47 3.466 ;
      RECT 53.455 3.027 53.46 3.473 ;
      RECT 53.425 3.06 53.455 3.487 ;
      RECT 53.415 3.095 53.425 3.502 ;
      RECT 53.41 3.102 53.415 3.508 ;
      RECT 53.39 3.117 53.41 3.515 ;
      RECT 53.385 3.132 53.39 3.523 ;
      RECT 53.38 3.141 53.385 3.528 ;
      RECT 53.365 3.147 53.38 3.535 ;
      RECT 53.36 3.153 53.365 3.543 ;
      RECT 53.355 3.157 53.36 3.55 ;
      RECT 53.35 3.161 53.355 3.56 ;
      RECT 53.34 3.166 53.35 3.57 ;
      RECT 53.32 3.177 53.34 3.598 ;
      RECT 53.305 3.189 53.32 3.625 ;
      RECT 53.285 3.202 53.305 3.65 ;
      RECT 53.265 3.217 53.285 3.674 ;
      RECT 53.25 3.232 53.265 3.689 ;
      RECT 53.245 3.243 53.25 3.698 ;
      RECT 53.18 3.288 53.245 3.708 ;
      RECT 53.145 3.347 53.18 3.721 ;
      RECT 53.14 3.37 53.145 3.727 ;
      RECT 53.135 3.377 53.14 3.729 ;
      RECT 53.12 3.387 53.135 3.732 ;
      RECT 53.09 3.412 53.12 3.736 ;
      RECT 53.085 3.43 53.09 3.74 ;
      RECT 53.08 3.437 53.085 3.741 ;
      RECT 53.06 3.445 53.08 3.745 ;
      RECT 53.05 3.452 53.06 3.749 ;
      RECT 53.006 3.463 53.05 3.756 ;
      RECT 52.92 3.491 53.006 3.772 ;
      RECT 52.86 3.515 52.92 3.79 ;
      RECT 52.815 3.525 52.86 3.804 ;
      RECT 52.756 3.533 52.815 3.818 ;
      RECT 52.67 3.54 52.756 3.837 ;
      RECT 52.645 3.545 52.67 3.852 ;
      RECT 52.565 3.548 52.645 3.855 ;
      RECT 52.485 3.552 52.565 3.842 ;
      RECT 52.476 3.555 52.485 3.827 ;
      RECT 52.39 3.555 52.476 3.812 ;
      RECT 52.33 3.557 52.39 3.789 ;
      RECT 52.326 3.56 52.33 3.779 ;
      RECT 52.24 3.56 52.326 3.764 ;
      RECT 52.165 3.56 52.24 3.74 ;
      RECT 53.48 2.569 53.49 2.745 ;
      RECT 53.435 2.536 53.48 2.745 ;
      RECT 53.39 2.487 53.435 2.745 ;
      RECT 53.36 2.457 53.39 2.746 ;
      RECT 53.355 2.44 53.36 2.747 ;
      RECT 53.33 2.42 53.355 2.748 ;
      RECT 53.315 2.395 53.33 2.749 ;
      RECT 53.31 2.382 53.315 2.75 ;
      RECT 53.305 2.376 53.31 2.748 ;
      RECT 53.3 2.368 53.305 2.742 ;
      RECT 53.275 2.36 53.3 2.722 ;
      RECT 53.255 2.349 53.275 2.693 ;
      RECT 53.225 2.334 53.255 2.664 ;
      RECT 53.205 2.32 53.225 2.636 ;
      RECT 53.195 2.314 53.205 2.615 ;
      RECT 53.19 2.311 53.195 2.598 ;
      RECT 53.185 2.308 53.19 2.583 ;
      RECT 53.17 2.303 53.185 2.548 ;
      RECT 53.165 2.299 53.17 2.515 ;
      RECT 53.145 2.294 53.165 2.491 ;
      RECT 53.115 2.286 53.145 2.456 ;
      RECT 53.1 2.28 53.115 2.433 ;
      RECT 53.06 2.273 53.1 2.418 ;
      RECT 53.035 2.265 53.06 2.398 ;
      RECT 53.015 2.26 53.035 2.388 ;
      RECT 52.98 2.254 53.015 2.383 ;
      RECT 52.935 2.245 52.98 2.382 ;
      RECT 52.905 2.241 52.935 2.384 ;
      RECT 52.82 2.249 52.905 2.388 ;
      RECT 52.75 2.26 52.82 2.41 ;
      RECT 52.737 2.266 52.75 2.433 ;
      RECT 52.651 2.273 52.737 2.455 ;
      RECT 52.565 2.285 52.651 2.492 ;
      RECT 52.565 2.662 52.575 2.9 ;
      RECT 52.56 2.291 52.565 2.515 ;
      RECT 52.555 2.547 52.565 2.9 ;
      RECT 52.555 2.292 52.56 2.52 ;
      RECT 52.55 2.293 52.555 2.9 ;
      RECT 52.526 2.295 52.55 2.901 ;
      RECT 52.44 2.303 52.526 2.903 ;
      RECT 52.42 2.317 52.44 2.906 ;
      RECT 52.415 2.345 52.42 2.907 ;
      RECT 52.41 2.357 52.415 2.908 ;
      RECT 52.405 2.372 52.41 2.909 ;
      RECT 52.395 2.402 52.405 2.91 ;
      RECT 52.39 2.44 52.395 2.908 ;
      RECT 52.385 2.46 52.39 2.903 ;
      RECT 52.37 2.495 52.385 2.888 ;
      RECT 52.36 2.547 52.37 2.868 ;
      RECT 52.355 2.577 52.36 2.856 ;
      RECT 52.34 2.59 52.355 2.839 ;
      RECT 52.315 2.594 52.34 2.806 ;
      RECT 52.3 2.592 52.315 2.783 ;
      RECT 52.285 2.591 52.3 2.78 ;
      RECT 52.225 2.589 52.285 2.778 ;
      RECT 52.215 2.587 52.225 2.773 ;
      RECT 52.175 2.586 52.215 2.77 ;
      RECT 52.105 2.583 52.175 2.768 ;
      RECT 52.05 2.581 52.105 2.763 ;
      RECT 51.98 2.575 52.05 2.758 ;
      RECT 51.971 2.575 51.98 2.755 ;
      RECT 51.885 2.575 51.971 2.75 ;
      RECT 51.88 2.575 51.885 2.745 ;
      RECT 53.185 1.81 53.36 2.16 ;
      RECT 53.185 1.825 53.37 2.158 ;
      RECT 53.16 1.775 53.305 2.155 ;
      RECT 53.14 1.776 53.305 2.148 ;
      RECT 53.13 1.777 53.315 2.143 ;
      RECT 53.1 1.778 53.315 2.13 ;
      RECT 53.05 1.779 53.315 2.106 ;
      RECT 53.045 1.781 53.315 2.091 ;
      RECT 53.045 1.847 53.375 2.085 ;
      RECT 53.025 1.788 53.33 2.065 ;
      RECT 53.015 1.797 53.34 1.92 ;
      RECT 53.025 1.792 53.34 2.065 ;
      RECT 53.045 1.782 53.33 2.091 ;
      RECT 52.63 3.107 52.8 3.395 ;
      RECT 52.625 3.125 52.81 3.39 ;
      RECT 52.59 3.133 52.875 3.31 ;
      RECT 52.59 3.133 52.961 3.3 ;
      RECT 52.59 3.133 53.015 3.246 ;
      RECT 52.875 3.03 53.045 3.214 ;
      RECT 52.59 3.185 53.05 3.202 ;
      RECT 52.575 3.155 53.045 3.198 ;
      RECT 52.835 3.037 52.875 3.349 ;
      RECT 52.715 3.074 53.045 3.214 ;
      RECT 52.81 3.049 52.835 3.375 ;
      RECT 52.8 3.056 53.045 3.214 ;
      RECT 52.931 2.52 53 2.779 ;
      RECT 52.931 2.575 53.005 2.778 ;
      RECT 52.845 2.575 53.005 2.777 ;
      RECT 52.84 2.575 53.01 2.77 ;
      RECT 52.83 2.52 53 2.765 ;
      RECT 52.21 1.819 52.385 2.12 ;
      RECT 52.195 1.807 52.21 2.105 ;
      RECT 52.165 1.806 52.195 2.058 ;
      RECT 52.165 1.824 52.39 2.053 ;
      RECT 52.15 1.808 52.21 2.018 ;
      RECT 52.145 1.83 52.4 1.918 ;
      RECT 52.145 1.813 52.296 1.918 ;
      RECT 52.145 1.815 52.3 1.918 ;
      RECT 52.15 1.811 52.296 2.018 ;
      RECT 52.255 3.047 52.26 3.395 ;
      RECT 52.245 3.037 52.255 3.401 ;
      RECT 52.21 3.027 52.245 3.403 ;
      RECT 52.172 3.022 52.21 3.407 ;
      RECT 52.086 3.015 52.172 3.414 ;
      RECT 52 3.005 52.086 3.424 ;
      RECT 51.955 3 52 3.432 ;
      RECT 51.951 3 51.955 3.436 ;
      RECT 51.865 3 51.951 3.443 ;
      RECT 51.85 3 51.865 3.443 ;
      RECT 51.84 2.998 51.85 3.415 ;
      RECT 51.83 2.994 51.84 3.358 ;
      RECT 51.81 2.988 51.83 3.29 ;
      RECT 51.805 2.984 51.81 3.238 ;
      RECT 51.795 2.983 51.805 3.205 ;
      RECT 51.745 2.981 51.795 3.19 ;
      RECT 51.72 2.979 51.745 3.185 ;
      RECT 51.677 2.977 51.72 3.181 ;
      RECT 51.591 2.973 51.677 3.169 ;
      RECT 51.505 2.968 51.591 3.153 ;
      RECT 51.475 2.965 51.505 3.14 ;
      RECT 51.45 2.964 51.475 3.128 ;
      RECT 51.445 2.964 51.45 3.118 ;
      RECT 51.405 2.963 51.445 3.11 ;
      RECT 51.39 2.962 51.405 3.103 ;
      RECT 51.34 2.961 51.39 3.095 ;
      RECT 51.338 2.96 51.34 3.09 ;
      RECT 51.252 2.958 51.338 3.09 ;
      RECT 51.166 2.953 51.252 3.09 ;
      RECT 51.08 2.949 51.166 3.09 ;
      RECT 51.031 2.945 51.08 3.088 ;
      RECT 50.945 2.942 51.031 3.083 ;
      RECT 50.922 2.939 50.945 3.079 ;
      RECT 50.836 2.936 50.922 3.074 ;
      RECT 50.75 2.932 50.836 3.065 ;
      RECT 50.725 2.925 50.75 3.06 ;
      RECT 50.665 2.89 50.725 3.057 ;
      RECT 50.645 2.815 50.665 3.054 ;
      RECT 50.64 2.757 50.645 3.053 ;
      RECT 50.615 2.697 50.64 3.052 ;
      RECT 50.54 2.575 50.615 3.048 ;
      RECT 50.53 2.575 50.54 3.04 ;
      RECT 50.515 2.575 50.53 3.03 ;
      RECT 50.5 2.575 50.515 3 ;
      RECT 50.485 2.575 50.5 2.945 ;
      RECT 50.47 2.575 50.485 2.883 ;
      RECT 50.445 2.575 50.47 2.808 ;
      RECT 50.44 2.575 50.445 2.758 ;
      RECT 51.785 2.12 51.805 2.429 ;
      RECT 51.771 2.122 51.82 2.426 ;
      RECT 51.771 2.127 51.84 2.417 ;
      RECT 51.685 2.125 51.82 2.411 ;
      RECT 51.685 2.133 51.875 2.394 ;
      RECT 51.65 2.135 51.875 2.393 ;
      RECT 51.62 2.143 51.875 2.384 ;
      RECT 51.61 2.148 51.895 2.37 ;
      RECT 51.65 2.138 51.895 2.37 ;
      RECT 51.65 2.141 51.905 2.358 ;
      RECT 51.62 2.143 51.915 2.345 ;
      RECT 51.62 2.147 51.925 2.288 ;
      RECT 51.61 2.152 51.93 2.203 ;
      RECT 51.771 2.12 51.805 2.426 ;
      RECT 51.65 7.855 51.82 8.305 ;
      RECT 51.705 6.075 51.875 8.025 ;
      RECT 51.65 5.015 51.82 6.245 ;
      RECT 51.21 2.223 51.215 2.435 ;
      RECT 51.085 2.22 51.1 2.435 ;
      RECT 50.55 2.25 50.62 2.435 ;
      RECT 50.435 2.25 50.47 2.43 ;
      RECT 51.556 2.552 51.575 2.746 ;
      RECT 51.47 2.507 51.556 2.747 ;
      RECT 51.46 2.46 51.47 2.749 ;
      RECT 51.455 2.44 51.46 2.75 ;
      RECT 51.435 2.405 51.455 2.751 ;
      RECT 51.42 2.355 51.435 2.752 ;
      RECT 51.4 2.292 51.42 2.753 ;
      RECT 51.39 2.255 51.4 2.754 ;
      RECT 51.375 2.244 51.39 2.755 ;
      RECT 51.37 2.236 51.375 2.753 ;
      RECT 51.36 2.235 51.37 2.745 ;
      RECT 51.33 2.232 51.36 2.724 ;
      RECT 51.255 2.227 51.33 2.669 ;
      RECT 51.24 2.223 51.255 2.615 ;
      RECT 51.23 2.223 51.24 2.51 ;
      RECT 51.215 2.223 51.23 2.443 ;
      RECT 51.2 2.223 51.21 2.433 ;
      RECT 51.145 2.222 51.2 2.43 ;
      RECT 51.1 2.22 51.145 2.433 ;
      RECT 51.072 2.22 51.085 2.436 ;
      RECT 50.986 2.224 51.072 2.438 ;
      RECT 50.9 2.23 50.986 2.443 ;
      RECT 50.88 2.234 50.9 2.445 ;
      RECT 50.878 2.235 50.88 2.444 ;
      RECT 50.792 2.237 50.878 2.443 ;
      RECT 50.706 2.242 50.792 2.44 ;
      RECT 50.62 2.247 50.706 2.437 ;
      RECT 50.47 2.25 50.55 2.433 ;
      RECT 51.13 5.015 51.3 8.305 ;
      RECT 51.13 7.315 51.535 7.645 ;
      RECT 51.13 6.475 51.535 6.805 ;
      RECT 51.246 3.225 51.295 3.559 ;
      RECT 51.246 3.225 51.3 3.558 ;
      RECT 51.16 3.225 51.3 3.557 ;
      RECT 50.935 3.333 51.305 3.555 ;
      RECT 51.16 3.225 51.33 3.548 ;
      RECT 51.13 3.237 51.335 3.539 ;
      RECT 51.115 3.255 51.34 3.536 ;
      RECT 50.93 3.339 51.34 3.463 ;
      RECT 50.925 3.346 51.34 3.423 ;
      RECT 50.94 3.312 51.34 3.536 ;
      RECT 51.101 3.258 51.305 3.555 ;
      RECT 51.015 3.278 51.34 3.536 ;
      RECT 51.115 3.252 51.335 3.539 ;
      RECT 50.885 2.576 51.075 2.77 ;
      RECT 50.88 2.578 51.075 2.769 ;
      RECT 50.875 2.582 51.09 2.766 ;
      RECT 50.89 2.575 51.09 2.766 ;
      RECT 50.875 2.685 51.095 2.761 ;
      RECT 50.17 3.185 50.261 3.483 ;
      RECT 50.165 3.187 50.34 3.478 ;
      RECT 50.17 3.185 50.34 3.478 ;
      RECT 50.165 3.191 50.36 3.476 ;
      RECT 50.165 3.246 50.4 3.475 ;
      RECT 50.165 3.281 50.415 3.469 ;
      RECT 50.165 3.315 50.425 3.459 ;
      RECT 50.155 3.195 50.36 3.31 ;
      RECT 50.155 3.215 50.375 3.31 ;
      RECT 50.155 3.198 50.365 3.31 ;
      RECT 50.38 1.966 50.385 2.028 ;
      RECT 50.375 1.888 50.38 2.051 ;
      RECT 50.37 1.845 50.375 2.062 ;
      RECT 50.365 1.835 50.37 2.074 ;
      RECT 50.36 1.835 50.365 2.083 ;
      RECT 50.335 1.835 50.36 2.115 ;
      RECT 50.33 1.835 50.335 2.148 ;
      RECT 50.315 1.835 50.33 2.173 ;
      RECT 50.305 1.835 50.315 2.2 ;
      RECT 50.3 1.835 50.305 2.213 ;
      RECT 50.295 1.835 50.3 2.228 ;
      RECT 50.285 1.835 50.295 2.243 ;
      RECT 50.28 1.835 50.285 2.263 ;
      RECT 50.255 1.835 50.28 2.298 ;
      RECT 50.21 1.835 50.255 2.343 ;
      RECT 50.2 1.835 50.21 2.356 ;
      RECT 50.115 1.92 50.2 2.363 ;
      RECT 50.08 2.042 50.115 2.372 ;
      RECT 50.075 2.082 50.08 2.376 ;
      RECT 50.055 2.105 50.075 2.378 ;
      RECT 50.05 2.135 50.055 2.381 ;
      RECT 50.04 2.147 50.05 2.382 ;
      RECT 49.995 2.17 50.04 2.387 ;
      RECT 49.955 2.2 49.995 2.395 ;
      RECT 49.92 2.212 49.955 2.401 ;
      RECT 49.915 2.217 49.92 2.405 ;
      RECT 49.845 2.227 49.915 2.412 ;
      RECT 49.805 2.237 49.845 2.422 ;
      RECT 49.785 2.242 49.805 2.428 ;
      RECT 49.775 2.246 49.785 2.433 ;
      RECT 49.77 2.249 49.775 2.436 ;
      RECT 49.76 2.25 49.77 2.437 ;
      RECT 49.735 2.252 49.76 2.441 ;
      RECT 49.725 2.257 49.735 2.444 ;
      RECT 49.68 2.265 49.725 2.445 ;
      RECT 49.555 2.27 49.68 2.445 ;
      RECT 50.11 2.567 50.13 2.749 ;
      RECT 50.061 2.552 50.11 2.748 ;
      RECT 49.975 2.567 50.13 2.746 ;
      RECT 49.96 2.567 50.13 2.745 ;
      RECT 49.925 2.545 50.095 2.73 ;
      RECT 49.995 3.565 50.01 3.774 ;
      RECT 49.995 3.573 50.015 3.773 ;
      RECT 49.94 3.573 50.015 3.772 ;
      RECT 49.92 3.577 50.02 3.77 ;
      RECT 49.9 3.527 49.94 3.769 ;
      RECT 49.845 3.585 50.025 3.767 ;
      RECT 49.81 3.542 49.94 3.765 ;
      RECT 49.806 3.545 49.995 3.764 ;
      RECT 49.72 3.553 49.995 3.762 ;
      RECT 49.72 3.597 50.03 3.755 ;
      RECT 49.71 3.69 50.03 3.753 ;
      RECT 49.72 3.609 50.035 3.738 ;
      RECT 49.72 3.63 50.05 3.708 ;
      RECT 49.72 3.657 50.055 3.678 ;
      RECT 49.845 3.535 49.94 3.767 ;
      RECT 49.475 2.58 49.48 3.118 ;
      RECT 49.28 2.91 49.285 3.105 ;
      RECT 47.58 2.575 47.595 2.955 ;
      RECT 49.645 2.575 49.65 2.745 ;
      RECT 49.64 2.575 49.645 2.755 ;
      RECT 49.635 2.575 49.64 2.768 ;
      RECT 49.61 2.575 49.635 2.81 ;
      RECT 49.585 2.575 49.61 2.883 ;
      RECT 49.57 2.575 49.585 2.935 ;
      RECT 49.565 2.575 49.57 2.965 ;
      RECT 49.54 2.575 49.565 3.005 ;
      RECT 49.525 2.575 49.54 3.06 ;
      RECT 49.52 2.575 49.525 3.093 ;
      RECT 49.495 2.575 49.52 3.113 ;
      RECT 49.48 2.575 49.495 3.119 ;
      RECT 49.41 2.61 49.475 3.115 ;
      RECT 49.36 2.665 49.41 3.11 ;
      RECT 49.35 2.697 49.36 3.108 ;
      RECT 49.345 2.722 49.35 3.108 ;
      RECT 49.325 2.795 49.345 3.108 ;
      RECT 49.315 2.875 49.325 3.107 ;
      RECT 49.3 2.905 49.315 3.107 ;
      RECT 49.285 2.91 49.3 3.106 ;
      RECT 49.225 2.912 49.28 3.103 ;
      RECT 49.195 2.917 49.225 3.099 ;
      RECT 49.193 2.92 49.195 3.098 ;
      RECT 49.107 2.922 49.193 3.095 ;
      RECT 49.021 2.928 49.107 3.089 ;
      RECT 48.935 2.933 49.021 3.083 ;
      RECT 48.862 2.938 48.935 3.084 ;
      RECT 48.776 2.944 48.862 3.092 ;
      RECT 48.69 2.95 48.776 3.101 ;
      RECT 48.67 2.954 48.69 3.106 ;
      RECT 48.623 2.956 48.67 3.109 ;
      RECT 48.537 2.961 48.623 3.115 ;
      RECT 48.451 2.966 48.537 3.124 ;
      RECT 48.365 2.972 48.451 3.132 ;
      RECT 48.28 2.97 48.365 3.141 ;
      RECT 48.276 2.965 48.28 3.145 ;
      RECT 48.19 2.96 48.276 3.137 ;
      RECT 48.126 2.951 48.19 3.125 ;
      RECT 48.04 2.942 48.126 3.112 ;
      RECT 48.016 2.935 48.04 3.103 ;
      RECT 47.93 2.929 48.016 3.09 ;
      RECT 47.89 2.922 47.93 3.076 ;
      RECT 47.885 2.912 47.89 3.072 ;
      RECT 47.875 2.9 47.885 3.071 ;
      RECT 47.855 2.87 47.875 3.068 ;
      RECT 47.8 2.79 47.855 3.062 ;
      RECT 47.78 2.709 47.8 3.057 ;
      RECT 47.76 2.667 47.78 3.053 ;
      RECT 47.735 2.62 47.76 3.047 ;
      RECT 47.73 2.595 47.735 3.044 ;
      RECT 47.695 2.575 47.73 3.039 ;
      RECT 47.686 2.575 47.695 3.032 ;
      RECT 47.6 2.575 47.686 3.002 ;
      RECT 47.595 2.575 47.6 2.965 ;
      RECT 47.56 2.575 47.58 2.887 ;
      RECT 47.555 2.617 47.56 2.852 ;
      RECT 47.55 2.692 47.555 2.808 ;
      RECT 49 2.497 49.175 2.745 ;
      RECT 49 2.497 49.18 2.743 ;
      RECT 48.995 2.529 49.18 2.703 ;
      RECT 49.025 2.47 49.195 2.69 ;
      RECT 48.99 2.547 49.195 2.623 ;
      RECT 48.3 2.01 48.47 2.185 ;
      RECT 48.3 2.01 48.642 2.177 ;
      RECT 48.3 2.01 48.725 2.171 ;
      RECT 48.3 2.01 48.76 2.167 ;
      RECT 48.3 2.01 48.78 2.166 ;
      RECT 48.3 2.01 48.866 2.162 ;
      RECT 48.76 1.835 48.93 2.157 ;
      RECT 48.335 1.942 48.96 2.155 ;
      RECT 48.325 1.997 48.965 2.153 ;
      RECT 48.3 2.033 48.975 2.148 ;
      RECT 48.3 2.06 48.98 2.078 ;
      RECT 48.365 1.885 48.94 2.155 ;
      RECT 48.556 1.87 48.94 2.155 ;
      RECT 48.39 1.873 48.94 2.155 ;
      RECT 48.47 1.871 48.556 2.182 ;
      RECT 48.556 1.868 48.935 2.155 ;
      RECT 48.74 1.845 48.935 2.155 ;
      RECT 48.642 1.866 48.935 2.155 ;
      RECT 48.725 1.86 48.74 2.168 ;
      RECT 48.875 3.225 48.88 3.425 ;
      RECT 48.34 3.29 48.385 3.425 ;
      RECT 48.91 3.225 48.93 3.398 ;
      RECT 48.88 3.225 48.91 3.413 ;
      RECT 48.815 3.225 48.875 3.45 ;
      RECT 48.8 3.225 48.815 3.48 ;
      RECT 48.785 3.225 48.8 3.493 ;
      RECT 48.765 3.225 48.785 3.508 ;
      RECT 48.76 3.225 48.765 3.517 ;
      RECT 48.75 3.229 48.76 3.522 ;
      RECT 48.735 3.239 48.75 3.533 ;
      RECT 48.71 3.255 48.735 3.543 ;
      RECT 48.7 3.269 48.71 3.545 ;
      RECT 48.68 3.281 48.7 3.542 ;
      RECT 48.65 3.302 48.68 3.536 ;
      RECT 48.64 3.314 48.65 3.531 ;
      RECT 48.63 3.312 48.64 3.528 ;
      RECT 48.615 3.311 48.63 3.523 ;
      RECT 48.61 3.31 48.615 3.518 ;
      RECT 48.575 3.308 48.61 3.508 ;
      RECT 48.555 3.305 48.575 3.49 ;
      RECT 48.545 3.303 48.555 3.485 ;
      RECT 48.535 3.302 48.545 3.48 ;
      RECT 48.5 3.3 48.535 3.468 ;
      RECT 48.445 3.296 48.5 3.448 ;
      RECT 48.435 3.294 48.445 3.433 ;
      RECT 48.43 3.294 48.435 3.428 ;
      RECT 48.385 3.292 48.43 3.425 ;
      RECT 48.29 3.29 48.34 3.429 ;
      RECT 48.28 3.291 48.29 3.434 ;
      RECT 48.22 3.298 48.28 3.448 ;
      RECT 48.195 3.306 48.22 3.468 ;
      RECT 48.185 3.31 48.195 3.48 ;
      RECT 48.18 3.311 48.185 3.485 ;
      RECT 48.165 3.313 48.18 3.488 ;
      RECT 48.15 3.315 48.165 3.493 ;
      RECT 48.145 3.315 48.15 3.496 ;
      RECT 48.1 3.32 48.145 3.507 ;
      RECT 48.095 3.324 48.1 3.519 ;
      RECT 48.07 3.32 48.095 3.523 ;
      RECT 48.06 3.316 48.07 3.527 ;
      RECT 48.05 3.315 48.06 3.531 ;
      RECT 48.035 3.305 48.05 3.537 ;
      RECT 48.03 3.293 48.035 3.541 ;
      RECT 48.025 3.29 48.03 3.542 ;
      RECT 48.02 3.287 48.025 3.544 ;
      RECT 48.005 3.275 48.02 3.543 ;
      RECT 47.99 3.257 48.005 3.54 ;
      RECT 47.97 3.236 47.99 3.533 ;
      RECT 47.905 3.225 47.97 3.505 ;
      RECT 47.901 3.225 47.905 3.484 ;
      RECT 47.815 3.225 47.901 3.454 ;
      RECT 47.8 3.225 47.815 3.41 ;
      RECT 48.375 2.325 48.38 2.56 ;
      RECT 47.505 2.241 47.51 2.445 ;
      RECT 48.085 2.27 48.09 2.425 ;
      RECT 48.005 2.25 48.01 2.425 ;
      RECT 48.675 2.392 48.69 2.745 ;
      RECT 48.601 2.377 48.675 2.745 ;
      RECT 48.515 2.36 48.601 2.745 ;
      RECT 48.505 2.35 48.515 2.743 ;
      RECT 48.5 2.348 48.505 2.738 ;
      RECT 48.485 2.346 48.5 2.724 ;
      RECT 48.415 2.338 48.485 2.664 ;
      RECT 48.395 2.329 48.415 2.598 ;
      RECT 48.39 2.326 48.395 2.578 ;
      RECT 48.38 2.325 48.39 2.568 ;
      RECT 48.37 2.325 48.375 2.552 ;
      RECT 48.36 2.324 48.37 2.542 ;
      RECT 48.35 2.322 48.36 2.53 ;
      RECT 48.335 2.319 48.35 2.51 ;
      RECT 48.325 2.317 48.335 2.495 ;
      RECT 48.305 2.314 48.325 2.483 ;
      RECT 48.3 2.312 48.305 2.473 ;
      RECT 48.275 2.31 48.3 2.46 ;
      RECT 48.245 2.305 48.275 2.445 ;
      RECT 48.165 2.296 48.245 2.436 ;
      RECT 48.12 2.285 48.165 2.429 ;
      RECT 48.1 2.276 48.12 2.426 ;
      RECT 48.09 2.271 48.1 2.425 ;
      RECT 48.045 2.265 48.085 2.425 ;
      RECT 48.03 2.257 48.045 2.425 ;
      RECT 48.01 2.252 48.03 2.425 ;
      RECT 47.99 2.249 48.005 2.425 ;
      RECT 47.907 2.248 47.99 2.424 ;
      RECT 47.821 2.247 47.907 2.42 ;
      RECT 47.735 2.245 47.821 2.417 ;
      RECT 47.682 2.244 47.735 2.419 ;
      RECT 47.596 2.243 47.682 2.428 ;
      RECT 47.51 2.242 47.596 2.44 ;
      RECT 47.49 2.241 47.505 2.448 ;
      RECT 47.41 2.24 47.49 2.46 ;
      RECT 47.385 2.24 47.41 2.473 ;
      RECT 47.36 2.24 47.385 2.488 ;
      RECT 47.355 2.24 47.36 2.51 ;
      RECT 47.35 2.24 47.355 2.528 ;
      RECT 47.345 2.24 47.35 2.545 ;
      RECT 47.34 2.24 47.345 2.558 ;
      RECT 47.335 2.24 47.34 2.568 ;
      RECT 47.295 2.24 47.335 2.653 ;
      RECT 47.28 2.24 47.295 2.738 ;
      RECT 47.27 2.241 47.28 2.75 ;
      RECT 47.235 2.246 47.27 2.755 ;
      RECT 47.195 2.255 47.235 2.755 ;
      RECT 47.18 2.265 47.195 2.755 ;
      RECT 47.175 2.275 47.18 2.755 ;
      RECT 47.155 2.302 47.175 2.755 ;
      RECT 47.105 2.385 47.155 2.755 ;
      RECT 47.1 2.447 47.105 2.755 ;
      RECT 47.09 2.46 47.1 2.755 ;
      RECT 47.08 2.482 47.09 2.755 ;
      RECT 47.07 2.507 47.08 2.75 ;
      RECT 47.065 2.545 47.07 2.743 ;
      RECT 47.055 2.655 47.065 2.738 ;
      RECT 48.45 3.576 48.465 3.835 ;
      RECT 48.45 3.591 48.47 3.834 ;
      RECT 48.366 3.591 48.47 3.832 ;
      RECT 48.366 3.605 48.475 3.831 ;
      RECT 48.28 3.647 48.48 3.828 ;
      RECT 48.275 3.59 48.465 3.823 ;
      RECT 48.275 3.661 48.485 3.82 ;
      RECT 48.27 3.692 48.485 3.818 ;
      RECT 48.275 3.689 48.5 3.808 ;
      RECT 48.27 3.735 48.515 3.793 ;
      RECT 48.27 3.763 48.52 3.778 ;
      RECT 48.28 3.565 48.45 3.828 ;
      RECT 48.04 2.575 48.21 2.745 ;
      RECT 48.005 2.575 48.21 2.74 ;
      RECT 47.995 2.575 48.21 2.733 ;
      RECT 47.99 2.56 48.16 2.73 ;
      RECT 46.82 3.097 47.085 3.54 ;
      RECT 46.815 3.068 47.03 3.538 ;
      RECT 46.81 3.222 47.09 3.533 ;
      RECT 46.815 3.117 47.09 3.533 ;
      RECT 46.815 3.128 47.1 3.52 ;
      RECT 46.815 3.075 47.06 3.538 ;
      RECT 46.82 3.062 47.03 3.54 ;
      RECT 46.82 3.06 46.98 3.54 ;
      RECT 46.921 3.052 46.98 3.54 ;
      RECT 46.835 3.053 46.98 3.54 ;
      RECT 46.921 3.051 46.97 3.54 ;
      RECT 46.725 1.866 46.9 2.165 ;
      RECT 46.775 1.828 46.9 2.165 ;
      RECT 46.76 1.83 46.986 2.157 ;
      RECT 46.76 1.833 47.025 2.144 ;
      RECT 46.76 1.834 47.035 2.13 ;
      RECT 46.715 1.885 47.035 2.12 ;
      RECT 46.76 1.835 47.04 2.115 ;
      RECT 46.715 2.045 47.045 2.105 ;
      RECT 46.7 1.905 47.04 2.045 ;
      RECT 46.695 1.921 47.04 1.985 ;
      RECT 46.74 1.845 47.04 2.115 ;
      RECT 46.775 1.826 46.861 2.165 ;
      RECT 44.87 1.74 45.04 2.935 ;
      RECT 44.87 1.74 45.335 1.91 ;
      RECT 44.87 6.97 45.335 7.14 ;
      RECT 44.87 5.945 45.04 7.14 ;
      RECT 43.88 1.74 44.05 2.935 ;
      RECT 43.88 1.74 44.345 1.91 ;
      RECT 43.88 6.97 44.345 7.14 ;
      RECT 43.88 5.945 44.05 7.14 ;
      RECT 42.025 2.635 42.195 3.865 ;
      RECT 42.08 0.855 42.25 2.805 ;
      RECT 42.025 0.575 42.195 1.025 ;
      RECT 42.025 7.855 42.195 8.305 ;
      RECT 42.08 6.075 42.25 8.025 ;
      RECT 42.025 5.015 42.195 6.245 ;
      RECT 41.505 0.575 41.675 3.865 ;
      RECT 41.505 2.075 41.91 2.405 ;
      RECT 41.505 1.235 41.91 1.565 ;
      RECT 41.505 5.015 41.675 8.305 ;
      RECT 41.505 7.315 41.91 7.645 ;
      RECT 41.505 6.475 41.91 6.805 ;
      RECT 39.43 3.126 39.435 3.298 ;
      RECT 39.425 3.119 39.43 3.388 ;
      RECT 39.42 3.113 39.425 3.407 ;
      RECT 39.4 3.107 39.42 3.417 ;
      RECT 39.385 3.102 39.4 3.425 ;
      RECT 39.348 3.096 39.385 3.423 ;
      RECT 39.262 3.082 39.348 3.419 ;
      RECT 39.176 3.064 39.262 3.414 ;
      RECT 39.09 3.045 39.176 3.408 ;
      RECT 39.06 3.033 39.09 3.404 ;
      RECT 39.04 3.027 39.06 3.403 ;
      RECT 38.975 3.025 39.04 3.401 ;
      RECT 38.96 3.025 38.975 3.393 ;
      RECT 38.945 3.025 38.96 3.38 ;
      RECT 38.94 3.025 38.945 3.37 ;
      RECT 38.925 3.025 38.94 3.348 ;
      RECT 38.91 3.025 38.925 3.315 ;
      RECT 38.905 3.025 38.91 3.293 ;
      RECT 38.895 3.025 38.905 3.275 ;
      RECT 38.88 3.025 38.895 3.253 ;
      RECT 38.86 3.025 38.88 3.215 ;
      RECT 39.21 2.31 39.245 2.749 ;
      RECT 39.21 2.31 39.25 2.748 ;
      RECT 39.155 2.37 39.25 2.747 ;
      RECT 39.02 2.542 39.25 2.746 ;
      RECT 39.13 2.42 39.25 2.746 ;
      RECT 39.02 2.542 39.275 2.736 ;
      RECT 39.075 2.487 39.355 2.653 ;
      RECT 39.25 2.281 39.255 2.744 ;
      RECT 39.105 2.457 39.395 2.53 ;
      RECT 39.12 2.44 39.25 2.746 ;
      RECT 39.255 2.28 39.425 2.468 ;
      RECT 39.245 2.283 39.425 2.468 ;
      RECT 38.75 2.16 38.92 2.47 ;
      RECT 38.75 2.16 38.925 2.443 ;
      RECT 38.75 2.16 38.93 2.42 ;
      RECT 38.75 2.16 38.94 2.37 ;
      RECT 38.745 2.265 38.94 2.34 ;
      RECT 38.78 1.835 38.95 2.313 ;
      RECT 38.78 1.835 38.965 2.234 ;
      RECT 38.77 2.045 38.965 2.234 ;
      RECT 38.78 1.845 38.975 2.149 ;
      RECT 38.71 2.587 38.715 2.79 ;
      RECT 38.7 2.575 38.71 2.9 ;
      RECT 38.675 2.575 38.7 2.94 ;
      RECT 38.595 2.575 38.675 3.025 ;
      RECT 38.585 2.575 38.595 3.095 ;
      RECT 38.56 2.575 38.585 3.118 ;
      RECT 38.54 2.575 38.56 3.153 ;
      RECT 38.495 2.585 38.54 3.196 ;
      RECT 38.485 2.597 38.495 3.233 ;
      RECT 38.465 2.611 38.485 3.253 ;
      RECT 38.455 2.629 38.465 3.269 ;
      RECT 38.44 2.655 38.455 3.279 ;
      RECT 38.425 2.696 38.44 3.293 ;
      RECT 38.415 2.731 38.425 3.303 ;
      RECT 38.41 2.747 38.415 3.308 ;
      RECT 38.4 2.762 38.41 3.313 ;
      RECT 38.38 2.805 38.4 3.323 ;
      RECT 38.36 2.842 38.38 3.336 ;
      RECT 38.325 2.865 38.36 3.354 ;
      RECT 38.315 2.879 38.325 3.37 ;
      RECT 38.295 2.889 38.315 3.38 ;
      RECT 38.29 2.898 38.295 3.388 ;
      RECT 38.28 2.905 38.29 3.395 ;
      RECT 38.27 2.912 38.28 3.403 ;
      RECT 38.255 2.922 38.27 3.411 ;
      RECT 38.245 2.936 38.255 3.421 ;
      RECT 38.235 2.948 38.245 3.433 ;
      RECT 38.22 2.97 38.235 3.446 ;
      RECT 38.21 2.992 38.22 3.457 ;
      RECT 38.2 3.012 38.21 3.466 ;
      RECT 38.195 3.027 38.2 3.473 ;
      RECT 38.165 3.06 38.195 3.487 ;
      RECT 38.155 3.095 38.165 3.502 ;
      RECT 38.15 3.102 38.155 3.508 ;
      RECT 38.13 3.117 38.15 3.515 ;
      RECT 38.125 3.132 38.13 3.523 ;
      RECT 38.12 3.141 38.125 3.528 ;
      RECT 38.105 3.147 38.12 3.535 ;
      RECT 38.1 3.153 38.105 3.543 ;
      RECT 38.095 3.157 38.1 3.55 ;
      RECT 38.09 3.161 38.095 3.56 ;
      RECT 38.08 3.166 38.09 3.57 ;
      RECT 38.06 3.177 38.08 3.598 ;
      RECT 38.045 3.189 38.06 3.625 ;
      RECT 38.025 3.202 38.045 3.65 ;
      RECT 38.005 3.217 38.025 3.674 ;
      RECT 37.99 3.232 38.005 3.689 ;
      RECT 37.985 3.243 37.99 3.698 ;
      RECT 37.92 3.288 37.985 3.708 ;
      RECT 37.885 3.347 37.92 3.721 ;
      RECT 37.88 3.37 37.885 3.727 ;
      RECT 37.875 3.377 37.88 3.729 ;
      RECT 37.86 3.387 37.875 3.732 ;
      RECT 37.83 3.412 37.86 3.736 ;
      RECT 37.825 3.43 37.83 3.74 ;
      RECT 37.82 3.437 37.825 3.741 ;
      RECT 37.8 3.445 37.82 3.745 ;
      RECT 37.79 3.452 37.8 3.749 ;
      RECT 37.746 3.463 37.79 3.756 ;
      RECT 37.66 3.491 37.746 3.772 ;
      RECT 37.6 3.515 37.66 3.79 ;
      RECT 37.555 3.525 37.6 3.804 ;
      RECT 37.496 3.533 37.555 3.818 ;
      RECT 37.41 3.54 37.496 3.837 ;
      RECT 37.385 3.545 37.41 3.852 ;
      RECT 37.305 3.548 37.385 3.855 ;
      RECT 37.225 3.552 37.305 3.842 ;
      RECT 37.216 3.555 37.225 3.827 ;
      RECT 37.13 3.555 37.216 3.812 ;
      RECT 37.07 3.557 37.13 3.789 ;
      RECT 37.066 3.56 37.07 3.779 ;
      RECT 36.98 3.56 37.066 3.764 ;
      RECT 36.905 3.56 36.98 3.74 ;
      RECT 38.22 2.569 38.23 2.745 ;
      RECT 38.175 2.536 38.22 2.745 ;
      RECT 38.13 2.487 38.175 2.745 ;
      RECT 38.1 2.457 38.13 2.746 ;
      RECT 38.095 2.44 38.1 2.747 ;
      RECT 38.07 2.42 38.095 2.748 ;
      RECT 38.055 2.395 38.07 2.749 ;
      RECT 38.05 2.382 38.055 2.75 ;
      RECT 38.045 2.376 38.05 2.748 ;
      RECT 38.04 2.368 38.045 2.742 ;
      RECT 38.015 2.36 38.04 2.722 ;
      RECT 37.995 2.349 38.015 2.693 ;
      RECT 37.965 2.334 37.995 2.664 ;
      RECT 37.945 2.32 37.965 2.636 ;
      RECT 37.935 2.314 37.945 2.615 ;
      RECT 37.93 2.311 37.935 2.598 ;
      RECT 37.925 2.308 37.93 2.583 ;
      RECT 37.91 2.303 37.925 2.548 ;
      RECT 37.905 2.299 37.91 2.515 ;
      RECT 37.885 2.294 37.905 2.491 ;
      RECT 37.855 2.286 37.885 2.456 ;
      RECT 37.84 2.28 37.855 2.433 ;
      RECT 37.8 2.273 37.84 2.418 ;
      RECT 37.775 2.265 37.8 2.398 ;
      RECT 37.755 2.26 37.775 2.388 ;
      RECT 37.72 2.254 37.755 2.383 ;
      RECT 37.675 2.245 37.72 2.382 ;
      RECT 37.645 2.241 37.675 2.384 ;
      RECT 37.56 2.249 37.645 2.388 ;
      RECT 37.49 2.26 37.56 2.41 ;
      RECT 37.477 2.266 37.49 2.433 ;
      RECT 37.391 2.273 37.477 2.455 ;
      RECT 37.305 2.285 37.391 2.492 ;
      RECT 37.305 2.662 37.315 2.9 ;
      RECT 37.3 2.291 37.305 2.515 ;
      RECT 37.295 2.547 37.305 2.9 ;
      RECT 37.295 2.292 37.3 2.52 ;
      RECT 37.29 2.293 37.295 2.9 ;
      RECT 37.266 2.295 37.29 2.901 ;
      RECT 37.18 2.303 37.266 2.903 ;
      RECT 37.16 2.317 37.18 2.906 ;
      RECT 37.155 2.345 37.16 2.907 ;
      RECT 37.15 2.357 37.155 2.908 ;
      RECT 37.145 2.372 37.15 2.909 ;
      RECT 37.135 2.402 37.145 2.91 ;
      RECT 37.13 2.44 37.135 2.908 ;
      RECT 37.125 2.46 37.13 2.903 ;
      RECT 37.11 2.495 37.125 2.888 ;
      RECT 37.1 2.547 37.11 2.868 ;
      RECT 37.095 2.577 37.1 2.856 ;
      RECT 37.08 2.59 37.095 2.839 ;
      RECT 37.055 2.594 37.08 2.806 ;
      RECT 37.04 2.592 37.055 2.783 ;
      RECT 37.025 2.591 37.04 2.78 ;
      RECT 36.965 2.589 37.025 2.778 ;
      RECT 36.955 2.587 36.965 2.773 ;
      RECT 36.915 2.586 36.955 2.77 ;
      RECT 36.845 2.583 36.915 2.768 ;
      RECT 36.79 2.581 36.845 2.763 ;
      RECT 36.72 2.575 36.79 2.758 ;
      RECT 36.711 2.575 36.72 2.755 ;
      RECT 36.625 2.575 36.711 2.75 ;
      RECT 36.62 2.575 36.625 2.745 ;
      RECT 37.925 1.81 38.1 2.16 ;
      RECT 37.925 1.825 38.11 2.158 ;
      RECT 37.9 1.775 38.045 2.155 ;
      RECT 37.88 1.776 38.045 2.148 ;
      RECT 37.87 1.777 38.055 2.143 ;
      RECT 37.84 1.778 38.055 2.13 ;
      RECT 37.79 1.779 38.055 2.106 ;
      RECT 37.785 1.781 38.055 2.091 ;
      RECT 37.785 1.847 38.115 2.085 ;
      RECT 37.765 1.788 38.07 2.065 ;
      RECT 37.755 1.797 38.08 1.92 ;
      RECT 37.765 1.792 38.08 2.065 ;
      RECT 37.785 1.782 38.07 2.091 ;
      RECT 37.37 3.107 37.54 3.395 ;
      RECT 37.365 3.125 37.55 3.39 ;
      RECT 37.33 3.133 37.615 3.31 ;
      RECT 37.33 3.133 37.701 3.3 ;
      RECT 37.33 3.133 37.755 3.246 ;
      RECT 37.615 3.03 37.785 3.214 ;
      RECT 37.33 3.185 37.79 3.202 ;
      RECT 37.315 3.155 37.785 3.198 ;
      RECT 37.575 3.037 37.615 3.349 ;
      RECT 37.455 3.074 37.785 3.214 ;
      RECT 37.55 3.049 37.575 3.375 ;
      RECT 37.54 3.056 37.785 3.214 ;
      RECT 37.671 2.52 37.74 2.779 ;
      RECT 37.671 2.575 37.745 2.778 ;
      RECT 37.585 2.575 37.745 2.777 ;
      RECT 37.58 2.575 37.75 2.77 ;
      RECT 37.57 2.52 37.74 2.765 ;
      RECT 36.95 1.819 37.125 2.12 ;
      RECT 36.935 1.807 36.95 2.105 ;
      RECT 36.905 1.806 36.935 2.058 ;
      RECT 36.905 1.824 37.13 2.053 ;
      RECT 36.89 1.808 36.95 2.018 ;
      RECT 36.885 1.83 37.14 1.918 ;
      RECT 36.885 1.813 37.036 1.918 ;
      RECT 36.885 1.815 37.04 1.918 ;
      RECT 36.89 1.811 37.036 2.018 ;
      RECT 36.995 3.047 37 3.395 ;
      RECT 36.985 3.037 36.995 3.401 ;
      RECT 36.95 3.027 36.985 3.403 ;
      RECT 36.912 3.022 36.95 3.407 ;
      RECT 36.826 3.015 36.912 3.414 ;
      RECT 36.74 3.005 36.826 3.424 ;
      RECT 36.695 3 36.74 3.432 ;
      RECT 36.691 3 36.695 3.436 ;
      RECT 36.605 3 36.691 3.443 ;
      RECT 36.59 3 36.605 3.443 ;
      RECT 36.58 2.998 36.59 3.415 ;
      RECT 36.57 2.994 36.58 3.358 ;
      RECT 36.55 2.988 36.57 3.29 ;
      RECT 36.545 2.984 36.55 3.238 ;
      RECT 36.535 2.983 36.545 3.205 ;
      RECT 36.485 2.981 36.535 3.19 ;
      RECT 36.46 2.979 36.485 3.185 ;
      RECT 36.417 2.977 36.46 3.181 ;
      RECT 36.331 2.973 36.417 3.169 ;
      RECT 36.245 2.968 36.331 3.153 ;
      RECT 36.215 2.965 36.245 3.14 ;
      RECT 36.19 2.964 36.215 3.128 ;
      RECT 36.185 2.964 36.19 3.118 ;
      RECT 36.145 2.963 36.185 3.11 ;
      RECT 36.13 2.962 36.145 3.103 ;
      RECT 36.08 2.961 36.13 3.095 ;
      RECT 36.078 2.96 36.08 3.09 ;
      RECT 35.992 2.958 36.078 3.09 ;
      RECT 35.906 2.953 35.992 3.09 ;
      RECT 35.82 2.949 35.906 3.09 ;
      RECT 35.771 2.945 35.82 3.088 ;
      RECT 35.685 2.942 35.771 3.083 ;
      RECT 35.662 2.939 35.685 3.079 ;
      RECT 35.576 2.936 35.662 3.074 ;
      RECT 35.49 2.932 35.576 3.065 ;
      RECT 35.465 2.925 35.49 3.06 ;
      RECT 35.405 2.89 35.465 3.057 ;
      RECT 35.385 2.815 35.405 3.054 ;
      RECT 35.38 2.757 35.385 3.053 ;
      RECT 35.355 2.697 35.38 3.052 ;
      RECT 35.28 2.575 35.355 3.048 ;
      RECT 35.27 2.575 35.28 3.04 ;
      RECT 35.255 2.575 35.27 3.03 ;
      RECT 35.24 2.575 35.255 3 ;
      RECT 35.225 2.575 35.24 2.945 ;
      RECT 35.21 2.575 35.225 2.883 ;
      RECT 35.185 2.575 35.21 2.808 ;
      RECT 35.18 2.575 35.185 2.758 ;
      RECT 36.525 2.12 36.545 2.429 ;
      RECT 36.511 2.122 36.56 2.426 ;
      RECT 36.511 2.127 36.58 2.417 ;
      RECT 36.425 2.125 36.56 2.411 ;
      RECT 36.425 2.133 36.615 2.394 ;
      RECT 36.39 2.135 36.615 2.393 ;
      RECT 36.36 2.143 36.615 2.384 ;
      RECT 36.35 2.148 36.635 2.37 ;
      RECT 36.39 2.138 36.635 2.37 ;
      RECT 36.39 2.141 36.645 2.358 ;
      RECT 36.36 2.143 36.655 2.345 ;
      RECT 36.36 2.147 36.665 2.288 ;
      RECT 36.35 2.152 36.67 2.203 ;
      RECT 36.511 2.12 36.545 2.426 ;
      RECT 36.39 7.855 36.56 8.305 ;
      RECT 36.445 6.075 36.615 8.025 ;
      RECT 36.39 5.015 36.56 6.245 ;
      RECT 35.95 2.223 35.955 2.435 ;
      RECT 35.825 2.22 35.84 2.435 ;
      RECT 35.29 2.25 35.36 2.435 ;
      RECT 35.175 2.25 35.21 2.43 ;
      RECT 36.296 2.552 36.315 2.746 ;
      RECT 36.21 2.507 36.296 2.747 ;
      RECT 36.2 2.46 36.21 2.749 ;
      RECT 36.195 2.44 36.2 2.75 ;
      RECT 36.175 2.405 36.195 2.751 ;
      RECT 36.16 2.355 36.175 2.752 ;
      RECT 36.14 2.292 36.16 2.753 ;
      RECT 36.13 2.255 36.14 2.754 ;
      RECT 36.115 2.244 36.13 2.755 ;
      RECT 36.11 2.236 36.115 2.753 ;
      RECT 36.1 2.235 36.11 2.745 ;
      RECT 36.07 2.232 36.1 2.724 ;
      RECT 35.995 2.227 36.07 2.669 ;
      RECT 35.98 2.223 35.995 2.615 ;
      RECT 35.97 2.223 35.98 2.51 ;
      RECT 35.955 2.223 35.97 2.443 ;
      RECT 35.94 2.223 35.95 2.433 ;
      RECT 35.885 2.222 35.94 2.43 ;
      RECT 35.84 2.22 35.885 2.433 ;
      RECT 35.812 2.22 35.825 2.436 ;
      RECT 35.726 2.224 35.812 2.438 ;
      RECT 35.64 2.23 35.726 2.443 ;
      RECT 35.62 2.234 35.64 2.445 ;
      RECT 35.618 2.235 35.62 2.444 ;
      RECT 35.532 2.237 35.618 2.443 ;
      RECT 35.446 2.242 35.532 2.44 ;
      RECT 35.36 2.247 35.446 2.437 ;
      RECT 35.21 2.25 35.29 2.433 ;
      RECT 35.87 5.015 36.04 8.305 ;
      RECT 35.87 7.315 36.275 7.645 ;
      RECT 35.87 6.475 36.275 6.805 ;
      RECT 35.986 3.225 36.035 3.559 ;
      RECT 35.986 3.225 36.04 3.558 ;
      RECT 35.9 3.225 36.04 3.557 ;
      RECT 35.675 3.333 36.045 3.555 ;
      RECT 35.9 3.225 36.07 3.548 ;
      RECT 35.87 3.237 36.075 3.539 ;
      RECT 35.855 3.255 36.08 3.536 ;
      RECT 35.67 3.339 36.08 3.463 ;
      RECT 35.665 3.346 36.08 3.423 ;
      RECT 35.68 3.312 36.08 3.536 ;
      RECT 35.841 3.258 36.045 3.555 ;
      RECT 35.755 3.278 36.08 3.536 ;
      RECT 35.855 3.252 36.075 3.539 ;
      RECT 35.625 2.576 35.815 2.77 ;
      RECT 35.62 2.578 35.815 2.769 ;
      RECT 35.615 2.582 35.83 2.766 ;
      RECT 35.63 2.575 35.83 2.766 ;
      RECT 35.615 2.685 35.835 2.761 ;
      RECT 34.91 3.185 35.001 3.483 ;
      RECT 34.905 3.187 35.08 3.478 ;
      RECT 34.91 3.185 35.08 3.478 ;
      RECT 34.905 3.191 35.1 3.476 ;
      RECT 34.905 3.246 35.14 3.475 ;
      RECT 34.905 3.281 35.155 3.469 ;
      RECT 34.905 3.315 35.165 3.459 ;
      RECT 34.895 3.195 35.1 3.31 ;
      RECT 34.895 3.215 35.115 3.31 ;
      RECT 34.895 3.198 35.105 3.31 ;
      RECT 35.12 1.966 35.125 2.028 ;
      RECT 35.115 1.888 35.12 2.051 ;
      RECT 35.11 1.845 35.115 2.062 ;
      RECT 35.105 1.835 35.11 2.074 ;
      RECT 35.1 1.835 35.105 2.083 ;
      RECT 35.075 1.835 35.1 2.115 ;
      RECT 35.07 1.835 35.075 2.148 ;
      RECT 35.055 1.835 35.07 2.173 ;
      RECT 35.045 1.835 35.055 2.2 ;
      RECT 35.04 1.835 35.045 2.213 ;
      RECT 35.035 1.835 35.04 2.228 ;
      RECT 35.025 1.835 35.035 2.243 ;
      RECT 35.02 1.835 35.025 2.263 ;
      RECT 34.995 1.835 35.02 2.298 ;
      RECT 34.95 1.835 34.995 2.343 ;
      RECT 34.94 1.835 34.95 2.356 ;
      RECT 34.855 1.92 34.94 2.363 ;
      RECT 34.82 2.042 34.855 2.372 ;
      RECT 34.815 2.082 34.82 2.376 ;
      RECT 34.795 2.105 34.815 2.378 ;
      RECT 34.79 2.135 34.795 2.381 ;
      RECT 34.78 2.147 34.79 2.382 ;
      RECT 34.735 2.17 34.78 2.387 ;
      RECT 34.695 2.2 34.735 2.395 ;
      RECT 34.66 2.212 34.695 2.401 ;
      RECT 34.655 2.217 34.66 2.405 ;
      RECT 34.585 2.227 34.655 2.412 ;
      RECT 34.545 2.237 34.585 2.422 ;
      RECT 34.525 2.242 34.545 2.428 ;
      RECT 34.515 2.246 34.525 2.433 ;
      RECT 34.51 2.249 34.515 2.436 ;
      RECT 34.5 2.25 34.51 2.437 ;
      RECT 34.475 2.252 34.5 2.441 ;
      RECT 34.465 2.257 34.475 2.444 ;
      RECT 34.42 2.265 34.465 2.445 ;
      RECT 34.295 2.27 34.42 2.445 ;
      RECT 34.85 2.567 34.87 2.749 ;
      RECT 34.801 2.552 34.85 2.748 ;
      RECT 34.715 2.567 34.87 2.746 ;
      RECT 34.7 2.567 34.87 2.745 ;
      RECT 34.665 2.545 34.835 2.73 ;
      RECT 34.735 3.565 34.75 3.774 ;
      RECT 34.735 3.573 34.755 3.773 ;
      RECT 34.68 3.573 34.755 3.772 ;
      RECT 34.66 3.577 34.76 3.77 ;
      RECT 34.64 3.527 34.68 3.769 ;
      RECT 34.585 3.585 34.765 3.767 ;
      RECT 34.55 3.542 34.68 3.765 ;
      RECT 34.546 3.545 34.735 3.764 ;
      RECT 34.46 3.553 34.735 3.762 ;
      RECT 34.46 3.597 34.77 3.755 ;
      RECT 34.45 3.69 34.77 3.753 ;
      RECT 34.46 3.609 34.775 3.738 ;
      RECT 34.46 3.63 34.79 3.708 ;
      RECT 34.46 3.657 34.795 3.678 ;
      RECT 34.585 3.535 34.68 3.767 ;
      RECT 34.215 2.58 34.22 3.118 ;
      RECT 34.02 2.91 34.025 3.105 ;
      RECT 32.32 2.575 32.335 2.955 ;
      RECT 34.385 2.575 34.39 2.745 ;
      RECT 34.38 2.575 34.385 2.755 ;
      RECT 34.375 2.575 34.38 2.768 ;
      RECT 34.35 2.575 34.375 2.81 ;
      RECT 34.325 2.575 34.35 2.883 ;
      RECT 34.31 2.575 34.325 2.935 ;
      RECT 34.305 2.575 34.31 2.965 ;
      RECT 34.28 2.575 34.305 3.005 ;
      RECT 34.265 2.575 34.28 3.06 ;
      RECT 34.26 2.575 34.265 3.093 ;
      RECT 34.235 2.575 34.26 3.113 ;
      RECT 34.22 2.575 34.235 3.119 ;
      RECT 34.15 2.61 34.215 3.115 ;
      RECT 34.1 2.665 34.15 3.11 ;
      RECT 34.09 2.697 34.1 3.108 ;
      RECT 34.085 2.722 34.09 3.108 ;
      RECT 34.065 2.795 34.085 3.108 ;
      RECT 34.055 2.875 34.065 3.107 ;
      RECT 34.04 2.905 34.055 3.107 ;
      RECT 34.025 2.91 34.04 3.106 ;
      RECT 33.965 2.912 34.02 3.103 ;
      RECT 33.935 2.917 33.965 3.099 ;
      RECT 33.933 2.92 33.935 3.098 ;
      RECT 33.847 2.922 33.933 3.095 ;
      RECT 33.761 2.928 33.847 3.089 ;
      RECT 33.675 2.933 33.761 3.083 ;
      RECT 33.602 2.938 33.675 3.084 ;
      RECT 33.516 2.944 33.602 3.092 ;
      RECT 33.43 2.95 33.516 3.101 ;
      RECT 33.41 2.954 33.43 3.106 ;
      RECT 33.363 2.956 33.41 3.109 ;
      RECT 33.277 2.961 33.363 3.115 ;
      RECT 33.191 2.966 33.277 3.124 ;
      RECT 33.105 2.972 33.191 3.132 ;
      RECT 33.02 2.97 33.105 3.141 ;
      RECT 33.016 2.965 33.02 3.145 ;
      RECT 32.93 2.96 33.016 3.137 ;
      RECT 32.866 2.951 32.93 3.125 ;
      RECT 32.78 2.942 32.866 3.112 ;
      RECT 32.756 2.935 32.78 3.103 ;
      RECT 32.67 2.929 32.756 3.09 ;
      RECT 32.63 2.922 32.67 3.076 ;
      RECT 32.625 2.912 32.63 3.072 ;
      RECT 32.615 2.9 32.625 3.071 ;
      RECT 32.595 2.87 32.615 3.068 ;
      RECT 32.54 2.79 32.595 3.062 ;
      RECT 32.52 2.709 32.54 3.057 ;
      RECT 32.5 2.667 32.52 3.053 ;
      RECT 32.475 2.62 32.5 3.047 ;
      RECT 32.47 2.595 32.475 3.044 ;
      RECT 32.435 2.575 32.47 3.039 ;
      RECT 32.426 2.575 32.435 3.032 ;
      RECT 32.34 2.575 32.426 3.002 ;
      RECT 32.335 2.575 32.34 2.965 ;
      RECT 32.3 2.575 32.32 2.887 ;
      RECT 32.295 2.617 32.3 2.852 ;
      RECT 32.29 2.692 32.295 2.808 ;
      RECT 33.74 2.497 33.915 2.745 ;
      RECT 33.74 2.497 33.92 2.743 ;
      RECT 33.735 2.529 33.92 2.703 ;
      RECT 33.765 2.47 33.935 2.69 ;
      RECT 33.73 2.547 33.935 2.623 ;
      RECT 33.04 2.01 33.21 2.185 ;
      RECT 33.04 2.01 33.382 2.177 ;
      RECT 33.04 2.01 33.465 2.171 ;
      RECT 33.04 2.01 33.5 2.167 ;
      RECT 33.04 2.01 33.52 2.166 ;
      RECT 33.04 2.01 33.606 2.162 ;
      RECT 33.5 1.835 33.67 2.157 ;
      RECT 33.075 1.942 33.7 2.155 ;
      RECT 33.065 1.997 33.705 2.153 ;
      RECT 33.04 2.033 33.715 2.148 ;
      RECT 33.04 2.06 33.72 2.078 ;
      RECT 33.105 1.885 33.68 2.155 ;
      RECT 33.296 1.87 33.68 2.155 ;
      RECT 33.13 1.873 33.68 2.155 ;
      RECT 33.21 1.871 33.296 2.182 ;
      RECT 33.296 1.868 33.675 2.155 ;
      RECT 33.48 1.845 33.675 2.155 ;
      RECT 33.382 1.866 33.675 2.155 ;
      RECT 33.465 1.86 33.48 2.168 ;
      RECT 33.615 3.225 33.62 3.425 ;
      RECT 33.08 3.29 33.125 3.425 ;
      RECT 33.65 3.225 33.67 3.398 ;
      RECT 33.62 3.225 33.65 3.413 ;
      RECT 33.555 3.225 33.615 3.45 ;
      RECT 33.54 3.225 33.555 3.48 ;
      RECT 33.525 3.225 33.54 3.493 ;
      RECT 33.505 3.225 33.525 3.508 ;
      RECT 33.5 3.225 33.505 3.517 ;
      RECT 33.49 3.229 33.5 3.522 ;
      RECT 33.475 3.239 33.49 3.533 ;
      RECT 33.45 3.255 33.475 3.543 ;
      RECT 33.44 3.269 33.45 3.545 ;
      RECT 33.42 3.281 33.44 3.542 ;
      RECT 33.39 3.302 33.42 3.536 ;
      RECT 33.38 3.314 33.39 3.531 ;
      RECT 33.37 3.312 33.38 3.528 ;
      RECT 33.355 3.311 33.37 3.523 ;
      RECT 33.35 3.31 33.355 3.518 ;
      RECT 33.315 3.308 33.35 3.508 ;
      RECT 33.295 3.305 33.315 3.49 ;
      RECT 33.285 3.303 33.295 3.485 ;
      RECT 33.275 3.302 33.285 3.48 ;
      RECT 33.24 3.3 33.275 3.468 ;
      RECT 33.185 3.296 33.24 3.448 ;
      RECT 33.175 3.294 33.185 3.433 ;
      RECT 33.17 3.294 33.175 3.428 ;
      RECT 33.125 3.292 33.17 3.425 ;
      RECT 33.03 3.29 33.08 3.429 ;
      RECT 33.02 3.291 33.03 3.434 ;
      RECT 32.96 3.298 33.02 3.448 ;
      RECT 32.935 3.306 32.96 3.468 ;
      RECT 32.925 3.31 32.935 3.48 ;
      RECT 32.92 3.311 32.925 3.485 ;
      RECT 32.905 3.313 32.92 3.488 ;
      RECT 32.89 3.315 32.905 3.493 ;
      RECT 32.885 3.315 32.89 3.496 ;
      RECT 32.84 3.32 32.885 3.507 ;
      RECT 32.835 3.324 32.84 3.519 ;
      RECT 32.81 3.32 32.835 3.523 ;
      RECT 32.8 3.316 32.81 3.527 ;
      RECT 32.79 3.315 32.8 3.531 ;
      RECT 32.775 3.305 32.79 3.537 ;
      RECT 32.77 3.293 32.775 3.541 ;
      RECT 32.765 3.29 32.77 3.542 ;
      RECT 32.76 3.287 32.765 3.544 ;
      RECT 32.745 3.275 32.76 3.543 ;
      RECT 32.73 3.257 32.745 3.54 ;
      RECT 32.71 3.236 32.73 3.533 ;
      RECT 32.645 3.225 32.71 3.505 ;
      RECT 32.641 3.225 32.645 3.484 ;
      RECT 32.555 3.225 32.641 3.454 ;
      RECT 32.54 3.225 32.555 3.41 ;
      RECT 33.115 2.325 33.12 2.56 ;
      RECT 32.245 2.241 32.25 2.445 ;
      RECT 32.825 2.27 32.83 2.425 ;
      RECT 32.745 2.25 32.75 2.425 ;
      RECT 33.415 2.392 33.43 2.745 ;
      RECT 33.341 2.377 33.415 2.745 ;
      RECT 33.255 2.36 33.341 2.745 ;
      RECT 33.245 2.35 33.255 2.743 ;
      RECT 33.24 2.348 33.245 2.738 ;
      RECT 33.225 2.346 33.24 2.724 ;
      RECT 33.155 2.338 33.225 2.664 ;
      RECT 33.135 2.329 33.155 2.598 ;
      RECT 33.13 2.326 33.135 2.578 ;
      RECT 33.12 2.325 33.13 2.568 ;
      RECT 33.11 2.325 33.115 2.552 ;
      RECT 33.1 2.324 33.11 2.542 ;
      RECT 33.09 2.322 33.1 2.53 ;
      RECT 33.075 2.319 33.09 2.51 ;
      RECT 33.065 2.317 33.075 2.495 ;
      RECT 33.045 2.314 33.065 2.483 ;
      RECT 33.04 2.312 33.045 2.473 ;
      RECT 33.015 2.31 33.04 2.46 ;
      RECT 32.985 2.305 33.015 2.445 ;
      RECT 32.905 2.296 32.985 2.436 ;
      RECT 32.86 2.285 32.905 2.429 ;
      RECT 32.84 2.276 32.86 2.426 ;
      RECT 32.83 2.271 32.84 2.425 ;
      RECT 32.785 2.265 32.825 2.425 ;
      RECT 32.77 2.257 32.785 2.425 ;
      RECT 32.75 2.252 32.77 2.425 ;
      RECT 32.73 2.249 32.745 2.425 ;
      RECT 32.647 2.248 32.73 2.424 ;
      RECT 32.561 2.247 32.647 2.42 ;
      RECT 32.475 2.245 32.561 2.417 ;
      RECT 32.422 2.244 32.475 2.419 ;
      RECT 32.336 2.243 32.422 2.428 ;
      RECT 32.25 2.242 32.336 2.44 ;
      RECT 32.23 2.241 32.245 2.448 ;
      RECT 32.15 2.24 32.23 2.46 ;
      RECT 32.125 2.24 32.15 2.473 ;
      RECT 32.1 2.24 32.125 2.488 ;
      RECT 32.095 2.24 32.1 2.51 ;
      RECT 32.09 2.24 32.095 2.528 ;
      RECT 32.085 2.24 32.09 2.545 ;
      RECT 32.08 2.24 32.085 2.558 ;
      RECT 32.075 2.24 32.08 2.568 ;
      RECT 32.035 2.24 32.075 2.653 ;
      RECT 32.02 2.24 32.035 2.738 ;
      RECT 32.01 2.241 32.02 2.75 ;
      RECT 31.975 2.246 32.01 2.755 ;
      RECT 31.935 2.255 31.975 2.755 ;
      RECT 31.92 2.265 31.935 2.755 ;
      RECT 31.915 2.275 31.92 2.755 ;
      RECT 31.895 2.302 31.915 2.755 ;
      RECT 31.845 2.385 31.895 2.755 ;
      RECT 31.84 2.447 31.845 2.755 ;
      RECT 31.83 2.46 31.84 2.755 ;
      RECT 31.82 2.482 31.83 2.755 ;
      RECT 31.81 2.507 31.82 2.75 ;
      RECT 31.805 2.545 31.81 2.743 ;
      RECT 31.795 2.655 31.805 2.738 ;
      RECT 33.19 3.576 33.205 3.835 ;
      RECT 33.19 3.591 33.21 3.834 ;
      RECT 33.106 3.591 33.21 3.832 ;
      RECT 33.106 3.605 33.215 3.831 ;
      RECT 33.02 3.647 33.22 3.828 ;
      RECT 33.015 3.59 33.205 3.823 ;
      RECT 33.015 3.661 33.225 3.82 ;
      RECT 33.01 3.692 33.225 3.818 ;
      RECT 33.015 3.689 33.24 3.808 ;
      RECT 33.01 3.735 33.255 3.793 ;
      RECT 33.01 3.763 33.26 3.778 ;
      RECT 33.02 3.565 33.19 3.828 ;
      RECT 32.78 2.575 32.95 2.745 ;
      RECT 32.745 2.575 32.95 2.74 ;
      RECT 32.735 2.575 32.95 2.733 ;
      RECT 32.73 2.56 32.9 2.73 ;
      RECT 31.56 3.097 31.825 3.54 ;
      RECT 31.555 3.068 31.77 3.538 ;
      RECT 31.55 3.222 31.83 3.533 ;
      RECT 31.555 3.117 31.83 3.533 ;
      RECT 31.555 3.128 31.84 3.52 ;
      RECT 31.555 3.075 31.8 3.538 ;
      RECT 31.56 3.062 31.77 3.54 ;
      RECT 31.56 3.06 31.72 3.54 ;
      RECT 31.661 3.052 31.72 3.54 ;
      RECT 31.575 3.053 31.72 3.54 ;
      RECT 31.661 3.051 31.71 3.54 ;
      RECT 31.465 1.866 31.64 2.165 ;
      RECT 31.515 1.828 31.64 2.165 ;
      RECT 31.5 1.83 31.726 2.157 ;
      RECT 31.5 1.833 31.765 2.144 ;
      RECT 31.5 1.834 31.775 2.13 ;
      RECT 31.455 1.885 31.775 2.12 ;
      RECT 31.5 1.835 31.78 2.115 ;
      RECT 31.455 2.045 31.785 2.105 ;
      RECT 31.44 1.905 31.78 2.045 ;
      RECT 31.435 1.921 31.78 1.985 ;
      RECT 31.48 1.845 31.78 2.115 ;
      RECT 31.515 1.826 31.601 2.165 ;
      RECT 29.61 1.74 29.78 2.935 ;
      RECT 29.61 1.74 30.075 1.91 ;
      RECT 29.61 6.97 30.075 7.14 ;
      RECT 29.61 5.945 29.78 7.14 ;
      RECT 28.62 1.74 28.79 2.935 ;
      RECT 28.62 1.74 29.085 1.91 ;
      RECT 28.62 6.97 29.085 7.14 ;
      RECT 28.62 5.945 28.79 7.14 ;
      RECT 26.765 2.635 26.935 3.865 ;
      RECT 26.82 0.855 26.99 2.805 ;
      RECT 26.765 0.575 26.935 1.025 ;
      RECT 26.765 7.855 26.935 8.305 ;
      RECT 26.82 6.075 26.99 8.025 ;
      RECT 26.765 5.015 26.935 6.245 ;
      RECT 26.245 0.575 26.415 3.865 ;
      RECT 26.245 2.075 26.65 2.405 ;
      RECT 26.245 1.235 26.65 1.565 ;
      RECT 26.245 5.015 26.415 8.305 ;
      RECT 26.245 7.315 26.65 7.645 ;
      RECT 26.245 6.475 26.65 6.805 ;
      RECT 24.17 3.126 24.175 3.298 ;
      RECT 24.165 3.119 24.17 3.388 ;
      RECT 24.16 3.113 24.165 3.407 ;
      RECT 24.14 3.107 24.16 3.417 ;
      RECT 24.125 3.102 24.14 3.425 ;
      RECT 24.088 3.096 24.125 3.423 ;
      RECT 24.002 3.082 24.088 3.419 ;
      RECT 23.916 3.064 24.002 3.414 ;
      RECT 23.83 3.045 23.916 3.408 ;
      RECT 23.8 3.033 23.83 3.404 ;
      RECT 23.78 3.027 23.8 3.403 ;
      RECT 23.715 3.025 23.78 3.401 ;
      RECT 23.7 3.025 23.715 3.393 ;
      RECT 23.685 3.025 23.7 3.38 ;
      RECT 23.68 3.025 23.685 3.37 ;
      RECT 23.665 3.025 23.68 3.348 ;
      RECT 23.65 3.025 23.665 3.315 ;
      RECT 23.645 3.025 23.65 3.293 ;
      RECT 23.635 3.025 23.645 3.275 ;
      RECT 23.62 3.025 23.635 3.253 ;
      RECT 23.6 3.025 23.62 3.215 ;
      RECT 23.95 2.31 23.985 2.749 ;
      RECT 23.95 2.31 23.99 2.748 ;
      RECT 23.895 2.37 23.99 2.747 ;
      RECT 23.76 2.542 23.99 2.746 ;
      RECT 23.87 2.42 23.99 2.746 ;
      RECT 23.76 2.542 24.015 2.736 ;
      RECT 23.815 2.487 24.095 2.653 ;
      RECT 23.99 2.281 23.995 2.744 ;
      RECT 23.845 2.457 24.135 2.53 ;
      RECT 23.86 2.44 23.99 2.746 ;
      RECT 23.995 2.28 24.165 2.468 ;
      RECT 23.985 2.283 24.165 2.468 ;
      RECT 23.49 2.16 23.66 2.47 ;
      RECT 23.49 2.16 23.665 2.443 ;
      RECT 23.49 2.16 23.67 2.42 ;
      RECT 23.49 2.16 23.68 2.37 ;
      RECT 23.485 2.265 23.68 2.34 ;
      RECT 23.52 1.835 23.69 2.313 ;
      RECT 23.52 1.835 23.705 2.234 ;
      RECT 23.51 2.045 23.705 2.234 ;
      RECT 23.52 1.845 23.715 2.149 ;
      RECT 23.45 2.587 23.455 2.79 ;
      RECT 23.44 2.575 23.45 2.9 ;
      RECT 23.415 2.575 23.44 2.94 ;
      RECT 23.335 2.575 23.415 3.025 ;
      RECT 23.325 2.575 23.335 3.095 ;
      RECT 23.3 2.575 23.325 3.118 ;
      RECT 23.28 2.575 23.3 3.153 ;
      RECT 23.235 2.585 23.28 3.196 ;
      RECT 23.225 2.597 23.235 3.233 ;
      RECT 23.205 2.611 23.225 3.253 ;
      RECT 23.195 2.629 23.205 3.269 ;
      RECT 23.18 2.655 23.195 3.279 ;
      RECT 23.165 2.696 23.18 3.293 ;
      RECT 23.155 2.731 23.165 3.303 ;
      RECT 23.15 2.747 23.155 3.308 ;
      RECT 23.14 2.762 23.15 3.313 ;
      RECT 23.12 2.805 23.14 3.323 ;
      RECT 23.1 2.842 23.12 3.336 ;
      RECT 23.065 2.865 23.1 3.354 ;
      RECT 23.055 2.879 23.065 3.37 ;
      RECT 23.035 2.889 23.055 3.38 ;
      RECT 23.03 2.898 23.035 3.388 ;
      RECT 23.02 2.905 23.03 3.395 ;
      RECT 23.01 2.912 23.02 3.403 ;
      RECT 22.995 2.922 23.01 3.411 ;
      RECT 22.985 2.936 22.995 3.421 ;
      RECT 22.975 2.948 22.985 3.433 ;
      RECT 22.96 2.97 22.975 3.446 ;
      RECT 22.95 2.992 22.96 3.457 ;
      RECT 22.94 3.012 22.95 3.466 ;
      RECT 22.935 3.027 22.94 3.473 ;
      RECT 22.905 3.06 22.935 3.487 ;
      RECT 22.895 3.095 22.905 3.502 ;
      RECT 22.89 3.102 22.895 3.508 ;
      RECT 22.87 3.117 22.89 3.515 ;
      RECT 22.865 3.132 22.87 3.523 ;
      RECT 22.86 3.141 22.865 3.528 ;
      RECT 22.845 3.147 22.86 3.535 ;
      RECT 22.84 3.153 22.845 3.543 ;
      RECT 22.835 3.157 22.84 3.55 ;
      RECT 22.83 3.161 22.835 3.56 ;
      RECT 22.82 3.166 22.83 3.57 ;
      RECT 22.8 3.177 22.82 3.598 ;
      RECT 22.785 3.189 22.8 3.625 ;
      RECT 22.765 3.202 22.785 3.65 ;
      RECT 22.745 3.217 22.765 3.674 ;
      RECT 22.73 3.232 22.745 3.689 ;
      RECT 22.725 3.243 22.73 3.698 ;
      RECT 22.66 3.288 22.725 3.708 ;
      RECT 22.625 3.347 22.66 3.721 ;
      RECT 22.62 3.37 22.625 3.727 ;
      RECT 22.615 3.377 22.62 3.729 ;
      RECT 22.6 3.387 22.615 3.732 ;
      RECT 22.57 3.412 22.6 3.736 ;
      RECT 22.565 3.43 22.57 3.74 ;
      RECT 22.56 3.437 22.565 3.741 ;
      RECT 22.54 3.445 22.56 3.745 ;
      RECT 22.53 3.452 22.54 3.749 ;
      RECT 22.486 3.463 22.53 3.756 ;
      RECT 22.4 3.491 22.486 3.772 ;
      RECT 22.34 3.515 22.4 3.79 ;
      RECT 22.295 3.525 22.34 3.804 ;
      RECT 22.236 3.533 22.295 3.818 ;
      RECT 22.15 3.54 22.236 3.837 ;
      RECT 22.125 3.545 22.15 3.852 ;
      RECT 22.045 3.548 22.125 3.855 ;
      RECT 21.965 3.552 22.045 3.842 ;
      RECT 21.956 3.555 21.965 3.827 ;
      RECT 21.87 3.555 21.956 3.812 ;
      RECT 21.81 3.557 21.87 3.789 ;
      RECT 21.806 3.56 21.81 3.779 ;
      RECT 21.72 3.56 21.806 3.764 ;
      RECT 21.645 3.56 21.72 3.74 ;
      RECT 22.96 2.569 22.97 2.745 ;
      RECT 22.915 2.536 22.96 2.745 ;
      RECT 22.87 2.487 22.915 2.745 ;
      RECT 22.84 2.457 22.87 2.746 ;
      RECT 22.835 2.44 22.84 2.747 ;
      RECT 22.81 2.42 22.835 2.748 ;
      RECT 22.795 2.395 22.81 2.749 ;
      RECT 22.79 2.382 22.795 2.75 ;
      RECT 22.785 2.376 22.79 2.748 ;
      RECT 22.78 2.368 22.785 2.742 ;
      RECT 22.755 2.36 22.78 2.722 ;
      RECT 22.735 2.349 22.755 2.693 ;
      RECT 22.705 2.334 22.735 2.664 ;
      RECT 22.685 2.32 22.705 2.636 ;
      RECT 22.675 2.314 22.685 2.615 ;
      RECT 22.67 2.311 22.675 2.598 ;
      RECT 22.665 2.308 22.67 2.583 ;
      RECT 22.65 2.303 22.665 2.548 ;
      RECT 22.645 2.299 22.65 2.515 ;
      RECT 22.625 2.294 22.645 2.491 ;
      RECT 22.595 2.286 22.625 2.456 ;
      RECT 22.58 2.28 22.595 2.433 ;
      RECT 22.54 2.273 22.58 2.418 ;
      RECT 22.515 2.265 22.54 2.398 ;
      RECT 22.495 2.26 22.515 2.388 ;
      RECT 22.46 2.254 22.495 2.383 ;
      RECT 22.415 2.245 22.46 2.382 ;
      RECT 22.385 2.241 22.415 2.384 ;
      RECT 22.3 2.249 22.385 2.388 ;
      RECT 22.23 2.26 22.3 2.41 ;
      RECT 22.217 2.266 22.23 2.433 ;
      RECT 22.131 2.273 22.217 2.455 ;
      RECT 22.045 2.285 22.131 2.492 ;
      RECT 22.045 2.662 22.055 2.9 ;
      RECT 22.04 2.291 22.045 2.515 ;
      RECT 22.035 2.547 22.045 2.9 ;
      RECT 22.035 2.292 22.04 2.52 ;
      RECT 22.03 2.293 22.035 2.9 ;
      RECT 22.006 2.295 22.03 2.901 ;
      RECT 21.92 2.303 22.006 2.903 ;
      RECT 21.9 2.317 21.92 2.906 ;
      RECT 21.895 2.345 21.9 2.907 ;
      RECT 21.89 2.357 21.895 2.908 ;
      RECT 21.885 2.372 21.89 2.909 ;
      RECT 21.875 2.402 21.885 2.91 ;
      RECT 21.87 2.44 21.875 2.908 ;
      RECT 21.865 2.46 21.87 2.903 ;
      RECT 21.85 2.495 21.865 2.888 ;
      RECT 21.84 2.547 21.85 2.868 ;
      RECT 21.835 2.577 21.84 2.856 ;
      RECT 21.82 2.59 21.835 2.839 ;
      RECT 21.795 2.594 21.82 2.806 ;
      RECT 21.78 2.592 21.795 2.783 ;
      RECT 21.765 2.591 21.78 2.78 ;
      RECT 21.705 2.589 21.765 2.778 ;
      RECT 21.695 2.587 21.705 2.773 ;
      RECT 21.655 2.586 21.695 2.77 ;
      RECT 21.585 2.583 21.655 2.768 ;
      RECT 21.53 2.581 21.585 2.763 ;
      RECT 21.46 2.575 21.53 2.758 ;
      RECT 21.451 2.575 21.46 2.755 ;
      RECT 21.365 2.575 21.451 2.75 ;
      RECT 21.36 2.575 21.365 2.745 ;
      RECT 22.665 1.81 22.84 2.16 ;
      RECT 22.665 1.825 22.85 2.158 ;
      RECT 22.64 1.775 22.785 2.155 ;
      RECT 22.62 1.776 22.785 2.148 ;
      RECT 22.61 1.777 22.795 2.143 ;
      RECT 22.58 1.778 22.795 2.13 ;
      RECT 22.53 1.779 22.795 2.106 ;
      RECT 22.525 1.781 22.795 2.091 ;
      RECT 22.525 1.847 22.855 2.085 ;
      RECT 22.505 1.788 22.81 2.065 ;
      RECT 22.495 1.797 22.82 1.92 ;
      RECT 22.505 1.792 22.82 2.065 ;
      RECT 22.525 1.782 22.81 2.091 ;
      RECT 22.11 3.107 22.28 3.395 ;
      RECT 22.105 3.125 22.29 3.39 ;
      RECT 22.07 3.133 22.355 3.31 ;
      RECT 22.07 3.133 22.441 3.3 ;
      RECT 22.07 3.133 22.495 3.246 ;
      RECT 22.355 3.03 22.525 3.214 ;
      RECT 22.07 3.185 22.53 3.202 ;
      RECT 22.055 3.155 22.525 3.198 ;
      RECT 22.315 3.037 22.355 3.349 ;
      RECT 22.195 3.074 22.525 3.214 ;
      RECT 22.29 3.049 22.315 3.375 ;
      RECT 22.28 3.056 22.525 3.214 ;
      RECT 22.411 2.52 22.48 2.779 ;
      RECT 22.411 2.575 22.485 2.778 ;
      RECT 22.325 2.575 22.485 2.777 ;
      RECT 22.32 2.575 22.49 2.77 ;
      RECT 22.31 2.52 22.48 2.765 ;
      RECT 21.69 1.819 21.865 2.12 ;
      RECT 21.675 1.807 21.69 2.105 ;
      RECT 21.645 1.806 21.675 2.058 ;
      RECT 21.645 1.824 21.87 2.053 ;
      RECT 21.63 1.808 21.69 2.018 ;
      RECT 21.625 1.83 21.88 1.918 ;
      RECT 21.625 1.813 21.776 1.918 ;
      RECT 21.625 1.815 21.78 1.918 ;
      RECT 21.63 1.811 21.776 2.018 ;
      RECT 21.735 3.047 21.74 3.395 ;
      RECT 21.725 3.037 21.735 3.401 ;
      RECT 21.69 3.027 21.725 3.403 ;
      RECT 21.652 3.022 21.69 3.407 ;
      RECT 21.566 3.015 21.652 3.414 ;
      RECT 21.48 3.005 21.566 3.424 ;
      RECT 21.435 3 21.48 3.432 ;
      RECT 21.431 3 21.435 3.436 ;
      RECT 21.345 3 21.431 3.443 ;
      RECT 21.33 3 21.345 3.443 ;
      RECT 21.32 2.998 21.33 3.415 ;
      RECT 21.31 2.994 21.32 3.358 ;
      RECT 21.29 2.988 21.31 3.29 ;
      RECT 21.285 2.984 21.29 3.238 ;
      RECT 21.275 2.983 21.285 3.205 ;
      RECT 21.225 2.981 21.275 3.19 ;
      RECT 21.2 2.979 21.225 3.185 ;
      RECT 21.157 2.977 21.2 3.181 ;
      RECT 21.071 2.973 21.157 3.169 ;
      RECT 20.985 2.968 21.071 3.153 ;
      RECT 20.955 2.965 20.985 3.14 ;
      RECT 20.93 2.964 20.955 3.128 ;
      RECT 20.925 2.964 20.93 3.118 ;
      RECT 20.885 2.963 20.925 3.11 ;
      RECT 20.87 2.962 20.885 3.103 ;
      RECT 20.82 2.961 20.87 3.095 ;
      RECT 20.818 2.96 20.82 3.09 ;
      RECT 20.732 2.958 20.818 3.09 ;
      RECT 20.646 2.953 20.732 3.09 ;
      RECT 20.56 2.949 20.646 3.09 ;
      RECT 20.511 2.945 20.56 3.088 ;
      RECT 20.425 2.942 20.511 3.083 ;
      RECT 20.402 2.939 20.425 3.079 ;
      RECT 20.316 2.936 20.402 3.074 ;
      RECT 20.23 2.932 20.316 3.065 ;
      RECT 20.205 2.925 20.23 3.06 ;
      RECT 20.145 2.89 20.205 3.057 ;
      RECT 20.125 2.815 20.145 3.054 ;
      RECT 20.12 2.757 20.125 3.053 ;
      RECT 20.095 2.697 20.12 3.052 ;
      RECT 20.02 2.575 20.095 3.048 ;
      RECT 20.01 2.575 20.02 3.04 ;
      RECT 19.995 2.575 20.01 3.03 ;
      RECT 19.98 2.575 19.995 3 ;
      RECT 19.965 2.575 19.98 2.945 ;
      RECT 19.95 2.575 19.965 2.883 ;
      RECT 19.925 2.575 19.95 2.808 ;
      RECT 19.92 2.575 19.925 2.758 ;
      RECT 21.265 2.12 21.285 2.429 ;
      RECT 21.251 2.122 21.3 2.426 ;
      RECT 21.251 2.127 21.32 2.417 ;
      RECT 21.165 2.125 21.3 2.411 ;
      RECT 21.165 2.133 21.355 2.394 ;
      RECT 21.13 2.135 21.355 2.393 ;
      RECT 21.1 2.143 21.355 2.384 ;
      RECT 21.09 2.148 21.375 2.37 ;
      RECT 21.13 2.138 21.375 2.37 ;
      RECT 21.13 2.141 21.385 2.358 ;
      RECT 21.1 2.143 21.395 2.345 ;
      RECT 21.1 2.147 21.405 2.288 ;
      RECT 21.09 2.152 21.41 2.203 ;
      RECT 21.251 2.12 21.285 2.426 ;
      RECT 21.13 7.855 21.3 8.305 ;
      RECT 21.185 6.075 21.355 8.025 ;
      RECT 21.13 5.015 21.3 6.245 ;
      RECT 20.69 2.223 20.695 2.435 ;
      RECT 20.565 2.22 20.58 2.435 ;
      RECT 20.03 2.25 20.1 2.435 ;
      RECT 19.915 2.25 19.95 2.43 ;
      RECT 21.036 2.552 21.055 2.746 ;
      RECT 20.95 2.507 21.036 2.747 ;
      RECT 20.94 2.46 20.95 2.749 ;
      RECT 20.935 2.44 20.94 2.75 ;
      RECT 20.915 2.405 20.935 2.751 ;
      RECT 20.9 2.355 20.915 2.752 ;
      RECT 20.88 2.292 20.9 2.753 ;
      RECT 20.87 2.255 20.88 2.754 ;
      RECT 20.855 2.244 20.87 2.755 ;
      RECT 20.85 2.236 20.855 2.753 ;
      RECT 20.84 2.235 20.85 2.745 ;
      RECT 20.81 2.232 20.84 2.724 ;
      RECT 20.735 2.227 20.81 2.669 ;
      RECT 20.72 2.223 20.735 2.615 ;
      RECT 20.71 2.223 20.72 2.51 ;
      RECT 20.695 2.223 20.71 2.443 ;
      RECT 20.68 2.223 20.69 2.433 ;
      RECT 20.625 2.222 20.68 2.43 ;
      RECT 20.58 2.22 20.625 2.433 ;
      RECT 20.552 2.22 20.565 2.436 ;
      RECT 20.466 2.224 20.552 2.438 ;
      RECT 20.38 2.23 20.466 2.443 ;
      RECT 20.36 2.234 20.38 2.445 ;
      RECT 20.358 2.235 20.36 2.444 ;
      RECT 20.272 2.237 20.358 2.443 ;
      RECT 20.186 2.242 20.272 2.44 ;
      RECT 20.1 2.247 20.186 2.437 ;
      RECT 19.95 2.25 20.03 2.433 ;
      RECT 20.61 5.015 20.78 8.305 ;
      RECT 20.61 7.315 21.015 7.645 ;
      RECT 20.61 6.475 21.015 6.805 ;
      RECT 20.726 3.225 20.775 3.559 ;
      RECT 20.726 3.225 20.78 3.558 ;
      RECT 20.64 3.225 20.78 3.557 ;
      RECT 20.415 3.333 20.785 3.555 ;
      RECT 20.64 3.225 20.81 3.548 ;
      RECT 20.61 3.237 20.815 3.539 ;
      RECT 20.595 3.255 20.82 3.536 ;
      RECT 20.41 3.339 20.82 3.463 ;
      RECT 20.405 3.346 20.82 3.423 ;
      RECT 20.42 3.312 20.82 3.536 ;
      RECT 20.581 3.258 20.785 3.555 ;
      RECT 20.495 3.278 20.82 3.536 ;
      RECT 20.595 3.252 20.815 3.539 ;
      RECT 20.365 2.576 20.555 2.77 ;
      RECT 20.36 2.578 20.555 2.769 ;
      RECT 20.355 2.582 20.57 2.766 ;
      RECT 20.37 2.575 20.57 2.766 ;
      RECT 20.355 2.685 20.575 2.761 ;
      RECT 19.65 3.185 19.741 3.483 ;
      RECT 19.645 3.187 19.82 3.478 ;
      RECT 19.65 3.185 19.82 3.478 ;
      RECT 19.645 3.191 19.84 3.476 ;
      RECT 19.645 3.246 19.88 3.475 ;
      RECT 19.645 3.281 19.895 3.469 ;
      RECT 19.645 3.315 19.905 3.459 ;
      RECT 19.635 3.195 19.84 3.31 ;
      RECT 19.635 3.215 19.855 3.31 ;
      RECT 19.635 3.198 19.845 3.31 ;
      RECT 19.86 1.966 19.865 2.028 ;
      RECT 19.855 1.888 19.86 2.051 ;
      RECT 19.85 1.845 19.855 2.062 ;
      RECT 19.845 1.835 19.85 2.074 ;
      RECT 19.84 1.835 19.845 2.083 ;
      RECT 19.815 1.835 19.84 2.115 ;
      RECT 19.81 1.835 19.815 2.148 ;
      RECT 19.795 1.835 19.81 2.173 ;
      RECT 19.785 1.835 19.795 2.2 ;
      RECT 19.78 1.835 19.785 2.213 ;
      RECT 19.775 1.835 19.78 2.228 ;
      RECT 19.765 1.835 19.775 2.243 ;
      RECT 19.76 1.835 19.765 2.263 ;
      RECT 19.735 1.835 19.76 2.298 ;
      RECT 19.69 1.835 19.735 2.343 ;
      RECT 19.68 1.835 19.69 2.356 ;
      RECT 19.595 1.92 19.68 2.363 ;
      RECT 19.56 2.042 19.595 2.372 ;
      RECT 19.555 2.082 19.56 2.376 ;
      RECT 19.535 2.105 19.555 2.378 ;
      RECT 19.53 2.135 19.535 2.381 ;
      RECT 19.52 2.147 19.53 2.382 ;
      RECT 19.475 2.17 19.52 2.387 ;
      RECT 19.435 2.2 19.475 2.395 ;
      RECT 19.4 2.212 19.435 2.401 ;
      RECT 19.395 2.217 19.4 2.405 ;
      RECT 19.325 2.227 19.395 2.412 ;
      RECT 19.285 2.237 19.325 2.422 ;
      RECT 19.265 2.242 19.285 2.428 ;
      RECT 19.255 2.246 19.265 2.433 ;
      RECT 19.25 2.249 19.255 2.436 ;
      RECT 19.24 2.25 19.25 2.437 ;
      RECT 19.215 2.252 19.24 2.441 ;
      RECT 19.205 2.257 19.215 2.444 ;
      RECT 19.16 2.265 19.205 2.445 ;
      RECT 19.035 2.27 19.16 2.445 ;
      RECT 19.59 2.567 19.61 2.749 ;
      RECT 19.541 2.552 19.59 2.748 ;
      RECT 19.455 2.567 19.61 2.746 ;
      RECT 19.44 2.567 19.61 2.745 ;
      RECT 19.405 2.545 19.575 2.73 ;
      RECT 19.475 3.565 19.49 3.774 ;
      RECT 19.475 3.573 19.495 3.773 ;
      RECT 19.42 3.573 19.495 3.772 ;
      RECT 19.4 3.577 19.5 3.77 ;
      RECT 19.38 3.527 19.42 3.769 ;
      RECT 19.325 3.585 19.505 3.767 ;
      RECT 19.29 3.542 19.42 3.765 ;
      RECT 19.286 3.545 19.475 3.764 ;
      RECT 19.2 3.553 19.475 3.762 ;
      RECT 19.2 3.597 19.51 3.755 ;
      RECT 19.19 3.69 19.51 3.753 ;
      RECT 19.2 3.609 19.515 3.738 ;
      RECT 19.2 3.63 19.53 3.708 ;
      RECT 19.2 3.657 19.535 3.678 ;
      RECT 19.325 3.535 19.42 3.767 ;
      RECT 18.955 2.58 18.96 3.118 ;
      RECT 18.76 2.91 18.765 3.105 ;
      RECT 17.06 2.575 17.075 2.955 ;
      RECT 19.125 2.575 19.13 2.745 ;
      RECT 19.12 2.575 19.125 2.755 ;
      RECT 19.115 2.575 19.12 2.768 ;
      RECT 19.09 2.575 19.115 2.81 ;
      RECT 19.065 2.575 19.09 2.883 ;
      RECT 19.05 2.575 19.065 2.935 ;
      RECT 19.045 2.575 19.05 2.965 ;
      RECT 19.02 2.575 19.045 3.005 ;
      RECT 19.005 2.575 19.02 3.06 ;
      RECT 19 2.575 19.005 3.093 ;
      RECT 18.975 2.575 19 3.113 ;
      RECT 18.96 2.575 18.975 3.119 ;
      RECT 18.89 2.61 18.955 3.115 ;
      RECT 18.84 2.665 18.89 3.11 ;
      RECT 18.83 2.697 18.84 3.108 ;
      RECT 18.825 2.722 18.83 3.108 ;
      RECT 18.805 2.795 18.825 3.108 ;
      RECT 18.795 2.875 18.805 3.107 ;
      RECT 18.78 2.905 18.795 3.107 ;
      RECT 18.765 2.91 18.78 3.106 ;
      RECT 18.705 2.912 18.76 3.103 ;
      RECT 18.675 2.917 18.705 3.099 ;
      RECT 18.673 2.92 18.675 3.098 ;
      RECT 18.587 2.922 18.673 3.095 ;
      RECT 18.501 2.928 18.587 3.089 ;
      RECT 18.415 2.933 18.501 3.083 ;
      RECT 18.342 2.938 18.415 3.084 ;
      RECT 18.256 2.944 18.342 3.092 ;
      RECT 18.17 2.95 18.256 3.101 ;
      RECT 18.15 2.954 18.17 3.106 ;
      RECT 18.103 2.956 18.15 3.109 ;
      RECT 18.017 2.961 18.103 3.115 ;
      RECT 17.931 2.966 18.017 3.124 ;
      RECT 17.845 2.972 17.931 3.132 ;
      RECT 17.76 2.97 17.845 3.141 ;
      RECT 17.756 2.965 17.76 3.145 ;
      RECT 17.67 2.96 17.756 3.137 ;
      RECT 17.606 2.951 17.67 3.125 ;
      RECT 17.52 2.942 17.606 3.112 ;
      RECT 17.496 2.935 17.52 3.103 ;
      RECT 17.41 2.929 17.496 3.09 ;
      RECT 17.37 2.922 17.41 3.076 ;
      RECT 17.365 2.912 17.37 3.072 ;
      RECT 17.355 2.9 17.365 3.071 ;
      RECT 17.335 2.87 17.355 3.068 ;
      RECT 17.28 2.79 17.335 3.062 ;
      RECT 17.26 2.709 17.28 3.057 ;
      RECT 17.24 2.667 17.26 3.053 ;
      RECT 17.215 2.62 17.24 3.047 ;
      RECT 17.21 2.595 17.215 3.044 ;
      RECT 17.175 2.575 17.21 3.039 ;
      RECT 17.166 2.575 17.175 3.032 ;
      RECT 17.08 2.575 17.166 3.002 ;
      RECT 17.075 2.575 17.08 2.965 ;
      RECT 17.04 2.575 17.06 2.887 ;
      RECT 17.035 2.617 17.04 2.852 ;
      RECT 17.03 2.692 17.035 2.808 ;
      RECT 18.48 2.497 18.655 2.745 ;
      RECT 18.48 2.497 18.66 2.743 ;
      RECT 18.475 2.529 18.66 2.703 ;
      RECT 18.505 2.47 18.675 2.69 ;
      RECT 18.47 2.547 18.675 2.623 ;
      RECT 17.78 2.01 17.95 2.185 ;
      RECT 17.78 2.01 18.122 2.177 ;
      RECT 17.78 2.01 18.205 2.171 ;
      RECT 17.78 2.01 18.24 2.167 ;
      RECT 17.78 2.01 18.26 2.166 ;
      RECT 17.78 2.01 18.346 2.162 ;
      RECT 18.24 1.835 18.41 2.157 ;
      RECT 17.815 1.942 18.44 2.155 ;
      RECT 17.805 1.997 18.445 2.153 ;
      RECT 17.78 2.033 18.455 2.148 ;
      RECT 17.78 2.06 18.46 2.078 ;
      RECT 17.845 1.885 18.42 2.155 ;
      RECT 18.036 1.87 18.42 2.155 ;
      RECT 17.87 1.873 18.42 2.155 ;
      RECT 17.95 1.871 18.036 2.182 ;
      RECT 18.036 1.868 18.415 2.155 ;
      RECT 18.22 1.845 18.415 2.155 ;
      RECT 18.122 1.866 18.415 2.155 ;
      RECT 18.205 1.86 18.22 2.168 ;
      RECT 18.355 3.225 18.36 3.425 ;
      RECT 17.82 3.29 17.865 3.425 ;
      RECT 18.39 3.225 18.41 3.398 ;
      RECT 18.36 3.225 18.39 3.413 ;
      RECT 18.295 3.225 18.355 3.45 ;
      RECT 18.28 3.225 18.295 3.48 ;
      RECT 18.265 3.225 18.28 3.493 ;
      RECT 18.245 3.225 18.265 3.508 ;
      RECT 18.24 3.225 18.245 3.517 ;
      RECT 18.23 3.229 18.24 3.522 ;
      RECT 18.215 3.239 18.23 3.533 ;
      RECT 18.19 3.255 18.215 3.543 ;
      RECT 18.18 3.269 18.19 3.545 ;
      RECT 18.16 3.281 18.18 3.542 ;
      RECT 18.13 3.302 18.16 3.536 ;
      RECT 18.12 3.314 18.13 3.531 ;
      RECT 18.11 3.312 18.12 3.528 ;
      RECT 18.095 3.311 18.11 3.523 ;
      RECT 18.09 3.31 18.095 3.518 ;
      RECT 18.055 3.308 18.09 3.508 ;
      RECT 18.035 3.305 18.055 3.49 ;
      RECT 18.025 3.303 18.035 3.485 ;
      RECT 18.015 3.302 18.025 3.48 ;
      RECT 17.98 3.3 18.015 3.468 ;
      RECT 17.925 3.296 17.98 3.448 ;
      RECT 17.915 3.294 17.925 3.433 ;
      RECT 17.91 3.294 17.915 3.428 ;
      RECT 17.865 3.292 17.91 3.425 ;
      RECT 17.77 3.29 17.82 3.429 ;
      RECT 17.76 3.291 17.77 3.434 ;
      RECT 17.7 3.298 17.76 3.448 ;
      RECT 17.675 3.306 17.7 3.468 ;
      RECT 17.665 3.31 17.675 3.48 ;
      RECT 17.66 3.311 17.665 3.485 ;
      RECT 17.645 3.313 17.66 3.488 ;
      RECT 17.63 3.315 17.645 3.493 ;
      RECT 17.625 3.315 17.63 3.496 ;
      RECT 17.58 3.32 17.625 3.507 ;
      RECT 17.575 3.324 17.58 3.519 ;
      RECT 17.55 3.32 17.575 3.523 ;
      RECT 17.54 3.316 17.55 3.527 ;
      RECT 17.53 3.315 17.54 3.531 ;
      RECT 17.515 3.305 17.53 3.537 ;
      RECT 17.51 3.293 17.515 3.541 ;
      RECT 17.505 3.29 17.51 3.542 ;
      RECT 17.5 3.287 17.505 3.544 ;
      RECT 17.485 3.275 17.5 3.543 ;
      RECT 17.47 3.257 17.485 3.54 ;
      RECT 17.45 3.236 17.47 3.533 ;
      RECT 17.385 3.225 17.45 3.505 ;
      RECT 17.381 3.225 17.385 3.484 ;
      RECT 17.295 3.225 17.381 3.454 ;
      RECT 17.28 3.225 17.295 3.41 ;
      RECT 17.855 2.325 17.86 2.56 ;
      RECT 16.985 2.241 16.99 2.445 ;
      RECT 17.565 2.27 17.57 2.425 ;
      RECT 17.485 2.25 17.49 2.425 ;
      RECT 18.155 2.392 18.17 2.745 ;
      RECT 18.081 2.377 18.155 2.745 ;
      RECT 17.995 2.36 18.081 2.745 ;
      RECT 17.985 2.35 17.995 2.743 ;
      RECT 17.98 2.348 17.985 2.738 ;
      RECT 17.965 2.346 17.98 2.724 ;
      RECT 17.895 2.338 17.965 2.664 ;
      RECT 17.875 2.329 17.895 2.598 ;
      RECT 17.87 2.326 17.875 2.578 ;
      RECT 17.86 2.325 17.87 2.568 ;
      RECT 17.85 2.325 17.855 2.552 ;
      RECT 17.84 2.324 17.85 2.542 ;
      RECT 17.83 2.322 17.84 2.53 ;
      RECT 17.815 2.319 17.83 2.51 ;
      RECT 17.805 2.317 17.815 2.495 ;
      RECT 17.785 2.314 17.805 2.483 ;
      RECT 17.78 2.312 17.785 2.473 ;
      RECT 17.755 2.31 17.78 2.46 ;
      RECT 17.725 2.305 17.755 2.445 ;
      RECT 17.645 2.296 17.725 2.436 ;
      RECT 17.6 2.285 17.645 2.429 ;
      RECT 17.58 2.276 17.6 2.426 ;
      RECT 17.57 2.271 17.58 2.425 ;
      RECT 17.525 2.265 17.565 2.425 ;
      RECT 17.51 2.257 17.525 2.425 ;
      RECT 17.49 2.252 17.51 2.425 ;
      RECT 17.47 2.249 17.485 2.425 ;
      RECT 17.387 2.248 17.47 2.424 ;
      RECT 17.301 2.247 17.387 2.42 ;
      RECT 17.215 2.245 17.301 2.417 ;
      RECT 17.162 2.244 17.215 2.419 ;
      RECT 17.076 2.243 17.162 2.428 ;
      RECT 16.99 2.242 17.076 2.44 ;
      RECT 16.97 2.241 16.985 2.448 ;
      RECT 16.89 2.24 16.97 2.46 ;
      RECT 16.865 2.24 16.89 2.473 ;
      RECT 16.84 2.24 16.865 2.488 ;
      RECT 16.835 2.24 16.84 2.51 ;
      RECT 16.83 2.24 16.835 2.528 ;
      RECT 16.825 2.24 16.83 2.545 ;
      RECT 16.82 2.24 16.825 2.558 ;
      RECT 16.815 2.24 16.82 2.568 ;
      RECT 16.775 2.24 16.815 2.653 ;
      RECT 16.76 2.24 16.775 2.738 ;
      RECT 16.75 2.241 16.76 2.75 ;
      RECT 16.715 2.246 16.75 2.755 ;
      RECT 16.675 2.255 16.715 2.755 ;
      RECT 16.66 2.265 16.675 2.755 ;
      RECT 16.655 2.275 16.66 2.755 ;
      RECT 16.635 2.302 16.655 2.755 ;
      RECT 16.585 2.385 16.635 2.755 ;
      RECT 16.58 2.447 16.585 2.755 ;
      RECT 16.57 2.46 16.58 2.755 ;
      RECT 16.56 2.482 16.57 2.755 ;
      RECT 16.55 2.507 16.56 2.75 ;
      RECT 16.545 2.545 16.55 2.743 ;
      RECT 16.535 2.655 16.545 2.738 ;
      RECT 17.93 3.576 17.945 3.835 ;
      RECT 17.93 3.591 17.95 3.834 ;
      RECT 17.846 3.591 17.95 3.832 ;
      RECT 17.846 3.605 17.955 3.831 ;
      RECT 17.76 3.647 17.96 3.828 ;
      RECT 17.755 3.59 17.945 3.823 ;
      RECT 17.755 3.661 17.965 3.82 ;
      RECT 17.75 3.692 17.965 3.818 ;
      RECT 17.755 3.689 17.98 3.808 ;
      RECT 17.75 3.735 17.995 3.793 ;
      RECT 17.75 3.763 18 3.778 ;
      RECT 17.76 3.565 17.93 3.828 ;
      RECT 17.52 2.575 17.69 2.745 ;
      RECT 17.485 2.575 17.69 2.74 ;
      RECT 17.475 2.575 17.69 2.733 ;
      RECT 17.47 2.56 17.64 2.73 ;
      RECT 16.3 3.097 16.565 3.54 ;
      RECT 16.295 3.068 16.51 3.538 ;
      RECT 16.29 3.222 16.57 3.533 ;
      RECT 16.295 3.117 16.57 3.533 ;
      RECT 16.295 3.128 16.58 3.52 ;
      RECT 16.295 3.075 16.54 3.538 ;
      RECT 16.3 3.062 16.51 3.54 ;
      RECT 16.3 3.06 16.46 3.54 ;
      RECT 16.401 3.052 16.46 3.54 ;
      RECT 16.315 3.053 16.46 3.54 ;
      RECT 16.401 3.051 16.45 3.54 ;
      RECT 16.205 1.866 16.38 2.165 ;
      RECT 16.255 1.828 16.38 2.165 ;
      RECT 16.24 1.83 16.466 2.157 ;
      RECT 16.24 1.833 16.505 2.144 ;
      RECT 16.24 1.834 16.515 2.13 ;
      RECT 16.195 1.885 16.515 2.12 ;
      RECT 16.24 1.835 16.52 2.115 ;
      RECT 16.195 2.045 16.525 2.105 ;
      RECT 16.18 1.905 16.52 2.045 ;
      RECT 16.175 1.921 16.52 1.985 ;
      RECT 16.22 1.845 16.52 2.115 ;
      RECT 16.255 1.826 16.341 2.165 ;
      RECT 14.35 1.74 14.52 2.935 ;
      RECT 14.35 1.74 14.815 1.91 ;
      RECT 14.35 6.97 14.815 7.14 ;
      RECT 14.35 5.945 14.52 7.14 ;
      RECT 13.36 1.74 13.53 2.935 ;
      RECT 13.36 1.74 13.825 1.91 ;
      RECT 13.36 6.97 13.825 7.14 ;
      RECT 13.36 5.945 13.53 7.14 ;
      RECT 11.505 2.635 11.675 3.865 ;
      RECT 11.56 0.855 11.73 2.805 ;
      RECT 11.505 0.575 11.675 1.025 ;
      RECT 11.505 7.855 11.675 8.305 ;
      RECT 11.56 6.075 11.73 8.025 ;
      RECT 11.505 5.015 11.675 6.245 ;
      RECT 10.985 0.575 11.155 3.865 ;
      RECT 10.985 2.075 11.39 2.405 ;
      RECT 10.985 1.235 11.39 1.565 ;
      RECT 10.985 5.015 11.155 8.305 ;
      RECT 10.985 7.315 11.39 7.645 ;
      RECT 10.985 6.475 11.39 6.805 ;
      RECT 8.91 3.126 8.915 3.298 ;
      RECT 8.905 3.119 8.91 3.388 ;
      RECT 8.9 3.113 8.905 3.407 ;
      RECT 8.88 3.107 8.9 3.417 ;
      RECT 8.865 3.102 8.88 3.425 ;
      RECT 8.828 3.096 8.865 3.423 ;
      RECT 8.742 3.082 8.828 3.419 ;
      RECT 8.656 3.064 8.742 3.414 ;
      RECT 8.57 3.045 8.656 3.408 ;
      RECT 8.54 3.033 8.57 3.404 ;
      RECT 8.52 3.027 8.54 3.403 ;
      RECT 8.455 3.025 8.52 3.401 ;
      RECT 8.44 3.025 8.455 3.393 ;
      RECT 8.425 3.025 8.44 3.38 ;
      RECT 8.42 3.025 8.425 3.37 ;
      RECT 8.405 3.025 8.42 3.348 ;
      RECT 8.39 3.025 8.405 3.315 ;
      RECT 8.385 3.025 8.39 3.293 ;
      RECT 8.375 3.025 8.385 3.275 ;
      RECT 8.36 3.025 8.375 3.253 ;
      RECT 8.34 3.025 8.36 3.215 ;
      RECT 8.69 2.31 8.725 2.749 ;
      RECT 8.69 2.31 8.73 2.748 ;
      RECT 8.635 2.37 8.73 2.747 ;
      RECT 8.5 2.542 8.73 2.746 ;
      RECT 8.61 2.42 8.73 2.746 ;
      RECT 8.5 2.542 8.755 2.736 ;
      RECT 8.555 2.487 8.835 2.653 ;
      RECT 8.73 2.281 8.735 2.744 ;
      RECT 8.585 2.457 8.875 2.53 ;
      RECT 8.6 2.44 8.73 2.746 ;
      RECT 8.735 2.28 8.905 2.468 ;
      RECT 8.725 2.283 8.905 2.468 ;
      RECT 8.23 2.16 8.4 2.47 ;
      RECT 8.23 2.16 8.405 2.443 ;
      RECT 8.23 2.16 8.41 2.42 ;
      RECT 8.23 2.16 8.42 2.37 ;
      RECT 8.225 2.265 8.42 2.34 ;
      RECT 8.26 1.835 8.43 2.313 ;
      RECT 8.26 1.835 8.445 2.234 ;
      RECT 8.25 2.045 8.445 2.234 ;
      RECT 8.26 1.845 8.455 2.149 ;
      RECT 8.19 2.587 8.195 2.79 ;
      RECT 8.18 2.575 8.19 2.9 ;
      RECT 8.155 2.575 8.18 2.94 ;
      RECT 8.075 2.575 8.155 3.025 ;
      RECT 8.065 2.575 8.075 3.095 ;
      RECT 8.04 2.575 8.065 3.118 ;
      RECT 8.02 2.575 8.04 3.153 ;
      RECT 7.975 2.585 8.02 3.196 ;
      RECT 7.965 2.597 7.975 3.233 ;
      RECT 7.945 2.611 7.965 3.253 ;
      RECT 7.935 2.629 7.945 3.269 ;
      RECT 7.92 2.655 7.935 3.279 ;
      RECT 7.905 2.696 7.92 3.293 ;
      RECT 7.895 2.731 7.905 3.303 ;
      RECT 7.89 2.747 7.895 3.308 ;
      RECT 7.88 2.762 7.89 3.313 ;
      RECT 7.86 2.805 7.88 3.323 ;
      RECT 7.84 2.842 7.86 3.336 ;
      RECT 7.805 2.865 7.84 3.354 ;
      RECT 7.795 2.879 7.805 3.37 ;
      RECT 7.775 2.889 7.795 3.38 ;
      RECT 7.77 2.898 7.775 3.388 ;
      RECT 7.76 2.905 7.77 3.395 ;
      RECT 7.75 2.912 7.76 3.403 ;
      RECT 7.735 2.922 7.75 3.411 ;
      RECT 7.725 2.936 7.735 3.421 ;
      RECT 7.715 2.948 7.725 3.433 ;
      RECT 7.7 2.97 7.715 3.446 ;
      RECT 7.69 2.992 7.7 3.457 ;
      RECT 7.68 3.012 7.69 3.466 ;
      RECT 7.675 3.027 7.68 3.473 ;
      RECT 7.645 3.06 7.675 3.487 ;
      RECT 7.635 3.095 7.645 3.502 ;
      RECT 7.63 3.102 7.635 3.508 ;
      RECT 7.61 3.117 7.63 3.515 ;
      RECT 7.605 3.132 7.61 3.523 ;
      RECT 7.6 3.141 7.605 3.528 ;
      RECT 7.585 3.147 7.6 3.535 ;
      RECT 7.58 3.153 7.585 3.543 ;
      RECT 7.575 3.157 7.58 3.55 ;
      RECT 7.57 3.161 7.575 3.56 ;
      RECT 7.56 3.166 7.57 3.57 ;
      RECT 7.54 3.177 7.56 3.598 ;
      RECT 7.525 3.189 7.54 3.625 ;
      RECT 7.505 3.202 7.525 3.65 ;
      RECT 7.485 3.217 7.505 3.674 ;
      RECT 7.47 3.232 7.485 3.689 ;
      RECT 7.465 3.243 7.47 3.698 ;
      RECT 7.4 3.288 7.465 3.708 ;
      RECT 7.365 3.347 7.4 3.721 ;
      RECT 7.36 3.37 7.365 3.727 ;
      RECT 7.355 3.377 7.36 3.729 ;
      RECT 7.34 3.387 7.355 3.732 ;
      RECT 7.31 3.412 7.34 3.736 ;
      RECT 7.305 3.43 7.31 3.74 ;
      RECT 7.3 3.437 7.305 3.741 ;
      RECT 7.28 3.445 7.3 3.745 ;
      RECT 7.27 3.452 7.28 3.749 ;
      RECT 7.226 3.463 7.27 3.756 ;
      RECT 7.14 3.491 7.226 3.772 ;
      RECT 7.08 3.515 7.14 3.79 ;
      RECT 7.035 3.525 7.08 3.804 ;
      RECT 6.976 3.533 7.035 3.818 ;
      RECT 6.89 3.54 6.976 3.837 ;
      RECT 6.865 3.545 6.89 3.852 ;
      RECT 6.785 3.548 6.865 3.855 ;
      RECT 6.705 3.552 6.785 3.842 ;
      RECT 6.696 3.555 6.705 3.827 ;
      RECT 6.61 3.555 6.696 3.812 ;
      RECT 6.55 3.557 6.61 3.789 ;
      RECT 6.546 3.56 6.55 3.779 ;
      RECT 6.46 3.56 6.546 3.764 ;
      RECT 6.385 3.56 6.46 3.74 ;
      RECT 7.7 2.569 7.71 2.745 ;
      RECT 7.655 2.536 7.7 2.745 ;
      RECT 7.61 2.487 7.655 2.745 ;
      RECT 7.58 2.457 7.61 2.746 ;
      RECT 7.575 2.44 7.58 2.747 ;
      RECT 7.55 2.42 7.575 2.748 ;
      RECT 7.535 2.395 7.55 2.749 ;
      RECT 7.53 2.382 7.535 2.75 ;
      RECT 7.525 2.376 7.53 2.748 ;
      RECT 7.52 2.368 7.525 2.742 ;
      RECT 7.495 2.36 7.52 2.722 ;
      RECT 7.475 2.349 7.495 2.693 ;
      RECT 7.445 2.334 7.475 2.664 ;
      RECT 7.425 2.32 7.445 2.636 ;
      RECT 7.415 2.314 7.425 2.615 ;
      RECT 7.41 2.311 7.415 2.598 ;
      RECT 7.405 2.308 7.41 2.583 ;
      RECT 7.39 2.303 7.405 2.548 ;
      RECT 7.385 2.299 7.39 2.515 ;
      RECT 7.365 2.294 7.385 2.491 ;
      RECT 7.335 2.286 7.365 2.456 ;
      RECT 7.32 2.28 7.335 2.433 ;
      RECT 7.28 2.273 7.32 2.418 ;
      RECT 7.255 2.265 7.28 2.398 ;
      RECT 7.235 2.26 7.255 2.388 ;
      RECT 7.2 2.254 7.235 2.383 ;
      RECT 7.155 2.245 7.2 2.382 ;
      RECT 7.125 2.241 7.155 2.384 ;
      RECT 7.04 2.249 7.125 2.388 ;
      RECT 6.97 2.26 7.04 2.41 ;
      RECT 6.957 2.266 6.97 2.433 ;
      RECT 6.871 2.273 6.957 2.455 ;
      RECT 6.785 2.285 6.871 2.492 ;
      RECT 6.785 2.662 6.795 2.9 ;
      RECT 6.78 2.291 6.785 2.515 ;
      RECT 6.775 2.547 6.785 2.9 ;
      RECT 6.775 2.292 6.78 2.52 ;
      RECT 6.77 2.293 6.775 2.9 ;
      RECT 6.746 2.295 6.77 2.901 ;
      RECT 6.66 2.303 6.746 2.903 ;
      RECT 6.64 2.317 6.66 2.906 ;
      RECT 6.635 2.345 6.64 2.907 ;
      RECT 6.63 2.357 6.635 2.908 ;
      RECT 6.625 2.372 6.63 2.909 ;
      RECT 6.615 2.402 6.625 2.91 ;
      RECT 6.61 2.44 6.615 2.908 ;
      RECT 6.605 2.46 6.61 2.903 ;
      RECT 6.59 2.495 6.605 2.888 ;
      RECT 6.58 2.547 6.59 2.868 ;
      RECT 6.575 2.577 6.58 2.856 ;
      RECT 6.56 2.59 6.575 2.839 ;
      RECT 6.535 2.594 6.56 2.806 ;
      RECT 6.52 2.592 6.535 2.783 ;
      RECT 6.505 2.591 6.52 2.78 ;
      RECT 6.445 2.589 6.505 2.778 ;
      RECT 6.435 2.587 6.445 2.773 ;
      RECT 6.395 2.586 6.435 2.77 ;
      RECT 6.325 2.583 6.395 2.768 ;
      RECT 6.27 2.581 6.325 2.763 ;
      RECT 6.2 2.575 6.27 2.758 ;
      RECT 6.191 2.575 6.2 2.755 ;
      RECT 6.105 2.575 6.191 2.75 ;
      RECT 6.1 2.575 6.105 2.745 ;
      RECT 7.405 1.81 7.58 2.16 ;
      RECT 7.405 1.825 7.59 2.158 ;
      RECT 7.38 1.775 7.525 2.155 ;
      RECT 7.36 1.776 7.525 2.148 ;
      RECT 7.35 1.777 7.535 2.143 ;
      RECT 7.32 1.778 7.535 2.13 ;
      RECT 7.27 1.779 7.535 2.106 ;
      RECT 7.265 1.781 7.535 2.091 ;
      RECT 7.265 1.847 7.595 2.085 ;
      RECT 7.245 1.788 7.55 2.065 ;
      RECT 7.235 1.797 7.56 1.92 ;
      RECT 7.245 1.792 7.56 2.065 ;
      RECT 7.265 1.782 7.55 2.091 ;
      RECT 6.85 3.107 7.02 3.395 ;
      RECT 6.845 3.125 7.03 3.39 ;
      RECT 6.81 3.133 7.095 3.31 ;
      RECT 6.81 3.133 7.181 3.3 ;
      RECT 6.81 3.133 7.235 3.246 ;
      RECT 7.095 3.03 7.265 3.214 ;
      RECT 6.81 3.185 7.27 3.202 ;
      RECT 6.795 3.155 7.265 3.198 ;
      RECT 7.055 3.037 7.095 3.349 ;
      RECT 6.935 3.074 7.265 3.214 ;
      RECT 7.03 3.049 7.055 3.375 ;
      RECT 7.02 3.056 7.265 3.214 ;
      RECT 7.151 2.52 7.22 2.779 ;
      RECT 7.151 2.575 7.225 2.778 ;
      RECT 7.065 2.575 7.225 2.777 ;
      RECT 7.06 2.575 7.23 2.77 ;
      RECT 7.05 2.52 7.22 2.765 ;
      RECT 6.43 1.819 6.605 2.12 ;
      RECT 6.415 1.807 6.43 2.105 ;
      RECT 6.385 1.806 6.415 2.058 ;
      RECT 6.385 1.824 6.61 2.053 ;
      RECT 6.37 1.808 6.43 2.018 ;
      RECT 6.365 1.83 6.62 1.918 ;
      RECT 6.365 1.813 6.516 1.918 ;
      RECT 6.365 1.815 6.52 1.918 ;
      RECT 6.37 1.811 6.516 2.018 ;
      RECT 6.475 3.047 6.48 3.395 ;
      RECT 6.465 3.037 6.475 3.401 ;
      RECT 6.43 3.027 6.465 3.403 ;
      RECT 6.392 3.022 6.43 3.407 ;
      RECT 6.306 3.015 6.392 3.414 ;
      RECT 6.22 3.005 6.306 3.424 ;
      RECT 6.175 3 6.22 3.432 ;
      RECT 6.171 3 6.175 3.436 ;
      RECT 6.085 3 6.171 3.443 ;
      RECT 6.07 3 6.085 3.443 ;
      RECT 6.06 2.998 6.07 3.415 ;
      RECT 6.05 2.994 6.06 3.358 ;
      RECT 6.03 2.988 6.05 3.29 ;
      RECT 6.025 2.984 6.03 3.238 ;
      RECT 6.015 2.983 6.025 3.205 ;
      RECT 5.965 2.981 6.015 3.19 ;
      RECT 5.94 2.979 5.965 3.185 ;
      RECT 5.897 2.977 5.94 3.181 ;
      RECT 5.811 2.973 5.897 3.169 ;
      RECT 5.725 2.968 5.811 3.153 ;
      RECT 5.695 2.965 5.725 3.14 ;
      RECT 5.67 2.964 5.695 3.128 ;
      RECT 5.665 2.964 5.67 3.118 ;
      RECT 5.625 2.963 5.665 3.11 ;
      RECT 5.61 2.962 5.625 3.103 ;
      RECT 5.56 2.961 5.61 3.095 ;
      RECT 5.558 2.96 5.56 3.09 ;
      RECT 5.472 2.958 5.558 3.09 ;
      RECT 5.386 2.953 5.472 3.09 ;
      RECT 5.3 2.949 5.386 3.09 ;
      RECT 5.251 2.945 5.3 3.088 ;
      RECT 5.165 2.942 5.251 3.083 ;
      RECT 5.142 2.939 5.165 3.079 ;
      RECT 5.056 2.936 5.142 3.074 ;
      RECT 4.97 2.932 5.056 3.065 ;
      RECT 4.945 2.925 4.97 3.06 ;
      RECT 4.885 2.89 4.945 3.057 ;
      RECT 4.865 2.815 4.885 3.054 ;
      RECT 4.86 2.757 4.865 3.053 ;
      RECT 4.835 2.697 4.86 3.052 ;
      RECT 4.76 2.575 4.835 3.048 ;
      RECT 4.75 2.575 4.76 3.04 ;
      RECT 4.735 2.575 4.75 3.03 ;
      RECT 4.72 2.575 4.735 3 ;
      RECT 4.705 2.575 4.72 2.945 ;
      RECT 4.69 2.575 4.705 2.883 ;
      RECT 4.665 2.575 4.69 2.808 ;
      RECT 4.66 2.575 4.665 2.758 ;
      RECT 6.005 2.12 6.025 2.429 ;
      RECT 5.991 2.122 6.04 2.426 ;
      RECT 5.991 2.127 6.06 2.417 ;
      RECT 5.905 2.125 6.04 2.411 ;
      RECT 5.905 2.133 6.095 2.394 ;
      RECT 5.87 2.135 6.095 2.393 ;
      RECT 5.84 2.143 6.095 2.384 ;
      RECT 5.83 2.148 6.115 2.37 ;
      RECT 5.87 2.138 6.115 2.37 ;
      RECT 5.87 2.141 6.125 2.358 ;
      RECT 5.84 2.143 6.135 2.345 ;
      RECT 5.84 2.147 6.145 2.288 ;
      RECT 5.83 2.152 6.15 2.203 ;
      RECT 5.991 2.12 6.025 2.426 ;
      RECT 5.87 7.855 6.04 8.305 ;
      RECT 5.925 6.075 6.095 8.025 ;
      RECT 5.87 5.015 6.04 6.245 ;
      RECT 5.43 2.223 5.435 2.435 ;
      RECT 5.305 2.22 5.32 2.435 ;
      RECT 4.77 2.25 4.84 2.435 ;
      RECT 4.655 2.25 4.69 2.43 ;
      RECT 5.776 2.552 5.795 2.746 ;
      RECT 5.69 2.507 5.776 2.747 ;
      RECT 5.68 2.46 5.69 2.749 ;
      RECT 5.675 2.44 5.68 2.75 ;
      RECT 5.655 2.405 5.675 2.751 ;
      RECT 5.64 2.355 5.655 2.752 ;
      RECT 5.62 2.292 5.64 2.753 ;
      RECT 5.61 2.255 5.62 2.754 ;
      RECT 5.595 2.244 5.61 2.755 ;
      RECT 5.59 2.236 5.595 2.753 ;
      RECT 5.58 2.235 5.59 2.745 ;
      RECT 5.55 2.232 5.58 2.724 ;
      RECT 5.475 2.227 5.55 2.669 ;
      RECT 5.46 2.223 5.475 2.615 ;
      RECT 5.45 2.223 5.46 2.51 ;
      RECT 5.435 2.223 5.45 2.443 ;
      RECT 5.42 2.223 5.43 2.433 ;
      RECT 5.365 2.222 5.42 2.43 ;
      RECT 5.32 2.22 5.365 2.433 ;
      RECT 5.292 2.22 5.305 2.436 ;
      RECT 5.206 2.224 5.292 2.438 ;
      RECT 5.12 2.23 5.206 2.443 ;
      RECT 5.1 2.234 5.12 2.445 ;
      RECT 5.098 2.235 5.1 2.444 ;
      RECT 5.012 2.237 5.098 2.443 ;
      RECT 4.926 2.242 5.012 2.44 ;
      RECT 4.84 2.247 4.926 2.437 ;
      RECT 4.69 2.25 4.77 2.433 ;
      RECT 5.35 5.015 5.52 8.305 ;
      RECT 5.35 7.315 5.755 7.645 ;
      RECT 5.35 6.475 5.755 6.805 ;
      RECT 5.466 3.225 5.515 3.559 ;
      RECT 5.466 3.225 5.52 3.558 ;
      RECT 5.38 3.225 5.52 3.557 ;
      RECT 5.155 3.333 5.525 3.555 ;
      RECT 5.38 3.225 5.55 3.548 ;
      RECT 5.35 3.237 5.555 3.539 ;
      RECT 5.335 3.255 5.56 3.536 ;
      RECT 5.15 3.339 5.56 3.463 ;
      RECT 5.145 3.346 5.56 3.423 ;
      RECT 5.16 3.312 5.56 3.536 ;
      RECT 5.321 3.258 5.525 3.555 ;
      RECT 5.235 3.278 5.56 3.536 ;
      RECT 5.335 3.252 5.555 3.539 ;
      RECT 5.105 2.576 5.295 2.77 ;
      RECT 5.1 2.578 5.295 2.769 ;
      RECT 5.095 2.582 5.31 2.766 ;
      RECT 5.11 2.575 5.31 2.766 ;
      RECT 5.095 2.685 5.315 2.761 ;
      RECT 4.39 3.185 4.481 3.483 ;
      RECT 4.385 3.187 4.56 3.478 ;
      RECT 4.39 3.185 4.56 3.478 ;
      RECT 4.385 3.191 4.58 3.476 ;
      RECT 4.385 3.246 4.62 3.475 ;
      RECT 4.385 3.281 4.635 3.469 ;
      RECT 4.385 3.315 4.645 3.459 ;
      RECT 4.375 3.195 4.58 3.31 ;
      RECT 4.375 3.215 4.595 3.31 ;
      RECT 4.375 3.198 4.585 3.31 ;
      RECT 4.6 1.966 4.605 2.028 ;
      RECT 4.595 1.888 4.6 2.051 ;
      RECT 4.59 1.845 4.595 2.062 ;
      RECT 4.585 1.835 4.59 2.074 ;
      RECT 4.58 1.835 4.585 2.083 ;
      RECT 4.555 1.835 4.58 2.115 ;
      RECT 4.55 1.835 4.555 2.148 ;
      RECT 4.535 1.835 4.55 2.173 ;
      RECT 4.525 1.835 4.535 2.2 ;
      RECT 4.52 1.835 4.525 2.213 ;
      RECT 4.515 1.835 4.52 2.228 ;
      RECT 4.505 1.835 4.515 2.243 ;
      RECT 4.5 1.835 4.505 2.263 ;
      RECT 4.475 1.835 4.5 2.298 ;
      RECT 4.43 1.835 4.475 2.343 ;
      RECT 4.42 1.835 4.43 2.356 ;
      RECT 4.335 1.92 4.42 2.363 ;
      RECT 4.3 2.042 4.335 2.372 ;
      RECT 4.295 2.082 4.3 2.376 ;
      RECT 4.275 2.105 4.295 2.378 ;
      RECT 4.27 2.135 4.275 2.381 ;
      RECT 4.26 2.147 4.27 2.382 ;
      RECT 4.215 2.17 4.26 2.387 ;
      RECT 4.175 2.2 4.215 2.395 ;
      RECT 4.14 2.212 4.175 2.401 ;
      RECT 4.135 2.217 4.14 2.405 ;
      RECT 4.065 2.227 4.135 2.412 ;
      RECT 4.025 2.237 4.065 2.422 ;
      RECT 4.005 2.242 4.025 2.428 ;
      RECT 3.995 2.246 4.005 2.433 ;
      RECT 3.99 2.249 3.995 2.436 ;
      RECT 3.98 2.25 3.99 2.437 ;
      RECT 3.955 2.252 3.98 2.441 ;
      RECT 3.945 2.257 3.955 2.444 ;
      RECT 3.9 2.265 3.945 2.445 ;
      RECT 3.775 2.27 3.9 2.445 ;
      RECT 4.33 2.567 4.35 2.749 ;
      RECT 4.281 2.552 4.33 2.748 ;
      RECT 4.195 2.567 4.35 2.746 ;
      RECT 4.18 2.567 4.35 2.745 ;
      RECT 4.145 2.545 4.315 2.73 ;
      RECT 4.215 3.565 4.23 3.774 ;
      RECT 4.215 3.573 4.235 3.773 ;
      RECT 4.16 3.573 4.235 3.772 ;
      RECT 4.14 3.577 4.24 3.77 ;
      RECT 4.12 3.527 4.16 3.769 ;
      RECT 4.065 3.585 4.245 3.767 ;
      RECT 4.03 3.542 4.16 3.765 ;
      RECT 4.026 3.545 4.215 3.764 ;
      RECT 3.94 3.553 4.215 3.762 ;
      RECT 3.94 3.597 4.25 3.755 ;
      RECT 3.93 3.69 4.25 3.753 ;
      RECT 3.94 3.609 4.255 3.738 ;
      RECT 3.94 3.63 4.27 3.708 ;
      RECT 3.94 3.657 4.275 3.678 ;
      RECT 4.065 3.535 4.16 3.767 ;
      RECT 3.695 2.58 3.7 3.118 ;
      RECT 3.5 2.91 3.505 3.105 ;
      RECT 1.8 2.575 1.815 2.955 ;
      RECT 3.865 2.575 3.87 2.745 ;
      RECT 3.86 2.575 3.865 2.755 ;
      RECT 3.855 2.575 3.86 2.768 ;
      RECT 3.83 2.575 3.855 2.81 ;
      RECT 3.805 2.575 3.83 2.883 ;
      RECT 3.79 2.575 3.805 2.935 ;
      RECT 3.785 2.575 3.79 2.965 ;
      RECT 3.76 2.575 3.785 3.005 ;
      RECT 3.745 2.575 3.76 3.06 ;
      RECT 3.74 2.575 3.745 3.093 ;
      RECT 3.715 2.575 3.74 3.113 ;
      RECT 3.7 2.575 3.715 3.119 ;
      RECT 3.63 2.61 3.695 3.115 ;
      RECT 3.58 2.665 3.63 3.11 ;
      RECT 3.57 2.697 3.58 3.108 ;
      RECT 3.565 2.722 3.57 3.108 ;
      RECT 3.545 2.795 3.565 3.108 ;
      RECT 3.535 2.875 3.545 3.107 ;
      RECT 3.52 2.905 3.535 3.107 ;
      RECT 3.505 2.91 3.52 3.106 ;
      RECT 3.445 2.912 3.5 3.103 ;
      RECT 3.415 2.917 3.445 3.099 ;
      RECT 3.413 2.92 3.415 3.098 ;
      RECT 3.327 2.922 3.413 3.095 ;
      RECT 3.241 2.928 3.327 3.089 ;
      RECT 3.155 2.933 3.241 3.083 ;
      RECT 3.082 2.938 3.155 3.084 ;
      RECT 2.996 2.944 3.082 3.092 ;
      RECT 2.91 2.95 2.996 3.101 ;
      RECT 2.89 2.954 2.91 3.106 ;
      RECT 2.843 2.956 2.89 3.109 ;
      RECT 2.757 2.961 2.843 3.115 ;
      RECT 2.671 2.966 2.757 3.124 ;
      RECT 2.585 2.972 2.671 3.132 ;
      RECT 2.5 2.97 2.585 3.141 ;
      RECT 2.496 2.965 2.5 3.145 ;
      RECT 2.41 2.96 2.496 3.137 ;
      RECT 2.346 2.951 2.41 3.125 ;
      RECT 2.26 2.942 2.346 3.112 ;
      RECT 2.236 2.935 2.26 3.103 ;
      RECT 2.15 2.929 2.236 3.09 ;
      RECT 2.11 2.922 2.15 3.076 ;
      RECT 2.105 2.912 2.11 3.072 ;
      RECT 2.095 2.9 2.105 3.071 ;
      RECT 2.075 2.87 2.095 3.068 ;
      RECT 2.02 2.79 2.075 3.062 ;
      RECT 2 2.709 2.02 3.057 ;
      RECT 1.98 2.667 2 3.053 ;
      RECT 1.955 2.62 1.98 3.047 ;
      RECT 1.95 2.595 1.955 3.044 ;
      RECT 1.915 2.575 1.95 3.039 ;
      RECT 1.906 2.575 1.915 3.032 ;
      RECT 1.82 2.575 1.906 3.002 ;
      RECT 1.815 2.575 1.82 2.965 ;
      RECT 1.78 2.575 1.8 2.887 ;
      RECT 1.775 2.617 1.78 2.852 ;
      RECT 1.77 2.692 1.775 2.808 ;
      RECT 3.22 2.497 3.395 2.745 ;
      RECT 3.22 2.497 3.4 2.743 ;
      RECT 3.215 2.529 3.4 2.703 ;
      RECT 3.245 2.47 3.415 2.69 ;
      RECT 3.21 2.547 3.415 2.623 ;
      RECT 2.52 2.01 2.69 2.185 ;
      RECT 2.52 2.01 2.862 2.177 ;
      RECT 2.52 2.01 2.945 2.171 ;
      RECT 2.52 2.01 2.98 2.167 ;
      RECT 2.52 2.01 3 2.166 ;
      RECT 2.52 2.01 3.086 2.162 ;
      RECT 2.98 1.835 3.15 2.157 ;
      RECT 2.555 1.942 3.18 2.155 ;
      RECT 2.545 1.997 3.185 2.153 ;
      RECT 2.52 2.033 3.195 2.148 ;
      RECT 2.52 2.06 3.2 2.078 ;
      RECT 2.585 1.885 3.16 2.155 ;
      RECT 2.776 1.87 3.16 2.155 ;
      RECT 2.61 1.873 3.16 2.155 ;
      RECT 2.69 1.871 2.776 2.182 ;
      RECT 2.776 1.868 3.155 2.155 ;
      RECT 2.96 1.845 3.155 2.155 ;
      RECT 2.862 1.866 3.155 2.155 ;
      RECT 2.945 1.86 2.96 2.168 ;
      RECT 3.095 3.225 3.1 3.425 ;
      RECT 2.56 3.29 2.605 3.425 ;
      RECT 3.13 3.225 3.15 3.398 ;
      RECT 3.1 3.225 3.13 3.413 ;
      RECT 3.035 3.225 3.095 3.45 ;
      RECT 3.02 3.225 3.035 3.48 ;
      RECT 3.005 3.225 3.02 3.493 ;
      RECT 2.985 3.225 3.005 3.508 ;
      RECT 2.98 3.225 2.985 3.517 ;
      RECT 2.97 3.229 2.98 3.522 ;
      RECT 2.955 3.239 2.97 3.533 ;
      RECT 2.93 3.255 2.955 3.543 ;
      RECT 2.92 3.269 2.93 3.545 ;
      RECT 2.9 3.281 2.92 3.542 ;
      RECT 2.87 3.302 2.9 3.536 ;
      RECT 2.86 3.314 2.87 3.531 ;
      RECT 2.85 3.312 2.86 3.528 ;
      RECT 2.835 3.311 2.85 3.523 ;
      RECT 2.83 3.31 2.835 3.518 ;
      RECT 2.795 3.308 2.83 3.508 ;
      RECT 2.775 3.305 2.795 3.49 ;
      RECT 2.765 3.303 2.775 3.485 ;
      RECT 2.755 3.302 2.765 3.48 ;
      RECT 2.72 3.3 2.755 3.468 ;
      RECT 2.665 3.296 2.72 3.448 ;
      RECT 2.655 3.294 2.665 3.433 ;
      RECT 2.65 3.294 2.655 3.428 ;
      RECT 2.605 3.292 2.65 3.425 ;
      RECT 2.51 3.29 2.56 3.429 ;
      RECT 2.5 3.291 2.51 3.434 ;
      RECT 2.44 3.298 2.5 3.448 ;
      RECT 2.415 3.306 2.44 3.468 ;
      RECT 2.405 3.31 2.415 3.48 ;
      RECT 2.4 3.311 2.405 3.485 ;
      RECT 2.385 3.313 2.4 3.488 ;
      RECT 2.37 3.315 2.385 3.493 ;
      RECT 2.365 3.315 2.37 3.496 ;
      RECT 2.32 3.32 2.365 3.507 ;
      RECT 2.315 3.324 2.32 3.519 ;
      RECT 2.29 3.32 2.315 3.523 ;
      RECT 2.28 3.316 2.29 3.527 ;
      RECT 2.27 3.315 2.28 3.531 ;
      RECT 2.255 3.305 2.27 3.537 ;
      RECT 2.25 3.293 2.255 3.541 ;
      RECT 2.245 3.29 2.25 3.542 ;
      RECT 2.24 3.287 2.245 3.544 ;
      RECT 2.225 3.275 2.24 3.543 ;
      RECT 2.21 3.257 2.225 3.54 ;
      RECT 2.19 3.236 2.21 3.533 ;
      RECT 2.125 3.225 2.19 3.505 ;
      RECT 2.121 3.225 2.125 3.484 ;
      RECT 2.035 3.225 2.121 3.454 ;
      RECT 2.02 3.225 2.035 3.41 ;
      RECT 2.595 2.325 2.6 2.56 ;
      RECT 1.725 2.241 1.73 2.445 ;
      RECT 2.305 2.27 2.31 2.425 ;
      RECT 2.225 2.25 2.23 2.425 ;
      RECT 2.895 2.392 2.91 2.745 ;
      RECT 2.821 2.377 2.895 2.745 ;
      RECT 2.735 2.36 2.821 2.745 ;
      RECT 2.725 2.35 2.735 2.743 ;
      RECT 2.72 2.348 2.725 2.738 ;
      RECT 2.705 2.346 2.72 2.724 ;
      RECT 2.635 2.338 2.705 2.664 ;
      RECT 2.615 2.329 2.635 2.598 ;
      RECT 2.61 2.326 2.615 2.578 ;
      RECT 2.6 2.325 2.61 2.568 ;
      RECT 2.59 2.325 2.595 2.552 ;
      RECT 2.58 2.324 2.59 2.542 ;
      RECT 2.57 2.322 2.58 2.53 ;
      RECT 2.555 2.319 2.57 2.51 ;
      RECT 2.545 2.317 2.555 2.495 ;
      RECT 2.525 2.314 2.545 2.483 ;
      RECT 2.52 2.312 2.525 2.473 ;
      RECT 2.495 2.31 2.52 2.46 ;
      RECT 2.465 2.305 2.495 2.445 ;
      RECT 2.385 2.296 2.465 2.436 ;
      RECT 2.34 2.285 2.385 2.429 ;
      RECT 2.32 2.276 2.34 2.426 ;
      RECT 2.31 2.271 2.32 2.425 ;
      RECT 2.265 2.265 2.305 2.425 ;
      RECT 2.25 2.257 2.265 2.425 ;
      RECT 2.23 2.252 2.25 2.425 ;
      RECT 2.21 2.249 2.225 2.425 ;
      RECT 2.127 2.248 2.21 2.424 ;
      RECT 2.041 2.247 2.127 2.42 ;
      RECT 1.955 2.245 2.041 2.417 ;
      RECT 1.902 2.244 1.955 2.419 ;
      RECT 1.816 2.243 1.902 2.428 ;
      RECT 1.73 2.242 1.816 2.44 ;
      RECT 1.71 2.241 1.725 2.448 ;
      RECT 1.63 2.24 1.71 2.46 ;
      RECT 1.605 2.24 1.63 2.473 ;
      RECT 1.58 2.24 1.605 2.488 ;
      RECT 1.575 2.24 1.58 2.51 ;
      RECT 1.57 2.24 1.575 2.528 ;
      RECT 1.565 2.24 1.57 2.545 ;
      RECT 1.56 2.24 1.565 2.558 ;
      RECT 1.555 2.24 1.56 2.568 ;
      RECT 1.515 2.24 1.555 2.653 ;
      RECT 1.5 2.24 1.515 2.738 ;
      RECT 1.49 2.241 1.5 2.75 ;
      RECT 1.455 2.246 1.49 2.755 ;
      RECT 1.415 2.255 1.455 2.755 ;
      RECT 1.4 2.265 1.415 2.755 ;
      RECT 1.395 2.275 1.4 2.755 ;
      RECT 1.375 2.302 1.395 2.755 ;
      RECT 1.325 2.385 1.375 2.755 ;
      RECT 1.32 2.447 1.325 2.755 ;
      RECT 1.31 2.46 1.32 2.755 ;
      RECT 1.3 2.482 1.31 2.755 ;
      RECT 1.29 2.507 1.3 2.75 ;
      RECT 1.285 2.545 1.29 2.743 ;
      RECT 1.275 2.655 1.285 2.738 ;
      RECT 2.67 3.576 2.685 3.835 ;
      RECT 2.67 3.591 2.69 3.834 ;
      RECT 2.586 3.591 2.69 3.832 ;
      RECT 2.586 3.605 2.695 3.831 ;
      RECT 2.5 3.647 2.7 3.828 ;
      RECT 2.495 3.59 2.685 3.823 ;
      RECT 2.495 3.661 2.705 3.82 ;
      RECT 2.49 3.692 2.705 3.818 ;
      RECT 2.495 3.689 2.72 3.808 ;
      RECT 2.49 3.735 2.735 3.793 ;
      RECT 2.49 3.763 2.74 3.778 ;
      RECT 2.5 3.565 2.67 3.828 ;
      RECT 2.26 2.575 2.43 2.745 ;
      RECT 2.225 2.575 2.43 2.74 ;
      RECT 2.215 2.575 2.43 2.733 ;
      RECT 2.21 2.56 2.38 2.73 ;
      RECT 1.04 3.097 1.305 3.54 ;
      RECT 1.035 3.068 1.25 3.538 ;
      RECT 1.03 3.222 1.31 3.533 ;
      RECT 1.035 3.117 1.31 3.533 ;
      RECT 1.035 3.128 1.32 3.52 ;
      RECT 1.035 3.075 1.28 3.538 ;
      RECT 1.04 3.062 1.25 3.54 ;
      RECT 1.04 3.06 1.2 3.54 ;
      RECT 1.141 3.052 1.2 3.54 ;
      RECT 1.055 3.053 1.2 3.54 ;
      RECT 1.141 3.051 1.19 3.54 ;
      RECT 0.945 1.866 1.12 2.165 ;
      RECT 0.995 1.828 1.12 2.165 ;
      RECT 0.98 1.83 1.206 2.157 ;
      RECT 0.98 1.833 1.245 2.144 ;
      RECT 0.98 1.834 1.255 2.13 ;
      RECT 0.935 1.885 1.255 2.12 ;
      RECT 0.98 1.835 1.26 2.115 ;
      RECT 0.935 2.045 1.265 2.105 ;
      RECT 0.92 1.905 1.26 2.045 ;
      RECT 0.915 1.921 1.26 1.985 ;
      RECT 0.96 1.845 1.26 2.115 ;
      RECT 0.995 1.826 1.081 2.165 ;
      RECT -1.625 7.855 -1.455 8.305 ;
      RECT -1.57 6.075 -1.4 8.025 ;
      RECT -1.625 5.015 -1.455 6.245 ;
      RECT -2.145 5.015 -1.975 8.305 ;
      RECT -2.145 7.315 -1.74 7.645 ;
      RECT -2.145 6.475 -1.74 6.805 ;
      RECT 75.76 0.575 75.93 1.085 ;
      RECT 75.76 2.395 75.93 3.865 ;
      RECT 75.76 5.015 75.93 6.485 ;
      RECT 75.76 7.795 75.93 8.305 ;
      RECT 74.77 0.575 74.94 1.085 ;
      RECT 74.77 2.395 74.94 3.865 ;
      RECT 74.77 5.015 74.94 6.485 ;
      RECT 74.77 7.795 74.94 8.305 ;
      RECT 73.405 0.575 73.575 3.865 ;
      RECT 73.405 5.015 73.575 8.305 ;
      RECT 72.975 0.575 73.145 1.085 ;
      RECT 72.975 1.655 73.145 3.865 ;
      RECT 72.975 5.015 73.145 7.225 ;
      RECT 72.975 7.795 73.145 8.305 ;
      RECT 71.605 1.66 71.775 2.935 ;
      RECT 71.605 5.945 71.775 7.22 ;
      RECT 67.77 5.015 67.94 8.305 ;
      RECT 67.34 5.015 67.51 7.225 ;
      RECT 67.34 7.795 67.51 8.305 ;
      RECT 65.97 5.945 66.14 7.22 ;
      RECT 60.5 0.575 60.67 1.085 ;
      RECT 60.5 2.395 60.67 3.865 ;
      RECT 60.5 5.015 60.67 6.485 ;
      RECT 60.5 7.795 60.67 8.305 ;
      RECT 59.51 0.575 59.68 1.085 ;
      RECT 59.51 2.395 59.68 3.865 ;
      RECT 59.51 5.015 59.68 6.485 ;
      RECT 59.51 7.795 59.68 8.305 ;
      RECT 58.145 0.575 58.315 3.865 ;
      RECT 58.145 5.015 58.315 8.305 ;
      RECT 57.715 0.575 57.885 1.085 ;
      RECT 57.715 1.655 57.885 3.865 ;
      RECT 57.715 5.015 57.885 7.225 ;
      RECT 57.715 7.795 57.885 8.305 ;
      RECT 56.345 1.66 56.515 2.935 ;
      RECT 56.345 5.945 56.515 7.22 ;
      RECT 52.51 5.015 52.68 8.305 ;
      RECT 52.08 5.015 52.25 7.225 ;
      RECT 52.08 7.795 52.25 8.305 ;
      RECT 50.71 5.945 50.88 7.22 ;
      RECT 45.24 0.575 45.41 1.085 ;
      RECT 45.24 2.395 45.41 3.865 ;
      RECT 45.24 5.015 45.41 6.485 ;
      RECT 45.24 7.795 45.41 8.305 ;
      RECT 44.25 0.575 44.42 1.085 ;
      RECT 44.25 2.395 44.42 3.865 ;
      RECT 44.25 5.015 44.42 6.485 ;
      RECT 44.25 7.795 44.42 8.305 ;
      RECT 42.885 0.575 43.055 3.865 ;
      RECT 42.885 5.015 43.055 8.305 ;
      RECT 42.455 0.575 42.625 1.085 ;
      RECT 42.455 1.655 42.625 3.865 ;
      RECT 42.455 5.015 42.625 7.225 ;
      RECT 42.455 7.795 42.625 8.305 ;
      RECT 41.085 1.66 41.255 2.935 ;
      RECT 41.085 5.945 41.255 7.22 ;
      RECT 37.25 5.015 37.42 8.305 ;
      RECT 36.82 5.015 36.99 7.225 ;
      RECT 36.82 7.795 36.99 8.305 ;
      RECT 35.45 5.945 35.62 7.22 ;
      RECT 29.98 0.575 30.15 1.085 ;
      RECT 29.98 2.395 30.15 3.865 ;
      RECT 29.98 5.015 30.15 6.485 ;
      RECT 29.98 7.795 30.15 8.305 ;
      RECT 28.99 0.575 29.16 1.085 ;
      RECT 28.99 2.395 29.16 3.865 ;
      RECT 28.99 5.015 29.16 6.485 ;
      RECT 28.99 7.795 29.16 8.305 ;
      RECT 27.625 0.575 27.795 3.865 ;
      RECT 27.625 5.015 27.795 8.305 ;
      RECT 27.195 0.575 27.365 1.085 ;
      RECT 27.195 1.655 27.365 3.865 ;
      RECT 27.195 5.015 27.365 7.225 ;
      RECT 27.195 7.795 27.365 8.305 ;
      RECT 25.825 1.66 25.995 2.935 ;
      RECT 25.825 5.945 25.995 7.22 ;
      RECT 21.99 5.015 22.16 8.305 ;
      RECT 21.56 5.015 21.73 7.225 ;
      RECT 21.56 7.795 21.73 8.305 ;
      RECT 20.19 5.945 20.36 7.22 ;
      RECT 14.72 0.575 14.89 1.085 ;
      RECT 14.72 2.395 14.89 3.865 ;
      RECT 14.72 5.015 14.89 6.485 ;
      RECT 14.72 7.795 14.89 8.305 ;
      RECT 13.73 0.575 13.9 1.085 ;
      RECT 13.73 2.395 13.9 3.865 ;
      RECT 13.73 5.015 13.9 6.485 ;
      RECT 13.73 7.795 13.9 8.305 ;
      RECT 12.365 0.575 12.535 3.865 ;
      RECT 12.365 5.015 12.535 8.305 ;
      RECT 11.935 0.575 12.105 1.085 ;
      RECT 11.935 1.655 12.105 3.865 ;
      RECT 11.935 5.015 12.105 7.225 ;
      RECT 11.935 7.795 12.105 8.305 ;
      RECT 10.565 1.66 10.735 2.935 ;
      RECT 10.565 5.945 10.735 7.22 ;
      RECT 6.73 5.015 6.9 8.305 ;
      RECT 6.3 5.015 6.47 7.225 ;
      RECT 6.3 7.795 6.47 8.305 ;
      RECT 4.93 5.945 5.1 7.22 ;
      RECT -1.195 5.015 -1.025 7.225 ;
      RECT -1.195 7.795 -1.025 8.305 ;
      RECT -2.565 5.945 -2.395 7.22 ;
  END
END sky130_osu_ring_oscillator_mpr2ya_8_b0r1

MACRO sky130_osu_ring_oscillator_mpr2ya_8_b0r2
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 2.795 0 ;
  SIZE 79.095 BY 8.88 ;
  SYMMETRY X Y R90 ;
  SITE CoreSite ;
  OBS
    LAYER met3 ;
      RECT 70.91 0.95 71.24 3.055 ;
      RECT 70.91 2.735 71.255 3.025 ;
      RECT 64.9 0.95 65.23 2.585 ;
      RECT 64.9 0.95 71.24 1.28 ;
      RECT 67.24 7.055 67.61 7.425 ;
      RECT 67.275 4.27 67.575 7.425 ;
      RECT 63.085 4.27 67.575 4.57 ;
      RECT 66.265 1.855 66.565 4.57 ;
      RECT 63.085 2.435 63.385 4.57 ;
      RECT 66.22 2.76 66.565 3.49 ;
      RECT 62.98 2.015 63.31 2.745 ;
      RECT 65.86 1.855 66.59 2.185 ;
      RECT 55.65 0.95 55.98 3.055 ;
      RECT 55.65 2.735 55.995 3.025 ;
      RECT 49.64 0.95 49.97 2.585 ;
      RECT 49.64 0.95 55.98 1.28 ;
      RECT 51.98 7.055 52.35 7.425 ;
      RECT 52.015 4.27 52.315 7.425 ;
      RECT 47.825 4.27 52.315 4.57 ;
      RECT 51.005 1.855 51.305 4.57 ;
      RECT 47.825 2.435 48.125 4.57 ;
      RECT 50.96 2.76 51.305 3.49 ;
      RECT 47.72 2.015 48.05 2.745 ;
      RECT 50.6 1.855 51.33 2.185 ;
      RECT 40.39 0.95 40.72 3.055 ;
      RECT 40.39 2.735 40.735 3.025 ;
      RECT 34.38 0.95 34.71 2.585 ;
      RECT 34.38 0.95 40.72 1.28 ;
      RECT 36.72 7.055 37.09 7.425 ;
      RECT 36.755 4.27 37.055 7.425 ;
      RECT 32.565 4.27 37.055 4.57 ;
      RECT 35.745 1.855 36.045 4.57 ;
      RECT 32.565 2.435 32.865 4.57 ;
      RECT 35.7 2.76 36.045 3.49 ;
      RECT 32.46 2.015 32.79 2.745 ;
      RECT 35.34 1.855 36.07 2.185 ;
      RECT 25.13 0.95 25.46 3.055 ;
      RECT 25.13 2.735 25.475 3.025 ;
      RECT 19.12 0.95 19.45 2.585 ;
      RECT 19.12 0.95 25.46 1.28 ;
      RECT 21.46 7.055 21.83 7.425 ;
      RECT 21.495 4.27 21.795 7.425 ;
      RECT 17.305 4.27 21.795 4.57 ;
      RECT 20.485 1.855 20.785 4.57 ;
      RECT 17.305 2.435 17.605 4.57 ;
      RECT 20.44 2.76 20.785 3.49 ;
      RECT 17.2 2.015 17.53 2.745 ;
      RECT 20.08 1.855 20.81 2.185 ;
      RECT 9.87 0.95 10.2 3.055 ;
      RECT 9.87 2.735 10.215 3.025 ;
      RECT 3.86 0.95 4.19 2.585 ;
      RECT 3.86 0.95 10.2 1.28 ;
      RECT 6.2 7.055 6.57 7.425 ;
      RECT 6.235 4.27 6.535 7.425 ;
      RECT 2.045 4.27 6.535 4.57 ;
      RECT 5.225 1.855 5.525 4.57 ;
      RECT 2.045 2.435 2.345 4.57 ;
      RECT 5.18 2.76 5.525 3.49 ;
      RECT 1.94 2.015 2.27 2.745 ;
      RECT 4.82 1.855 5.55 2.185 ;
      RECT 69.34 2.015 69.67 2.745 ;
      RECT 68.14 2.88 68.47 3.61 ;
      RECT 67.3 1.855 68.03 2.185 ;
      RECT 63.7 2.015 64.03 2.745 ;
      RECT 54.08 2.015 54.41 2.745 ;
      RECT 52.88 2.88 53.21 3.61 ;
      RECT 52.04 1.855 52.77 2.185 ;
      RECT 48.44 2.015 48.77 2.745 ;
      RECT 38.82 2.015 39.15 2.745 ;
      RECT 37.62 2.88 37.95 3.61 ;
      RECT 36.78 1.855 37.51 2.185 ;
      RECT 33.18 2.015 33.51 2.745 ;
      RECT 23.56 2.015 23.89 2.745 ;
      RECT 22.36 2.88 22.69 3.61 ;
      RECT 21.52 1.855 22.25 2.185 ;
      RECT 17.92 2.015 18.25 2.745 ;
      RECT 8.3 2.015 8.63 2.745 ;
      RECT 7.1 2.88 7.43 3.61 ;
      RECT 6.26 1.855 6.99 2.185 ;
      RECT 2.66 2.015 2.99 2.745 ;
    LAYER via2 ;
      RECT 71.01 2.78 71.21 2.98 ;
      RECT 69.405 2.48 69.605 2.68 ;
      RECT 68.205 3.04 68.405 3.24 ;
      RECT 67.365 1.92 67.565 2.12 ;
      RECT 67.325 7.14 67.525 7.34 ;
      RECT 66.285 2.825 66.485 3.025 ;
      RECT 65.925 1.92 66.125 2.12 ;
      RECT 64.965 1.92 65.165 2.12 ;
      RECT 63.765 2.48 63.965 2.68 ;
      RECT 63.045 2.48 63.245 2.68 ;
      RECT 55.75 2.78 55.95 2.98 ;
      RECT 54.145 2.48 54.345 2.68 ;
      RECT 52.945 3.04 53.145 3.24 ;
      RECT 52.105 1.92 52.305 2.12 ;
      RECT 52.065 7.14 52.265 7.34 ;
      RECT 51.025 2.825 51.225 3.025 ;
      RECT 50.665 1.92 50.865 2.12 ;
      RECT 49.705 1.92 49.905 2.12 ;
      RECT 48.505 2.48 48.705 2.68 ;
      RECT 47.785 2.48 47.985 2.68 ;
      RECT 40.49 2.78 40.69 2.98 ;
      RECT 38.885 2.48 39.085 2.68 ;
      RECT 37.685 3.04 37.885 3.24 ;
      RECT 36.845 1.92 37.045 2.12 ;
      RECT 36.805 7.14 37.005 7.34 ;
      RECT 35.765 2.825 35.965 3.025 ;
      RECT 35.405 1.92 35.605 2.12 ;
      RECT 34.445 1.92 34.645 2.12 ;
      RECT 33.245 2.48 33.445 2.68 ;
      RECT 32.525 2.48 32.725 2.68 ;
      RECT 25.23 2.78 25.43 2.98 ;
      RECT 23.625 2.48 23.825 2.68 ;
      RECT 22.425 3.04 22.625 3.24 ;
      RECT 21.585 1.92 21.785 2.12 ;
      RECT 21.545 7.14 21.745 7.34 ;
      RECT 20.505 2.825 20.705 3.025 ;
      RECT 20.145 1.92 20.345 2.12 ;
      RECT 19.185 1.92 19.385 2.12 ;
      RECT 17.985 2.48 18.185 2.68 ;
      RECT 17.265 2.48 17.465 2.68 ;
      RECT 9.97 2.78 10.17 2.98 ;
      RECT 8.365 2.48 8.565 2.68 ;
      RECT 7.165 3.04 7.365 3.24 ;
      RECT 6.325 1.92 6.525 2.12 ;
      RECT 6.285 7.14 6.485 7.34 ;
      RECT 5.245 2.825 5.445 3.025 ;
      RECT 4.885 1.92 5.085 2.12 ;
      RECT 3.925 1.92 4.125 2.12 ;
      RECT 2.725 2.48 2.925 2.68 ;
      RECT 2.005 2.48 2.205 2.68 ;
    LAYER met2 ;
      RECT -1.57 8.4 75.93 8.57 ;
      RECT 75.76 7.275 75.93 8.57 ;
      RECT -1.57 6.255 -1.4 8.57 ;
      RECT 75.73 7.275 76.08 7.625 ;
      RECT -1.63 6.255 -1.34 6.605 ;
      RECT 72.57 6.22 72.89 6.545 ;
      RECT 72.6 5.695 72.77 6.545 ;
      RECT 72.6 5.695 72.775 6.045 ;
      RECT 72.6 5.695 73.575 5.87 ;
      RECT 73.4 1.965 73.575 5.87 ;
      RECT 73.345 1.965 73.695 2.315 ;
      RECT 73.37 6.655 73.695 6.98 ;
      RECT 72.255 6.745 73.695 6.915 ;
      RECT 72.255 2.395 72.415 6.915 ;
      RECT 72.57 2.365 72.89 2.685 ;
      RECT 72.255 2.395 72.89 2.565 ;
      RECT 71.52 5.86 71.86 6.21 ;
      RECT 71.6 2.705 71.775 6.21 ;
      RECT 71.525 2.705 71.865 3.055 ;
      RECT 70.92 2.705 71.305 3.055 ;
      RECT 70.91 2.77 71.305 2.97 ;
      RECT 71.055 2.7 71.225 3.055 ;
      RECT 69.365 2.44 69.645 2.72 ;
      RECT 69.36 2.44 69.645 2.673 ;
      RECT 69.34 2.44 69.645 2.65 ;
      RECT 69.33 2.44 69.645 2.63 ;
      RECT 69.32 2.44 69.645 2.615 ;
      RECT 69.295 2.44 69.645 2.588 ;
      RECT 69.285 2.44 69.645 2.563 ;
      RECT 69.24 2.295 69.52 2.555 ;
      RECT 69.24 2.39 69.62 2.555 ;
      RECT 69.24 2.335 69.565 2.555 ;
      RECT 69.24 2.327 69.56 2.555 ;
      RECT 69.24 2.317 69.555 2.555 ;
      RECT 69.24 2.305 69.55 2.555 ;
      RECT 68.165 3 68.445 3.28 ;
      RECT 68.165 3 68.48 3.26 ;
      RECT 60.445 6.655 60.795 7.005 ;
      RECT 67.91 6.61 68.26 6.96 ;
      RECT 60.445 6.685 68.26 6.885 ;
      RECT 68.2 2.42 68.25 2.68 ;
      RECT 67.99 2.42 67.995 2.68 ;
      RECT 67.185 1.975 67.215 2.235 ;
      RECT 66.955 1.975 67.03 2.235 ;
      RECT 68.175 2.37 68.2 2.68 ;
      RECT 68.17 2.327 68.175 2.68 ;
      RECT 68.165 2.31 68.17 2.68 ;
      RECT 68.16 2.297 68.165 2.68 ;
      RECT 68.085 2.18 68.16 2.68 ;
      RECT 68.04 1.997 68.085 2.68 ;
      RECT 68.035 1.925 68.04 2.68 ;
      RECT 68.02 1.9 68.035 2.68 ;
      RECT 67.995 1.862 68.02 2.68 ;
      RECT 67.985 1.842 67.995 2.402 ;
      RECT 67.97 1.834 67.985 2.357 ;
      RECT 67.965 1.826 67.97 2.328 ;
      RECT 67.96 1.823 67.965 2.308 ;
      RECT 67.955 1.82 67.96 2.288 ;
      RECT 67.95 1.817 67.955 2.268 ;
      RECT 67.92 1.806 67.95 2.205 ;
      RECT 67.9 1.791 67.92 2.12 ;
      RECT 67.895 1.783 67.9 2.083 ;
      RECT 67.885 1.777 67.895 2.05 ;
      RECT 67.87 1.769 67.885 2.01 ;
      RECT 67.865 1.762 67.87 1.97 ;
      RECT 67.86 1.759 67.865 1.948 ;
      RECT 67.855 1.756 67.86 1.935 ;
      RECT 67.85 1.755 67.855 1.925 ;
      RECT 67.835 1.749 67.85 1.915 ;
      RECT 67.81 1.736 67.835 1.9 ;
      RECT 67.76 1.711 67.81 1.871 ;
      RECT 67.745 1.69 67.76 1.846 ;
      RECT 67.735 1.683 67.745 1.835 ;
      RECT 67.68 1.664 67.735 1.808 ;
      RECT 67.655 1.642 67.68 1.781 ;
      RECT 67.65 1.635 67.655 1.776 ;
      RECT 67.635 1.635 67.65 1.774 ;
      RECT 67.61 1.627 67.635 1.77 ;
      RECT 67.595 1.625 67.61 1.766 ;
      RECT 67.565 1.625 67.595 1.763 ;
      RECT 67.555 1.625 67.565 1.758 ;
      RECT 67.51 1.625 67.555 1.756 ;
      RECT 67.481 1.625 67.51 1.757 ;
      RECT 67.395 1.625 67.481 1.759 ;
      RECT 67.381 1.626 67.395 1.761 ;
      RECT 67.295 1.627 67.381 1.763 ;
      RECT 67.28 1.628 67.295 1.773 ;
      RECT 67.275 1.629 67.28 1.782 ;
      RECT 67.255 1.632 67.275 1.792 ;
      RECT 67.24 1.64 67.255 1.807 ;
      RECT 67.22 1.658 67.24 1.822 ;
      RECT 67.21 1.67 67.22 1.845 ;
      RECT 67.2 1.679 67.21 1.875 ;
      RECT 67.185 1.691 67.2 1.92 ;
      RECT 67.13 1.724 67.185 2.235 ;
      RECT 67.125 1.752 67.13 2.235 ;
      RECT 67.105 1.767 67.125 2.235 ;
      RECT 67.07 1.827 67.105 2.235 ;
      RECT 67.068 1.877 67.07 2.235 ;
      RECT 67.065 1.885 67.068 2.235 ;
      RECT 67.055 1.9 67.065 2.235 ;
      RECT 67.05 1.912 67.055 2.235 ;
      RECT 67.04 1.937 67.05 2.235 ;
      RECT 67.03 1.965 67.04 2.235 ;
      RECT 64.935 3.47 64.985 3.73 ;
      RECT 67.845 3.02 67.905 3.28 ;
      RECT 67.83 3.02 67.845 3.29 ;
      RECT 67.811 3.02 67.83 3.323 ;
      RECT 67.725 3.02 67.811 3.448 ;
      RECT 67.645 3.02 67.725 3.63 ;
      RECT 67.64 3.257 67.645 3.715 ;
      RECT 67.615 3.327 67.64 3.743 ;
      RECT 67.61 3.397 67.615 3.77 ;
      RECT 67.59 3.469 67.61 3.792 ;
      RECT 67.585 3.536 67.59 3.815 ;
      RECT 67.575 3.565 67.585 3.83 ;
      RECT 67.565 3.587 67.575 3.847 ;
      RECT 67.56 3.597 67.565 3.858 ;
      RECT 67.555 3.605 67.56 3.866 ;
      RECT 67.545 3.613 67.555 3.878 ;
      RECT 67.54 3.625 67.545 3.888 ;
      RECT 67.535 3.633 67.54 3.893 ;
      RECT 67.515 3.651 67.535 3.903 ;
      RECT 67.51 3.668 67.515 3.91 ;
      RECT 67.505 3.676 67.51 3.911 ;
      RECT 67.5 3.687 67.505 3.913 ;
      RECT 67.46 3.725 67.5 3.923 ;
      RECT 67.455 3.76 67.46 3.934 ;
      RECT 67.45 3.765 67.455 3.937 ;
      RECT 67.425 3.775 67.45 3.944 ;
      RECT 67.415 3.789 67.425 3.953 ;
      RECT 67.395 3.801 67.415 3.956 ;
      RECT 67.345 3.82 67.395 3.96 ;
      RECT 67.3 3.835 67.345 3.965 ;
      RECT 67.235 3.838 67.3 3.971 ;
      RECT 67.22 3.836 67.235 3.978 ;
      RECT 67.19 3.835 67.22 3.978 ;
      RECT 67.151 3.834 67.19 3.974 ;
      RECT 67.065 3.831 67.151 3.97 ;
      RECT 67.048 3.829 67.065 3.967 ;
      RECT 66.962 3.827 67.048 3.964 ;
      RECT 66.876 3.824 66.962 3.958 ;
      RECT 66.79 3.82 66.876 3.953 ;
      RECT 66.712 3.817 66.79 3.949 ;
      RECT 66.626 3.814 66.712 3.947 ;
      RECT 66.54 3.811 66.626 3.944 ;
      RECT 66.482 3.809 66.54 3.941 ;
      RECT 66.396 3.806 66.482 3.939 ;
      RECT 66.31 3.802 66.396 3.937 ;
      RECT 66.224 3.799 66.31 3.934 ;
      RECT 66.138 3.795 66.224 3.932 ;
      RECT 66.052 3.791 66.138 3.929 ;
      RECT 65.966 3.788 66.052 3.927 ;
      RECT 65.88 3.784 65.966 3.924 ;
      RECT 65.794 3.781 65.88 3.922 ;
      RECT 65.708 3.777 65.794 3.919 ;
      RECT 65.622 3.774 65.708 3.917 ;
      RECT 65.536 3.77 65.622 3.914 ;
      RECT 65.45 3.767 65.536 3.912 ;
      RECT 65.44 3.765 65.45 3.908 ;
      RECT 65.435 3.765 65.44 3.906 ;
      RECT 65.395 3.76 65.435 3.9 ;
      RECT 65.381 3.751 65.395 3.893 ;
      RECT 65.295 3.721 65.381 3.878 ;
      RECT 65.275 3.687 65.295 3.863 ;
      RECT 65.205 3.656 65.275 3.85 ;
      RECT 65.2 3.631 65.205 3.839 ;
      RECT 65.195 3.625 65.2 3.837 ;
      RECT 65.126 3.47 65.195 3.825 ;
      RECT 65.04 3.47 65.126 3.799 ;
      RECT 65.015 3.47 65.04 3.778 ;
      RECT 65.01 3.47 65.015 3.768 ;
      RECT 65.005 3.47 65.01 3.76 ;
      RECT 64.985 3.47 65.005 3.743 ;
      RECT 67.405 2.04 67.665 2.3 ;
      RECT 67.39 2.04 67.665 2.203 ;
      RECT 67.36 2.04 67.665 2.178 ;
      RECT 67.325 1.88 67.605 2.16 ;
      RECT 67.295 3.37 67.355 3.63 ;
      RECT 66.32 2.06 66.375 2.32 ;
      RECT 67.255 3.327 67.295 3.63 ;
      RECT 67.226 3.248 67.255 3.63 ;
      RECT 67.14 3.12 67.226 3.63 ;
      RECT 67.12 3 67.14 3.63 ;
      RECT 67.095 2.951 67.12 3.63 ;
      RECT 67.09 2.916 67.095 3.48 ;
      RECT 67.06 2.876 67.09 3.418 ;
      RECT 67.035 2.813 67.06 3.333 ;
      RECT 67.025 2.775 67.035 3.27 ;
      RECT 67.01 2.75 67.025 3.231 ;
      RECT 66.967 2.708 67.01 3.137 ;
      RECT 66.965 2.681 66.967 3.064 ;
      RECT 66.96 2.676 66.965 3.055 ;
      RECT 66.955 2.669 66.96 3.03 ;
      RECT 66.95 2.663 66.955 3.015 ;
      RECT 66.945 2.657 66.95 3.003 ;
      RECT 66.935 2.648 66.945 2.985 ;
      RECT 66.93 2.639 66.935 2.963 ;
      RECT 66.905 2.62 66.93 2.913 ;
      RECT 66.9 2.601 66.905 2.863 ;
      RECT 66.885 2.587 66.9 2.823 ;
      RECT 66.88 2.573 66.885 2.79 ;
      RECT 66.875 2.566 66.88 2.783 ;
      RECT 66.86 2.553 66.875 2.775 ;
      RECT 66.815 2.515 66.86 2.748 ;
      RECT 66.785 2.468 66.815 2.713 ;
      RECT 66.765 2.437 66.785 2.69 ;
      RECT 66.685 2.37 66.765 2.643 ;
      RECT 66.655 2.3 66.685 2.59 ;
      RECT 66.65 2.277 66.655 2.573 ;
      RECT 66.62 2.255 66.65 2.558 ;
      RECT 66.59 2.214 66.62 2.53 ;
      RECT 66.585 2.189 66.59 2.515 ;
      RECT 66.58 2.183 66.585 2.508 ;
      RECT 66.57 2.06 66.58 2.5 ;
      RECT 66.56 2.06 66.57 2.493 ;
      RECT 66.555 2.06 66.56 2.485 ;
      RECT 66.535 2.06 66.555 2.473 ;
      RECT 66.485 2.06 66.535 2.443 ;
      RECT 66.43 2.06 66.485 2.393 ;
      RECT 66.4 2.06 66.43 2.353 ;
      RECT 66.375 2.06 66.4 2.33 ;
      RECT 66.245 2.785 66.525 3.065 ;
      RECT 66.21 2.7 66.47 2.96 ;
      RECT 66.21 2.782 66.48 2.96 ;
      RECT 64.41 2.155 64.415 2.64 ;
      RECT 64.3 2.34 64.305 2.64 ;
      RECT 64.21 2.38 64.275 2.64 ;
      RECT 65.885 1.88 65.975 2.51 ;
      RECT 65.85 1.93 65.855 2.51 ;
      RECT 65.795 1.955 65.805 2.51 ;
      RECT 65.75 1.955 65.76 2.51 ;
      RECT 66.12 1.88 66.165 2.16 ;
      RECT 64.97 1.61 65.17 1.75 ;
      RECT 66.086 1.88 66.12 2.172 ;
      RECT 66 1.88 66.086 2.212 ;
      RECT 65.985 1.88 66 2.253 ;
      RECT 65.98 1.88 65.985 2.273 ;
      RECT 65.975 1.88 65.98 2.293 ;
      RECT 65.855 1.922 65.885 2.51 ;
      RECT 65.805 1.942 65.85 2.51 ;
      RECT 65.79 1.957 65.795 2.51 ;
      RECT 65.76 1.957 65.79 2.51 ;
      RECT 65.715 1.942 65.75 2.51 ;
      RECT 65.71 1.93 65.715 2.29 ;
      RECT 65.705 1.927 65.71 2.27 ;
      RECT 65.69 1.917 65.705 2.223 ;
      RECT 65.685 1.91 65.69 2.186 ;
      RECT 65.68 1.907 65.685 2.169 ;
      RECT 65.665 1.897 65.68 2.125 ;
      RECT 65.66 1.888 65.665 2.085 ;
      RECT 65.655 1.884 65.66 2.07 ;
      RECT 65.645 1.878 65.655 2.053 ;
      RECT 65.605 1.859 65.645 2.028 ;
      RECT 65.6 1.841 65.605 2.008 ;
      RECT 65.59 1.835 65.6 2.003 ;
      RECT 65.56 1.819 65.59 1.99 ;
      RECT 65.545 1.801 65.56 1.973 ;
      RECT 65.53 1.789 65.545 1.96 ;
      RECT 65.525 1.781 65.53 1.953 ;
      RECT 65.495 1.767 65.525 1.94 ;
      RECT 65.49 1.752 65.495 1.928 ;
      RECT 65.48 1.746 65.49 1.92 ;
      RECT 65.46 1.734 65.48 1.908 ;
      RECT 65.45 1.722 65.46 1.895 ;
      RECT 65.42 1.706 65.45 1.88 ;
      RECT 65.4 1.686 65.42 1.863 ;
      RECT 65.395 1.676 65.4 1.853 ;
      RECT 65.37 1.664 65.395 1.84 ;
      RECT 65.365 1.652 65.37 1.828 ;
      RECT 65.36 1.647 65.365 1.824 ;
      RECT 65.345 1.64 65.36 1.816 ;
      RECT 65.335 1.627 65.345 1.806 ;
      RECT 65.33 1.625 65.335 1.8 ;
      RECT 65.305 1.618 65.33 1.789 ;
      RECT 65.3 1.611 65.305 1.778 ;
      RECT 65.275 1.61 65.3 1.765 ;
      RECT 65.256 1.61 65.275 1.755 ;
      RECT 65.17 1.61 65.256 1.752 ;
      RECT 64.94 1.61 64.97 1.755 ;
      RECT 64.9 1.617 64.94 1.768 ;
      RECT 64.875 1.627 64.9 1.781 ;
      RECT 64.86 1.636 64.875 1.791 ;
      RECT 64.83 1.641 64.86 1.81 ;
      RECT 64.825 1.647 64.83 1.828 ;
      RECT 64.805 1.657 64.825 1.843 ;
      RECT 64.795 1.67 64.805 1.863 ;
      RECT 64.78 1.682 64.795 1.88 ;
      RECT 64.775 1.692 64.78 1.89 ;
      RECT 64.77 1.697 64.775 1.895 ;
      RECT 64.76 1.705 64.77 1.908 ;
      RECT 64.71 1.737 64.76 1.945 ;
      RECT 64.695 1.772 64.71 1.986 ;
      RECT 64.69 1.782 64.695 2.001 ;
      RECT 64.685 1.787 64.69 2.008 ;
      RECT 64.66 1.803 64.685 2.028 ;
      RECT 64.645 1.824 64.66 2.053 ;
      RECT 64.62 1.845 64.645 2.078 ;
      RECT 64.61 1.864 64.62 2.101 ;
      RECT 64.585 1.882 64.61 2.124 ;
      RECT 64.57 1.902 64.585 2.148 ;
      RECT 64.565 1.912 64.57 2.16 ;
      RECT 64.55 1.924 64.565 2.18 ;
      RECT 64.54 1.939 64.55 2.22 ;
      RECT 64.535 1.947 64.54 2.248 ;
      RECT 64.525 1.957 64.535 2.268 ;
      RECT 64.52 1.97 64.525 2.293 ;
      RECT 64.515 1.983 64.52 2.313 ;
      RECT 64.51 1.989 64.515 2.335 ;
      RECT 64.5 1.998 64.51 2.355 ;
      RECT 64.495 2.018 64.5 2.378 ;
      RECT 64.49 2.024 64.495 2.398 ;
      RECT 64.485 2.031 64.49 2.42 ;
      RECT 64.48 2.042 64.485 2.433 ;
      RECT 64.47 2.052 64.48 2.458 ;
      RECT 64.45 2.077 64.47 2.64 ;
      RECT 64.42 2.117 64.45 2.64 ;
      RECT 64.415 2.147 64.42 2.64 ;
      RECT 64.39 2.175 64.41 2.64 ;
      RECT 64.36 2.22 64.39 2.64 ;
      RECT 64.355 2.247 64.36 2.64 ;
      RECT 64.335 2.265 64.355 2.64 ;
      RECT 64.325 2.29 64.335 2.64 ;
      RECT 64.32 2.302 64.325 2.64 ;
      RECT 64.305 2.325 64.32 2.64 ;
      RECT 64.285 2.352 64.3 2.64 ;
      RECT 64.275 2.375 64.285 2.64 ;
      RECT 66.065 3.26 66.145 3.52 ;
      RECT 65.3 2.48 65.37 2.74 ;
      RECT 66.031 3.227 66.065 3.52 ;
      RECT 65.945 3.13 66.031 3.52 ;
      RECT 65.925 3.042 65.945 3.52 ;
      RECT 65.915 3.012 65.925 3.52 ;
      RECT 65.905 2.992 65.915 3.52 ;
      RECT 65.885 2.979 65.905 3.52 ;
      RECT 65.87 2.969 65.885 3.348 ;
      RECT 65.865 2.962 65.87 3.303 ;
      RECT 65.855 2.956 65.865 3.293 ;
      RECT 65.845 2.948 65.855 3.275 ;
      RECT 65.84 2.942 65.845 3.263 ;
      RECT 65.83 2.937 65.84 3.25 ;
      RECT 65.81 2.927 65.83 3.223 ;
      RECT 65.77 2.906 65.81 3.175 ;
      RECT 65.755 2.887 65.77 3.133 ;
      RECT 65.73 2.873 65.755 3.103 ;
      RECT 65.72 2.861 65.73 3.07 ;
      RECT 65.715 2.856 65.72 3.06 ;
      RECT 65.685 2.842 65.715 3.04 ;
      RECT 65.675 2.826 65.685 3.013 ;
      RECT 65.67 2.821 65.675 3.003 ;
      RECT 65.645 2.812 65.67 2.983 ;
      RECT 65.635 2.8 65.645 2.963 ;
      RECT 65.565 2.768 65.635 2.938 ;
      RECT 65.56 2.737 65.565 2.915 ;
      RECT 65.511 2.48 65.56 2.898 ;
      RECT 65.425 2.48 65.511 2.857 ;
      RECT 65.37 2.48 65.425 2.785 ;
      RECT 65.46 3.265 65.62 3.525 ;
      RECT 64.985 1.88 65.035 2.565 ;
      RECT 64.775 2.305 64.81 2.565 ;
      RECT 65.09 1.88 65.095 2.34 ;
      RECT 65.18 1.88 65.205 2.16 ;
      RECT 65.455 3.262 65.46 3.525 ;
      RECT 65.42 3.25 65.455 3.525 ;
      RECT 65.36 3.223 65.42 3.525 ;
      RECT 65.355 3.206 65.36 3.379 ;
      RECT 65.35 3.203 65.355 3.366 ;
      RECT 65.33 3.196 65.35 3.353 ;
      RECT 65.295 3.179 65.33 3.335 ;
      RECT 65.255 3.158 65.295 3.315 ;
      RECT 65.25 3.146 65.255 3.303 ;
      RECT 65.21 3.132 65.25 3.289 ;
      RECT 65.19 3.115 65.21 3.271 ;
      RECT 65.18 3.107 65.19 3.263 ;
      RECT 65.165 1.88 65.18 2.178 ;
      RECT 65.15 3.097 65.18 3.25 ;
      RECT 65.135 1.88 65.165 2.223 ;
      RECT 65.14 3.087 65.15 3.237 ;
      RECT 65.11 3.072 65.14 3.224 ;
      RECT 65.095 1.88 65.135 2.29 ;
      RECT 65.095 3.04 65.11 3.21 ;
      RECT 65.09 3.012 65.095 3.204 ;
      RECT 65.085 1.88 65.09 2.345 ;
      RECT 65.075 2.982 65.09 3.198 ;
      RECT 65.08 1.88 65.085 2.358 ;
      RECT 65.07 1.88 65.08 2.378 ;
      RECT 65.035 2.895 65.075 3.183 ;
      RECT 65.035 1.88 65.07 2.418 ;
      RECT 65.03 2.827 65.035 3.171 ;
      RECT 65.015 2.782 65.03 3.166 ;
      RECT 65.01 2.72 65.015 3.161 ;
      RECT 64.985 2.627 65.01 3.154 ;
      RECT 64.98 1.88 64.985 3.146 ;
      RECT 64.965 1.88 64.98 3.133 ;
      RECT 64.945 1.88 64.965 3.09 ;
      RECT 64.935 1.88 64.945 3.04 ;
      RECT 64.93 1.88 64.935 3.013 ;
      RECT 64.925 1.88 64.93 2.991 ;
      RECT 64.92 2.106 64.925 2.974 ;
      RECT 64.915 2.128 64.92 2.952 ;
      RECT 64.91 2.17 64.915 2.935 ;
      RECT 64.88 2.22 64.91 2.879 ;
      RECT 64.875 2.247 64.88 2.821 ;
      RECT 64.86 2.265 64.875 2.785 ;
      RECT 64.855 2.283 64.86 2.749 ;
      RECT 64.849 2.29 64.855 2.73 ;
      RECT 64.845 2.297 64.849 2.713 ;
      RECT 64.84 2.302 64.845 2.682 ;
      RECT 64.83 2.305 64.84 2.657 ;
      RECT 64.82 2.305 64.83 2.623 ;
      RECT 64.815 2.305 64.82 2.6 ;
      RECT 64.81 2.305 64.815 2.58 ;
      RECT 63.725 2.44 64.005 2.72 ;
      RECT 63.725 2.44 64.025 2.615 ;
      RECT 63.815 2.33 64.075 2.59 ;
      RECT 63.78 2.425 64.075 2.59 ;
      RECT 63.905 0.945 64.07 2.59 ;
      RECT 63.805 0.945 64.175 1.315 ;
      RECT 63.43 3.47 63.69 3.73 ;
      RECT 63.45 3.397 63.63 3.73 ;
      RECT 63.45 3.14 63.625 3.73 ;
      RECT 63.45 2.932 63.615 3.73 ;
      RECT 63.455 2.85 63.615 3.73 ;
      RECT 63.455 2.615 63.605 3.73 ;
      RECT 63.455 2.462 63.6 3.73 ;
      RECT 63.46 2.447 63.6 3.73 ;
      RECT 63.51 2.162 63.6 3.73 ;
      RECT 63.465 2.397 63.6 3.73 ;
      RECT 63.495 2.215 63.6 3.73 ;
      RECT 63.48 2.327 63.6 3.73 ;
      RECT 63.485 2.285 63.6 3.73 ;
      RECT 63.48 2.327 63.615 2.39 ;
      RECT 63.515 1.915 63.62 2.335 ;
      RECT 63.515 1.915 63.635 2.318 ;
      RECT 63.515 1.915 63.67 2.28 ;
      RECT 63.51 2.162 63.72 2.213 ;
      RECT 63.515 1.915 63.775 2.175 ;
      RECT 62.775 2.62 63.035 2.88 ;
      RECT 62.775 2.62 63.045 2.838 ;
      RECT 62.775 2.62 63.131 2.809 ;
      RECT 62.775 2.62 63.2 2.761 ;
      RECT 62.775 2.62 63.235 2.73 ;
      RECT 63.005 2.44 63.285 2.72 ;
      RECT 62.84 2.605 63.285 2.72 ;
      RECT 62.93 2.482 63.035 2.88 ;
      RECT 62.86 2.545 63.285 2.72 ;
      RECT 57.31 6.22 57.63 6.545 ;
      RECT 57.34 5.695 57.51 6.545 ;
      RECT 57.34 5.695 57.515 6.045 ;
      RECT 57.34 5.695 58.315 5.87 ;
      RECT 58.14 1.965 58.315 5.87 ;
      RECT 58.085 1.965 58.435 2.315 ;
      RECT 58.11 6.655 58.435 6.98 ;
      RECT 56.995 6.745 58.435 6.915 ;
      RECT 56.995 2.395 57.155 6.915 ;
      RECT 57.31 2.365 57.63 2.685 ;
      RECT 56.995 2.395 57.63 2.565 ;
      RECT 56.26 5.86 56.6 6.21 ;
      RECT 56.34 2.705 56.515 6.21 ;
      RECT 56.265 2.705 56.605 3.055 ;
      RECT 55.66 2.705 56.045 3.055 ;
      RECT 55.65 2.77 56.045 2.97 ;
      RECT 55.795 2.7 55.965 3.055 ;
      RECT 54.105 2.44 54.385 2.72 ;
      RECT 54.1 2.44 54.385 2.673 ;
      RECT 54.08 2.44 54.385 2.65 ;
      RECT 54.07 2.44 54.385 2.63 ;
      RECT 54.06 2.44 54.385 2.615 ;
      RECT 54.035 2.44 54.385 2.588 ;
      RECT 54.025 2.44 54.385 2.563 ;
      RECT 53.98 2.295 54.26 2.555 ;
      RECT 53.98 2.39 54.36 2.555 ;
      RECT 53.98 2.335 54.305 2.555 ;
      RECT 53.98 2.327 54.3 2.555 ;
      RECT 53.98 2.317 54.295 2.555 ;
      RECT 53.98 2.305 54.29 2.555 ;
      RECT 52.905 3 53.185 3.28 ;
      RECT 52.905 3 53.22 3.26 ;
      RECT 45.185 6.655 45.535 7.005 ;
      RECT 52.65 6.61 53 6.96 ;
      RECT 45.185 6.685 53 6.885 ;
      RECT 52.94 2.42 52.99 2.68 ;
      RECT 52.73 2.42 52.735 2.68 ;
      RECT 51.925 1.975 51.955 2.235 ;
      RECT 51.695 1.975 51.77 2.235 ;
      RECT 52.915 2.37 52.94 2.68 ;
      RECT 52.91 2.327 52.915 2.68 ;
      RECT 52.905 2.31 52.91 2.68 ;
      RECT 52.9 2.297 52.905 2.68 ;
      RECT 52.825 2.18 52.9 2.68 ;
      RECT 52.78 1.997 52.825 2.68 ;
      RECT 52.775 1.925 52.78 2.68 ;
      RECT 52.76 1.9 52.775 2.68 ;
      RECT 52.735 1.862 52.76 2.68 ;
      RECT 52.725 1.842 52.735 2.402 ;
      RECT 52.71 1.834 52.725 2.357 ;
      RECT 52.705 1.826 52.71 2.328 ;
      RECT 52.7 1.823 52.705 2.308 ;
      RECT 52.695 1.82 52.7 2.288 ;
      RECT 52.69 1.817 52.695 2.268 ;
      RECT 52.66 1.806 52.69 2.205 ;
      RECT 52.64 1.791 52.66 2.12 ;
      RECT 52.635 1.783 52.64 2.083 ;
      RECT 52.625 1.777 52.635 2.05 ;
      RECT 52.61 1.769 52.625 2.01 ;
      RECT 52.605 1.762 52.61 1.97 ;
      RECT 52.6 1.759 52.605 1.948 ;
      RECT 52.595 1.756 52.6 1.935 ;
      RECT 52.59 1.755 52.595 1.925 ;
      RECT 52.575 1.749 52.59 1.915 ;
      RECT 52.55 1.736 52.575 1.9 ;
      RECT 52.5 1.711 52.55 1.871 ;
      RECT 52.485 1.69 52.5 1.846 ;
      RECT 52.475 1.683 52.485 1.835 ;
      RECT 52.42 1.664 52.475 1.808 ;
      RECT 52.395 1.642 52.42 1.781 ;
      RECT 52.39 1.635 52.395 1.776 ;
      RECT 52.375 1.635 52.39 1.774 ;
      RECT 52.35 1.627 52.375 1.77 ;
      RECT 52.335 1.625 52.35 1.766 ;
      RECT 52.305 1.625 52.335 1.763 ;
      RECT 52.295 1.625 52.305 1.758 ;
      RECT 52.25 1.625 52.295 1.756 ;
      RECT 52.221 1.625 52.25 1.757 ;
      RECT 52.135 1.625 52.221 1.759 ;
      RECT 52.121 1.626 52.135 1.761 ;
      RECT 52.035 1.627 52.121 1.763 ;
      RECT 52.02 1.628 52.035 1.773 ;
      RECT 52.015 1.629 52.02 1.782 ;
      RECT 51.995 1.632 52.015 1.792 ;
      RECT 51.98 1.64 51.995 1.807 ;
      RECT 51.96 1.658 51.98 1.822 ;
      RECT 51.95 1.67 51.96 1.845 ;
      RECT 51.94 1.679 51.95 1.875 ;
      RECT 51.925 1.691 51.94 1.92 ;
      RECT 51.87 1.724 51.925 2.235 ;
      RECT 51.865 1.752 51.87 2.235 ;
      RECT 51.845 1.767 51.865 2.235 ;
      RECT 51.81 1.827 51.845 2.235 ;
      RECT 51.808 1.877 51.81 2.235 ;
      RECT 51.805 1.885 51.808 2.235 ;
      RECT 51.795 1.9 51.805 2.235 ;
      RECT 51.79 1.912 51.795 2.235 ;
      RECT 51.78 1.937 51.79 2.235 ;
      RECT 51.77 1.965 51.78 2.235 ;
      RECT 49.675 3.47 49.725 3.73 ;
      RECT 52.585 3.02 52.645 3.28 ;
      RECT 52.57 3.02 52.585 3.29 ;
      RECT 52.551 3.02 52.57 3.323 ;
      RECT 52.465 3.02 52.551 3.448 ;
      RECT 52.385 3.02 52.465 3.63 ;
      RECT 52.38 3.257 52.385 3.715 ;
      RECT 52.355 3.327 52.38 3.743 ;
      RECT 52.35 3.397 52.355 3.77 ;
      RECT 52.33 3.469 52.35 3.792 ;
      RECT 52.325 3.536 52.33 3.815 ;
      RECT 52.315 3.565 52.325 3.83 ;
      RECT 52.305 3.587 52.315 3.847 ;
      RECT 52.3 3.597 52.305 3.858 ;
      RECT 52.295 3.605 52.3 3.866 ;
      RECT 52.285 3.613 52.295 3.878 ;
      RECT 52.28 3.625 52.285 3.888 ;
      RECT 52.275 3.633 52.28 3.893 ;
      RECT 52.255 3.651 52.275 3.903 ;
      RECT 52.25 3.668 52.255 3.91 ;
      RECT 52.245 3.676 52.25 3.911 ;
      RECT 52.24 3.687 52.245 3.913 ;
      RECT 52.2 3.725 52.24 3.923 ;
      RECT 52.195 3.76 52.2 3.934 ;
      RECT 52.19 3.765 52.195 3.937 ;
      RECT 52.165 3.775 52.19 3.944 ;
      RECT 52.155 3.789 52.165 3.953 ;
      RECT 52.135 3.801 52.155 3.956 ;
      RECT 52.085 3.82 52.135 3.96 ;
      RECT 52.04 3.835 52.085 3.965 ;
      RECT 51.975 3.838 52.04 3.971 ;
      RECT 51.96 3.836 51.975 3.978 ;
      RECT 51.93 3.835 51.96 3.978 ;
      RECT 51.891 3.834 51.93 3.974 ;
      RECT 51.805 3.831 51.891 3.97 ;
      RECT 51.788 3.829 51.805 3.967 ;
      RECT 51.702 3.827 51.788 3.964 ;
      RECT 51.616 3.824 51.702 3.958 ;
      RECT 51.53 3.82 51.616 3.953 ;
      RECT 51.452 3.817 51.53 3.949 ;
      RECT 51.366 3.814 51.452 3.947 ;
      RECT 51.28 3.811 51.366 3.944 ;
      RECT 51.222 3.809 51.28 3.941 ;
      RECT 51.136 3.806 51.222 3.939 ;
      RECT 51.05 3.802 51.136 3.937 ;
      RECT 50.964 3.799 51.05 3.934 ;
      RECT 50.878 3.795 50.964 3.932 ;
      RECT 50.792 3.791 50.878 3.929 ;
      RECT 50.706 3.788 50.792 3.927 ;
      RECT 50.62 3.784 50.706 3.924 ;
      RECT 50.534 3.781 50.62 3.922 ;
      RECT 50.448 3.777 50.534 3.919 ;
      RECT 50.362 3.774 50.448 3.917 ;
      RECT 50.276 3.77 50.362 3.914 ;
      RECT 50.19 3.767 50.276 3.912 ;
      RECT 50.18 3.765 50.19 3.908 ;
      RECT 50.175 3.765 50.18 3.906 ;
      RECT 50.135 3.76 50.175 3.9 ;
      RECT 50.121 3.751 50.135 3.893 ;
      RECT 50.035 3.721 50.121 3.878 ;
      RECT 50.015 3.687 50.035 3.863 ;
      RECT 49.945 3.656 50.015 3.85 ;
      RECT 49.94 3.631 49.945 3.839 ;
      RECT 49.935 3.625 49.94 3.837 ;
      RECT 49.866 3.47 49.935 3.825 ;
      RECT 49.78 3.47 49.866 3.799 ;
      RECT 49.755 3.47 49.78 3.778 ;
      RECT 49.75 3.47 49.755 3.768 ;
      RECT 49.745 3.47 49.75 3.76 ;
      RECT 49.725 3.47 49.745 3.743 ;
      RECT 52.145 2.04 52.405 2.3 ;
      RECT 52.13 2.04 52.405 2.203 ;
      RECT 52.1 2.04 52.405 2.178 ;
      RECT 52.065 1.88 52.345 2.16 ;
      RECT 52.035 3.37 52.095 3.63 ;
      RECT 51.06 2.06 51.115 2.32 ;
      RECT 51.995 3.327 52.035 3.63 ;
      RECT 51.966 3.248 51.995 3.63 ;
      RECT 51.88 3.12 51.966 3.63 ;
      RECT 51.86 3 51.88 3.63 ;
      RECT 51.835 2.951 51.86 3.63 ;
      RECT 51.83 2.916 51.835 3.48 ;
      RECT 51.8 2.876 51.83 3.418 ;
      RECT 51.775 2.813 51.8 3.333 ;
      RECT 51.765 2.775 51.775 3.27 ;
      RECT 51.75 2.75 51.765 3.231 ;
      RECT 51.707 2.708 51.75 3.137 ;
      RECT 51.705 2.681 51.707 3.064 ;
      RECT 51.7 2.676 51.705 3.055 ;
      RECT 51.695 2.669 51.7 3.03 ;
      RECT 51.69 2.663 51.695 3.015 ;
      RECT 51.685 2.657 51.69 3.003 ;
      RECT 51.675 2.648 51.685 2.985 ;
      RECT 51.67 2.639 51.675 2.963 ;
      RECT 51.645 2.62 51.67 2.913 ;
      RECT 51.64 2.601 51.645 2.863 ;
      RECT 51.625 2.587 51.64 2.823 ;
      RECT 51.62 2.573 51.625 2.79 ;
      RECT 51.615 2.566 51.62 2.783 ;
      RECT 51.6 2.553 51.615 2.775 ;
      RECT 51.555 2.515 51.6 2.748 ;
      RECT 51.525 2.468 51.555 2.713 ;
      RECT 51.505 2.437 51.525 2.69 ;
      RECT 51.425 2.37 51.505 2.643 ;
      RECT 51.395 2.3 51.425 2.59 ;
      RECT 51.39 2.277 51.395 2.573 ;
      RECT 51.36 2.255 51.39 2.558 ;
      RECT 51.33 2.214 51.36 2.53 ;
      RECT 51.325 2.189 51.33 2.515 ;
      RECT 51.32 2.183 51.325 2.508 ;
      RECT 51.31 2.06 51.32 2.5 ;
      RECT 51.3 2.06 51.31 2.493 ;
      RECT 51.295 2.06 51.3 2.485 ;
      RECT 51.275 2.06 51.295 2.473 ;
      RECT 51.225 2.06 51.275 2.443 ;
      RECT 51.17 2.06 51.225 2.393 ;
      RECT 51.14 2.06 51.17 2.353 ;
      RECT 51.115 2.06 51.14 2.33 ;
      RECT 50.985 2.785 51.265 3.065 ;
      RECT 50.95 2.7 51.21 2.96 ;
      RECT 50.95 2.782 51.22 2.96 ;
      RECT 49.15 2.155 49.155 2.64 ;
      RECT 49.04 2.34 49.045 2.64 ;
      RECT 48.95 2.38 49.015 2.64 ;
      RECT 50.625 1.88 50.715 2.51 ;
      RECT 50.59 1.93 50.595 2.51 ;
      RECT 50.535 1.955 50.545 2.51 ;
      RECT 50.49 1.955 50.5 2.51 ;
      RECT 50.86 1.88 50.905 2.16 ;
      RECT 49.71 1.61 49.91 1.75 ;
      RECT 50.826 1.88 50.86 2.172 ;
      RECT 50.74 1.88 50.826 2.212 ;
      RECT 50.725 1.88 50.74 2.253 ;
      RECT 50.72 1.88 50.725 2.273 ;
      RECT 50.715 1.88 50.72 2.293 ;
      RECT 50.595 1.922 50.625 2.51 ;
      RECT 50.545 1.942 50.59 2.51 ;
      RECT 50.53 1.957 50.535 2.51 ;
      RECT 50.5 1.957 50.53 2.51 ;
      RECT 50.455 1.942 50.49 2.51 ;
      RECT 50.45 1.93 50.455 2.29 ;
      RECT 50.445 1.927 50.45 2.27 ;
      RECT 50.43 1.917 50.445 2.223 ;
      RECT 50.425 1.91 50.43 2.186 ;
      RECT 50.42 1.907 50.425 2.169 ;
      RECT 50.405 1.897 50.42 2.125 ;
      RECT 50.4 1.888 50.405 2.085 ;
      RECT 50.395 1.884 50.4 2.07 ;
      RECT 50.385 1.878 50.395 2.053 ;
      RECT 50.345 1.859 50.385 2.028 ;
      RECT 50.34 1.841 50.345 2.008 ;
      RECT 50.33 1.835 50.34 2.003 ;
      RECT 50.3 1.819 50.33 1.99 ;
      RECT 50.285 1.801 50.3 1.973 ;
      RECT 50.27 1.789 50.285 1.96 ;
      RECT 50.265 1.781 50.27 1.953 ;
      RECT 50.235 1.767 50.265 1.94 ;
      RECT 50.23 1.752 50.235 1.928 ;
      RECT 50.22 1.746 50.23 1.92 ;
      RECT 50.2 1.734 50.22 1.908 ;
      RECT 50.19 1.722 50.2 1.895 ;
      RECT 50.16 1.706 50.19 1.88 ;
      RECT 50.14 1.686 50.16 1.863 ;
      RECT 50.135 1.676 50.14 1.853 ;
      RECT 50.11 1.664 50.135 1.84 ;
      RECT 50.105 1.652 50.11 1.828 ;
      RECT 50.1 1.647 50.105 1.824 ;
      RECT 50.085 1.64 50.1 1.816 ;
      RECT 50.075 1.627 50.085 1.806 ;
      RECT 50.07 1.625 50.075 1.8 ;
      RECT 50.045 1.618 50.07 1.789 ;
      RECT 50.04 1.611 50.045 1.778 ;
      RECT 50.015 1.61 50.04 1.765 ;
      RECT 49.996 1.61 50.015 1.755 ;
      RECT 49.91 1.61 49.996 1.752 ;
      RECT 49.68 1.61 49.71 1.755 ;
      RECT 49.64 1.617 49.68 1.768 ;
      RECT 49.615 1.627 49.64 1.781 ;
      RECT 49.6 1.636 49.615 1.791 ;
      RECT 49.57 1.641 49.6 1.81 ;
      RECT 49.565 1.647 49.57 1.828 ;
      RECT 49.545 1.657 49.565 1.843 ;
      RECT 49.535 1.67 49.545 1.863 ;
      RECT 49.52 1.682 49.535 1.88 ;
      RECT 49.515 1.692 49.52 1.89 ;
      RECT 49.51 1.697 49.515 1.895 ;
      RECT 49.5 1.705 49.51 1.908 ;
      RECT 49.45 1.737 49.5 1.945 ;
      RECT 49.435 1.772 49.45 1.986 ;
      RECT 49.43 1.782 49.435 2.001 ;
      RECT 49.425 1.787 49.43 2.008 ;
      RECT 49.4 1.803 49.425 2.028 ;
      RECT 49.385 1.824 49.4 2.053 ;
      RECT 49.36 1.845 49.385 2.078 ;
      RECT 49.35 1.864 49.36 2.101 ;
      RECT 49.325 1.882 49.35 2.124 ;
      RECT 49.31 1.902 49.325 2.148 ;
      RECT 49.305 1.912 49.31 2.16 ;
      RECT 49.29 1.924 49.305 2.18 ;
      RECT 49.28 1.939 49.29 2.22 ;
      RECT 49.275 1.947 49.28 2.248 ;
      RECT 49.265 1.957 49.275 2.268 ;
      RECT 49.26 1.97 49.265 2.293 ;
      RECT 49.255 1.983 49.26 2.313 ;
      RECT 49.25 1.989 49.255 2.335 ;
      RECT 49.24 1.998 49.25 2.355 ;
      RECT 49.235 2.018 49.24 2.378 ;
      RECT 49.23 2.024 49.235 2.398 ;
      RECT 49.225 2.031 49.23 2.42 ;
      RECT 49.22 2.042 49.225 2.433 ;
      RECT 49.21 2.052 49.22 2.458 ;
      RECT 49.19 2.077 49.21 2.64 ;
      RECT 49.16 2.117 49.19 2.64 ;
      RECT 49.155 2.147 49.16 2.64 ;
      RECT 49.13 2.175 49.15 2.64 ;
      RECT 49.1 2.22 49.13 2.64 ;
      RECT 49.095 2.247 49.1 2.64 ;
      RECT 49.075 2.265 49.095 2.64 ;
      RECT 49.065 2.29 49.075 2.64 ;
      RECT 49.06 2.302 49.065 2.64 ;
      RECT 49.045 2.325 49.06 2.64 ;
      RECT 49.025 2.352 49.04 2.64 ;
      RECT 49.015 2.375 49.025 2.64 ;
      RECT 50.805 3.26 50.885 3.52 ;
      RECT 50.04 2.48 50.11 2.74 ;
      RECT 50.771 3.227 50.805 3.52 ;
      RECT 50.685 3.13 50.771 3.52 ;
      RECT 50.665 3.042 50.685 3.52 ;
      RECT 50.655 3.012 50.665 3.52 ;
      RECT 50.645 2.992 50.655 3.52 ;
      RECT 50.625 2.979 50.645 3.52 ;
      RECT 50.61 2.969 50.625 3.348 ;
      RECT 50.605 2.962 50.61 3.303 ;
      RECT 50.595 2.956 50.605 3.293 ;
      RECT 50.585 2.948 50.595 3.275 ;
      RECT 50.58 2.942 50.585 3.263 ;
      RECT 50.57 2.937 50.58 3.25 ;
      RECT 50.55 2.927 50.57 3.223 ;
      RECT 50.51 2.906 50.55 3.175 ;
      RECT 50.495 2.887 50.51 3.133 ;
      RECT 50.47 2.873 50.495 3.103 ;
      RECT 50.46 2.861 50.47 3.07 ;
      RECT 50.455 2.856 50.46 3.06 ;
      RECT 50.425 2.842 50.455 3.04 ;
      RECT 50.415 2.826 50.425 3.013 ;
      RECT 50.41 2.821 50.415 3.003 ;
      RECT 50.385 2.812 50.41 2.983 ;
      RECT 50.375 2.8 50.385 2.963 ;
      RECT 50.305 2.768 50.375 2.938 ;
      RECT 50.3 2.737 50.305 2.915 ;
      RECT 50.251 2.48 50.3 2.898 ;
      RECT 50.165 2.48 50.251 2.857 ;
      RECT 50.11 2.48 50.165 2.785 ;
      RECT 50.2 3.265 50.36 3.525 ;
      RECT 49.725 1.88 49.775 2.565 ;
      RECT 49.515 2.305 49.55 2.565 ;
      RECT 49.83 1.88 49.835 2.34 ;
      RECT 49.92 1.88 49.945 2.16 ;
      RECT 50.195 3.262 50.2 3.525 ;
      RECT 50.16 3.25 50.195 3.525 ;
      RECT 50.1 3.223 50.16 3.525 ;
      RECT 50.095 3.206 50.1 3.379 ;
      RECT 50.09 3.203 50.095 3.366 ;
      RECT 50.07 3.196 50.09 3.353 ;
      RECT 50.035 3.179 50.07 3.335 ;
      RECT 49.995 3.158 50.035 3.315 ;
      RECT 49.99 3.146 49.995 3.303 ;
      RECT 49.95 3.132 49.99 3.289 ;
      RECT 49.93 3.115 49.95 3.271 ;
      RECT 49.92 3.107 49.93 3.263 ;
      RECT 49.905 1.88 49.92 2.178 ;
      RECT 49.89 3.097 49.92 3.25 ;
      RECT 49.875 1.88 49.905 2.223 ;
      RECT 49.88 3.087 49.89 3.237 ;
      RECT 49.85 3.072 49.88 3.224 ;
      RECT 49.835 1.88 49.875 2.29 ;
      RECT 49.835 3.04 49.85 3.21 ;
      RECT 49.83 3.012 49.835 3.204 ;
      RECT 49.825 1.88 49.83 2.345 ;
      RECT 49.815 2.982 49.83 3.198 ;
      RECT 49.82 1.88 49.825 2.358 ;
      RECT 49.81 1.88 49.82 2.378 ;
      RECT 49.775 2.895 49.815 3.183 ;
      RECT 49.775 1.88 49.81 2.418 ;
      RECT 49.77 2.827 49.775 3.171 ;
      RECT 49.755 2.782 49.77 3.166 ;
      RECT 49.75 2.72 49.755 3.161 ;
      RECT 49.725 2.627 49.75 3.154 ;
      RECT 49.72 1.88 49.725 3.146 ;
      RECT 49.705 1.88 49.72 3.133 ;
      RECT 49.685 1.88 49.705 3.09 ;
      RECT 49.675 1.88 49.685 3.04 ;
      RECT 49.67 1.88 49.675 3.013 ;
      RECT 49.665 1.88 49.67 2.991 ;
      RECT 49.66 2.106 49.665 2.974 ;
      RECT 49.655 2.128 49.66 2.952 ;
      RECT 49.65 2.17 49.655 2.935 ;
      RECT 49.62 2.22 49.65 2.879 ;
      RECT 49.615 2.247 49.62 2.821 ;
      RECT 49.6 2.265 49.615 2.785 ;
      RECT 49.595 2.283 49.6 2.749 ;
      RECT 49.589 2.29 49.595 2.73 ;
      RECT 49.585 2.297 49.589 2.713 ;
      RECT 49.58 2.302 49.585 2.682 ;
      RECT 49.57 2.305 49.58 2.657 ;
      RECT 49.56 2.305 49.57 2.623 ;
      RECT 49.555 2.305 49.56 2.6 ;
      RECT 49.55 2.305 49.555 2.58 ;
      RECT 48.465 2.44 48.745 2.72 ;
      RECT 48.465 2.44 48.765 2.615 ;
      RECT 48.555 2.33 48.815 2.59 ;
      RECT 48.52 2.425 48.815 2.59 ;
      RECT 48.645 0.945 48.81 2.59 ;
      RECT 48.545 0.945 48.915 1.315 ;
      RECT 48.17 3.47 48.43 3.73 ;
      RECT 48.19 3.397 48.37 3.73 ;
      RECT 48.19 3.14 48.365 3.73 ;
      RECT 48.19 2.932 48.355 3.73 ;
      RECT 48.195 2.85 48.355 3.73 ;
      RECT 48.195 2.615 48.345 3.73 ;
      RECT 48.195 2.462 48.34 3.73 ;
      RECT 48.2 2.447 48.34 3.73 ;
      RECT 48.25 2.162 48.34 3.73 ;
      RECT 48.205 2.397 48.34 3.73 ;
      RECT 48.235 2.215 48.34 3.73 ;
      RECT 48.22 2.327 48.34 3.73 ;
      RECT 48.225 2.285 48.34 3.73 ;
      RECT 48.22 2.327 48.355 2.39 ;
      RECT 48.255 1.915 48.36 2.335 ;
      RECT 48.255 1.915 48.375 2.318 ;
      RECT 48.255 1.915 48.41 2.28 ;
      RECT 48.25 2.162 48.46 2.213 ;
      RECT 48.255 1.915 48.515 2.175 ;
      RECT 47.515 2.62 47.775 2.88 ;
      RECT 47.515 2.62 47.785 2.838 ;
      RECT 47.515 2.62 47.871 2.809 ;
      RECT 47.515 2.62 47.94 2.761 ;
      RECT 47.515 2.62 47.975 2.73 ;
      RECT 47.745 2.44 48.025 2.72 ;
      RECT 47.58 2.605 48.025 2.72 ;
      RECT 47.67 2.482 47.775 2.88 ;
      RECT 47.6 2.545 48.025 2.72 ;
      RECT 42.05 6.22 42.37 6.545 ;
      RECT 42.08 5.695 42.25 6.545 ;
      RECT 42.08 5.695 42.255 6.045 ;
      RECT 42.08 5.695 43.055 5.87 ;
      RECT 42.88 1.965 43.055 5.87 ;
      RECT 42.825 1.965 43.175 2.315 ;
      RECT 42.85 6.655 43.175 6.98 ;
      RECT 41.735 6.745 43.175 6.915 ;
      RECT 41.735 2.395 41.895 6.915 ;
      RECT 42.05 2.365 42.37 2.685 ;
      RECT 41.735 2.395 42.37 2.565 ;
      RECT 41 5.86 41.34 6.21 ;
      RECT 41.08 2.705 41.255 6.21 ;
      RECT 41.005 2.705 41.345 3.055 ;
      RECT 40.4 2.705 40.785 3.055 ;
      RECT 40.39 2.77 40.785 2.97 ;
      RECT 40.535 2.7 40.705 3.055 ;
      RECT 38.845 2.44 39.125 2.72 ;
      RECT 38.84 2.44 39.125 2.673 ;
      RECT 38.82 2.44 39.125 2.65 ;
      RECT 38.81 2.44 39.125 2.63 ;
      RECT 38.8 2.44 39.125 2.615 ;
      RECT 38.775 2.44 39.125 2.588 ;
      RECT 38.765 2.44 39.125 2.563 ;
      RECT 38.72 2.295 39 2.555 ;
      RECT 38.72 2.39 39.1 2.555 ;
      RECT 38.72 2.335 39.045 2.555 ;
      RECT 38.72 2.327 39.04 2.555 ;
      RECT 38.72 2.317 39.035 2.555 ;
      RECT 38.72 2.305 39.03 2.555 ;
      RECT 37.645 3 37.925 3.28 ;
      RECT 37.645 3 37.96 3.26 ;
      RECT 29.97 6.66 30.32 7.01 ;
      RECT 37.39 6.615 37.74 6.965 ;
      RECT 29.97 6.69 37.74 6.89 ;
      RECT 37.68 2.42 37.73 2.68 ;
      RECT 37.47 2.42 37.475 2.68 ;
      RECT 36.665 1.975 36.695 2.235 ;
      RECT 36.435 1.975 36.51 2.235 ;
      RECT 37.655 2.37 37.68 2.68 ;
      RECT 37.65 2.327 37.655 2.68 ;
      RECT 37.645 2.31 37.65 2.68 ;
      RECT 37.64 2.297 37.645 2.68 ;
      RECT 37.565 2.18 37.64 2.68 ;
      RECT 37.52 1.997 37.565 2.68 ;
      RECT 37.515 1.925 37.52 2.68 ;
      RECT 37.5 1.9 37.515 2.68 ;
      RECT 37.475 1.862 37.5 2.68 ;
      RECT 37.465 1.842 37.475 2.402 ;
      RECT 37.45 1.834 37.465 2.357 ;
      RECT 37.445 1.826 37.45 2.328 ;
      RECT 37.44 1.823 37.445 2.308 ;
      RECT 37.435 1.82 37.44 2.288 ;
      RECT 37.43 1.817 37.435 2.268 ;
      RECT 37.4 1.806 37.43 2.205 ;
      RECT 37.38 1.791 37.4 2.12 ;
      RECT 37.375 1.783 37.38 2.083 ;
      RECT 37.365 1.777 37.375 2.05 ;
      RECT 37.35 1.769 37.365 2.01 ;
      RECT 37.345 1.762 37.35 1.97 ;
      RECT 37.34 1.759 37.345 1.948 ;
      RECT 37.335 1.756 37.34 1.935 ;
      RECT 37.33 1.755 37.335 1.925 ;
      RECT 37.315 1.749 37.33 1.915 ;
      RECT 37.29 1.736 37.315 1.9 ;
      RECT 37.24 1.711 37.29 1.871 ;
      RECT 37.225 1.69 37.24 1.846 ;
      RECT 37.215 1.683 37.225 1.835 ;
      RECT 37.16 1.664 37.215 1.808 ;
      RECT 37.135 1.642 37.16 1.781 ;
      RECT 37.13 1.635 37.135 1.776 ;
      RECT 37.115 1.635 37.13 1.774 ;
      RECT 37.09 1.627 37.115 1.77 ;
      RECT 37.075 1.625 37.09 1.766 ;
      RECT 37.045 1.625 37.075 1.763 ;
      RECT 37.035 1.625 37.045 1.758 ;
      RECT 36.99 1.625 37.035 1.756 ;
      RECT 36.961 1.625 36.99 1.757 ;
      RECT 36.875 1.625 36.961 1.759 ;
      RECT 36.861 1.626 36.875 1.761 ;
      RECT 36.775 1.627 36.861 1.763 ;
      RECT 36.76 1.628 36.775 1.773 ;
      RECT 36.755 1.629 36.76 1.782 ;
      RECT 36.735 1.632 36.755 1.792 ;
      RECT 36.72 1.64 36.735 1.807 ;
      RECT 36.7 1.658 36.72 1.822 ;
      RECT 36.69 1.67 36.7 1.845 ;
      RECT 36.68 1.679 36.69 1.875 ;
      RECT 36.665 1.691 36.68 1.92 ;
      RECT 36.61 1.724 36.665 2.235 ;
      RECT 36.605 1.752 36.61 2.235 ;
      RECT 36.585 1.767 36.605 2.235 ;
      RECT 36.55 1.827 36.585 2.235 ;
      RECT 36.548 1.877 36.55 2.235 ;
      RECT 36.545 1.885 36.548 2.235 ;
      RECT 36.535 1.9 36.545 2.235 ;
      RECT 36.53 1.912 36.535 2.235 ;
      RECT 36.52 1.937 36.53 2.235 ;
      RECT 36.51 1.965 36.52 2.235 ;
      RECT 34.415 3.47 34.465 3.73 ;
      RECT 37.325 3.02 37.385 3.28 ;
      RECT 37.31 3.02 37.325 3.29 ;
      RECT 37.291 3.02 37.31 3.323 ;
      RECT 37.205 3.02 37.291 3.448 ;
      RECT 37.125 3.02 37.205 3.63 ;
      RECT 37.12 3.257 37.125 3.715 ;
      RECT 37.095 3.327 37.12 3.743 ;
      RECT 37.09 3.397 37.095 3.77 ;
      RECT 37.07 3.469 37.09 3.792 ;
      RECT 37.065 3.536 37.07 3.815 ;
      RECT 37.055 3.565 37.065 3.83 ;
      RECT 37.045 3.587 37.055 3.847 ;
      RECT 37.04 3.597 37.045 3.858 ;
      RECT 37.035 3.605 37.04 3.866 ;
      RECT 37.025 3.613 37.035 3.878 ;
      RECT 37.02 3.625 37.025 3.888 ;
      RECT 37.015 3.633 37.02 3.893 ;
      RECT 36.995 3.651 37.015 3.903 ;
      RECT 36.99 3.668 36.995 3.91 ;
      RECT 36.985 3.676 36.99 3.911 ;
      RECT 36.98 3.687 36.985 3.913 ;
      RECT 36.94 3.725 36.98 3.923 ;
      RECT 36.935 3.76 36.94 3.934 ;
      RECT 36.93 3.765 36.935 3.937 ;
      RECT 36.905 3.775 36.93 3.944 ;
      RECT 36.895 3.789 36.905 3.953 ;
      RECT 36.875 3.801 36.895 3.956 ;
      RECT 36.825 3.82 36.875 3.96 ;
      RECT 36.78 3.835 36.825 3.965 ;
      RECT 36.715 3.838 36.78 3.971 ;
      RECT 36.7 3.836 36.715 3.978 ;
      RECT 36.67 3.835 36.7 3.978 ;
      RECT 36.631 3.834 36.67 3.974 ;
      RECT 36.545 3.831 36.631 3.97 ;
      RECT 36.528 3.829 36.545 3.967 ;
      RECT 36.442 3.827 36.528 3.964 ;
      RECT 36.356 3.824 36.442 3.958 ;
      RECT 36.27 3.82 36.356 3.953 ;
      RECT 36.192 3.817 36.27 3.949 ;
      RECT 36.106 3.814 36.192 3.947 ;
      RECT 36.02 3.811 36.106 3.944 ;
      RECT 35.962 3.809 36.02 3.941 ;
      RECT 35.876 3.806 35.962 3.939 ;
      RECT 35.79 3.802 35.876 3.937 ;
      RECT 35.704 3.799 35.79 3.934 ;
      RECT 35.618 3.795 35.704 3.932 ;
      RECT 35.532 3.791 35.618 3.929 ;
      RECT 35.446 3.788 35.532 3.927 ;
      RECT 35.36 3.784 35.446 3.924 ;
      RECT 35.274 3.781 35.36 3.922 ;
      RECT 35.188 3.777 35.274 3.919 ;
      RECT 35.102 3.774 35.188 3.917 ;
      RECT 35.016 3.77 35.102 3.914 ;
      RECT 34.93 3.767 35.016 3.912 ;
      RECT 34.92 3.765 34.93 3.908 ;
      RECT 34.915 3.765 34.92 3.906 ;
      RECT 34.875 3.76 34.915 3.9 ;
      RECT 34.861 3.751 34.875 3.893 ;
      RECT 34.775 3.721 34.861 3.878 ;
      RECT 34.755 3.687 34.775 3.863 ;
      RECT 34.685 3.656 34.755 3.85 ;
      RECT 34.68 3.631 34.685 3.839 ;
      RECT 34.675 3.625 34.68 3.837 ;
      RECT 34.606 3.47 34.675 3.825 ;
      RECT 34.52 3.47 34.606 3.799 ;
      RECT 34.495 3.47 34.52 3.778 ;
      RECT 34.49 3.47 34.495 3.768 ;
      RECT 34.485 3.47 34.49 3.76 ;
      RECT 34.465 3.47 34.485 3.743 ;
      RECT 36.885 2.04 37.145 2.3 ;
      RECT 36.87 2.04 37.145 2.203 ;
      RECT 36.84 2.04 37.145 2.178 ;
      RECT 36.805 1.88 37.085 2.16 ;
      RECT 36.775 3.37 36.835 3.63 ;
      RECT 35.8 2.06 35.855 2.32 ;
      RECT 36.735 3.327 36.775 3.63 ;
      RECT 36.706 3.248 36.735 3.63 ;
      RECT 36.62 3.12 36.706 3.63 ;
      RECT 36.6 3 36.62 3.63 ;
      RECT 36.575 2.951 36.6 3.63 ;
      RECT 36.57 2.916 36.575 3.48 ;
      RECT 36.54 2.876 36.57 3.418 ;
      RECT 36.515 2.813 36.54 3.333 ;
      RECT 36.505 2.775 36.515 3.27 ;
      RECT 36.49 2.75 36.505 3.231 ;
      RECT 36.447 2.708 36.49 3.137 ;
      RECT 36.445 2.681 36.447 3.064 ;
      RECT 36.44 2.676 36.445 3.055 ;
      RECT 36.435 2.669 36.44 3.03 ;
      RECT 36.43 2.663 36.435 3.015 ;
      RECT 36.425 2.657 36.43 3.003 ;
      RECT 36.415 2.648 36.425 2.985 ;
      RECT 36.41 2.639 36.415 2.963 ;
      RECT 36.385 2.62 36.41 2.913 ;
      RECT 36.38 2.601 36.385 2.863 ;
      RECT 36.365 2.587 36.38 2.823 ;
      RECT 36.36 2.573 36.365 2.79 ;
      RECT 36.355 2.566 36.36 2.783 ;
      RECT 36.34 2.553 36.355 2.775 ;
      RECT 36.295 2.515 36.34 2.748 ;
      RECT 36.265 2.468 36.295 2.713 ;
      RECT 36.245 2.437 36.265 2.69 ;
      RECT 36.165 2.37 36.245 2.643 ;
      RECT 36.135 2.3 36.165 2.59 ;
      RECT 36.13 2.277 36.135 2.573 ;
      RECT 36.1 2.255 36.13 2.558 ;
      RECT 36.07 2.214 36.1 2.53 ;
      RECT 36.065 2.189 36.07 2.515 ;
      RECT 36.06 2.183 36.065 2.508 ;
      RECT 36.05 2.06 36.06 2.5 ;
      RECT 36.04 2.06 36.05 2.493 ;
      RECT 36.035 2.06 36.04 2.485 ;
      RECT 36.015 2.06 36.035 2.473 ;
      RECT 35.965 2.06 36.015 2.443 ;
      RECT 35.91 2.06 35.965 2.393 ;
      RECT 35.88 2.06 35.91 2.353 ;
      RECT 35.855 2.06 35.88 2.33 ;
      RECT 35.725 2.785 36.005 3.065 ;
      RECT 35.69 2.7 35.95 2.96 ;
      RECT 35.69 2.782 35.96 2.96 ;
      RECT 33.89 2.155 33.895 2.64 ;
      RECT 33.78 2.34 33.785 2.64 ;
      RECT 33.69 2.38 33.755 2.64 ;
      RECT 35.365 1.88 35.455 2.51 ;
      RECT 35.33 1.93 35.335 2.51 ;
      RECT 35.275 1.955 35.285 2.51 ;
      RECT 35.23 1.955 35.24 2.51 ;
      RECT 35.6 1.88 35.645 2.16 ;
      RECT 34.45 1.61 34.65 1.75 ;
      RECT 35.566 1.88 35.6 2.172 ;
      RECT 35.48 1.88 35.566 2.212 ;
      RECT 35.465 1.88 35.48 2.253 ;
      RECT 35.46 1.88 35.465 2.273 ;
      RECT 35.455 1.88 35.46 2.293 ;
      RECT 35.335 1.922 35.365 2.51 ;
      RECT 35.285 1.942 35.33 2.51 ;
      RECT 35.27 1.957 35.275 2.51 ;
      RECT 35.24 1.957 35.27 2.51 ;
      RECT 35.195 1.942 35.23 2.51 ;
      RECT 35.19 1.93 35.195 2.29 ;
      RECT 35.185 1.927 35.19 2.27 ;
      RECT 35.17 1.917 35.185 2.223 ;
      RECT 35.165 1.91 35.17 2.186 ;
      RECT 35.16 1.907 35.165 2.169 ;
      RECT 35.145 1.897 35.16 2.125 ;
      RECT 35.14 1.888 35.145 2.085 ;
      RECT 35.135 1.884 35.14 2.07 ;
      RECT 35.125 1.878 35.135 2.053 ;
      RECT 35.085 1.859 35.125 2.028 ;
      RECT 35.08 1.841 35.085 2.008 ;
      RECT 35.07 1.835 35.08 2.003 ;
      RECT 35.04 1.819 35.07 1.99 ;
      RECT 35.025 1.801 35.04 1.973 ;
      RECT 35.01 1.789 35.025 1.96 ;
      RECT 35.005 1.781 35.01 1.953 ;
      RECT 34.975 1.767 35.005 1.94 ;
      RECT 34.97 1.752 34.975 1.928 ;
      RECT 34.96 1.746 34.97 1.92 ;
      RECT 34.94 1.734 34.96 1.908 ;
      RECT 34.93 1.722 34.94 1.895 ;
      RECT 34.9 1.706 34.93 1.88 ;
      RECT 34.88 1.686 34.9 1.863 ;
      RECT 34.875 1.676 34.88 1.853 ;
      RECT 34.85 1.664 34.875 1.84 ;
      RECT 34.845 1.652 34.85 1.828 ;
      RECT 34.84 1.647 34.845 1.824 ;
      RECT 34.825 1.64 34.84 1.816 ;
      RECT 34.815 1.627 34.825 1.806 ;
      RECT 34.81 1.625 34.815 1.8 ;
      RECT 34.785 1.618 34.81 1.789 ;
      RECT 34.78 1.611 34.785 1.778 ;
      RECT 34.755 1.61 34.78 1.765 ;
      RECT 34.736 1.61 34.755 1.755 ;
      RECT 34.65 1.61 34.736 1.752 ;
      RECT 34.42 1.61 34.45 1.755 ;
      RECT 34.38 1.617 34.42 1.768 ;
      RECT 34.355 1.627 34.38 1.781 ;
      RECT 34.34 1.636 34.355 1.791 ;
      RECT 34.31 1.641 34.34 1.81 ;
      RECT 34.305 1.647 34.31 1.828 ;
      RECT 34.285 1.657 34.305 1.843 ;
      RECT 34.275 1.67 34.285 1.863 ;
      RECT 34.26 1.682 34.275 1.88 ;
      RECT 34.255 1.692 34.26 1.89 ;
      RECT 34.25 1.697 34.255 1.895 ;
      RECT 34.24 1.705 34.25 1.908 ;
      RECT 34.19 1.737 34.24 1.945 ;
      RECT 34.175 1.772 34.19 1.986 ;
      RECT 34.17 1.782 34.175 2.001 ;
      RECT 34.165 1.787 34.17 2.008 ;
      RECT 34.14 1.803 34.165 2.028 ;
      RECT 34.125 1.824 34.14 2.053 ;
      RECT 34.1 1.845 34.125 2.078 ;
      RECT 34.09 1.864 34.1 2.101 ;
      RECT 34.065 1.882 34.09 2.124 ;
      RECT 34.05 1.902 34.065 2.148 ;
      RECT 34.045 1.912 34.05 2.16 ;
      RECT 34.03 1.924 34.045 2.18 ;
      RECT 34.02 1.939 34.03 2.22 ;
      RECT 34.015 1.947 34.02 2.248 ;
      RECT 34.005 1.957 34.015 2.268 ;
      RECT 34 1.97 34.005 2.293 ;
      RECT 33.995 1.983 34 2.313 ;
      RECT 33.99 1.989 33.995 2.335 ;
      RECT 33.98 1.998 33.99 2.355 ;
      RECT 33.975 2.018 33.98 2.378 ;
      RECT 33.97 2.024 33.975 2.398 ;
      RECT 33.965 2.031 33.97 2.42 ;
      RECT 33.96 2.042 33.965 2.433 ;
      RECT 33.95 2.052 33.96 2.458 ;
      RECT 33.93 2.077 33.95 2.64 ;
      RECT 33.9 2.117 33.93 2.64 ;
      RECT 33.895 2.147 33.9 2.64 ;
      RECT 33.87 2.175 33.89 2.64 ;
      RECT 33.84 2.22 33.87 2.64 ;
      RECT 33.835 2.247 33.84 2.64 ;
      RECT 33.815 2.265 33.835 2.64 ;
      RECT 33.805 2.29 33.815 2.64 ;
      RECT 33.8 2.302 33.805 2.64 ;
      RECT 33.785 2.325 33.8 2.64 ;
      RECT 33.765 2.352 33.78 2.64 ;
      RECT 33.755 2.375 33.765 2.64 ;
      RECT 35.545 3.26 35.625 3.52 ;
      RECT 34.78 2.48 34.85 2.74 ;
      RECT 35.511 3.227 35.545 3.52 ;
      RECT 35.425 3.13 35.511 3.52 ;
      RECT 35.405 3.042 35.425 3.52 ;
      RECT 35.395 3.012 35.405 3.52 ;
      RECT 35.385 2.992 35.395 3.52 ;
      RECT 35.365 2.979 35.385 3.52 ;
      RECT 35.35 2.969 35.365 3.348 ;
      RECT 35.345 2.962 35.35 3.303 ;
      RECT 35.335 2.956 35.345 3.293 ;
      RECT 35.325 2.948 35.335 3.275 ;
      RECT 35.32 2.942 35.325 3.263 ;
      RECT 35.31 2.937 35.32 3.25 ;
      RECT 35.29 2.927 35.31 3.223 ;
      RECT 35.25 2.906 35.29 3.175 ;
      RECT 35.235 2.887 35.25 3.133 ;
      RECT 35.21 2.873 35.235 3.103 ;
      RECT 35.2 2.861 35.21 3.07 ;
      RECT 35.195 2.856 35.2 3.06 ;
      RECT 35.165 2.842 35.195 3.04 ;
      RECT 35.155 2.826 35.165 3.013 ;
      RECT 35.15 2.821 35.155 3.003 ;
      RECT 35.125 2.812 35.15 2.983 ;
      RECT 35.115 2.8 35.125 2.963 ;
      RECT 35.045 2.768 35.115 2.938 ;
      RECT 35.04 2.737 35.045 2.915 ;
      RECT 34.991 2.48 35.04 2.898 ;
      RECT 34.905 2.48 34.991 2.857 ;
      RECT 34.85 2.48 34.905 2.785 ;
      RECT 34.94 3.265 35.1 3.525 ;
      RECT 34.465 1.88 34.515 2.565 ;
      RECT 34.255 2.305 34.29 2.565 ;
      RECT 34.57 1.88 34.575 2.34 ;
      RECT 34.66 1.88 34.685 2.16 ;
      RECT 34.935 3.262 34.94 3.525 ;
      RECT 34.9 3.25 34.935 3.525 ;
      RECT 34.84 3.223 34.9 3.525 ;
      RECT 34.835 3.206 34.84 3.379 ;
      RECT 34.83 3.203 34.835 3.366 ;
      RECT 34.81 3.196 34.83 3.353 ;
      RECT 34.775 3.179 34.81 3.335 ;
      RECT 34.735 3.158 34.775 3.315 ;
      RECT 34.73 3.146 34.735 3.303 ;
      RECT 34.69 3.132 34.73 3.289 ;
      RECT 34.67 3.115 34.69 3.271 ;
      RECT 34.66 3.107 34.67 3.263 ;
      RECT 34.645 1.88 34.66 2.178 ;
      RECT 34.63 3.097 34.66 3.25 ;
      RECT 34.615 1.88 34.645 2.223 ;
      RECT 34.62 3.087 34.63 3.237 ;
      RECT 34.59 3.072 34.62 3.224 ;
      RECT 34.575 1.88 34.615 2.29 ;
      RECT 34.575 3.04 34.59 3.21 ;
      RECT 34.57 3.012 34.575 3.204 ;
      RECT 34.565 1.88 34.57 2.345 ;
      RECT 34.555 2.982 34.57 3.198 ;
      RECT 34.56 1.88 34.565 2.358 ;
      RECT 34.55 1.88 34.56 2.378 ;
      RECT 34.515 2.895 34.555 3.183 ;
      RECT 34.515 1.88 34.55 2.418 ;
      RECT 34.51 2.827 34.515 3.171 ;
      RECT 34.495 2.782 34.51 3.166 ;
      RECT 34.49 2.72 34.495 3.161 ;
      RECT 34.465 2.627 34.49 3.154 ;
      RECT 34.46 1.88 34.465 3.146 ;
      RECT 34.445 1.88 34.46 3.133 ;
      RECT 34.425 1.88 34.445 3.09 ;
      RECT 34.415 1.88 34.425 3.04 ;
      RECT 34.41 1.88 34.415 3.013 ;
      RECT 34.405 1.88 34.41 2.991 ;
      RECT 34.4 2.106 34.405 2.974 ;
      RECT 34.395 2.128 34.4 2.952 ;
      RECT 34.39 2.17 34.395 2.935 ;
      RECT 34.36 2.22 34.39 2.879 ;
      RECT 34.355 2.247 34.36 2.821 ;
      RECT 34.34 2.265 34.355 2.785 ;
      RECT 34.335 2.283 34.34 2.749 ;
      RECT 34.329 2.29 34.335 2.73 ;
      RECT 34.325 2.297 34.329 2.713 ;
      RECT 34.32 2.302 34.325 2.682 ;
      RECT 34.31 2.305 34.32 2.657 ;
      RECT 34.3 2.305 34.31 2.623 ;
      RECT 34.295 2.305 34.3 2.6 ;
      RECT 34.29 2.305 34.295 2.58 ;
      RECT 33.205 2.44 33.485 2.72 ;
      RECT 33.205 2.44 33.505 2.615 ;
      RECT 33.295 2.33 33.555 2.59 ;
      RECT 33.26 2.425 33.555 2.59 ;
      RECT 33.385 0.945 33.55 2.59 ;
      RECT 33.285 0.945 33.655 1.315 ;
      RECT 32.91 3.47 33.17 3.73 ;
      RECT 32.93 3.397 33.11 3.73 ;
      RECT 32.93 3.14 33.105 3.73 ;
      RECT 32.93 2.932 33.095 3.73 ;
      RECT 32.935 2.85 33.095 3.73 ;
      RECT 32.935 2.615 33.085 3.73 ;
      RECT 32.935 2.462 33.08 3.73 ;
      RECT 32.94 2.447 33.08 3.73 ;
      RECT 32.99 2.162 33.08 3.73 ;
      RECT 32.945 2.397 33.08 3.73 ;
      RECT 32.975 2.215 33.08 3.73 ;
      RECT 32.96 2.327 33.08 3.73 ;
      RECT 32.965 2.285 33.08 3.73 ;
      RECT 32.96 2.327 33.095 2.39 ;
      RECT 32.995 1.915 33.1 2.335 ;
      RECT 32.995 1.915 33.115 2.318 ;
      RECT 32.995 1.915 33.15 2.28 ;
      RECT 32.99 2.162 33.2 2.213 ;
      RECT 32.995 1.915 33.255 2.175 ;
      RECT 32.255 2.62 32.515 2.88 ;
      RECT 32.255 2.62 32.525 2.838 ;
      RECT 32.255 2.62 32.611 2.809 ;
      RECT 32.255 2.62 32.68 2.761 ;
      RECT 32.255 2.62 32.715 2.73 ;
      RECT 32.485 2.44 32.765 2.72 ;
      RECT 32.32 2.605 32.765 2.72 ;
      RECT 32.41 2.482 32.515 2.88 ;
      RECT 32.34 2.545 32.765 2.72 ;
      RECT 26.79 6.22 27.11 6.545 ;
      RECT 26.82 5.695 26.99 6.545 ;
      RECT 26.82 5.695 26.995 6.045 ;
      RECT 26.82 5.695 27.795 5.87 ;
      RECT 27.62 1.965 27.795 5.87 ;
      RECT 27.565 1.965 27.915 2.315 ;
      RECT 27.59 6.655 27.915 6.98 ;
      RECT 26.475 6.745 27.915 6.915 ;
      RECT 26.475 2.395 26.635 6.915 ;
      RECT 26.79 2.365 27.11 2.685 ;
      RECT 26.475 2.395 27.11 2.565 ;
      RECT 25.74 5.86 26.08 6.21 ;
      RECT 25.82 2.705 25.995 6.21 ;
      RECT 25.745 2.705 26.085 3.055 ;
      RECT 25.14 2.705 25.525 3.055 ;
      RECT 25.13 2.77 25.525 2.97 ;
      RECT 25.275 2.7 25.445 3.055 ;
      RECT 23.585 2.44 23.865 2.72 ;
      RECT 23.58 2.44 23.865 2.673 ;
      RECT 23.56 2.44 23.865 2.65 ;
      RECT 23.55 2.44 23.865 2.63 ;
      RECT 23.54 2.44 23.865 2.615 ;
      RECT 23.515 2.44 23.865 2.588 ;
      RECT 23.505 2.44 23.865 2.563 ;
      RECT 23.46 2.295 23.74 2.555 ;
      RECT 23.46 2.39 23.84 2.555 ;
      RECT 23.46 2.335 23.785 2.555 ;
      RECT 23.46 2.327 23.78 2.555 ;
      RECT 23.46 2.317 23.775 2.555 ;
      RECT 23.46 2.305 23.77 2.555 ;
      RECT 22.385 3 22.665 3.28 ;
      RECT 22.385 3 22.7 3.26 ;
      RECT 14.71 6.655 15.06 7.005 ;
      RECT 22.13 6.61 22.48 6.96 ;
      RECT 14.71 6.685 22.48 6.885 ;
      RECT 22.42 2.42 22.47 2.68 ;
      RECT 22.21 2.42 22.215 2.68 ;
      RECT 21.405 1.975 21.435 2.235 ;
      RECT 21.175 1.975 21.25 2.235 ;
      RECT 22.395 2.37 22.42 2.68 ;
      RECT 22.39 2.327 22.395 2.68 ;
      RECT 22.385 2.31 22.39 2.68 ;
      RECT 22.38 2.297 22.385 2.68 ;
      RECT 22.305 2.18 22.38 2.68 ;
      RECT 22.26 1.997 22.305 2.68 ;
      RECT 22.255 1.925 22.26 2.68 ;
      RECT 22.24 1.9 22.255 2.68 ;
      RECT 22.215 1.862 22.24 2.68 ;
      RECT 22.205 1.842 22.215 2.402 ;
      RECT 22.19 1.834 22.205 2.357 ;
      RECT 22.185 1.826 22.19 2.328 ;
      RECT 22.18 1.823 22.185 2.308 ;
      RECT 22.175 1.82 22.18 2.288 ;
      RECT 22.17 1.817 22.175 2.268 ;
      RECT 22.14 1.806 22.17 2.205 ;
      RECT 22.12 1.791 22.14 2.12 ;
      RECT 22.115 1.783 22.12 2.083 ;
      RECT 22.105 1.777 22.115 2.05 ;
      RECT 22.09 1.769 22.105 2.01 ;
      RECT 22.085 1.762 22.09 1.97 ;
      RECT 22.08 1.759 22.085 1.948 ;
      RECT 22.075 1.756 22.08 1.935 ;
      RECT 22.07 1.755 22.075 1.925 ;
      RECT 22.055 1.749 22.07 1.915 ;
      RECT 22.03 1.736 22.055 1.9 ;
      RECT 21.98 1.711 22.03 1.871 ;
      RECT 21.965 1.69 21.98 1.846 ;
      RECT 21.955 1.683 21.965 1.835 ;
      RECT 21.9 1.664 21.955 1.808 ;
      RECT 21.875 1.642 21.9 1.781 ;
      RECT 21.87 1.635 21.875 1.776 ;
      RECT 21.855 1.635 21.87 1.774 ;
      RECT 21.83 1.627 21.855 1.77 ;
      RECT 21.815 1.625 21.83 1.766 ;
      RECT 21.785 1.625 21.815 1.763 ;
      RECT 21.775 1.625 21.785 1.758 ;
      RECT 21.73 1.625 21.775 1.756 ;
      RECT 21.701 1.625 21.73 1.757 ;
      RECT 21.615 1.625 21.701 1.759 ;
      RECT 21.601 1.626 21.615 1.761 ;
      RECT 21.515 1.627 21.601 1.763 ;
      RECT 21.5 1.628 21.515 1.773 ;
      RECT 21.495 1.629 21.5 1.782 ;
      RECT 21.475 1.632 21.495 1.792 ;
      RECT 21.46 1.64 21.475 1.807 ;
      RECT 21.44 1.658 21.46 1.822 ;
      RECT 21.43 1.67 21.44 1.845 ;
      RECT 21.42 1.679 21.43 1.875 ;
      RECT 21.405 1.691 21.42 1.92 ;
      RECT 21.35 1.724 21.405 2.235 ;
      RECT 21.345 1.752 21.35 2.235 ;
      RECT 21.325 1.767 21.345 2.235 ;
      RECT 21.29 1.827 21.325 2.235 ;
      RECT 21.288 1.877 21.29 2.235 ;
      RECT 21.285 1.885 21.288 2.235 ;
      RECT 21.275 1.9 21.285 2.235 ;
      RECT 21.27 1.912 21.275 2.235 ;
      RECT 21.26 1.937 21.27 2.235 ;
      RECT 21.25 1.965 21.26 2.235 ;
      RECT 19.155 3.47 19.205 3.73 ;
      RECT 22.065 3.02 22.125 3.28 ;
      RECT 22.05 3.02 22.065 3.29 ;
      RECT 22.031 3.02 22.05 3.323 ;
      RECT 21.945 3.02 22.031 3.448 ;
      RECT 21.865 3.02 21.945 3.63 ;
      RECT 21.86 3.257 21.865 3.715 ;
      RECT 21.835 3.327 21.86 3.743 ;
      RECT 21.83 3.397 21.835 3.77 ;
      RECT 21.81 3.469 21.83 3.792 ;
      RECT 21.805 3.536 21.81 3.815 ;
      RECT 21.795 3.565 21.805 3.83 ;
      RECT 21.785 3.587 21.795 3.847 ;
      RECT 21.78 3.597 21.785 3.858 ;
      RECT 21.775 3.605 21.78 3.866 ;
      RECT 21.765 3.613 21.775 3.878 ;
      RECT 21.76 3.625 21.765 3.888 ;
      RECT 21.755 3.633 21.76 3.893 ;
      RECT 21.735 3.651 21.755 3.903 ;
      RECT 21.73 3.668 21.735 3.91 ;
      RECT 21.725 3.676 21.73 3.911 ;
      RECT 21.72 3.687 21.725 3.913 ;
      RECT 21.68 3.725 21.72 3.923 ;
      RECT 21.675 3.76 21.68 3.934 ;
      RECT 21.67 3.765 21.675 3.937 ;
      RECT 21.645 3.775 21.67 3.944 ;
      RECT 21.635 3.789 21.645 3.953 ;
      RECT 21.615 3.801 21.635 3.956 ;
      RECT 21.565 3.82 21.615 3.96 ;
      RECT 21.52 3.835 21.565 3.965 ;
      RECT 21.455 3.838 21.52 3.971 ;
      RECT 21.44 3.836 21.455 3.978 ;
      RECT 21.41 3.835 21.44 3.978 ;
      RECT 21.371 3.834 21.41 3.974 ;
      RECT 21.285 3.831 21.371 3.97 ;
      RECT 21.268 3.829 21.285 3.967 ;
      RECT 21.182 3.827 21.268 3.964 ;
      RECT 21.096 3.824 21.182 3.958 ;
      RECT 21.01 3.82 21.096 3.953 ;
      RECT 20.932 3.817 21.01 3.949 ;
      RECT 20.846 3.814 20.932 3.947 ;
      RECT 20.76 3.811 20.846 3.944 ;
      RECT 20.702 3.809 20.76 3.941 ;
      RECT 20.616 3.806 20.702 3.939 ;
      RECT 20.53 3.802 20.616 3.937 ;
      RECT 20.444 3.799 20.53 3.934 ;
      RECT 20.358 3.795 20.444 3.932 ;
      RECT 20.272 3.791 20.358 3.929 ;
      RECT 20.186 3.788 20.272 3.927 ;
      RECT 20.1 3.784 20.186 3.924 ;
      RECT 20.014 3.781 20.1 3.922 ;
      RECT 19.928 3.777 20.014 3.919 ;
      RECT 19.842 3.774 19.928 3.917 ;
      RECT 19.756 3.77 19.842 3.914 ;
      RECT 19.67 3.767 19.756 3.912 ;
      RECT 19.66 3.765 19.67 3.908 ;
      RECT 19.655 3.765 19.66 3.906 ;
      RECT 19.615 3.76 19.655 3.9 ;
      RECT 19.601 3.751 19.615 3.893 ;
      RECT 19.515 3.721 19.601 3.878 ;
      RECT 19.495 3.687 19.515 3.863 ;
      RECT 19.425 3.656 19.495 3.85 ;
      RECT 19.42 3.631 19.425 3.839 ;
      RECT 19.415 3.625 19.42 3.837 ;
      RECT 19.346 3.47 19.415 3.825 ;
      RECT 19.26 3.47 19.346 3.799 ;
      RECT 19.235 3.47 19.26 3.778 ;
      RECT 19.23 3.47 19.235 3.768 ;
      RECT 19.225 3.47 19.23 3.76 ;
      RECT 19.205 3.47 19.225 3.743 ;
      RECT 21.625 2.04 21.885 2.3 ;
      RECT 21.61 2.04 21.885 2.203 ;
      RECT 21.58 2.04 21.885 2.178 ;
      RECT 21.545 1.88 21.825 2.16 ;
      RECT 21.515 3.37 21.575 3.63 ;
      RECT 20.54 2.06 20.595 2.32 ;
      RECT 21.475 3.327 21.515 3.63 ;
      RECT 21.446 3.248 21.475 3.63 ;
      RECT 21.36 3.12 21.446 3.63 ;
      RECT 21.34 3 21.36 3.63 ;
      RECT 21.315 2.951 21.34 3.63 ;
      RECT 21.31 2.916 21.315 3.48 ;
      RECT 21.28 2.876 21.31 3.418 ;
      RECT 21.255 2.813 21.28 3.333 ;
      RECT 21.245 2.775 21.255 3.27 ;
      RECT 21.23 2.75 21.245 3.231 ;
      RECT 21.187 2.708 21.23 3.137 ;
      RECT 21.185 2.681 21.187 3.064 ;
      RECT 21.18 2.676 21.185 3.055 ;
      RECT 21.175 2.669 21.18 3.03 ;
      RECT 21.17 2.663 21.175 3.015 ;
      RECT 21.165 2.657 21.17 3.003 ;
      RECT 21.155 2.648 21.165 2.985 ;
      RECT 21.15 2.639 21.155 2.963 ;
      RECT 21.125 2.62 21.15 2.913 ;
      RECT 21.12 2.601 21.125 2.863 ;
      RECT 21.105 2.587 21.12 2.823 ;
      RECT 21.1 2.573 21.105 2.79 ;
      RECT 21.095 2.566 21.1 2.783 ;
      RECT 21.08 2.553 21.095 2.775 ;
      RECT 21.035 2.515 21.08 2.748 ;
      RECT 21.005 2.468 21.035 2.713 ;
      RECT 20.985 2.437 21.005 2.69 ;
      RECT 20.905 2.37 20.985 2.643 ;
      RECT 20.875 2.3 20.905 2.59 ;
      RECT 20.87 2.277 20.875 2.573 ;
      RECT 20.84 2.255 20.87 2.558 ;
      RECT 20.81 2.214 20.84 2.53 ;
      RECT 20.805 2.189 20.81 2.515 ;
      RECT 20.8 2.183 20.805 2.508 ;
      RECT 20.79 2.06 20.8 2.5 ;
      RECT 20.78 2.06 20.79 2.493 ;
      RECT 20.775 2.06 20.78 2.485 ;
      RECT 20.755 2.06 20.775 2.473 ;
      RECT 20.705 2.06 20.755 2.443 ;
      RECT 20.65 2.06 20.705 2.393 ;
      RECT 20.62 2.06 20.65 2.353 ;
      RECT 20.595 2.06 20.62 2.33 ;
      RECT 20.465 2.785 20.745 3.065 ;
      RECT 20.43 2.7 20.69 2.96 ;
      RECT 20.43 2.782 20.7 2.96 ;
      RECT 18.63 2.155 18.635 2.64 ;
      RECT 18.52 2.34 18.525 2.64 ;
      RECT 18.43 2.38 18.495 2.64 ;
      RECT 20.105 1.88 20.195 2.51 ;
      RECT 20.07 1.93 20.075 2.51 ;
      RECT 20.015 1.955 20.025 2.51 ;
      RECT 19.97 1.955 19.98 2.51 ;
      RECT 20.34 1.88 20.385 2.16 ;
      RECT 19.19 1.61 19.39 1.75 ;
      RECT 20.306 1.88 20.34 2.172 ;
      RECT 20.22 1.88 20.306 2.212 ;
      RECT 20.205 1.88 20.22 2.253 ;
      RECT 20.2 1.88 20.205 2.273 ;
      RECT 20.195 1.88 20.2 2.293 ;
      RECT 20.075 1.922 20.105 2.51 ;
      RECT 20.025 1.942 20.07 2.51 ;
      RECT 20.01 1.957 20.015 2.51 ;
      RECT 19.98 1.957 20.01 2.51 ;
      RECT 19.935 1.942 19.97 2.51 ;
      RECT 19.93 1.93 19.935 2.29 ;
      RECT 19.925 1.927 19.93 2.27 ;
      RECT 19.91 1.917 19.925 2.223 ;
      RECT 19.905 1.91 19.91 2.186 ;
      RECT 19.9 1.907 19.905 2.169 ;
      RECT 19.885 1.897 19.9 2.125 ;
      RECT 19.88 1.888 19.885 2.085 ;
      RECT 19.875 1.884 19.88 2.07 ;
      RECT 19.865 1.878 19.875 2.053 ;
      RECT 19.825 1.859 19.865 2.028 ;
      RECT 19.82 1.841 19.825 2.008 ;
      RECT 19.81 1.835 19.82 2.003 ;
      RECT 19.78 1.819 19.81 1.99 ;
      RECT 19.765 1.801 19.78 1.973 ;
      RECT 19.75 1.789 19.765 1.96 ;
      RECT 19.745 1.781 19.75 1.953 ;
      RECT 19.715 1.767 19.745 1.94 ;
      RECT 19.71 1.752 19.715 1.928 ;
      RECT 19.7 1.746 19.71 1.92 ;
      RECT 19.68 1.734 19.7 1.908 ;
      RECT 19.67 1.722 19.68 1.895 ;
      RECT 19.64 1.706 19.67 1.88 ;
      RECT 19.62 1.686 19.64 1.863 ;
      RECT 19.615 1.676 19.62 1.853 ;
      RECT 19.59 1.664 19.615 1.84 ;
      RECT 19.585 1.652 19.59 1.828 ;
      RECT 19.58 1.647 19.585 1.824 ;
      RECT 19.565 1.64 19.58 1.816 ;
      RECT 19.555 1.627 19.565 1.806 ;
      RECT 19.55 1.625 19.555 1.8 ;
      RECT 19.525 1.618 19.55 1.789 ;
      RECT 19.52 1.611 19.525 1.778 ;
      RECT 19.495 1.61 19.52 1.765 ;
      RECT 19.476 1.61 19.495 1.755 ;
      RECT 19.39 1.61 19.476 1.752 ;
      RECT 19.16 1.61 19.19 1.755 ;
      RECT 19.12 1.617 19.16 1.768 ;
      RECT 19.095 1.627 19.12 1.781 ;
      RECT 19.08 1.636 19.095 1.791 ;
      RECT 19.05 1.641 19.08 1.81 ;
      RECT 19.045 1.647 19.05 1.828 ;
      RECT 19.025 1.657 19.045 1.843 ;
      RECT 19.015 1.67 19.025 1.863 ;
      RECT 19 1.682 19.015 1.88 ;
      RECT 18.995 1.692 19 1.89 ;
      RECT 18.99 1.697 18.995 1.895 ;
      RECT 18.98 1.705 18.99 1.908 ;
      RECT 18.93 1.737 18.98 1.945 ;
      RECT 18.915 1.772 18.93 1.986 ;
      RECT 18.91 1.782 18.915 2.001 ;
      RECT 18.905 1.787 18.91 2.008 ;
      RECT 18.88 1.803 18.905 2.028 ;
      RECT 18.865 1.824 18.88 2.053 ;
      RECT 18.84 1.845 18.865 2.078 ;
      RECT 18.83 1.864 18.84 2.101 ;
      RECT 18.805 1.882 18.83 2.124 ;
      RECT 18.79 1.902 18.805 2.148 ;
      RECT 18.785 1.912 18.79 2.16 ;
      RECT 18.77 1.924 18.785 2.18 ;
      RECT 18.76 1.939 18.77 2.22 ;
      RECT 18.755 1.947 18.76 2.248 ;
      RECT 18.745 1.957 18.755 2.268 ;
      RECT 18.74 1.97 18.745 2.293 ;
      RECT 18.735 1.983 18.74 2.313 ;
      RECT 18.73 1.989 18.735 2.335 ;
      RECT 18.72 1.998 18.73 2.355 ;
      RECT 18.715 2.018 18.72 2.378 ;
      RECT 18.71 2.024 18.715 2.398 ;
      RECT 18.705 2.031 18.71 2.42 ;
      RECT 18.7 2.042 18.705 2.433 ;
      RECT 18.69 2.052 18.7 2.458 ;
      RECT 18.67 2.077 18.69 2.64 ;
      RECT 18.64 2.117 18.67 2.64 ;
      RECT 18.635 2.147 18.64 2.64 ;
      RECT 18.61 2.175 18.63 2.64 ;
      RECT 18.58 2.22 18.61 2.64 ;
      RECT 18.575 2.247 18.58 2.64 ;
      RECT 18.555 2.265 18.575 2.64 ;
      RECT 18.545 2.29 18.555 2.64 ;
      RECT 18.54 2.302 18.545 2.64 ;
      RECT 18.525 2.325 18.54 2.64 ;
      RECT 18.505 2.352 18.52 2.64 ;
      RECT 18.495 2.375 18.505 2.64 ;
      RECT 20.285 3.26 20.365 3.52 ;
      RECT 19.52 2.48 19.59 2.74 ;
      RECT 20.251 3.227 20.285 3.52 ;
      RECT 20.165 3.13 20.251 3.52 ;
      RECT 20.145 3.042 20.165 3.52 ;
      RECT 20.135 3.012 20.145 3.52 ;
      RECT 20.125 2.992 20.135 3.52 ;
      RECT 20.105 2.979 20.125 3.52 ;
      RECT 20.09 2.969 20.105 3.348 ;
      RECT 20.085 2.962 20.09 3.303 ;
      RECT 20.075 2.956 20.085 3.293 ;
      RECT 20.065 2.948 20.075 3.275 ;
      RECT 20.06 2.942 20.065 3.263 ;
      RECT 20.05 2.937 20.06 3.25 ;
      RECT 20.03 2.927 20.05 3.223 ;
      RECT 19.99 2.906 20.03 3.175 ;
      RECT 19.975 2.887 19.99 3.133 ;
      RECT 19.95 2.873 19.975 3.103 ;
      RECT 19.94 2.861 19.95 3.07 ;
      RECT 19.935 2.856 19.94 3.06 ;
      RECT 19.905 2.842 19.935 3.04 ;
      RECT 19.895 2.826 19.905 3.013 ;
      RECT 19.89 2.821 19.895 3.003 ;
      RECT 19.865 2.812 19.89 2.983 ;
      RECT 19.855 2.8 19.865 2.963 ;
      RECT 19.785 2.768 19.855 2.938 ;
      RECT 19.78 2.737 19.785 2.915 ;
      RECT 19.731 2.48 19.78 2.898 ;
      RECT 19.645 2.48 19.731 2.857 ;
      RECT 19.59 2.48 19.645 2.785 ;
      RECT 19.68 3.265 19.84 3.525 ;
      RECT 19.205 1.88 19.255 2.565 ;
      RECT 18.995 2.305 19.03 2.565 ;
      RECT 19.31 1.88 19.315 2.34 ;
      RECT 19.4 1.88 19.425 2.16 ;
      RECT 19.675 3.262 19.68 3.525 ;
      RECT 19.64 3.25 19.675 3.525 ;
      RECT 19.58 3.223 19.64 3.525 ;
      RECT 19.575 3.206 19.58 3.379 ;
      RECT 19.57 3.203 19.575 3.366 ;
      RECT 19.55 3.196 19.57 3.353 ;
      RECT 19.515 3.179 19.55 3.335 ;
      RECT 19.475 3.158 19.515 3.315 ;
      RECT 19.47 3.146 19.475 3.303 ;
      RECT 19.43 3.132 19.47 3.289 ;
      RECT 19.41 3.115 19.43 3.271 ;
      RECT 19.4 3.107 19.41 3.263 ;
      RECT 19.385 1.88 19.4 2.178 ;
      RECT 19.37 3.097 19.4 3.25 ;
      RECT 19.355 1.88 19.385 2.223 ;
      RECT 19.36 3.087 19.37 3.237 ;
      RECT 19.33 3.072 19.36 3.224 ;
      RECT 19.315 1.88 19.355 2.29 ;
      RECT 19.315 3.04 19.33 3.21 ;
      RECT 19.31 3.012 19.315 3.204 ;
      RECT 19.305 1.88 19.31 2.345 ;
      RECT 19.295 2.982 19.31 3.198 ;
      RECT 19.3 1.88 19.305 2.358 ;
      RECT 19.29 1.88 19.3 2.378 ;
      RECT 19.255 2.895 19.295 3.183 ;
      RECT 19.255 1.88 19.29 2.418 ;
      RECT 19.25 2.827 19.255 3.171 ;
      RECT 19.235 2.782 19.25 3.166 ;
      RECT 19.23 2.72 19.235 3.161 ;
      RECT 19.205 2.627 19.23 3.154 ;
      RECT 19.2 1.88 19.205 3.146 ;
      RECT 19.185 1.88 19.2 3.133 ;
      RECT 19.165 1.88 19.185 3.09 ;
      RECT 19.155 1.88 19.165 3.04 ;
      RECT 19.15 1.88 19.155 3.013 ;
      RECT 19.145 1.88 19.15 2.991 ;
      RECT 19.14 2.106 19.145 2.974 ;
      RECT 19.135 2.128 19.14 2.952 ;
      RECT 19.13 2.17 19.135 2.935 ;
      RECT 19.1 2.22 19.13 2.879 ;
      RECT 19.095 2.247 19.1 2.821 ;
      RECT 19.08 2.265 19.095 2.785 ;
      RECT 19.075 2.283 19.08 2.749 ;
      RECT 19.069 2.29 19.075 2.73 ;
      RECT 19.065 2.297 19.069 2.713 ;
      RECT 19.06 2.302 19.065 2.682 ;
      RECT 19.05 2.305 19.06 2.657 ;
      RECT 19.04 2.305 19.05 2.623 ;
      RECT 19.035 2.305 19.04 2.6 ;
      RECT 19.03 2.305 19.035 2.58 ;
      RECT 17.945 2.44 18.225 2.72 ;
      RECT 17.945 2.44 18.245 2.615 ;
      RECT 18.035 2.33 18.295 2.59 ;
      RECT 18 2.425 18.295 2.59 ;
      RECT 18.125 0.945 18.29 2.59 ;
      RECT 18.025 0.945 18.395 1.315 ;
      RECT 17.65 3.47 17.91 3.73 ;
      RECT 17.67 3.397 17.85 3.73 ;
      RECT 17.67 3.14 17.845 3.73 ;
      RECT 17.67 2.932 17.835 3.73 ;
      RECT 17.675 2.85 17.835 3.73 ;
      RECT 17.675 2.615 17.825 3.73 ;
      RECT 17.675 2.462 17.82 3.73 ;
      RECT 17.68 2.447 17.82 3.73 ;
      RECT 17.73 2.162 17.82 3.73 ;
      RECT 17.685 2.397 17.82 3.73 ;
      RECT 17.715 2.215 17.82 3.73 ;
      RECT 17.7 2.327 17.82 3.73 ;
      RECT 17.705 2.285 17.82 3.73 ;
      RECT 17.7 2.327 17.835 2.39 ;
      RECT 17.735 1.915 17.84 2.335 ;
      RECT 17.735 1.915 17.855 2.318 ;
      RECT 17.735 1.915 17.89 2.28 ;
      RECT 17.73 2.162 17.94 2.213 ;
      RECT 17.735 1.915 17.995 2.175 ;
      RECT 16.995 2.62 17.255 2.88 ;
      RECT 16.995 2.62 17.265 2.838 ;
      RECT 16.995 2.62 17.351 2.809 ;
      RECT 16.995 2.62 17.42 2.761 ;
      RECT 16.995 2.62 17.455 2.73 ;
      RECT 17.225 2.44 17.505 2.72 ;
      RECT 17.06 2.605 17.505 2.72 ;
      RECT 17.15 2.482 17.255 2.88 ;
      RECT 17.08 2.545 17.505 2.72 ;
      RECT 11.53 6.22 11.85 6.545 ;
      RECT 11.56 5.695 11.73 6.545 ;
      RECT 11.56 5.695 11.735 6.045 ;
      RECT 11.56 5.695 12.535 5.87 ;
      RECT 12.36 1.965 12.535 5.87 ;
      RECT 12.305 1.965 12.655 2.315 ;
      RECT 12.33 6.655 12.655 6.98 ;
      RECT 11.215 6.745 12.655 6.915 ;
      RECT 11.215 2.395 11.375 6.915 ;
      RECT 11.53 2.365 11.85 2.685 ;
      RECT 11.215 2.395 11.85 2.565 ;
      RECT 10.48 5.86 10.82 6.21 ;
      RECT 10.56 2.705 10.735 6.21 ;
      RECT 10.485 2.705 10.825 3.055 ;
      RECT 9.88 2.705 10.265 3.055 ;
      RECT 9.87 2.77 10.265 2.97 ;
      RECT 10.015 2.7 10.185 3.055 ;
      RECT 8.325 2.44 8.605 2.72 ;
      RECT 8.32 2.44 8.605 2.673 ;
      RECT 8.3 2.44 8.605 2.65 ;
      RECT 8.29 2.44 8.605 2.63 ;
      RECT 8.28 2.44 8.605 2.615 ;
      RECT 8.255 2.44 8.605 2.588 ;
      RECT 8.245 2.44 8.605 2.563 ;
      RECT 8.2 2.295 8.48 2.555 ;
      RECT 8.2 2.39 8.58 2.555 ;
      RECT 8.2 2.335 8.525 2.555 ;
      RECT 8.2 2.327 8.52 2.555 ;
      RECT 8.2 2.317 8.515 2.555 ;
      RECT 8.2 2.305 8.51 2.555 ;
      RECT 7.125 3 7.405 3.28 ;
      RECT 7.125 3 7.44 3.26 ;
      RECT -1.255 6.995 -0.965 7.345 ;
      RECT -1.255 7.07 0.11 7.24 ;
      RECT -0.06 6.685 0.11 7.24 ;
      RECT 6.87 6.605 7.22 6.955 ;
      RECT -0.06 6.685 7.22 6.855 ;
      RECT 7.16 2.42 7.21 2.68 ;
      RECT 6.95 2.42 6.955 2.68 ;
      RECT 6.145 1.975 6.175 2.235 ;
      RECT 5.915 1.975 5.99 2.235 ;
      RECT 7.135 2.37 7.16 2.68 ;
      RECT 7.13 2.327 7.135 2.68 ;
      RECT 7.125 2.31 7.13 2.68 ;
      RECT 7.12 2.297 7.125 2.68 ;
      RECT 7.045 2.18 7.12 2.68 ;
      RECT 7 1.997 7.045 2.68 ;
      RECT 6.995 1.925 7 2.68 ;
      RECT 6.98 1.9 6.995 2.68 ;
      RECT 6.955 1.862 6.98 2.68 ;
      RECT 6.945 1.842 6.955 2.402 ;
      RECT 6.93 1.834 6.945 2.357 ;
      RECT 6.925 1.826 6.93 2.328 ;
      RECT 6.92 1.823 6.925 2.308 ;
      RECT 6.915 1.82 6.92 2.288 ;
      RECT 6.91 1.817 6.915 2.268 ;
      RECT 6.88 1.806 6.91 2.205 ;
      RECT 6.86 1.791 6.88 2.12 ;
      RECT 6.855 1.783 6.86 2.083 ;
      RECT 6.845 1.777 6.855 2.05 ;
      RECT 6.83 1.769 6.845 2.01 ;
      RECT 6.825 1.762 6.83 1.97 ;
      RECT 6.82 1.759 6.825 1.948 ;
      RECT 6.815 1.756 6.82 1.935 ;
      RECT 6.81 1.755 6.815 1.925 ;
      RECT 6.795 1.749 6.81 1.915 ;
      RECT 6.77 1.736 6.795 1.9 ;
      RECT 6.72 1.711 6.77 1.871 ;
      RECT 6.705 1.69 6.72 1.846 ;
      RECT 6.695 1.683 6.705 1.835 ;
      RECT 6.64 1.664 6.695 1.808 ;
      RECT 6.615 1.642 6.64 1.781 ;
      RECT 6.61 1.635 6.615 1.776 ;
      RECT 6.595 1.635 6.61 1.774 ;
      RECT 6.57 1.627 6.595 1.77 ;
      RECT 6.555 1.625 6.57 1.766 ;
      RECT 6.525 1.625 6.555 1.763 ;
      RECT 6.515 1.625 6.525 1.758 ;
      RECT 6.47 1.625 6.515 1.756 ;
      RECT 6.441 1.625 6.47 1.757 ;
      RECT 6.355 1.625 6.441 1.759 ;
      RECT 6.341 1.626 6.355 1.761 ;
      RECT 6.255 1.627 6.341 1.763 ;
      RECT 6.24 1.628 6.255 1.773 ;
      RECT 6.235 1.629 6.24 1.782 ;
      RECT 6.215 1.632 6.235 1.792 ;
      RECT 6.2 1.64 6.215 1.807 ;
      RECT 6.18 1.658 6.2 1.822 ;
      RECT 6.17 1.67 6.18 1.845 ;
      RECT 6.16 1.679 6.17 1.875 ;
      RECT 6.145 1.691 6.16 1.92 ;
      RECT 6.09 1.724 6.145 2.235 ;
      RECT 6.085 1.752 6.09 2.235 ;
      RECT 6.065 1.767 6.085 2.235 ;
      RECT 6.03 1.827 6.065 2.235 ;
      RECT 6.028 1.877 6.03 2.235 ;
      RECT 6.025 1.885 6.028 2.235 ;
      RECT 6.015 1.9 6.025 2.235 ;
      RECT 6.01 1.912 6.015 2.235 ;
      RECT 6 1.937 6.01 2.235 ;
      RECT 5.99 1.965 6 2.235 ;
      RECT 3.895 3.47 3.945 3.73 ;
      RECT 6.805 3.02 6.865 3.28 ;
      RECT 6.79 3.02 6.805 3.29 ;
      RECT 6.771 3.02 6.79 3.323 ;
      RECT 6.685 3.02 6.771 3.448 ;
      RECT 6.605 3.02 6.685 3.63 ;
      RECT 6.6 3.257 6.605 3.715 ;
      RECT 6.575 3.327 6.6 3.743 ;
      RECT 6.57 3.397 6.575 3.77 ;
      RECT 6.55 3.469 6.57 3.792 ;
      RECT 6.545 3.536 6.55 3.815 ;
      RECT 6.535 3.565 6.545 3.83 ;
      RECT 6.525 3.587 6.535 3.847 ;
      RECT 6.52 3.597 6.525 3.858 ;
      RECT 6.515 3.605 6.52 3.866 ;
      RECT 6.505 3.613 6.515 3.878 ;
      RECT 6.5 3.625 6.505 3.888 ;
      RECT 6.495 3.633 6.5 3.893 ;
      RECT 6.475 3.651 6.495 3.903 ;
      RECT 6.47 3.668 6.475 3.91 ;
      RECT 6.465 3.676 6.47 3.911 ;
      RECT 6.46 3.687 6.465 3.913 ;
      RECT 6.42 3.725 6.46 3.923 ;
      RECT 6.415 3.76 6.42 3.934 ;
      RECT 6.41 3.765 6.415 3.937 ;
      RECT 6.385 3.775 6.41 3.944 ;
      RECT 6.375 3.789 6.385 3.953 ;
      RECT 6.355 3.801 6.375 3.956 ;
      RECT 6.305 3.82 6.355 3.96 ;
      RECT 6.26 3.835 6.305 3.965 ;
      RECT 6.195 3.838 6.26 3.971 ;
      RECT 6.18 3.836 6.195 3.978 ;
      RECT 6.15 3.835 6.18 3.978 ;
      RECT 6.111 3.834 6.15 3.974 ;
      RECT 6.025 3.831 6.111 3.97 ;
      RECT 6.008 3.829 6.025 3.967 ;
      RECT 5.922 3.827 6.008 3.964 ;
      RECT 5.836 3.824 5.922 3.958 ;
      RECT 5.75 3.82 5.836 3.953 ;
      RECT 5.672 3.817 5.75 3.949 ;
      RECT 5.586 3.814 5.672 3.947 ;
      RECT 5.5 3.811 5.586 3.944 ;
      RECT 5.442 3.809 5.5 3.941 ;
      RECT 5.356 3.806 5.442 3.939 ;
      RECT 5.27 3.802 5.356 3.937 ;
      RECT 5.184 3.799 5.27 3.934 ;
      RECT 5.098 3.795 5.184 3.932 ;
      RECT 5.012 3.791 5.098 3.929 ;
      RECT 4.926 3.788 5.012 3.927 ;
      RECT 4.84 3.784 4.926 3.924 ;
      RECT 4.754 3.781 4.84 3.922 ;
      RECT 4.668 3.777 4.754 3.919 ;
      RECT 4.582 3.774 4.668 3.917 ;
      RECT 4.496 3.77 4.582 3.914 ;
      RECT 4.41 3.767 4.496 3.912 ;
      RECT 4.4 3.765 4.41 3.908 ;
      RECT 4.395 3.765 4.4 3.906 ;
      RECT 4.355 3.76 4.395 3.9 ;
      RECT 4.341 3.751 4.355 3.893 ;
      RECT 4.255 3.721 4.341 3.878 ;
      RECT 4.235 3.687 4.255 3.863 ;
      RECT 4.165 3.656 4.235 3.85 ;
      RECT 4.16 3.631 4.165 3.839 ;
      RECT 4.155 3.625 4.16 3.837 ;
      RECT 4.086 3.47 4.155 3.825 ;
      RECT 4 3.47 4.086 3.799 ;
      RECT 3.975 3.47 4 3.778 ;
      RECT 3.97 3.47 3.975 3.768 ;
      RECT 3.965 3.47 3.97 3.76 ;
      RECT 3.945 3.47 3.965 3.743 ;
      RECT 6.365 2.04 6.625 2.3 ;
      RECT 6.35 2.04 6.625 2.203 ;
      RECT 6.32 2.04 6.625 2.178 ;
      RECT 6.285 1.88 6.565 2.16 ;
      RECT 6.255 3.37 6.315 3.63 ;
      RECT 5.28 2.06 5.335 2.32 ;
      RECT 6.215 3.327 6.255 3.63 ;
      RECT 6.186 3.248 6.215 3.63 ;
      RECT 6.1 3.12 6.186 3.63 ;
      RECT 6.08 3 6.1 3.63 ;
      RECT 6.055 2.951 6.08 3.63 ;
      RECT 6.05 2.916 6.055 3.48 ;
      RECT 6.02 2.876 6.05 3.418 ;
      RECT 5.995 2.813 6.02 3.333 ;
      RECT 5.985 2.775 5.995 3.27 ;
      RECT 5.97 2.75 5.985 3.231 ;
      RECT 5.927 2.708 5.97 3.137 ;
      RECT 5.925 2.681 5.927 3.064 ;
      RECT 5.92 2.676 5.925 3.055 ;
      RECT 5.915 2.669 5.92 3.03 ;
      RECT 5.91 2.663 5.915 3.015 ;
      RECT 5.905 2.657 5.91 3.003 ;
      RECT 5.895 2.648 5.905 2.985 ;
      RECT 5.89 2.639 5.895 2.963 ;
      RECT 5.865 2.62 5.89 2.913 ;
      RECT 5.86 2.601 5.865 2.863 ;
      RECT 5.845 2.587 5.86 2.823 ;
      RECT 5.84 2.573 5.845 2.79 ;
      RECT 5.835 2.566 5.84 2.783 ;
      RECT 5.82 2.553 5.835 2.775 ;
      RECT 5.775 2.515 5.82 2.748 ;
      RECT 5.745 2.468 5.775 2.713 ;
      RECT 5.725 2.437 5.745 2.69 ;
      RECT 5.645 2.37 5.725 2.643 ;
      RECT 5.615 2.3 5.645 2.59 ;
      RECT 5.61 2.277 5.615 2.573 ;
      RECT 5.58 2.255 5.61 2.558 ;
      RECT 5.55 2.214 5.58 2.53 ;
      RECT 5.545 2.189 5.55 2.515 ;
      RECT 5.54 2.183 5.545 2.508 ;
      RECT 5.53 2.06 5.54 2.5 ;
      RECT 5.52 2.06 5.53 2.493 ;
      RECT 5.515 2.06 5.52 2.485 ;
      RECT 5.495 2.06 5.515 2.473 ;
      RECT 5.445 2.06 5.495 2.443 ;
      RECT 5.39 2.06 5.445 2.393 ;
      RECT 5.36 2.06 5.39 2.353 ;
      RECT 5.335 2.06 5.36 2.33 ;
      RECT 5.205 2.785 5.485 3.065 ;
      RECT 5.17 2.7 5.43 2.96 ;
      RECT 5.17 2.782 5.44 2.96 ;
      RECT 3.37 2.155 3.375 2.64 ;
      RECT 3.26 2.34 3.265 2.64 ;
      RECT 3.17 2.38 3.235 2.64 ;
      RECT 4.845 1.88 4.935 2.51 ;
      RECT 4.81 1.93 4.815 2.51 ;
      RECT 4.755 1.955 4.765 2.51 ;
      RECT 4.71 1.955 4.72 2.51 ;
      RECT 5.08 1.88 5.125 2.16 ;
      RECT 3.93 1.61 4.13 1.75 ;
      RECT 5.046 1.88 5.08 2.172 ;
      RECT 4.96 1.88 5.046 2.212 ;
      RECT 4.945 1.88 4.96 2.253 ;
      RECT 4.94 1.88 4.945 2.273 ;
      RECT 4.935 1.88 4.94 2.293 ;
      RECT 4.815 1.922 4.845 2.51 ;
      RECT 4.765 1.942 4.81 2.51 ;
      RECT 4.75 1.957 4.755 2.51 ;
      RECT 4.72 1.957 4.75 2.51 ;
      RECT 4.675 1.942 4.71 2.51 ;
      RECT 4.67 1.93 4.675 2.29 ;
      RECT 4.665 1.927 4.67 2.27 ;
      RECT 4.65 1.917 4.665 2.223 ;
      RECT 4.645 1.91 4.65 2.186 ;
      RECT 4.64 1.907 4.645 2.169 ;
      RECT 4.625 1.897 4.64 2.125 ;
      RECT 4.62 1.888 4.625 2.085 ;
      RECT 4.615 1.884 4.62 2.07 ;
      RECT 4.605 1.878 4.615 2.053 ;
      RECT 4.565 1.859 4.605 2.028 ;
      RECT 4.56 1.841 4.565 2.008 ;
      RECT 4.55 1.835 4.56 2.003 ;
      RECT 4.52 1.819 4.55 1.99 ;
      RECT 4.505 1.801 4.52 1.973 ;
      RECT 4.49 1.789 4.505 1.96 ;
      RECT 4.485 1.781 4.49 1.953 ;
      RECT 4.455 1.767 4.485 1.94 ;
      RECT 4.45 1.752 4.455 1.928 ;
      RECT 4.44 1.746 4.45 1.92 ;
      RECT 4.42 1.734 4.44 1.908 ;
      RECT 4.41 1.722 4.42 1.895 ;
      RECT 4.38 1.706 4.41 1.88 ;
      RECT 4.36 1.686 4.38 1.863 ;
      RECT 4.355 1.676 4.36 1.853 ;
      RECT 4.33 1.664 4.355 1.84 ;
      RECT 4.325 1.652 4.33 1.828 ;
      RECT 4.32 1.647 4.325 1.824 ;
      RECT 4.305 1.64 4.32 1.816 ;
      RECT 4.295 1.627 4.305 1.806 ;
      RECT 4.29 1.625 4.295 1.8 ;
      RECT 4.265 1.618 4.29 1.789 ;
      RECT 4.26 1.611 4.265 1.778 ;
      RECT 4.235 1.61 4.26 1.765 ;
      RECT 4.216 1.61 4.235 1.755 ;
      RECT 4.13 1.61 4.216 1.752 ;
      RECT 3.9 1.61 3.93 1.755 ;
      RECT 3.86 1.617 3.9 1.768 ;
      RECT 3.835 1.627 3.86 1.781 ;
      RECT 3.82 1.636 3.835 1.791 ;
      RECT 3.79 1.641 3.82 1.81 ;
      RECT 3.785 1.647 3.79 1.828 ;
      RECT 3.765 1.657 3.785 1.843 ;
      RECT 3.755 1.67 3.765 1.863 ;
      RECT 3.74 1.682 3.755 1.88 ;
      RECT 3.735 1.692 3.74 1.89 ;
      RECT 3.73 1.697 3.735 1.895 ;
      RECT 3.72 1.705 3.73 1.908 ;
      RECT 3.67 1.737 3.72 1.945 ;
      RECT 3.655 1.772 3.67 1.986 ;
      RECT 3.65 1.782 3.655 2.001 ;
      RECT 3.645 1.787 3.65 2.008 ;
      RECT 3.62 1.803 3.645 2.028 ;
      RECT 3.605 1.824 3.62 2.053 ;
      RECT 3.58 1.845 3.605 2.078 ;
      RECT 3.57 1.864 3.58 2.101 ;
      RECT 3.545 1.882 3.57 2.124 ;
      RECT 3.53 1.902 3.545 2.148 ;
      RECT 3.525 1.912 3.53 2.16 ;
      RECT 3.51 1.924 3.525 2.18 ;
      RECT 3.5 1.939 3.51 2.22 ;
      RECT 3.495 1.947 3.5 2.248 ;
      RECT 3.485 1.957 3.495 2.268 ;
      RECT 3.48 1.97 3.485 2.293 ;
      RECT 3.475 1.983 3.48 2.313 ;
      RECT 3.47 1.989 3.475 2.335 ;
      RECT 3.46 1.998 3.47 2.355 ;
      RECT 3.455 2.018 3.46 2.378 ;
      RECT 3.45 2.024 3.455 2.398 ;
      RECT 3.445 2.031 3.45 2.42 ;
      RECT 3.44 2.042 3.445 2.433 ;
      RECT 3.43 2.052 3.44 2.458 ;
      RECT 3.41 2.077 3.43 2.64 ;
      RECT 3.38 2.117 3.41 2.64 ;
      RECT 3.375 2.147 3.38 2.64 ;
      RECT 3.35 2.175 3.37 2.64 ;
      RECT 3.32 2.22 3.35 2.64 ;
      RECT 3.315 2.247 3.32 2.64 ;
      RECT 3.295 2.265 3.315 2.64 ;
      RECT 3.285 2.29 3.295 2.64 ;
      RECT 3.28 2.302 3.285 2.64 ;
      RECT 3.265 2.325 3.28 2.64 ;
      RECT 3.245 2.352 3.26 2.64 ;
      RECT 3.235 2.375 3.245 2.64 ;
      RECT 5.025 3.26 5.105 3.52 ;
      RECT 4.26 2.48 4.33 2.74 ;
      RECT 4.991 3.227 5.025 3.52 ;
      RECT 4.905 3.13 4.991 3.52 ;
      RECT 4.885 3.042 4.905 3.52 ;
      RECT 4.875 3.012 4.885 3.52 ;
      RECT 4.865 2.992 4.875 3.52 ;
      RECT 4.845 2.979 4.865 3.52 ;
      RECT 4.83 2.969 4.845 3.348 ;
      RECT 4.825 2.962 4.83 3.303 ;
      RECT 4.815 2.956 4.825 3.293 ;
      RECT 4.805 2.948 4.815 3.275 ;
      RECT 4.8 2.942 4.805 3.263 ;
      RECT 4.79 2.937 4.8 3.25 ;
      RECT 4.77 2.927 4.79 3.223 ;
      RECT 4.73 2.906 4.77 3.175 ;
      RECT 4.715 2.887 4.73 3.133 ;
      RECT 4.69 2.873 4.715 3.103 ;
      RECT 4.68 2.861 4.69 3.07 ;
      RECT 4.675 2.856 4.68 3.06 ;
      RECT 4.645 2.842 4.675 3.04 ;
      RECT 4.635 2.826 4.645 3.013 ;
      RECT 4.63 2.821 4.635 3.003 ;
      RECT 4.605 2.812 4.63 2.983 ;
      RECT 4.595 2.8 4.605 2.963 ;
      RECT 4.525 2.768 4.595 2.938 ;
      RECT 4.52 2.737 4.525 2.915 ;
      RECT 4.471 2.48 4.52 2.898 ;
      RECT 4.385 2.48 4.471 2.857 ;
      RECT 4.33 2.48 4.385 2.785 ;
      RECT 4.42 3.265 4.58 3.525 ;
      RECT 3.945 1.88 3.995 2.565 ;
      RECT 3.735 2.305 3.77 2.565 ;
      RECT 4.05 1.88 4.055 2.34 ;
      RECT 4.14 1.88 4.165 2.16 ;
      RECT 4.415 3.262 4.42 3.525 ;
      RECT 4.38 3.25 4.415 3.525 ;
      RECT 4.32 3.223 4.38 3.525 ;
      RECT 4.315 3.206 4.32 3.379 ;
      RECT 4.31 3.203 4.315 3.366 ;
      RECT 4.29 3.196 4.31 3.353 ;
      RECT 4.255 3.179 4.29 3.335 ;
      RECT 4.215 3.158 4.255 3.315 ;
      RECT 4.21 3.146 4.215 3.303 ;
      RECT 4.17 3.132 4.21 3.289 ;
      RECT 4.15 3.115 4.17 3.271 ;
      RECT 4.14 3.107 4.15 3.263 ;
      RECT 4.125 1.88 4.14 2.178 ;
      RECT 4.11 3.097 4.14 3.25 ;
      RECT 4.095 1.88 4.125 2.223 ;
      RECT 4.1 3.087 4.11 3.237 ;
      RECT 4.07 3.072 4.1 3.224 ;
      RECT 4.055 1.88 4.095 2.29 ;
      RECT 4.055 3.04 4.07 3.21 ;
      RECT 4.05 3.012 4.055 3.204 ;
      RECT 4.045 1.88 4.05 2.345 ;
      RECT 4.035 2.982 4.05 3.198 ;
      RECT 4.04 1.88 4.045 2.358 ;
      RECT 4.03 1.88 4.04 2.378 ;
      RECT 3.995 2.895 4.035 3.183 ;
      RECT 3.995 1.88 4.03 2.418 ;
      RECT 3.99 2.827 3.995 3.171 ;
      RECT 3.975 2.782 3.99 3.166 ;
      RECT 3.97 2.72 3.975 3.161 ;
      RECT 3.945 2.627 3.97 3.154 ;
      RECT 3.94 1.88 3.945 3.146 ;
      RECT 3.925 1.88 3.94 3.133 ;
      RECT 3.905 1.88 3.925 3.09 ;
      RECT 3.895 1.88 3.905 3.04 ;
      RECT 3.89 1.88 3.895 3.013 ;
      RECT 3.885 1.88 3.89 2.991 ;
      RECT 3.88 2.106 3.885 2.974 ;
      RECT 3.875 2.128 3.88 2.952 ;
      RECT 3.87 2.17 3.875 2.935 ;
      RECT 3.84 2.22 3.87 2.879 ;
      RECT 3.835 2.247 3.84 2.821 ;
      RECT 3.82 2.265 3.835 2.785 ;
      RECT 3.815 2.283 3.82 2.749 ;
      RECT 3.809 2.29 3.815 2.73 ;
      RECT 3.805 2.297 3.809 2.713 ;
      RECT 3.8 2.302 3.805 2.682 ;
      RECT 3.79 2.305 3.8 2.657 ;
      RECT 3.78 2.305 3.79 2.623 ;
      RECT 3.775 2.305 3.78 2.6 ;
      RECT 3.77 2.305 3.775 2.58 ;
      RECT 2.685 2.44 2.965 2.72 ;
      RECT 2.685 2.44 2.985 2.615 ;
      RECT 2.775 2.33 3.035 2.59 ;
      RECT 2.74 2.425 3.035 2.59 ;
      RECT 2.865 0.945 3.03 2.59 ;
      RECT 2.765 0.945 3.135 1.315 ;
      RECT 2.39 3.47 2.65 3.73 ;
      RECT 2.41 3.397 2.59 3.73 ;
      RECT 2.41 3.14 2.585 3.73 ;
      RECT 2.41 2.932 2.575 3.73 ;
      RECT 2.415 2.85 2.575 3.73 ;
      RECT 2.415 2.615 2.565 3.73 ;
      RECT 2.415 2.462 2.56 3.73 ;
      RECT 2.42 2.447 2.56 3.73 ;
      RECT 2.47 2.162 2.56 3.73 ;
      RECT 2.425 2.397 2.56 3.73 ;
      RECT 2.455 2.215 2.56 3.73 ;
      RECT 2.44 2.327 2.56 3.73 ;
      RECT 2.445 2.285 2.56 3.73 ;
      RECT 2.44 2.327 2.575 2.39 ;
      RECT 2.475 1.915 2.58 2.335 ;
      RECT 2.475 1.915 2.595 2.318 ;
      RECT 2.475 1.915 2.63 2.28 ;
      RECT 2.47 2.162 2.68 2.213 ;
      RECT 2.475 1.915 2.735 2.175 ;
      RECT 1.735 2.62 1.995 2.88 ;
      RECT 1.735 2.62 2.005 2.838 ;
      RECT 1.735 2.62 2.091 2.809 ;
      RECT 1.735 2.62 2.16 2.761 ;
      RECT 1.735 2.62 2.195 2.73 ;
      RECT 1.965 2.44 2.245 2.72 ;
      RECT 1.8 2.605 2.245 2.72 ;
      RECT 1.89 2.482 1.995 2.88 ;
      RECT 1.82 2.545 2.245 2.72 ;
      RECT 67.24 7.055 67.61 7.425 ;
      RECT 51.98 7.055 52.35 7.425 ;
      RECT 36.72 7.055 37.09 7.425 ;
      RECT 21.46 7.055 21.83 7.425 ;
      RECT 6.2 7.055 6.57 7.425 ;
    LAYER via1 ;
      RECT 75.83 7.375 75.98 7.525 ;
      RECT 73.46 6.74 73.61 6.89 ;
      RECT 73.445 2.065 73.595 2.215 ;
      RECT 72.655 2.45 72.805 2.6 ;
      RECT 72.655 6.325 72.805 6.475 ;
      RECT 71.625 2.805 71.775 2.955 ;
      RECT 71.62 5.96 71.77 6.11 ;
      RECT 71.065 2.805 71.215 2.955 ;
      RECT 69.295 2.35 69.445 2.5 ;
      RECT 68.275 3.055 68.425 3.205 ;
      RECT 68.045 2.475 68.195 2.625 ;
      RECT 68.01 6.71 68.16 6.86 ;
      RECT 67.7 3.075 67.85 3.225 ;
      RECT 67.46 2.095 67.61 2.245 ;
      RECT 67.35 7.165 67.5 7.315 ;
      RECT 67.15 3.425 67.3 3.575 ;
      RECT 67.01 2.03 67.16 2.18 ;
      RECT 66.375 2.115 66.525 2.265 ;
      RECT 66.265 2.755 66.415 2.905 ;
      RECT 65.94 3.315 66.09 3.465 ;
      RECT 65.77 2.305 65.92 2.455 ;
      RECT 65.415 3.32 65.565 3.47 ;
      RECT 65.355 2.535 65.505 2.685 ;
      RECT 64.99 3.525 65.14 3.675 ;
      RECT 64.83 2.36 64.98 2.51 ;
      RECT 64.265 2.435 64.415 2.585 ;
      RECT 63.915 1.055 64.065 1.205 ;
      RECT 63.87 2.385 64.02 2.535 ;
      RECT 63.57 1.97 63.72 2.12 ;
      RECT 63.485 3.525 63.635 3.675 ;
      RECT 62.83 2.675 62.98 2.825 ;
      RECT 60.545 6.755 60.695 6.905 ;
      RECT 58.2 6.74 58.35 6.89 ;
      RECT 58.185 2.065 58.335 2.215 ;
      RECT 57.395 2.45 57.545 2.6 ;
      RECT 57.395 6.325 57.545 6.475 ;
      RECT 56.365 2.805 56.515 2.955 ;
      RECT 56.36 5.96 56.51 6.11 ;
      RECT 55.805 2.805 55.955 2.955 ;
      RECT 54.035 2.35 54.185 2.5 ;
      RECT 53.015 3.055 53.165 3.205 ;
      RECT 52.785 2.475 52.935 2.625 ;
      RECT 52.75 6.71 52.9 6.86 ;
      RECT 52.44 3.075 52.59 3.225 ;
      RECT 52.2 2.095 52.35 2.245 ;
      RECT 52.09 7.165 52.24 7.315 ;
      RECT 51.89 3.425 52.04 3.575 ;
      RECT 51.75 2.03 51.9 2.18 ;
      RECT 51.115 2.115 51.265 2.265 ;
      RECT 51.005 2.755 51.155 2.905 ;
      RECT 50.68 3.315 50.83 3.465 ;
      RECT 50.51 2.305 50.66 2.455 ;
      RECT 50.155 3.32 50.305 3.47 ;
      RECT 50.095 2.535 50.245 2.685 ;
      RECT 49.73 3.525 49.88 3.675 ;
      RECT 49.57 2.36 49.72 2.51 ;
      RECT 49.005 2.435 49.155 2.585 ;
      RECT 48.655 1.055 48.805 1.205 ;
      RECT 48.61 2.385 48.76 2.535 ;
      RECT 48.31 1.97 48.46 2.12 ;
      RECT 48.225 3.525 48.375 3.675 ;
      RECT 47.57 2.675 47.72 2.825 ;
      RECT 45.285 6.755 45.435 6.905 ;
      RECT 42.94 6.74 43.09 6.89 ;
      RECT 42.925 2.065 43.075 2.215 ;
      RECT 42.135 2.45 42.285 2.6 ;
      RECT 42.135 6.325 42.285 6.475 ;
      RECT 41.105 2.805 41.255 2.955 ;
      RECT 41.1 5.96 41.25 6.11 ;
      RECT 40.545 2.805 40.695 2.955 ;
      RECT 38.775 2.35 38.925 2.5 ;
      RECT 37.755 3.055 37.905 3.205 ;
      RECT 37.525 2.475 37.675 2.625 ;
      RECT 37.49 6.715 37.64 6.865 ;
      RECT 37.18 3.075 37.33 3.225 ;
      RECT 36.94 2.095 37.09 2.245 ;
      RECT 36.83 7.165 36.98 7.315 ;
      RECT 36.63 3.425 36.78 3.575 ;
      RECT 36.49 2.03 36.64 2.18 ;
      RECT 35.855 2.115 36.005 2.265 ;
      RECT 35.745 2.755 35.895 2.905 ;
      RECT 35.42 3.315 35.57 3.465 ;
      RECT 35.25 2.305 35.4 2.455 ;
      RECT 34.895 3.32 35.045 3.47 ;
      RECT 34.835 2.535 34.985 2.685 ;
      RECT 34.47 3.525 34.62 3.675 ;
      RECT 34.31 2.36 34.46 2.51 ;
      RECT 33.745 2.435 33.895 2.585 ;
      RECT 33.395 1.055 33.545 1.205 ;
      RECT 33.35 2.385 33.5 2.535 ;
      RECT 33.05 1.97 33.2 2.12 ;
      RECT 32.965 3.525 33.115 3.675 ;
      RECT 32.31 2.675 32.46 2.825 ;
      RECT 30.07 6.76 30.22 6.91 ;
      RECT 27.68 6.74 27.83 6.89 ;
      RECT 27.665 2.065 27.815 2.215 ;
      RECT 26.875 2.45 27.025 2.6 ;
      RECT 26.875 6.325 27.025 6.475 ;
      RECT 25.845 2.805 25.995 2.955 ;
      RECT 25.84 5.96 25.99 6.11 ;
      RECT 25.285 2.805 25.435 2.955 ;
      RECT 23.515 2.35 23.665 2.5 ;
      RECT 22.495 3.055 22.645 3.205 ;
      RECT 22.265 2.475 22.415 2.625 ;
      RECT 22.23 6.71 22.38 6.86 ;
      RECT 21.92 3.075 22.07 3.225 ;
      RECT 21.68 2.095 21.83 2.245 ;
      RECT 21.57 7.165 21.72 7.315 ;
      RECT 21.37 3.425 21.52 3.575 ;
      RECT 21.23 2.03 21.38 2.18 ;
      RECT 20.595 2.115 20.745 2.265 ;
      RECT 20.485 2.755 20.635 2.905 ;
      RECT 20.16 3.315 20.31 3.465 ;
      RECT 19.99 2.305 20.14 2.455 ;
      RECT 19.635 3.32 19.785 3.47 ;
      RECT 19.575 2.535 19.725 2.685 ;
      RECT 19.21 3.525 19.36 3.675 ;
      RECT 19.05 2.36 19.2 2.51 ;
      RECT 18.485 2.435 18.635 2.585 ;
      RECT 18.135 1.055 18.285 1.205 ;
      RECT 18.09 2.385 18.24 2.535 ;
      RECT 17.79 1.97 17.94 2.12 ;
      RECT 17.705 3.525 17.855 3.675 ;
      RECT 17.05 2.675 17.2 2.825 ;
      RECT 14.81 6.755 14.96 6.905 ;
      RECT 12.42 6.74 12.57 6.89 ;
      RECT 12.405 2.065 12.555 2.215 ;
      RECT 11.615 2.45 11.765 2.6 ;
      RECT 11.615 6.325 11.765 6.475 ;
      RECT 10.585 2.805 10.735 2.955 ;
      RECT 10.58 5.96 10.73 6.11 ;
      RECT 10.025 2.805 10.175 2.955 ;
      RECT 8.255 2.35 8.405 2.5 ;
      RECT 7.235 3.055 7.385 3.205 ;
      RECT 7.005 2.475 7.155 2.625 ;
      RECT 6.97 6.705 7.12 6.855 ;
      RECT 6.66 3.075 6.81 3.225 ;
      RECT 6.42 2.095 6.57 2.245 ;
      RECT 6.31 7.165 6.46 7.315 ;
      RECT 6.11 3.425 6.26 3.575 ;
      RECT 5.97 2.03 6.12 2.18 ;
      RECT 5.335 2.115 5.485 2.265 ;
      RECT 5.225 2.755 5.375 2.905 ;
      RECT 4.9 3.315 5.05 3.465 ;
      RECT 4.73 2.305 4.88 2.455 ;
      RECT 4.375 3.32 4.525 3.47 ;
      RECT 4.315 2.535 4.465 2.685 ;
      RECT 3.95 3.525 4.1 3.675 ;
      RECT 3.79 2.36 3.94 2.51 ;
      RECT 3.225 2.435 3.375 2.585 ;
      RECT 2.875 1.055 3.025 1.205 ;
      RECT 2.83 2.385 2.98 2.535 ;
      RECT 2.53 1.97 2.68 2.12 ;
      RECT 2.445 3.525 2.595 3.675 ;
      RECT 1.79 2.675 1.94 2.825 ;
      RECT -1.185 7.095 -1.035 7.245 ;
      RECT -1.56 6.355 -1.41 6.505 ;
    LAYER met1 ;
      RECT 61.79 0 70.53 1.74 ;
      RECT 46.53 0 55.27 1.74 ;
      RECT 31.27 0 40.01 1.74 ;
      RECT 16.01 0 24.75 1.74 ;
      RECT 0.75 0 9.49 1.74 ;
      RECT -2.75 0 76.3 0.305 ;
      RECT -2.75 4.14 76.3 4.745 ;
      RECT 61.79 4.135 76.3 4.745 ;
      RECT 46.53 4.135 61.04 4.745 ;
      RECT 31.27 4.135 45.78 4.745 ;
      RECT 16.01 4.135 30.52 4.745 ;
      RECT 0.75 4.135 15.26 4.745 ;
      RECT 61.79 3.98 70.53 4.745 ;
      RECT 46.53 3.98 55.27 4.745 ;
      RECT 31.27 3.98 40.01 4.745 ;
      RECT 16.01 3.98 24.75 4.745 ;
      RECT 0.75 3.98 9.49 4.745 ;
      RECT -2.75 8.575 76.3 8.88 ;
      RECT 66.735 6.315 66.905 8.88 ;
      RECT 51.475 6.315 51.645 8.88 ;
      RECT 36.215 6.315 36.385 8.88 ;
      RECT 20.955 6.315 21.125 8.88 ;
      RECT 5.695 6.315 5.865 8.88 ;
      RECT 66.905 6.285 67.195 6.515 ;
      RECT 51.645 6.285 51.935 6.515 ;
      RECT 36.385 6.285 36.675 6.515 ;
      RECT 21.125 6.285 21.415 6.515 ;
      RECT 5.865 6.285 6.155 6.515 ;
      RECT 75.7 7.765 75.99 7.995 ;
      RECT 75.76 6.285 75.93 7.995 ;
      RECT 75.73 7.275 76.08 7.625 ;
      RECT 75.7 6.285 75.99 6.515 ;
      RECT 75.7 2.365 75.99 2.595 ;
      RECT 75.76 0.885 75.93 2.595 ;
      RECT 75.7 0.885 75.99 1.115 ;
      RECT 75.29 2.735 75.62 2.965 ;
      RECT 75.29 2.765 75.79 2.935 ;
      RECT 75.29 2.395 75.48 2.965 ;
      RECT 74.71 2.365 75 2.595 ;
      RECT 74.71 2.395 75.48 2.565 ;
      RECT 74.77 0.885 74.94 2.595 ;
      RECT 74.71 0.885 75 1.115 ;
      RECT 74.71 7.765 75 7.995 ;
      RECT 74.77 6.285 74.94 7.995 ;
      RECT 74.71 6.285 75 6.515 ;
      RECT 74.71 6.325 75.56 6.485 ;
      RECT 75.39 5.915 75.56 6.485 ;
      RECT 74.71 6.32 75.1 6.485 ;
      RECT 75.33 5.915 75.62 6.145 ;
      RECT 75.33 5.945 75.79 6.115 ;
      RECT 74.34 2.735 74.63 2.965 ;
      RECT 74.34 2.765 74.8 2.935 ;
      RECT 74.4 1.655 74.565 2.965 ;
      RECT 72.915 1.625 73.205 1.855 ;
      RECT 72.915 1.655 74.565 1.825 ;
      RECT 72.975 0.885 73.145 1.855 ;
      RECT 72.915 0.885 73.205 1.115 ;
      RECT 72.915 7.765 73.205 7.995 ;
      RECT 72.975 7.025 73.145 7.995 ;
      RECT 72.975 7.12 74.565 7.29 ;
      RECT 74.395 5.915 74.565 7.29 ;
      RECT 72.915 7.025 73.205 7.255 ;
      RECT 74.34 5.915 74.63 6.145 ;
      RECT 74.34 5.945 74.8 6.115 ;
      RECT 70.965 2.705 71.305 3.055 ;
      RECT 71.055 2.025 71.225 3.055 ;
      RECT 73.345 1.965 73.695 2.315 ;
      RECT 71.055 2.025 73.695 2.195 ;
      RECT 73.37 6.655 73.695 6.98 ;
      RECT 67.91 6.61 68.26 6.96 ;
      RECT 73.345 6.655 73.695 6.885 ;
      RECT 67.71 6.655 68.26 6.885 ;
      RECT 67.54 6.685 73.695 6.855 ;
      RECT 72.57 2.365 72.89 2.685 ;
      RECT 72.54 2.365 72.89 2.595 ;
      RECT 72.37 2.395 72.89 2.565 ;
      RECT 72.57 6.255 72.89 6.545 ;
      RECT 72.54 6.285 72.89 6.515 ;
      RECT 72.37 6.315 72.89 6.485 ;
      RECT 71.525 2.705 71.865 3.055 ;
      RECT 71.525 2.765 72.005 2.935 ;
      RECT 71.52 5.86 71.86 6.21 ;
      RECT 65.91 5.915 66.2 6.145 ;
      RECT 65.91 5.945 72.005 6.115 ;
      RECT 68.26 2.985 68.41 3.26 ;
      RECT 68.8 2.065 68.805 2.285 ;
      RECT 69.95 2.265 69.965 2.463 ;
      RECT 69.915 2.257 69.95 2.47 ;
      RECT 69.885 2.25 69.915 2.47 ;
      RECT 69.83 2.215 69.885 2.47 ;
      RECT 69.765 2.152 69.83 2.47 ;
      RECT 69.76 2.117 69.765 2.468 ;
      RECT 69.755 2.112 69.76 2.46 ;
      RECT 69.75 2.107 69.755 2.446 ;
      RECT 69.745 2.104 69.75 2.439 ;
      RECT 69.7 2.094 69.745 2.39 ;
      RECT 69.68 2.081 69.7 2.325 ;
      RECT 69.675 2.076 69.68 2.298 ;
      RECT 69.67 2.075 69.675 2.291 ;
      RECT 69.665 2.074 69.67 2.284 ;
      RECT 69.58 2.059 69.665 2.23 ;
      RECT 69.55 2.04 69.58 2.18 ;
      RECT 69.47 2.023 69.55 2.165 ;
      RECT 69.435 2.01 69.47 2.15 ;
      RECT 69.427 2.01 69.435 2.145 ;
      RECT 69.341 2.011 69.427 2.145 ;
      RECT 69.255 2.013 69.341 2.145 ;
      RECT 69.23 2.014 69.255 2.149 ;
      RECT 69.155 2.02 69.23 2.164 ;
      RECT 69.072 2.032 69.155 2.188 ;
      RECT 68.986 2.045 69.072 2.214 ;
      RECT 68.9 2.058 68.986 2.24 ;
      RECT 68.865 2.067 68.9 2.259 ;
      RECT 68.815 2.067 68.865 2.272 ;
      RECT 68.805 2.065 68.815 2.283 ;
      RECT 68.79 2.062 68.8 2.285 ;
      RECT 68.775 2.054 68.79 2.293 ;
      RECT 68.76 2.046 68.775 2.313 ;
      RECT 68.755 2.041 68.76 2.37 ;
      RECT 68.74 2.036 68.755 2.443 ;
      RECT 68.735 2.031 68.74 2.485 ;
      RECT 68.73 2.029 68.735 2.513 ;
      RECT 68.725 2.027 68.73 2.535 ;
      RECT 68.715 2.023 68.725 2.578 ;
      RECT 68.71 2.02 68.715 2.603 ;
      RECT 68.705 2.018 68.71 2.623 ;
      RECT 68.7 2.016 68.705 2.647 ;
      RECT 68.695 2.012 68.7 2.67 ;
      RECT 68.69 2.008 68.695 2.693 ;
      RECT 68.655 1.998 68.69 2.8 ;
      RECT 68.65 1.988 68.655 2.898 ;
      RECT 68.645 1.986 68.65 2.925 ;
      RECT 68.64 1.985 68.645 2.945 ;
      RECT 68.635 1.977 68.64 2.965 ;
      RECT 68.63 1.972 68.635 3 ;
      RECT 68.625 1.97 68.63 3.018 ;
      RECT 68.62 1.97 68.625 3.043 ;
      RECT 68.615 1.97 68.62 3.065 ;
      RECT 68.58 1.97 68.615 3.108 ;
      RECT 68.555 1.97 68.58 3.137 ;
      RECT 68.545 1.97 68.555 2.323 ;
      RECT 68.548 2.38 68.555 3.147 ;
      RECT 68.545 2.437 68.548 3.15 ;
      RECT 68.54 1.97 68.545 2.295 ;
      RECT 68.54 2.487 68.545 3.153 ;
      RECT 68.53 1.97 68.54 2.285 ;
      RECT 68.535 2.54 68.54 3.156 ;
      RECT 68.53 2.625 68.535 3.16 ;
      RECT 68.52 1.97 68.53 2.273 ;
      RECT 68.525 2.672 68.53 3.164 ;
      RECT 68.52 2.747 68.525 3.168 ;
      RECT 68.485 1.97 68.52 2.248 ;
      RECT 68.51 2.83 68.52 3.173 ;
      RECT 68.5 2.897 68.51 3.18 ;
      RECT 68.495 2.925 68.5 3.185 ;
      RECT 68.485 2.938 68.495 3.191 ;
      RECT 68.44 1.97 68.485 2.205 ;
      RECT 68.48 2.943 68.485 3.198 ;
      RECT 68.44 2.96 68.48 3.26 ;
      RECT 68.435 1.972 68.44 2.178 ;
      RECT 68.41 2.98 68.44 3.26 ;
      RECT 68.43 1.977 68.435 2.15 ;
      RECT 68.22 2.989 68.26 3.26 ;
      RECT 68.195 2.997 68.22 3.23 ;
      RECT 68.15 3.005 68.195 3.23 ;
      RECT 68.135 3.01 68.15 3.225 ;
      RECT 68.125 3.01 68.135 3.219 ;
      RECT 68.115 3.017 68.125 3.216 ;
      RECT 68.11 3.055 68.115 3.205 ;
      RECT 68.105 3.117 68.11 3.183 ;
      RECT 69.375 2.992 69.56 3.215 ;
      RECT 69.375 3.007 69.565 3.211 ;
      RECT 69.365 2.28 69.45 3.21 ;
      RECT 69.365 3.007 69.57 3.204 ;
      RECT 69.36 3.015 69.57 3.203 ;
      RECT 69.565 2.735 69.885 3.055 ;
      RECT 69.36 2.907 69.53 2.998 ;
      RECT 69.355 2.907 69.53 2.98 ;
      RECT 69.345 2.715 69.48 2.955 ;
      RECT 69.34 2.715 69.48 2.9 ;
      RECT 69.3 2.295 69.47 2.8 ;
      RECT 69.285 2.295 69.47 2.67 ;
      RECT 69.28 2.295 69.47 2.623 ;
      RECT 69.275 2.295 69.47 2.603 ;
      RECT 69.27 2.295 69.47 2.578 ;
      RECT 69.24 2.295 69.5 2.555 ;
      RECT 69.25 2.292 69.46 2.555 ;
      RECT 69.375 2.287 69.46 3.215 ;
      RECT 69.26 2.28 69.45 2.555 ;
      RECT 69.255 2.285 69.45 2.555 ;
      RECT 68.085 2.497 68.27 2.71 ;
      RECT 68.085 2.505 68.28 2.703 ;
      RECT 68.065 2.505 68.28 2.7 ;
      RECT 68.06 2.505 68.28 2.685 ;
      RECT 67.99 2.42 68.25 2.68 ;
      RECT 67.99 2.565 68.285 2.593 ;
      RECT 67.645 3.02 67.905 3.28 ;
      RECT 67.67 2.965 67.865 3.28 ;
      RECT 67.665 2.714 67.845 3.008 ;
      RECT 67.665 2.72 67.855 3.008 ;
      RECT 67.645 2.722 67.855 2.953 ;
      RECT 67.64 2.732 67.855 2.82 ;
      RECT 67.67 2.712 67.845 3.28 ;
      RECT 67.756 2.71 67.845 3.28 ;
      RECT 67.615 1.93 67.65 2.3 ;
      RECT 67.405 2.04 67.41 2.3 ;
      RECT 67.65 1.937 67.665 2.3 ;
      RECT 67.54 1.93 67.615 2.378 ;
      RECT 67.53 1.93 67.54 2.463 ;
      RECT 67.505 1.93 67.53 2.498 ;
      RECT 67.465 1.93 67.505 2.566 ;
      RECT 67.455 1.937 67.465 2.618 ;
      RECT 67.425 2.04 67.455 2.659 ;
      RECT 67.42 2.04 67.425 2.698 ;
      RECT 67.41 2.04 67.42 2.718 ;
      RECT 67.405 2.335 67.41 2.755 ;
      RECT 67.4 2.352 67.405 2.775 ;
      RECT 67.385 2.415 67.4 2.815 ;
      RECT 67.38 2.458 67.385 2.85 ;
      RECT 67.375 2.466 67.38 2.863 ;
      RECT 67.365 2.48 67.375 2.885 ;
      RECT 67.34 2.515 67.365 2.95 ;
      RECT 67.33 2.55 67.34 3.013 ;
      RECT 67.31 2.58 67.33 3.074 ;
      RECT 67.295 2.616 67.31 3.141 ;
      RECT 67.285 2.644 67.295 3.18 ;
      RECT 67.275 2.666 67.285 3.2 ;
      RECT 67.27 2.676 67.275 3.211 ;
      RECT 67.265 2.685 67.27 3.214 ;
      RECT 67.255 2.703 67.265 3.218 ;
      RECT 67.245 2.721 67.255 3.219 ;
      RECT 67.22 2.76 67.245 3.216 ;
      RECT 67.2 2.802 67.22 3.213 ;
      RECT 67.185 2.84 67.2 3.212 ;
      RECT 67.15 2.875 67.185 3.209 ;
      RECT 67.145 2.897 67.15 3.207 ;
      RECT 67.08 2.937 67.145 3.204 ;
      RECT 67.075 2.977 67.08 3.2 ;
      RECT 67.06 2.987 67.075 3.191 ;
      RECT 67.05 3.107 67.06 3.176 ;
      RECT 67.53 3.52 67.54 3.78 ;
      RECT 67.53 3.523 67.55 3.779 ;
      RECT 67.52 3.513 67.53 3.778 ;
      RECT 67.51 3.528 67.59 3.774 ;
      RECT 67.495 3.507 67.51 3.772 ;
      RECT 67.47 3.532 67.595 3.768 ;
      RECT 67.455 3.492 67.47 3.763 ;
      RECT 67.455 3.534 67.605 3.762 ;
      RECT 67.455 3.542 67.62 3.755 ;
      RECT 67.395 3.479 67.455 3.745 ;
      RECT 67.385 3.466 67.395 3.727 ;
      RECT 67.36 3.456 67.385 3.717 ;
      RECT 67.355 3.446 67.36 3.709 ;
      RECT 67.29 3.542 67.62 3.691 ;
      RECT 67.205 3.542 67.62 3.653 ;
      RECT 67.095 3.37 67.355 3.63 ;
      RECT 67.47 3.5 67.495 3.768 ;
      RECT 67.51 3.51 67.52 3.774 ;
      RECT 67.095 3.518 67.535 3.63 ;
      RECT 67.28 7.765 67.57 7.995 ;
      RECT 67.34 7.025 67.51 7.995 ;
      RECT 67.24 7.055 67.61 7.425 ;
      RECT 67.28 7.025 67.57 7.425 ;
      RECT 66.31 3.275 66.34 3.575 ;
      RECT 66.085 3.26 66.09 3.535 ;
      RECT 65.885 3.26 66.04 3.52 ;
      RECT 67.185 1.975 67.215 2.235 ;
      RECT 67.175 1.975 67.185 2.343 ;
      RECT 67.155 1.975 67.175 2.353 ;
      RECT 67.14 1.975 67.155 2.365 ;
      RECT 67.085 1.975 67.14 2.415 ;
      RECT 67.07 1.975 67.085 2.463 ;
      RECT 67.04 1.975 67.07 2.498 ;
      RECT 66.985 1.975 67.04 2.56 ;
      RECT 66.965 1.975 66.985 2.628 ;
      RECT 66.96 1.975 66.965 2.658 ;
      RECT 66.955 1.975 66.96 2.67 ;
      RECT 66.95 2.092 66.955 2.688 ;
      RECT 66.93 2.11 66.95 2.713 ;
      RECT 66.91 2.137 66.93 2.763 ;
      RECT 66.905 2.157 66.91 2.794 ;
      RECT 66.9 2.165 66.905 2.811 ;
      RECT 66.885 2.191 66.9 2.84 ;
      RECT 66.87 2.233 66.885 2.875 ;
      RECT 66.865 2.262 66.87 2.898 ;
      RECT 66.86 2.277 66.865 2.911 ;
      RECT 66.855 2.3 66.86 2.922 ;
      RECT 66.845 2.32 66.855 2.94 ;
      RECT 66.835 2.35 66.845 2.963 ;
      RECT 66.83 2.372 66.835 2.983 ;
      RECT 66.825 2.387 66.83 2.998 ;
      RECT 66.81 2.417 66.825 3.025 ;
      RECT 66.805 2.447 66.81 3.051 ;
      RECT 66.8 2.465 66.805 3.063 ;
      RECT 66.79 2.495 66.8 3.082 ;
      RECT 66.78 2.52 66.79 3.107 ;
      RECT 66.775 2.54 66.78 3.126 ;
      RECT 66.77 2.557 66.775 3.139 ;
      RECT 66.76 2.583 66.77 3.158 ;
      RECT 66.75 2.621 66.76 3.185 ;
      RECT 66.745 2.647 66.75 3.205 ;
      RECT 66.74 2.657 66.745 3.215 ;
      RECT 66.735 2.67 66.74 3.23 ;
      RECT 66.73 2.685 66.735 3.24 ;
      RECT 66.725 2.707 66.73 3.255 ;
      RECT 66.72 2.725 66.725 3.266 ;
      RECT 66.715 2.735 66.72 3.277 ;
      RECT 66.71 2.743 66.715 3.289 ;
      RECT 66.705 2.751 66.71 3.3 ;
      RECT 66.7 2.777 66.705 3.313 ;
      RECT 66.69 2.805 66.7 3.326 ;
      RECT 66.685 2.835 66.69 3.335 ;
      RECT 66.68 2.85 66.685 3.342 ;
      RECT 66.665 2.875 66.68 3.349 ;
      RECT 66.66 2.897 66.665 3.355 ;
      RECT 66.655 2.922 66.66 3.358 ;
      RECT 66.646 2.95 66.655 3.362 ;
      RECT 66.64 2.967 66.646 3.367 ;
      RECT 66.635 2.985 66.64 3.371 ;
      RECT 66.63 2.997 66.635 3.374 ;
      RECT 66.625 3.018 66.63 3.378 ;
      RECT 66.62 3.036 66.625 3.381 ;
      RECT 66.615 3.05 66.62 3.384 ;
      RECT 66.61 3.067 66.615 3.387 ;
      RECT 66.605 3.08 66.61 3.39 ;
      RECT 66.58 3.117 66.605 3.398 ;
      RECT 66.575 3.162 66.58 3.407 ;
      RECT 66.57 3.19 66.575 3.41 ;
      RECT 66.56 3.21 66.57 3.414 ;
      RECT 66.555 3.23 66.56 3.419 ;
      RECT 66.55 3.245 66.555 3.422 ;
      RECT 66.53 3.255 66.55 3.429 ;
      RECT 66.465 3.262 66.53 3.455 ;
      RECT 66.43 3.265 66.465 3.483 ;
      RECT 66.415 3.268 66.43 3.498 ;
      RECT 66.405 3.269 66.415 3.513 ;
      RECT 66.395 3.27 66.405 3.53 ;
      RECT 66.39 3.27 66.395 3.545 ;
      RECT 66.385 3.27 66.39 3.553 ;
      RECT 66.37 3.271 66.385 3.568 ;
      RECT 66.34 3.273 66.37 3.575 ;
      RECT 66.23 3.28 66.31 3.575 ;
      RECT 66.185 3.285 66.23 3.575 ;
      RECT 66.175 3.286 66.185 3.565 ;
      RECT 66.165 3.287 66.175 3.558 ;
      RECT 66.145 3.289 66.165 3.553 ;
      RECT 66.135 3.26 66.145 3.548 ;
      RECT 66.09 3.26 66.135 3.54 ;
      RECT 66.06 3.26 66.085 3.53 ;
      RECT 66.04 3.26 66.06 3.523 ;
      RECT 66.32 2.06 66.58 2.32 ;
      RECT 66.2 2.075 66.21 2.24 ;
      RECT 66.185 2.075 66.19 2.235 ;
      RECT 63.55 1.915 63.735 2.205 ;
      RECT 65.365 2.04 65.38 2.195 ;
      RECT 63.515 1.915 63.54 2.175 ;
      RECT 65.93 1.965 65.935 2.107 ;
      RECT 65.845 1.96 65.87 2.1 ;
      RECT 66.245 2.077 66.32 2.27 ;
      RECT 66.23 2.075 66.245 2.253 ;
      RECT 66.21 2.075 66.23 2.245 ;
      RECT 66.19 2.075 66.2 2.238 ;
      RECT 66.145 2.07 66.185 2.228 ;
      RECT 66.105 2.045 66.145 2.213 ;
      RECT 66.09 2.02 66.105 2.203 ;
      RECT 66.085 2.014 66.09 2.201 ;
      RECT 66.05 2.006 66.085 2.184 ;
      RECT 66.045 1.999 66.05 2.172 ;
      RECT 66.025 1.994 66.045 2.16 ;
      RECT 66.015 1.988 66.025 2.145 ;
      RECT 65.995 1.983 66.015 2.13 ;
      RECT 65.985 1.978 65.995 2.123 ;
      RECT 65.98 1.976 65.985 2.118 ;
      RECT 65.975 1.975 65.98 2.115 ;
      RECT 65.935 1.97 65.975 2.111 ;
      RECT 65.915 1.964 65.93 2.106 ;
      RECT 65.88 1.961 65.915 2.103 ;
      RECT 65.87 1.96 65.88 2.101 ;
      RECT 65.81 1.96 65.845 2.098 ;
      RECT 65.765 1.96 65.81 2.098 ;
      RECT 65.715 1.96 65.765 2.101 ;
      RECT 65.7 1.962 65.715 2.103 ;
      RECT 65.685 1.965 65.7 2.104 ;
      RECT 65.675 1.97 65.685 2.105 ;
      RECT 65.645 1.975 65.675 2.11 ;
      RECT 65.635 1.981 65.645 2.118 ;
      RECT 65.625 1.983 65.635 2.122 ;
      RECT 65.615 1.987 65.625 2.126 ;
      RECT 65.59 1.993 65.615 2.134 ;
      RECT 65.58 1.998 65.59 2.142 ;
      RECT 65.565 2.002 65.58 2.146 ;
      RECT 65.53 2.008 65.565 2.154 ;
      RECT 65.51 2.013 65.53 2.164 ;
      RECT 65.48 2.02 65.51 2.173 ;
      RECT 65.435 2.029 65.48 2.187 ;
      RECT 65.43 2.034 65.435 2.198 ;
      RECT 65.41 2.037 65.43 2.199 ;
      RECT 65.38 2.04 65.41 2.197 ;
      RECT 65.345 2.04 65.365 2.193 ;
      RECT 65.275 2.04 65.345 2.184 ;
      RECT 65.26 2.037 65.275 2.176 ;
      RECT 65.22 2.03 65.26 2.171 ;
      RECT 65.195 2.02 65.22 2.164 ;
      RECT 65.19 2.014 65.195 2.161 ;
      RECT 65.15 2.008 65.19 2.158 ;
      RECT 65.135 2.001 65.15 2.153 ;
      RECT 65.115 1.997 65.135 2.148 ;
      RECT 65.1 1.992 65.115 2.144 ;
      RECT 65.085 1.987 65.1 2.142 ;
      RECT 65.07 1.983 65.085 2.141 ;
      RECT 65.055 1.981 65.07 2.137 ;
      RECT 65.045 1.979 65.055 2.132 ;
      RECT 65.03 1.976 65.045 2.128 ;
      RECT 65.02 1.974 65.03 2.123 ;
      RECT 65 1.971 65.02 2.119 ;
      RECT 64.955 1.97 65 2.117 ;
      RECT 64.895 1.972 64.955 2.118 ;
      RECT 64.875 1.974 64.895 2.12 ;
      RECT 64.845 1.977 64.875 2.121 ;
      RECT 64.795 1.982 64.845 2.123 ;
      RECT 64.79 1.985 64.795 2.125 ;
      RECT 64.78 1.987 64.79 2.128 ;
      RECT 64.775 1.989 64.78 2.131 ;
      RECT 64.725 1.992 64.775 2.138 ;
      RECT 64.705 1.996 64.725 2.15 ;
      RECT 64.695 1.999 64.705 2.156 ;
      RECT 64.685 2 64.695 2.159 ;
      RECT 64.646 2.003 64.685 2.161 ;
      RECT 64.56 2.01 64.646 2.164 ;
      RECT 64.486 2.02 64.56 2.168 ;
      RECT 64.4 2.031 64.486 2.173 ;
      RECT 64.385 2.038 64.4 2.175 ;
      RECT 64.33 2.042 64.385 2.176 ;
      RECT 64.316 2.045 64.33 2.178 ;
      RECT 64.23 2.045 64.316 2.18 ;
      RECT 64.19 2.042 64.23 2.183 ;
      RECT 64.166 2.038 64.19 2.185 ;
      RECT 64.08 2.028 64.166 2.188 ;
      RECT 64.05 2.017 64.08 2.189 ;
      RECT 64.031 2.013 64.05 2.188 ;
      RECT 63.945 2.006 64.031 2.185 ;
      RECT 63.885 1.995 63.945 2.182 ;
      RECT 63.865 1.987 63.885 2.18 ;
      RECT 63.83 1.982 63.865 2.179 ;
      RECT 63.805 1.977 63.83 2.178 ;
      RECT 63.775 1.972 63.805 2.177 ;
      RECT 63.75 1.915 63.775 2.176 ;
      RECT 63.735 1.915 63.75 2.2 ;
      RECT 63.54 1.915 63.55 2.2 ;
      RECT 65.315 2.935 65.32 3.075 ;
      RECT 64.975 2.935 65.01 3.073 ;
      RECT 64.55 2.92 64.565 3.065 ;
      RECT 66.38 2.7 66.47 2.96 ;
      RECT 66.21 2.565 66.31 2.96 ;
      RECT 63.245 2.54 63.325 2.75 ;
      RECT 66.335 2.677 66.38 2.96 ;
      RECT 66.325 2.647 66.335 2.96 ;
      RECT 66.31 2.57 66.325 2.96 ;
      RECT 66.125 2.565 66.21 2.925 ;
      RECT 66.12 2.567 66.125 2.92 ;
      RECT 66.115 2.572 66.12 2.92 ;
      RECT 66.08 2.672 66.115 2.92 ;
      RECT 66.07 2.7 66.08 2.92 ;
      RECT 66.06 2.715 66.07 2.92 ;
      RECT 66.05 2.727 66.06 2.92 ;
      RECT 66.045 2.737 66.05 2.92 ;
      RECT 66.03 2.747 66.045 2.922 ;
      RECT 66.025 2.762 66.03 2.924 ;
      RECT 66.01 2.775 66.025 2.926 ;
      RECT 66.005 2.79 66.01 2.929 ;
      RECT 65.985 2.8 66.005 2.933 ;
      RECT 65.97 2.81 65.985 2.936 ;
      RECT 65.935 2.817 65.97 2.941 ;
      RECT 65.891 2.824 65.935 2.949 ;
      RECT 65.805 2.836 65.891 2.962 ;
      RECT 65.78 2.847 65.805 2.973 ;
      RECT 65.75 2.852 65.78 2.978 ;
      RECT 65.715 2.857 65.75 2.986 ;
      RECT 65.685 2.862 65.715 2.993 ;
      RECT 65.66 2.867 65.685 2.998 ;
      RECT 65.595 2.874 65.66 3.007 ;
      RECT 65.525 2.887 65.595 3.023 ;
      RECT 65.495 2.897 65.525 3.035 ;
      RECT 65.47 2.902 65.495 3.042 ;
      RECT 65.415 2.909 65.47 3.05 ;
      RECT 65.41 2.916 65.415 3.055 ;
      RECT 65.405 2.918 65.41 3.056 ;
      RECT 65.39 2.92 65.405 3.058 ;
      RECT 65.385 2.92 65.39 3.061 ;
      RECT 65.32 2.927 65.385 3.068 ;
      RECT 65.285 2.937 65.315 3.078 ;
      RECT 65.268 2.94 65.285 3.08 ;
      RECT 65.182 2.939 65.268 3.079 ;
      RECT 65.096 2.937 65.182 3.076 ;
      RECT 65.01 2.936 65.096 3.074 ;
      RECT 64.909 2.934 64.975 3.073 ;
      RECT 64.823 2.931 64.909 3.071 ;
      RECT 64.737 2.927 64.823 3.069 ;
      RECT 64.651 2.924 64.737 3.068 ;
      RECT 64.565 2.921 64.651 3.066 ;
      RECT 64.465 2.92 64.55 3.063 ;
      RECT 64.415 2.918 64.465 3.061 ;
      RECT 64.395 2.915 64.415 3.059 ;
      RECT 64.375 2.913 64.395 3.056 ;
      RECT 64.35 2.909 64.375 3.053 ;
      RECT 64.305 2.903 64.35 3.048 ;
      RECT 64.265 2.897 64.305 3.04 ;
      RECT 64.24 2.892 64.265 3.033 ;
      RECT 64.185 2.885 64.24 3.025 ;
      RECT 64.161 2.878 64.185 3.018 ;
      RECT 64.075 2.869 64.161 3.008 ;
      RECT 64.045 2.861 64.075 2.998 ;
      RECT 64.015 2.857 64.045 2.993 ;
      RECT 64.01 2.854 64.015 2.99 ;
      RECT 64.005 2.853 64.01 2.99 ;
      RECT 63.93 2.846 64.005 2.983 ;
      RECT 63.891 2.837 63.93 2.972 ;
      RECT 63.805 2.827 63.891 2.96 ;
      RECT 63.765 2.817 63.805 2.948 ;
      RECT 63.726 2.812 63.765 2.941 ;
      RECT 63.64 2.802 63.726 2.93 ;
      RECT 63.6 2.79 63.64 2.919 ;
      RECT 63.565 2.775 63.6 2.912 ;
      RECT 63.555 2.765 63.565 2.909 ;
      RECT 63.535 2.75 63.555 2.907 ;
      RECT 63.505 2.72 63.535 2.903 ;
      RECT 63.495 2.7 63.505 2.898 ;
      RECT 63.49 2.692 63.495 2.895 ;
      RECT 63.485 2.685 63.49 2.893 ;
      RECT 63.47 2.672 63.485 2.886 ;
      RECT 63.465 2.662 63.47 2.878 ;
      RECT 63.46 2.655 63.465 2.873 ;
      RECT 63.455 2.65 63.46 2.869 ;
      RECT 63.44 2.637 63.455 2.861 ;
      RECT 63.435 2.547 63.44 2.85 ;
      RECT 63.43 2.542 63.435 2.843 ;
      RECT 63.355 2.54 63.43 2.803 ;
      RECT 63.325 2.54 63.355 2.758 ;
      RECT 63.23 2.545 63.245 2.745 ;
      RECT 65.715 2.25 65.975 2.51 ;
      RECT 65.7 2.238 65.88 2.475 ;
      RECT 65.695 2.239 65.88 2.473 ;
      RECT 65.68 2.243 65.89 2.463 ;
      RECT 65.675 2.248 65.895 2.433 ;
      RECT 65.68 2.245 65.895 2.463 ;
      RECT 65.695 2.24 65.89 2.473 ;
      RECT 65.715 2.237 65.88 2.51 ;
      RECT 65.715 2.236 65.87 2.51 ;
      RECT 65.74 2.235 65.87 2.51 ;
      RECT 65.3 2.48 65.56 2.74 ;
      RECT 65.175 2.525 65.56 2.735 ;
      RECT 65.165 2.53 65.56 2.73 ;
      RECT 65.18 3.47 65.195 3.78 ;
      RECT 63.775 3.24 63.785 3.37 ;
      RECT 63.555 3.235 63.66 3.37 ;
      RECT 63.47 3.24 63.52 3.37 ;
      RECT 62.02 1.975 62.025 3.08 ;
      RECT 65.275 3.562 65.28 3.698 ;
      RECT 65.27 3.557 65.275 3.758 ;
      RECT 65.265 3.555 65.27 3.771 ;
      RECT 65.25 3.552 65.265 3.773 ;
      RECT 65.245 3.547 65.25 3.775 ;
      RECT 65.24 3.543 65.245 3.778 ;
      RECT 65.225 3.538 65.24 3.78 ;
      RECT 65.195 3.53 65.225 3.78 ;
      RECT 65.156 3.47 65.18 3.78 ;
      RECT 65.07 3.47 65.156 3.777 ;
      RECT 65.04 3.47 65.07 3.77 ;
      RECT 65.015 3.47 65.04 3.763 ;
      RECT 64.99 3.47 65.015 3.755 ;
      RECT 64.975 3.47 64.99 3.748 ;
      RECT 64.95 3.47 64.975 3.74 ;
      RECT 64.935 3.47 64.95 3.733 ;
      RECT 64.895 3.48 64.935 3.722 ;
      RECT 64.885 3.475 64.895 3.712 ;
      RECT 64.881 3.474 64.885 3.709 ;
      RECT 64.795 3.466 64.881 3.692 ;
      RECT 64.762 3.455 64.795 3.669 ;
      RECT 64.676 3.444 64.762 3.647 ;
      RECT 64.59 3.428 64.676 3.616 ;
      RECT 64.52 3.413 64.59 3.588 ;
      RECT 64.51 3.406 64.52 3.575 ;
      RECT 64.48 3.403 64.51 3.565 ;
      RECT 64.455 3.399 64.48 3.558 ;
      RECT 64.44 3.396 64.455 3.553 ;
      RECT 64.435 3.395 64.44 3.548 ;
      RECT 64.405 3.39 64.435 3.541 ;
      RECT 64.4 3.385 64.405 3.536 ;
      RECT 64.385 3.382 64.4 3.531 ;
      RECT 64.38 3.377 64.385 3.526 ;
      RECT 64.36 3.372 64.38 3.523 ;
      RECT 64.345 3.367 64.36 3.515 ;
      RECT 64.33 3.361 64.345 3.51 ;
      RECT 64.3 3.352 64.33 3.503 ;
      RECT 64.295 3.345 64.3 3.495 ;
      RECT 64.29 3.343 64.295 3.493 ;
      RECT 64.285 3.342 64.29 3.49 ;
      RECT 64.245 3.335 64.285 3.483 ;
      RECT 64.231 3.325 64.245 3.473 ;
      RECT 64.18 3.314 64.231 3.461 ;
      RECT 64.155 3.3 64.18 3.447 ;
      RECT 64.13 3.289 64.155 3.439 ;
      RECT 64.11 3.278 64.13 3.433 ;
      RECT 64.1 3.272 64.11 3.428 ;
      RECT 64.095 3.27 64.1 3.424 ;
      RECT 64.075 3.265 64.095 3.419 ;
      RECT 64.045 3.255 64.075 3.409 ;
      RECT 64.04 3.247 64.045 3.402 ;
      RECT 64.025 3.245 64.04 3.398 ;
      RECT 64.005 3.245 64.025 3.393 ;
      RECT 64 3.244 64.005 3.391 ;
      RECT 63.995 3.244 64 3.388 ;
      RECT 63.955 3.243 63.995 3.383 ;
      RECT 63.93 3.242 63.955 3.378 ;
      RECT 63.87 3.241 63.93 3.375 ;
      RECT 63.785 3.24 63.87 3.373 ;
      RECT 63.746 3.239 63.775 3.37 ;
      RECT 63.66 3.237 63.746 3.37 ;
      RECT 63.52 3.237 63.555 3.37 ;
      RECT 63.43 3.241 63.47 3.373 ;
      RECT 63.415 3.244 63.43 3.38 ;
      RECT 63.405 3.245 63.415 3.387 ;
      RECT 63.38 3.248 63.405 3.392 ;
      RECT 63.375 3.25 63.38 3.395 ;
      RECT 63.325 3.252 63.375 3.396 ;
      RECT 63.286 3.256 63.325 3.398 ;
      RECT 63.2 3.258 63.286 3.401 ;
      RECT 63.182 3.26 63.2 3.403 ;
      RECT 63.096 3.263 63.182 3.405 ;
      RECT 63.01 3.267 63.096 3.408 ;
      RECT 62.973 3.271 63.01 3.411 ;
      RECT 62.887 3.274 62.973 3.414 ;
      RECT 62.801 3.278 62.887 3.417 ;
      RECT 62.715 3.283 62.801 3.421 ;
      RECT 62.695 3.285 62.715 3.424 ;
      RECT 62.675 3.284 62.695 3.425 ;
      RECT 62.626 3.281 62.675 3.426 ;
      RECT 62.54 3.276 62.626 3.429 ;
      RECT 62.49 3.271 62.54 3.431 ;
      RECT 62.466 3.269 62.49 3.432 ;
      RECT 62.38 3.264 62.466 3.434 ;
      RECT 62.355 3.26 62.38 3.433 ;
      RECT 62.345 3.257 62.355 3.431 ;
      RECT 62.335 3.25 62.345 3.428 ;
      RECT 62.33 3.23 62.335 3.423 ;
      RECT 62.32 3.2 62.33 3.418 ;
      RECT 62.305 3.07 62.32 3.409 ;
      RECT 62.3 3.062 62.305 3.402 ;
      RECT 62.28 3.055 62.3 3.394 ;
      RECT 62.275 3.037 62.28 3.386 ;
      RECT 62.265 3.017 62.275 3.381 ;
      RECT 62.26 2.99 62.265 3.377 ;
      RECT 62.255 2.967 62.26 3.374 ;
      RECT 62.235 2.925 62.255 3.366 ;
      RECT 62.2 2.84 62.235 3.35 ;
      RECT 62.195 2.772 62.2 3.338 ;
      RECT 62.18 2.742 62.195 3.332 ;
      RECT 62.175 1.987 62.18 2.233 ;
      RECT 62.165 2.712 62.18 3.323 ;
      RECT 62.17 1.982 62.175 2.265 ;
      RECT 62.165 1.977 62.17 2.308 ;
      RECT 62.16 1.975 62.165 2.343 ;
      RECT 62.145 2.675 62.165 3.313 ;
      RECT 62.155 1.975 62.16 2.38 ;
      RECT 62.14 1.975 62.155 2.478 ;
      RECT 62.14 2.648 62.145 3.306 ;
      RECT 62.135 1.975 62.14 2.553 ;
      RECT 62.135 2.636 62.14 3.303 ;
      RECT 62.13 1.975 62.135 2.585 ;
      RECT 62.13 2.615 62.135 3.3 ;
      RECT 62.125 1.975 62.13 3.297 ;
      RECT 62.09 1.975 62.125 3.283 ;
      RECT 62.075 1.975 62.09 3.265 ;
      RECT 62.055 1.975 62.075 3.255 ;
      RECT 62.03 1.975 62.055 3.238 ;
      RECT 62.025 1.975 62.03 3.188 ;
      RECT 62.015 1.975 62.02 3.018 ;
      RECT 62.01 1.975 62.015 2.925 ;
      RECT 62.005 1.975 62.01 2.838 ;
      RECT 62 1.975 62.005 2.77 ;
      RECT 61.995 1.975 62 2.713 ;
      RECT 61.985 1.975 61.995 2.608 ;
      RECT 61.98 1.975 61.985 2.48 ;
      RECT 61.975 1.975 61.98 2.398 ;
      RECT 61.97 1.977 61.975 2.315 ;
      RECT 61.965 1.982 61.97 2.248 ;
      RECT 61.96 1.987 61.965 2.175 ;
      RECT 64.775 2.305 65.035 2.565 ;
      RECT 64.795 2.272 65.005 2.565 ;
      RECT 64.795 2.27 64.995 2.565 ;
      RECT 64.805 2.257 64.995 2.565 ;
      RECT 64.805 2.255 64.92 2.565 ;
      RECT 64.28 2.38 64.455 2.66 ;
      RECT 64.275 2.38 64.455 2.658 ;
      RECT 64.275 2.38 64.47 2.655 ;
      RECT 64.265 2.38 64.47 2.653 ;
      RECT 64.21 2.38 64.47 2.64 ;
      RECT 64.21 2.455 64.475 2.618 ;
      RECT 63.755 2.392 63.775 2.635 ;
      RECT 63.755 2.392 63.815 2.634 ;
      RECT 63.75 2.394 63.815 2.633 ;
      RECT 63.75 2.394 63.901 2.632 ;
      RECT 63.75 2.394 63.97 2.631 ;
      RECT 63.75 2.394 63.99 2.623 ;
      RECT 63.73 2.397 63.99 2.621 ;
      RECT 63.715 2.407 63.99 2.606 ;
      RECT 63.715 2.407 64.005 2.605 ;
      RECT 63.71 2.416 64.005 2.597 ;
      RECT 63.71 2.416 64.01 2.593 ;
      RECT 63.815 2.33 64.075 2.59 ;
      RECT 63.705 2.418 64.075 2.475 ;
      RECT 63.775 2.385 64.075 2.59 ;
      RECT 63.74 3.578 63.745 3.785 ;
      RECT 63.69 3.572 63.74 3.784 ;
      RECT 63.657 3.586 63.75 3.783 ;
      RECT 63.571 3.586 63.75 3.782 ;
      RECT 63.485 3.586 63.75 3.781 ;
      RECT 63.485 3.685 63.755 3.778 ;
      RECT 63.48 3.685 63.755 3.773 ;
      RECT 63.475 3.685 63.755 3.755 ;
      RECT 63.47 3.685 63.755 3.738 ;
      RECT 63.43 3.47 63.69 3.73 ;
      RECT 62.89 2.62 62.976 3.034 ;
      RECT 62.89 2.62 63.015 3.031 ;
      RECT 62.89 2.62 63.035 3.021 ;
      RECT 62.845 2.62 63.035 3.018 ;
      RECT 62.845 2.772 63.045 3.008 ;
      RECT 62.845 2.793 63.05 3.002 ;
      RECT 62.845 2.811 63.055 2.998 ;
      RECT 62.845 2.831 63.065 2.993 ;
      RECT 62.82 2.831 63.065 2.99 ;
      RECT 62.81 2.831 63.065 2.968 ;
      RECT 62.81 2.847 63.07 2.938 ;
      RECT 62.775 2.62 63.035 2.925 ;
      RECT 62.775 2.859 63.075 2.88 ;
      RECT 60.44 7.765 60.73 7.995 ;
      RECT 60.5 6.285 60.67 7.995 ;
      RECT 60.445 6.655 60.795 7.005 ;
      RECT 60.44 6.285 60.73 6.515 ;
      RECT 60.44 2.365 60.73 2.595 ;
      RECT 60.5 0.885 60.67 2.595 ;
      RECT 60.44 0.885 60.73 1.115 ;
      RECT 60.03 2.735 60.36 2.965 ;
      RECT 60.03 2.765 60.53 2.935 ;
      RECT 60.03 2.395 60.22 2.965 ;
      RECT 59.45 2.365 59.74 2.595 ;
      RECT 59.45 2.395 60.22 2.565 ;
      RECT 59.51 0.885 59.68 2.595 ;
      RECT 59.45 0.885 59.74 1.115 ;
      RECT 59.45 7.765 59.74 7.995 ;
      RECT 59.51 6.285 59.68 7.995 ;
      RECT 59.45 6.285 59.74 6.515 ;
      RECT 59.45 6.325 60.3 6.485 ;
      RECT 60.13 5.915 60.3 6.485 ;
      RECT 59.45 6.32 59.84 6.485 ;
      RECT 60.07 5.915 60.36 6.145 ;
      RECT 60.07 5.945 60.53 6.115 ;
      RECT 59.08 2.735 59.37 2.965 ;
      RECT 59.08 2.765 59.54 2.935 ;
      RECT 59.14 1.655 59.305 2.965 ;
      RECT 57.655 1.625 57.945 1.855 ;
      RECT 57.655 1.655 59.305 1.825 ;
      RECT 57.715 0.885 57.885 1.855 ;
      RECT 57.655 0.885 57.945 1.115 ;
      RECT 57.655 7.765 57.945 7.995 ;
      RECT 57.715 7.025 57.885 7.995 ;
      RECT 57.715 7.12 59.305 7.29 ;
      RECT 59.135 5.915 59.305 7.29 ;
      RECT 57.655 7.025 57.945 7.255 ;
      RECT 59.08 5.915 59.37 6.145 ;
      RECT 59.08 5.945 59.54 6.115 ;
      RECT 55.705 2.705 56.045 3.055 ;
      RECT 55.795 2.025 55.965 3.055 ;
      RECT 58.085 1.965 58.435 2.315 ;
      RECT 55.795 2.025 58.435 2.195 ;
      RECT 58.11 6.655 58.435 6.98 ;
      RECT 52.65 6.61 53 6.96 ;
      RECT 58.085 6.655 58.435 6.885 ;
      RECT 52.45 6.655 53 6.885 ;
      RECT 52.28 6.685 58.435 6.855 ;
      RECT 57.31 2.365 57.63 2.685 ;
      RECT 57.28 2.365 57.63 2.595 ;
      RECT 57.11 2.395 57.63 2.565 ;
      RECT 57.31 6.255 57.63 6.545 ;
      RECT 57.28 6.285 57.63 6.515 ;
      RECT 57.11 6.315 57.63 6.485 ;
      RECT 56.265 2.705 56.605 3.055 ;
      RECT 56.265 2.765 56.745 2.935 ;
      RECT 56.26 5.86 56.6 6.21 ;
      RECT 50.65 5.915 50.94 6.145 ;
      RECT 50.65 5.945 56.745 6.115 ;
      RECT 53 2.985 53.15 3.26 ;
      RECT 53.54 2.065 53.545 2.285 ;
      RECT 54.69 2.265 54.705 2.463 ;
      RECT 54.655 2.257 54.69 2.47 ;
      RECT 54.625 2.25 54.655 2.47 ;
      RECT 54.57 2.215 54.625 2.47 ;
      RECT 54.505 2.152 54.57 2.47 ;
      RECT 54.5 2.117 54.505 2.468 ;
      RECT 54.495 2.112 54.5 2.46 ;
      RECT 54.49 2.107 54.495 2.446 ;
      RECT 54.485 2.104 54.49 2.439 ;
      RECT 54.44 2.094 54.485 2.39 ;
      RECT 54.42 2.081 54.44 2.325 ;
      RECT 54.415 2.076 54.42 2.298 ;
      RECT 54.41 2.075 54.415 2.291 ;
      RECT 54.405 2.074 54.41 2.284 ;
      RECT 54.32 2.059 54.405 2.23 ;
      RECT 54.29 2.04 54.32 2.18 ;
      RECT 54.21 2.023 54.29 2.165 ;
      RECT 54.175 2.01 54.21 2.15 ;
      RECT 54.167 2.01 54.175 2.145 ;
      RECT 54.081 2.011 54.167 2.145 ;
      RECT 53.995 2.013 54.081 2.145 ;
      RECT 53.97 2.014 53.995 2.149 ;
      RECT 53.895 2.02 53.97 2.164 ;
      RECT 53.812 2.032 53.895 2.188 ;
      RECT 53.726 2.045 53.812 2.214 ;
      RECT 53.64 2.058 53.726 2.24 ;
      RECT 53.605 2.067 53.64 2.259 ;
      RECT 53.555 2.067 53.605 2.272 ;
      RECT 53.545 2.065 53.555 2.283 ;
      RECT 53.53 2.062 53.54 2.285 ;
      RECT 53.515 2.054 53.53 2.293 ;
      RECT 53.5 2.046 53.515 2.313 ;
      RECT 53.495 2.041 53.5 2.37 ;
      RECT 53.48 2.036 53.495 2.443 ;
      RECT 53.475 2.031 53.48 2.485 ;
      RECT 53.47 2.029 53.475 2.513 ;
      RECT 53.465 2.027 53.47 2.535 ;
      RECT 53.455 2.023 53.465 2.578 ;
      RECT 53.45 2.02 53.455 2.603 ;
      RECT 53.445 2.018 53.45 2.623 ;
      RECT 53.44 2.016 53.445 2.647 ;
      RECT 53.435 2.012 53.44 2.67 ;
      RECT 53.43 2.008 53.435 2.693 ;
      RECT 53.395 1.998 53.43 2.8 ;
      RECT 53.39 1.988 53.395 2.898 ;
      RECT 53.385 1.986 53.39 2.925 ;
      RECT 53.38 1.985 53.385 2.945 ;
      RECT 53.375 1.977 53.38 2.965 ;
      RECT 53.37 1.972 53.375 3 ;
      RECT 53.365 1.97 53.37 3.018 ;
      RECT 53.36 1.97 53.365 3.043 ;
      RECT 53.355 1.97 53.36 3.065 ;
      RECT 53.32 1.97 53.355 3.108 ;
      RECT 53.295 1.97 53.32 3.137 ;
      RECT 53.285 1.97 53.295 2.323 ;
      RECT 53.288 2.38 53.295 3.147 ;
      RECT 53.285 2.437 53.288 3.15 ;
      RECT 53.28 1.97 53.285 2.295 ;
      RECT 53.28 2.487 53.285 3.153 ;
      RECT 53.27 1.97 53.28 2.285 ;
      RECT 53.275 2.54 53.28 3.156 ;
      RECT 53.27 2.625 53.275 3.16 ;
      RECT 53.26 1.97 53.27 2.273 ;
      RECT 53.265 2.672 53.27 3.164 ;
      RECT 53.26 2.747 53.265 3.168 ;
      RECT 53.225 1.97 53.26 2.248 ;
      RECT 53.25 2.83 53.26 3.173 ;
      RECT 53.24 2.897 53.25 3.18 ;
      RECT 53.235 2.925 53.24 3.185 ;
      RECT 53.225 2.938 53.235 3.191 ;
      RECT 53.18 1.97 53.225 2.205 ;
      RECT 53.22 2.943 53.225 3.198 ;
      RECT 53.18 2.96 53.22 3.26 ;
      RECT 53.175 1.972 53.18 2.178 ;
      RECT 53.15 2.98 53.18 3.26 ;
      RECT 53.17 1.977 53.175 2.15 ;
      RECT 52.96 2.989 53 3.26 ;
      RECT 52.935 2.997 52.96 3.23 ;
      RECT 52.89 3.005 52.935 3.23 ;
      RECT 52.875 3.01 52.89 3.225 ;
      RECT 52.865 3.01 52.875 3.219 ;
      RECT 52.855 3.017 52.865 3.216 ;
      RECT 52.85 3.055 52.855 3.205 ;
      RECT 52.845 3.117 52.85 3.183 ;
      RECT 54.115 2.992 54.3 3.215 ;
      RECT 54.115 3.007 54.305 3.211 ;
      RECT 54.105 2.28 54.19 3.21 ;
      RECT 54.105 3.007 54.31 3.204 ;
      RECT 54.1 3.015 54.31 3.203 ;
      RECT 54.305 2.735 54.625 3.055 ;
      RECT 54.1 2.907 54.27 2.998 ;
      RECT 54.095 2.907 54.27 2.98 ;
      RECT 54.085 2.715 54.22 2.955 ;
      RECT 54.08 2.715 54.22 2.9 ;
      RECT 54.04 2.295 54.21 2.8 ;
      RECT 54.025 2.295 54.21 2.67 ;
      RECT 54.02 2.295 54.21 2.623 ;
      RECT 54.015 2.295 54.21 2.603 ;
      RECT 54.01 2.295 54.21 2.578 ;
      RECT 53.98 2.295 54.24 2.555 ;
      RECT 53.99 2.292 54.2 2.555 ;
      RECT 54.115 2.287 54.2 3.215 ;
      RECT 54 2.28 54.19 2.555 ;
      RECT 53.995 2.285 54.19 2.555 ;
      RECT 52.825 2.497 53.01 2.71 ;
      RECT 52.825 2.505 53.02 2.703 ;
      RECT 52.805 2.505 53.02 2.7 ;
      RECT 52.8 2.505 53.02 2.685 ;
      RECT 52.73 2.42 52.99 2.68 ;
      RECT 52.73 2.565 53.025 2.593 ;
      RECT 52.385 3.02 52.645 3.28 ;
      RECT 52.41 2.965 52.605 3.28 ;
      RECT 52.405 2.714 52.585 3.008 ;
      RECT 52.405 2.72 52.595 3.008 ;
      RECT 52.385 2.722 52.595 2.953 ;
      RECT 52.38 2.732 52.595 2.82 ;
      RECT 52.41 2.712 52.585 3.28 ;
      RECT 52.496 2.71 52.585 3.28 ;
      RECT 52.355 1.93 52.39 2.3 ;
      RECT 52.145 2.04 52.15 2.3 ;
      RECT 52.39 1.937 52.405 2.3 ;
      RECT 52.28 1.93 52.355 2.378 ;
      RECT 52.27 1.93 52.28 2.463 ;
      RECT 52.245 1.93 52.27 2.498 ;
      RECT 52.205 1.93 52.245 2.566 ;
      RECT 52.195 1.937 52.205 2.618 ;
      RECT 52.165 2.04 52.195 2.659 ;
      RECT 52.16 2.04 52.165 2.698 ;
      RECT 52.15 2.04 52.16 2.718 ;
      RECT 52.145 2.335 52.15 2.755 ;
      RECT 52.14 2.352 52.145 2.775 ;
      RECT 52.125 2.415 52.14 2.815 ;
      RECT 52.12 2.458 52.125 2.85 ;
      RECT 52.115 2.466 52.12 2.863 ;
      RECT 52.105 2.48 52.115 2.885 ;
      RECT 52.08 2.515 52.105 2.95 ;
      RECT 52.07 2.55 52.08 3.013 ;
      RECT 52.05 2.58 52.07 3.074 ;
      RECT 52.035 2.616 52.05 3.141 ;
      RECT 52.025 2.644 52.035 3.18 ;
      RECT 52.015 2.666 52.025 3.2 ;
      RECT 52.01 2.676 52.015 3.211 ;
      RECT 52.005 2.685 52.01 3.214 ;
      RECT 51.995 2.703 52.005 3.218 ;
      RECT 51.985 2.721 51.995 3.219 ;
      RECT 51.96 2.76 51.985 3.216 ;
      RECT 51.94 2.802 51.96 3.213 ;
      RECT 51.925 2.84 51.94 3.212 ;
      RECT 51.89 2.875 51.925 3.209 ;
      RECT 51.885 2.897 51.89 3.207 ;
      RECT 51.82 2.937 51.885 3.204 ;
      RECT 51.815 2.977 51.82 3.2 ;
      RECT 51.8 2.987 51.815 3.191 ;
      RECT 51.79 3.107 51.8 3.176 ;
      RECT 52.27 3.52 52.28 3.78 ;
      RECT 52.27 3.523 52.29 3.779 ;
      RECT 52.26 3.513 52.27 3.778 ;
      RECT 52.25 3.528 52.33 3.774 ;
      RECT 52.235 3.507 52.25 3.772 ;
      RECT 52.21 3.532 52.335 3.768 ;
      RECT 52.195 3.492 52.21 3.763 ;
      RECT 52.195 3.534 52.345 3.762 ;
      RECT 52.195 3.542 52.36 3.755 ;
      RECT 52.135 3.479 52.195 3.745 ;
      RECT 52.125 3.466 52.135 3.727 ;
      RECT 52.1 3.456 52.125 3.717 ;
      RECT 52.095 3.446 52.1 3.709 ;
      RECT 52.03 3.542 52.36 3.691 ;
      RECT 51.945 3.542 52.36 3.653 ;
      RECT 51.835 3.37 52.095 3.63 ;
      RECT 52.21 3.5 52.235 3.768 ;
      RECT 52.25 3.51 52.26 3.774 ;
      RECT 51.835 3.518 52.275 3.63 ;
      RECT 52.02 7.765 52.31 7.995 ;
      RECT 52.08 7.025 52.25 7.995 ;
      RECT 51.98 7.055 52.35 7.425 ;
      RECT 52.02 7.025 52.31 7.425 ;
      RECT 51.05 3.275 51.08 3.575 ;
      RECT 50.825 3.26 50.83 3.535 ;
      RECT 50.625 3.26 50.78 3.52 ;
      RECT 51.925 1.975 51.955 2.235 ;
      RECT 51.915 1.975 51.925 2.343 ;
      RECT 51.895 1.975 51.915 2.353 ;
      RECT 51.88 1.975 51.895 2.365 ;
      RECT 51.825 1.975 51.88 2.415 ;
      RECT 51.81 1.975 51.825 2.463 ;
      RECT 51.78 1.975 51.81 2.498 ;
      RECT 51.725 1.975 51.78 2.56 ;
      RECT 51.705 1.975 51.725 2.628 ;
      RECT 51.7 1.975 51.705 2.658 ;
      RECT 51.695 1.975 51.7 2.67 ;
      RECT 51.69 2.092 51.695 2.688 ;
      RECT 51.67 2.11 51.69 2.713 ;
      RECT 51.65 2.137 51.67 2.763 ;
      RECT 51.645 2.157 51.65 2.794 ;
      RECT 51.64 2.165 51.645 2.811 ;
      RECT 51.625 2.191 51.64 2.84 ;
      RECT 51.61 2.233 51.625 2.875 ;
      RECT 51.605 2.262 51.61 2.898 ;
      RECT 51.6 2.277 51.605 2.911 ;
      RECT 51.595 2.3 51.6 2.922 ;
      RECT 51.585 2.32 51.595 2.94 ;
      RECT 51.575 2.35 51.585 2.963 ;
      RECT 51.57 2.372 51.575 2.983 ;
      RECT 51.565 2.387 51.57 2.998 ;
      RECT 51.55 2.417 51.565 3.025 ;
      RECT 51.545 2.447 51.55 3.051 ;
      RECT 51.54 2.465 51.545 3.063 ;
      RECT 51.53 2.495 51.54 3.082 ;
      RECT 51.52 2.52 51.53 3.107 ;
      RECT 51.515 2.54 51.52 3.126 ;
      RECT 51.51 2.557 51.515 3.139 ;
      RECT 51.5 2.583 51.51 3.158 ;
      RECT 51.49 2.621 51.5 3.185 ;
      RECT 51.485 2.647 51.49 3.205 ;
      RECT 51.48 2.657 51.485 3.215 ;
      RECT 51.475 2.67 51.48 3.23 ;
      RECT 51.47 2.685 51.475 3.24 ;
      RECT 51.465 2.707 51.47 3.255 ;
      RECT 51.46 2.725 51.465 3.266 ;
      RECT 51.455 2.735 51.46 3.277 ;
      RECT 51.45 2.743 51.455 3.289 ;
      RECT 51.445 2.751 51.45 3.3 ;
      RECT 51.44 2.777 51.445 3.313 ;
      RECT 51.43 2.805 51.44 3.326 ;
      RECT 51.425 2.835 51.43 3.335 ;
      RECT 51.42 2.85 51.425 3.342 ;
      RECT 51.405 2.875 51.42 3.349 ;
      RECT 51.4 2.897 51.405 3.355 ;
      RECT 51.395 2.922 51.4 3.358 ;
      RECT 51.386 2.95 51.395 3.362 ;
      RECT 51.38 2.967 51.386 3.367 ;
      RECT 51.375 2.985 51.38 3.371 ;
      RECT 51.37 2.997 51.375 3.374 ;
      RECT 51.365 3.018 51.37 3.378 ;
      RECT 51.36 3.036 51.365 3.381 ;
      RECT 51.355 3.05 51.36 3.384 ;
      RECT 51.35 3.067 51.355 3.387 ;
      RECT 51.345 3.08 51.35 3.39 ;
      RECT 51.32 3.117 51.345 3.398 ;
      RECT 51.315 3.162 51.32 3.407 ;
      RECT 51.31 3.19 51.315 3.41 ;
      RECT 51.3 3.21 51.31 3.414 ;
      RECT 51.295 3.23 51.3 3.419 ;
      RECT 51.29 3.245 51.295 3.422 ;
      RECT 51.27 3.255 51.29 3.429 ;
      RECT 51.205 3.262 51.27 3.455 ;
      RECT 51.17 3.265 51.205 3.483 ;
      RECT 51.155 3.268 51.17 3.498 ;
      RECT 51.145 3.269 51.155 3.513 ;
      RECT 51.135 3.27 51.145 3.53 ;
      RECT 51.13 3.27 51.135 3.545 ;
      RECT 51.125 3.27 51.13 3.553 ;
      RECT 51.11 3.271 51.125 3.568 ;
      RECT 51.08 3.273 51.11 3.575 ;
      RECT 50.97 3.28 51.05 3.575 ;
      RECT 50.925 3.285 50.97 3.575 ;
      RECT 50.915 3.286 50.925 3.565 ;
      RECT 50.905 3.287 50.915 3.558 ;
      RECT 50.885 3.289 50.905 3.553 ;
      RECT 50.875 3.26 50.885 3.548 ;
      RECT 50.83 3.26 50.875 3.54 ;
      RECT 50.8 3.26 50.825 3.53 ;
      RECT 50.78 3.26 50.8 3.523 ;
      RECT 51.06 2.06 51.32 2.32 ;
      RECT 50.94 2.075 50.95 2.24 ;
      RECT 50.925 2.075 50.93 2.235 ;
      RECT 48.29 1.915 48.475 2.205 ;
      RECT 50.105 2.04 50.12 2.195 ;
      RECT 48.255 1.915 48.28 2.175 ;
      RECT 50.67 1.965 50.675 2.107 ;
      RECT 50.585 1.96 50.61 2.1 ;
      RECT 50.985 2.077 51.06 2.27 ;
      RECT 50.97 2.075 50.985 2.253 ;
      RECT 50.95 2.075 50.97 2.245 ;
      RECT 50.93 2.075 50.94 2.238 ;
      RECT 50.885 2.07 50.925 2.228 ;
      RECT 50.845 2.045 50.885 2.213 ;
      RECT 50.83 2.02 50.845 2.203 ;
      RECT 50.825 2.014 50.83 2.201 ;
      RECT 50.79 2.006 50.825 2.184 ;
      RECT 50.785 1.999 50.79 2.172 ;
      RECT 50.765 1.994 50.785 2.16 ;
      RECT 50.755 1.988 50.765 2.145 ;
      RECT 50.735 1.983 50.755 2.13 ;
      RECT 50.725 1.978 50.735 2.123 ;
      RECT 50.72 1.976 50.725 2.118 ;
      RECT 50.715 1.975 50.72 2.115 ;
      RECT 50.675 1.97 50.715 2.111 ;
      RECT 50.655 1.964 50.67 2.106 ;
      RECT 50.62 1.961 50.655 2.103 ;
      RECT 50.61 1.96 50.62 2.101 ;
      RECT 50.55 1.96 50.585 2.098 ;
      RECT 50.505 1.96 50.55 2.098 ;
      RECT 50.455 1.96 50.505 2.101 ;
      RECT 50.44 1.962 50.455 2.103 ;
      RECT 50.425 1.965 50.44 2.104 ;
      RECT 50.415 1.97 50.425 2.105 ;
      RECT 50.385 1.975 50.415 2.11 ;
      RECT 50.375 1.981 50.385 2.118 ;
      RECT 50.365 1.983 50.375 2.122 ;
      RECT 50.355 1.987 50.365 2.126 ;
      RECT 50.33 1.993 50.355 2.134 ;
      RECT 50.32 1.998 50.33 2.142 ;
      RECT 50.305 2.002 50.32 2.146 ;
      RECT 50.27 2.008 50.305 2.154 ;
      RECT 50.25 2.013 50.27 2.164 ;
      RECT 50.22 2.02 50.25 2.173 ;
      RECT 50.175 2.029 50.22 2.187 ;
      RECT 50.17 2.034 50.175 2.198 ;
      RECT 50.15 2.037 50.17 2.199 ;
      RECT 50.12 2.04 50.15 2.197 ;
      RECT 50.085 2.04 50.105 2.193 ;
      RECT 50.015 2.04 50.085 2.184 ;
      RECT 50 2.037 50.015 2.176 ;
      RECT 49.96 2.03 50 2.171 ;
      RECT 49.935 2.02 49.96 2.164 ;
      RECT 49.93 2.014 49.935 2.161 ;
      RECT 49.89 2.008 49.93 2.158 ;
      RECT 49.875 2.001 49.89 2.153 ;
      RECT 49.855 1.997 49.875 2.148 ;
      RECT 49.84 1.992 49.855 2.144 ;
      RECT 49.825 1.987 49.84 2.142 ;
      RECT 49.81 1.983 49.825 2.141 ;
      RECT 49.795 1.981 49.81 2.137 ;
      RECT 49.785 1.979 49.795 2.132 ;
      RECT 49.77 1.976 49.785 2.128 ;
      RECT 49.76 1.974 49.77 2.123 ;
      RECT 49.74 1.971 49.76 2.119 ;
      RECT 49.695 1.97 49.74 2.117 ;
      RECT 49.635 1.972 49.695 2.118 ;
      RECT 49.615 1.974 49.635 2.12 ;
      RECT 49.585 1.977 49.615 2.121 ;
      RECT 49.535 1.982 49.585 2.123 ;
      RECT 49.53 1.985 49.535 2.125 ;
      RECT 49.52 1.987 49.53 2.128 ;
      RECT 49.515 1.989 49.52 2.131 ;
      RECT 49.465 1.992 49.515 2.138 ;
      RECT 49.445 1.996 49.465 2.15 ;
      RECT 49.435 1.999 49.445 2.156 ;
      RECT 49.425 2 49.435 2.159 ;
      RECT 49.386 2.003 49.425 2.161 ;
      RECT 49.3 2.01 49.386 2.164 ;
      RECT 49.226 2.02 49.3 2.168 ;
      RECT 49.14 2.031 49.226 2.173 ;
      RECT 49.125 2.038 49.14 2.175 ;
      RECT 49.07 2.042 49.125 2.176 ;
      RECT 49.056 2.045 49.07 2.178 ;
      RECT 48.97 2.045 49.056 2.18 ;
      RECT 48.93 2.042 48.97 2.183 ;
      RECT 48.906 2.038 48.93 2.185 ;
      RECT 48.82 2.028 48.906 2.188 ;
      RECT 48.79 2.017 48.82 2.189 ;
      RECT 48.771 2.013 48.79 2.188 ;
      RECT 48.685 2.006 48.771 2.185 ;
      RECT 48.625 1.995 48.685 2.182 ;
      RECT 48.605 1.987 48.625 2.18 ;
      RECT 48.57 1.982 48.605 2.179 ;
      RECT 48.545 1.977 48.57 2.178 ;
      RECT 48.515 1.972 48.545 2.177 ;
      RECT 48.49 1.915 48.515 2.176 ;
      RECT 48.475 1.915 48.49 2.2 ;
      RECT 48.28 1.915 48.29 2.2 ;
      RECT 50.055 2.935 50.06 3.075 ;
      RECT 49.715 2.935 49.75 3.073 ;
      RECT 49.29 2.92 49.305 3.065 ;
      RECT 51.12 2.7 51.21 2.96 ;
      RECT 50.95 2.565 51.05 2.96 ;
      RECT 47.985 2.54 48.065 2.75 ;
      RECT 51.075 2.677 51.12 2.96 ;
      RECT 51.065 2.647 51.075 2.96 ;
      RECT 51.05 2.57 51.065 2.96 ;
      RECT 50.865 2.565 50.95 2.925 ;
      RECT 50.86 2.567 50.865 2.92 ;
      RECT 50.855 2.572 50.86 2.92 ;
      RECT 50.82 2.672 50.855 2.92 ;
      RECT 50.81 2.7 50.82 2.92 ;
      RECT 50.8 2.715 50.81 2.92 ;
      RECT 50.79 2.727 50.8 2.92 ;
      RECT 50.785 2.737 50.79 2.92 ;
      RECT 50.77 2.747 50.785 2.922 ;
      RECT 50.765 2.762 50.77 2.924 ;
      RECT 50.75 2.775 50.765 2.926 ;
      RECT 50.745 2.79 50.75 2.929 ;
      RECT 50.725 2.8 50.745 2.933 ;
      RECT 50.71 2.81 50.725 2.936 ;
      RECT 50.675 2.817 50.71 2.941 ;
      RECT 50.631 2.824 50.675 2.949 ;
      RECT 50.545 2.836 50.631 2.962 ;
      RECT 50.52 2.847 50.545 2.973 ;
      RECT 50.49 2.852 50.52 2.978 ;
      RECT 50.455 2.857 50.49 2.986 ;
      RECT 50.425 2.862 50.455 2.993 ;
      RECT 50.4 2.867 50.425 2.998 ;
      RECT 50.335 2.874 50.4 3.007 ;
      RECT 50.265 2.887 50.335 3.023 ;
      RECT 50.235 2.897 50.265 3.035 ;
      RECT 50.21 2.902 50.235 3.042 ;
      RECT 50.155 2.909 50.21 3.05 ;
      RECT 50.15 2.916 50.155 3.055 ;
      RECT 50.145 2.918 50.15 3.056 ;
      RECT 50.13 2.92 50.145 3.058 ;
      RECT 50.125 2.92 50.13 3.061 ;
      RECT 50.06 2.927 50.125 3.068 ;
      RECT 50.025 2.937 50.055 3.078 ;
      RECT 50.008 2.94 50.025 3.08 ;
      RECT 49.922 2.939 50.008 3.079 ;
      RECT 49.836 2.937 49.922 3.076 ;
      RECT 49.75 2.936 49.836 3.074 ;
      RECT 49.649 2.934 49.715 3.073 ;
      RECT 49.563 2.931 49.649 3.071 ;
      RECT 49.477 2.927 49.563 3.069 ;
      RECT 49.391 2.924 49.477 3.068 ;
      RECT 49.305 2.921 49.391 3.066 ;
      RECT 49.205 2.92 49.29 3.063 ;
      RECT 49.155 2.918 49.205 3.061 ;
      RECT 49.135 2.915 49.155 3.059 ;
      RECT 49.115 2.913 49.135 3.056 ;
      RECT 49.09 2.909 49.115 3.053 ;
      RECT 49.045 2.903 49.09 3.048 ;
      RECT 49.005 2.897 49.045 3.04 ;
      RECT 48.98 2.892 49.005 3.033 ;
      RECT 48.925 2.885 48.98 3.025 ;
      RECT 48.901 2.878 48.925 3.018 ;
      RECT 48.815 2.869 48.901 3.008 ;
      RECT 48.785 2.861 48.815 2.998 ;
      RECT 48.755 2.857 48.785 2.993 ;
      RECT 48.75 2.854 48.755 2.99 ;
      RECT 48.745 2.853 48.75 2.99 ;
      RECT 48.67 2.846 48.745 2.983 ;
      RECT 48.631 2.837 48.67 2.972 ;
      RECT 48.545 2.827 48.631 2.96 ;
      RECT 48.505 2.817 48.545 2.948 ;
      RECT 48.466 2.812 48.505 2.941 ;
      RECT 48.38 2.802 48.466 2.93 ;
      RECT 48.34 2.79 48.38 2.919 ;
      RECT 48.305 2.775 48.34 2.912 ;
      RECT 48.295 2.765 48.305 2.909 ;
      RECT 48.275 2.75 48.295 2.907 ;
      RECT 48.245 2.72 48.275 2.903 ;
      RECT 48.235 2.7 48.245 2.898 ;
      RECT 48.23 2.692 48.235 2.895 ;
      RECT 48.225 2.685 48.23 2.893 ;
      RECT 48.21 2.672 48.225 2.886 ;
      RECT 48.205 2.662 48.21 2.878 ;
      RECT 48.2 2.655 48.205 2.873 ;
      RECT 48.195 2.65 48.2 2.869 ;
      RECT 48.18 2.637 48.195 2.861 ;
      RECT 48.175 2.547 48.18 2.85 ;
      RECT 48.17 2.542 48.175 2.843 ;
      RECT 48.095 2.54 48.17 2.803 ;
      RECT 48.065 2.54 48.095 2.758 ;
      RECT 47.97 2.545 47.985 2.745 ;
      RECT 50.455 2.25 50.715 2.51 ;
      RECT 50.44 2.238 50.62 2.475 ;
      RECT 50.435 2.239 50.62 2.473 ;
      RECT 50.42 2.243 50.63 2.463 ;
      RECT 50.415 2.248 50.635 2.433 ;
      RECT 50.42 2.245 50.635 2.463 ;
      RECT 50.435 2.24 50.63 2.473 ;
      RECT 50.455 2.237 50.62 2.51 ;
      RECT 50.455 2.236 50.61 2.51 ;
      RECT 50.48 2.235 50.61 2.51 ;
      RECT 50.04 2.48 50.3 2.74 ;
      RECT 49.915 2.525 50.3 2.735 ;
      RECT 49.905 2.53 50.3 2.73 ;
      RECT 49.92 3.47 49.935 3.78 ;
      RECT 48.515 3.24 48.525 3.37 ;
      RECT 48.295 3.235 48.4 3.37 ;
      RECT 48.21 3.24 48.26 3.37 ;
      RECT 46.76 1.975 46.765 3.08 ;
      RECT 50.015 3.562 50.02 3.698 ;
      RECT 50.01 3.557 50.015 3.758 ;
      RECT 50.005 3.555 50.01 3.771 ;
      RECT 49.99 3.552 50.005 3.773 ;
      RECT 49.985 3.547 49.99 3.775 ;
      RECT 49.98 3.543 49.985 3.778 ;
      RECT 49.965 3.538 49.98 3.78 ;
      RECT 49.935 3.53 49.965 3.78 ;
      RECT 49.896 3.47 49.92 3.78 ;
      RECT 49.81 3.47 49.896 3.777 ;
      RECT 49.78 3.47 49.81 3.77 ;
      RECT 49.755 3.47 49.78 3.763 ;
      RECT 49.73 3.47 49.755 3.755 ;
      RECT 49.715 3.47 49.73 3.748 ;
      RECT 49.69 3.47 49.715 3.74 ;
      RECT 49.675 3.47 49.69 3.733 ;
      RECT 49.635 3.48 49.675 3.722 ;
      RECT 49.625 3.475 49.635 3.712 ;
      RECT 49.621 3.474 49.625 3.709 ;
      RECT 49.535 3.466 49.621 3.692 ;
      RECT 49.502 3.455 49.535 3.669 ;
      RECT 49.416 3.444 49.502 3.647 ;
      RECT 49.33 3.428 49.416 3.616 ;
      RECT 49.26 3.413 49.33 3.588 ;
      RECT 49.25 3.406 49.26 3.575 ;
      RECT 49.22 3.403 49.25 3.565 ;
      RECT 49.195 3.399 49.22 3.558 ;
      RECT 49.18 3.396 49.195 3.553 ;
      RECT 49.175 3.395 49.18 3.548 ;
      RECT 49.145 3.39 49.175 3.541 ;
      RECT 49.14 3.385 49.145 3.536 ;
      RECT 49.125 3.382 49.14 3.531 ;
      RECT 49.12 3.377 49.125 3.526 ;
      RECT 49.1 3.372 49.12 3.523 ;
      RECT 49.085 3.367 49.1 3.515 ;
      RECT 49.07 3.361 49.085 3.51 ;
      RECT 49.04 3.352 49.07 3.503 ;
      RECT 49.035 3.345 49.04 3.495 ;
      RECT 49.03 3.343 49.035 3.493 ;
      RECT 49.025 3.342 49.03 3.49 ;
      RECT 48.985 3.335 49.025 3.483 ;
      RECT 48.971 3.325 48.985 3.473 ;
      RECT 48.92 3.314 48.971 3.461 ;
      RECT 48.895 3.3 48.92 3.447 ;
      RECT 48.87 3.289 48.895 3.439 ;
      RECT 48.85 3.278 48.87 3.433 ;
      RECT 48.84 3.272 48.85 3.428 ;
      RECT 48.835 3.27 48.84 3.424 ;
      RECT 48.815 3.265 48.835 3.419 ;
      RECT 48.785 3.255 48.815 3.409 ;
      RECT 48.78 3.247 48.785 3.402 ;
      RECT 48.765 3.245 48.78 3.398 ;
      RECT 48.745 3.245 48.765 3.393 ;
      RECT 48.74 3.244 48.745 3.391 ;
      RECT 48.735 3.244 48.74 3.388 ;
      RECT 48.695 3.243 48.735 3.383 ;
      RECT 48.67 3.242 48.695 3.378 ;
      RECT 48.61 3.241 48.67 3.375 ;
      RECT 48.525 3.24 48.61 3.373 ;
      RECT 48.486 3.239 48.515 3.37 ;
      RECT 48.4 3.237 48.486 3.37 ;
      RECT 48.26 3.237 48.295 3.37 ;
      RECT 48.17 3.241 48.21 3.373 ;
      RECT 48.155 3.244 48.17 3.38 ;
      RECT 48.145 3.245 48.155 3.387 ;
      RECT 48.12 3.248 48.145 3.392 ;
      RECT 48.115 3.25 48.12 3.395 ;
      RECT 48.065 3.252 48.115 3.396 ;
      RECT 48.026 3.256 48.065 3.398 ;
      RECT 47.94 3.258 48.026 3.401 ;
      RECT 47.922 3.26 47.94 3.403 ;
      RECT 47.836 3.263 47.922 3.405 ;
      RECT 47.75 3.267 47.836 3.408 ;
      RECT 47.713 3.271 47.75 3.411 ;
      RECT 47.627 3.274 47.713 3.414 ;
      RECT 47.541 3.278 47.627 3.417 ;
      RECT 47.455 3.283 47.541 3.421 ;
      RECT 47.435 3.285 47.455 3.424 ;
      RECT 47.415 3.284 47.435 3.425 ;
      RECT 47.366 3.281 47.415 3.426 ;
      RECT 47.28 3.276 47.366 3.429 ;
      RECT 47.23 3.271 47.28 3.431 ;
      RECT 47.206 3.269 47.23 3.432 ;
      RECT 47.12 3.264 47.206 3.434 ;
      RECT 47.095 3.26 47.12 3.433 ;
      RECT 47.085 3.257 47.095 3.431 ;
      RECT 47.075 3.25 47.085 3.428 ;
      RECT 47.07 3.23 47.075 3.423 ;
      RECT 47.06 3.2 47.07 3.418 ;
      RECT 47.045 3.07 47.06 3.409 ;
      RECT 47.04 3.062 47.045 3.402 ;
      RECT 47.02 3.055 47.04 3.394 ;
      RECT 47.015 3.037 47.02 3.386 ;
      RECT 47.005 3.017 47.015 3.381 ;
      RECT 47 2.99 47.005 3.377 ;
      RECT 46.995 2.967 47 3.374 ;
      RECT 46.975 2.925 46.995 3.366 ;
      RECT 46.94 2.84 46.975 3.35 ;
      RECT 46.935 2.772 46.94 3.338 ;
      RECT 46.92 2.742 46.935 3.332 ;
      RECT 46.915 1.987 46.92 2.233 ;
      RECT 46.905 2.712 46.92 3.323 ;
      RECT 46.91 1.982 46.915 2.265 ;
      RECT 46.905 1.977 46.91 2.308 ;
      RECT 46.9 1.975 46.905 2.343 ;
      RECT 46.885 2.675 46.905 3.313 ;
      RECT 46.895 1.975 46.9 2.38 ;
      RECT 46.88 1.975 46.895 2.478 ;
      RECT 46.88 2.648 46.885 3.306 ;
      RECT 46.875 1.975 46.88 2.553 ;
      RECT 46.875 2.636 46.88 3.303 ;
      RECT 46.87 1.975 46.875 2.585 ;
      RECT 46.87 2.615 46.875 3.3 ;
      RECT 46.865 1.975 46.87 3.297 ;
      RECT 46.83 1.975 46.865 3.283 ;
      RECT 46.815 1.975 46.83 3.265 ;
      RECT 46.795 1.975 46.815 3.255 ;
      RECT 46.77 1.975 46.795 3.238 ;
      RECT 46.765 1.975 46.77 3.188 ;
      RECT 46.755 1.975 46.76 3.018 ;
      RECT 46.75 1.975 46.755 2.925 ;
      RECT 46.745 1.975 46.75 2.838 ;
      RECT 46.74 1.975 46.745 2.77 ;
      RECT 46.735 1.975 46.74 2.713 ;
      RECT 46.725 1.975 46.735 2.608 ;
      RECT 46.72 1.975 46.725 2.48 ;
      RECT 46.715 1.975 46.72 2.398 ;
      RECT 46.71 1.977 46.715 2.315 ;
      RECT 46.705 1.982 46.71 2.248 ;
      RECT 46.7 1.987 46.705 2.175 ;
      RECT 49.515 2.305 49.775 2.565 ;
      RECT 49.535 2.272 49.745 2.565 ;
      RECT 49.535 2.27 49.735 2.565 ;
      RECT 49.545 2.257 49.735 2.565 ;
      RECT 49.545 2.255 49.66 2.565 ;
      RECT 49.02 2.38 49.195 2.66 ;
      RECT 49.015 2.38 49.195 2.658 ;
      RECT 49.015 2.38 49.21 2.655 ;
      RECT 49.005 2.38 49.21 2.653 ;
      RECT 48.95 2.38 49.21 2.64 ;
      RECT 48.95 2.455 49.215 2.618 ;
      RECT 48.495 2.392 48.515 2.635 ;
      RECT 48.495 2.392 48.555 2.634 ;
      RECT 48.49 2.394 48.555 2.633 ;
      RECT 48.49 2.394 48.641 2.632 ;
      RECT 48.49 2.394 48.71 2.631 ;
      RECT 48.49 2.394 48.73 2.623 ;
      RECT 48.47 2.397 48.73 2.621 ;
      RECT 48.455 2.407 48.73 2.606 ;
      RECT 48.455 2.407 48.745 2.605 ;
      RECT 48.45 2.416 48.745 2.597 ;
      RECT 48.45 2.416 48.75 2.593 ;
      RECT 48.555 2.33 48.815 2.59 ;
      RECT 48.445 2.418 48.815 2.475 ;
      RECT 48.515 2.385 48.815 2.59 ;
      RECT 48.48 3.578 48.485 3.785 ;
      RECT 48.43 3.572 48.48 3.784 ;
      RECT 48.397 3.586 48.49 3.783 ;
      RECT 48.311 3.586 48.49 3.782 ;
      RECT 48.225 3.586 48.49 3.781 ;
      RECT 48.225 3.685 48.495 3.778 ;
      RECT 48.22 3.685 48.495 3.773 ;
      RECT 48.215 3.685 48.495 3.755 ;
      RECT 48.21 3.685 48.495 3.738 ;
      RECT 48.17 3.47 48.43 3.73 ;
      RECT 47.63 2.62 47.716 3.034 ;
      RECT 47.63 2.62 47.755 3.031 ;
      RECT 47.63 2.62 47.775 3.021 ;
      RECT 47.585 2.62 47.775 3.018 ;
      RECT 47.585 2.772 47.785 3.008 ;
      RECT 47.585 2.793 47.79 3.002 ;
      RECT 47.585 2.811 47.795 2.998 ;
      RECT 47.585 2.831 47.805 2.993 ;
      RECT 47.56 2.831 47.805 2.99 ;
      RECT 47.55 2.831 47.805 2.968 ;
      RECT 47.55 2.847 47.81 2.938 ;
      RECT 47.515 2.62 47.775 2.925 ;
      RECT 47.515 2.859 47.815 2.88 ;
      RECT 45.18 7.765 45.47 7.995 ;
      RECT 45.24 6.285 45.41 7.995 ;
      RECT 45.185 6.655 45.535 7.005 ;
      RECT 45.18 6.285 45.47 6.515 ;
      RECT 45.18 2.365 45.47 2.595 ;
      RECT 45.24 0.885 45.41 2.595 ;
      RECT 45.18 0.885 45.47 1.115 ;
      RECT 44.77 2.735 45.1 2.965 ;
      RECT 44.77 2.765 45.27 2.935 ;
      RECT 44.77 2.395 44.96 2.965 ;
      RECT 44.19 2.365 44.48 2.595 ;
      RECT 44.19 2.395 44.96 2.565 ;
      RECT 44.25 0.885 44.42 2.595 ;
      RECT 44.19 0.885 44.48 1.115 ;
      RECT 44.19 7.765 44.48 7.995 ;
      RECT 44.25 6.285 44.42 7.995 ;
      RECT 44.19 6.285 44.48 6.515 ;
      RECT 44.19 6.325 45.04 6.485 ;
      RECT 44.87 5.915 45.04 6.485 ;
      RECT 44.19 6.32 44.58 6.485 ;
      RECT 44.81 5.915 45.1 6.145 ;
      RECT 44.81 5.945 45.27 6.115 ;
      RECT 43.82 2.735 44.11 2.965 ;
      RECT 43.82 2.765 44.28 2.935 ;
      RECT 43.88 1.655 44.045 2.965 ;
      RECT 42.395 1.625 42.685 1.855 ;
      RECT 42.395 1.655 44.045 1.825 ;
      RECT 42.455 0.885 42.625 1.855 ;
      RECT 42.395 0.885 42.685 1.115 ;
      RECT 42.395 7.765 42.685 7.995 ;
      RECT 42.455 7.025 42.625 7.995 ;
      RECT 42.455 7.12 44.045 7.29 ;
      RECT 43.875 5.915 44.045 7.29 ;
      RECT 42.395 7.025 42.685 7.255 ;
      RECT 43.82 5.915 44.11 6.145 ;
      RECT 43.82 5.945 44.28 6.115 ;
      RECT 40.445 2.705 40.785 3.055 ;
      RECT 40.535 2.025 40.705 3.055 ;
      RECT 42.825 1.965 43.175 2.315 ;
      RECT 40.535 2.025 43.175 2.195 ;
      RECT 42.85 6.655 43.175 6.98 ;
      RECT 37.39 6.615 37.74 6.965 ;
      RECT 42.825 6.655 43.175 6.885 ;
      RECT 37.19 6.655 37.74 6.885 ;
      RECT 37.02 6.685 43.175 6.855 ;
      RECT 42.05 2.365 42.37 2.685 ;
      RECT 42.02 2.365 42.37 2.595 ;
      RECT 41.85 2.395 42.37 2.565 ;
      RECT 42.05 6.255 42.37 6.545 ;
      RECT 42.02 6.285 42.37 6.515 ;
      RECT 41.85 6.315 42.37 6.485 ;
      RECT 41.005 2.705 41.345 3.055 ;
      RECT 41.005 2.765 41.485 2.935 ;
      RECT 41 5.86 41.34 6.21 ;
      RECT 35.39 5.915 35.68 6.145 ;
      RECT 35.39 5.945 41.485 6.115 ;
      RECT 37.74 2.985 37.89 3.26 ;
      RECT 38.28 2.065 38.285 2.285 ;
      RECT 39.43 2.265 39.445 2.463 ;
      RECT 39.395 2.257 39.43 2.47 ;
      RECT 39.365 2.25 39.395 2.47 ;
      RECT 39.31 2.215 39.365 2.47 ;
      RECT 39.245 2.152 39.31 2.47 ;
      RECT 39.24 2.117 39.245 2.468 ;
      RECT 39.235 2.112 39.24 2.46 ;
      RECT 39.23 2.107 39.235 2.446 ;
      RECT 39.225 2.104 39.23 2.439 ;
      RECT 39.18 2.094 39.225 2.39 ;
      RECT 39.16 2.081 39.18 2.325 ;
      RECT 39.155 2.076 39.16 2.298 ;
      RECT 39.15 2.075 39.155 2.291 ;
      RECT 39.145 2.074 39.15 2.284 ;
      RECT 39.06 2.059 39.145 2.23 ;
      RECT 39.03 2.04 39.06 2.18 ;
      RECT 38.95 2.023 39.03 2.165 ;
      RECT 38.915 2.01 38.95 2.15 ;
      RECT 38.907 2.01 38.915 2.145 ;
      RECT 38.821 2.011 38.907 2.145 ;
      RECT 38.735 2.013 38.821 2.145 ;
      RECT 38.71 2.014 38.735 2.149 ;
      RECT 38.635 2.02 38.71 2.164 ;
      RECT 38.552 2.032 38.635 2.188 ;
      RECT 38.466 2.045 38.552 2.214 ;
      RECT 38.38 2.058 38.466 2.24 ;
      RECT 38.345 2.067 38.38 2.259 ;
      RECT 38.295 2.067 38.345 2.272 ;
      RECT 38.285 2.065 38.295 2.283 ;
      RECT 38.27 2.062 38.28 2.285 ;
      RECT 38.255 2.054 38.27 2.293 ;
      RECT 38.24 2.046 38.255 2.313 ;
      RECT 38.235 2.041 38.24 2.37 ;
      RECT 38.22 2.036 38.235 2.443 ;
      RECT 38.215 2.031 38.22 2.485 ;
      RECT 38.21 2.029 38.215 2.513 ;
      RECT 38.205 2.027 38.21 2.535 ;
      RECT 38.195 2.023 38.205 2.578 ;
      RECT 38.19 2.02 38.195 2.603 ;
      RECT 38.185 2.018 38.19 2.623 ;
      RECT 38.18 2.016 38.185 2.647 ;
      RECT 38.175 2.012 38.18 2.67 ;
      RECT 38.17 2.008 38.175 2.693 ;
      RECT 38.135 1.998 38.17 2.8 ;
      RECT 38.13 1.988 38.135 2.898 ;
      RECT 38.125 1.986 38.13 2.925 ;
      RECT 38.12 1.985 38.125 2.945 ;
      RECT 38.115 1.977 38.12 2.965 ;
      RECT 38.11 1.972 38.115 3 ;
      RECT 38.105 1.97 38.11 3.018 ;
      RECT 38.1 1.97 38.105 3.043 ;
      RECT 38.095 1.97 38.1 3.065 ;
      RECT 38.06 1.97 38.095 3.108 ;
      RECT 38.035 1.97 38.06 3.137 ;
      RECT 38.025 1.97 38.035 2.323 ;
      RECT 38.028 2.38 38.035 3.147 ;
      RECT 38.025 2.437 38.028 3.15 ;
      RECT 38.02 1.97 38.025 2.295 ;
      RECT 38.02 2.487 38.025 3.153 ;
      RECT 38.01 1.97 38.02 2.285 ;
      RECT 38.015 2.54 38.02 3.156 ;
      RECT 38.01 2.625 38.015 3.16 ;
      RECT 38 1.97 38.01 2.273 ;
      RECT 38.005 2.672 38.01 3.164 ;
      RECT 38 2.747 38.005 3.168 ;
      RECT 37.965 1.97 38 2.248 ;
      RECT 37.99 2.83 38 3.173 ;
      RECT 37.98 2.897 37.99 3.18 ;
      RECT 37.975 2.925 37.98 3.185 ;
      RECT 37.965 2.938 37.975 3.191 ;
      RECT 37.92 1.97 37.965 2.205 ;
      RECT 37.96 2.943 37.965 3.198 ;
      RECT 37.92 2.96 37.96 3.26 ;
      RECT 37.915 1.972 37.92 2.178 ;
      RECT 37.89 2.98 37.92 3.26 ;
      RECT 37.91 1.977 37.915 2.15 ;
      RECT 37.7 2.989 37.74 3.26 ;
      RECT 37.675 2.997 37.7 3.23 ;
      RECT 37.63 3.005 37.675 3.23 ;
      RECT 37.615 3.01 37.63 3.225 ;
      RECT 37.605 3.01 37.615 3.219 ;
      RECT 37.595 3.017 37.605 3.216 ;
      RECT 37.59 3.055 37.595 3.205 ;
      RECT 37.585 3.117 37.59 3.183 ;
      RECT 38.855 2.992 39.04 3.215 ;
      RECT 38.855 3.007 39.045 3.211 ;
      RECT 38.845 2.28 38.93 3.21 ;
      RECT 38.845 3.007 39.05 3.204 ;
      RECT 38.84 3.015 39.05 3.203 ;
      RECT 39.045 2.735 39.365 3.055 ;
      RECT 38.84 2.907 39.01 2.998 ;
      RECT 38.835 2.907 39.01 2.98 ;
      RECT 38.825 2.715 38.96 2.955 ;
      RECT 38.82 2.715 38.96 2.9 ;
      RECT 38.78 2.295 38.95 2.8 ;
      RECT 38.765 2.295 38.95 2.67 ;
      RECT 38.76 2.295 38.95 2.623 ;
      RECT 38.755 2.295 38.95 2.603 ;
      RECT 38.75 2.295 38.95 2.578 ;
      RECT 38.72 2.295 38.98 2.555 ;
      RECT 38.73 2.292 38.94 2.555 ;
      RECT 38.855 2.287 38.94 3.215 ;
      RECT 38.74 2.28 38.93 2.555 ;
      RECT 38.735 2.285 38.93 2.555 ;
      RECT 37.565 2.497 37.75 2.71 ;
      RECT 37.565 2.505 37.76 2.703 ;
      RECT 37.545 2.505 37.76 2.7 ;
      RECT 37.54 2.505 37.76 2.685 ;
      RECT 37.47 2.42 37.73 2.68 ;
      RECT 37.47 2.565 37.765 2.593 ;
      RECT 37.125 3.02 37.385 3.28 ;
      RECT 37.15 2.965 37.345 3.28 ;
      RECT 37.145 2.714 37.325 3.008 ;
      RECT 37.145 2.72 37.335 3.008 ;
      RECT 37.125 2.722 37.335 2.953 ;
      RECT 37.12 2.732 37.335 2.82 ;
      RECT 37.15 2.712 37.325 3.28 ;
      RECT 37.236 2.71 37.325 3.28 ;
      RECT 37.095 1.93 37.13 2.3 ;
      RECT 36.885 2.04 36.89 2.3 ;
      RECT 37.13 1.937 37.145 2.3 ;
      RECT 37.02 1.93 37.095 2.378 ;
      RECT 37.01 1.93 37.02 2.463 ;
      RECT 36.985 1.93 37.01 2.498 ;
      RECT 36.945 1.93 36.985 2.566 ;
      RECT 36.935 1.937 36.945 2.618 ;
      RECT 36.905 2.04 36.935 2.659 ;
      RECT 36.9 2.04 36.905 2.698 ;
      RECT 36.89 2.04 36.9 2.718 ;
      RECT 36.885 2.335 36.89 2.755 ;
      RECT 36.88 2.352 36.885 2.775 ;
      RECT 36.865 2.415 36.88 2.815 ;
      RECT 36.86 2.458 36.865 2.85 ;
      RECT 36.855 2.466 36.86 2.863 ;
      RECT 36.845 2.48 36.855 2.885 ;
      RECT 36.82 2.515 36.845 2.95 ;
      RECT 36.81 2.55 36.82 3.013 ;
      RECT 36.79 2.58 36.81 3.074 ;
      RECT 36.775 2.616 36.79 3.141 ;
      RECT 36.765 2.644 36.775 3.18 ;
      RECT 36.755 2.666 36.765 3.2 ;
      RECT 36.75 2.676 36.755 3.211 ;
      RECT 36.745 2.685 36.75 3.214 ;
      RECT 36.735 2.703 36.745 3.218 ;
      RECT 36.725 2.721 36.735 3.219 ;
      RECT 36.7 2.76 36.725 3.216 ;
      RECT 36.68 2.802 36.7 3.213 ;
      RECT 36.665 2.84 36.68 3.212 ;
      RECT 36.63 2.875 36.665 3.209 ;
      RECT 36.625 2.897 36.63 3.207 ;
      RECT 36.56 2.937 36.625 3.204 ;
      RECT 36.555 2.977 36.56 3.2 ;
      RECT 36.54 2.987 36.555 3.191 ;
      RECT 36.53 3.107 36.54 3.176 ;
      RECT 37.01 3.52 37.02 3.78 ;
      RECT 37.01 3.523 37.03 3.779 ;
      RECT 37 3.513 37.01 3.778 ;
      RECT 36.99 3.528 37.07 3.774 ;
      RECT 36.975 3.507 36.99 3.772 ;
      RECT 36.95 3.532 37.075 3.768 ;
      RECT 36.935 3.492 36.95 3.763 ;
      RECT 36.935 3.534 37.085 3.762 ;
      RECT 36.935 3.542 37.1 3.755 ;
      RECT 36.875 3.479 36.935 3.745 ;
      RECT 36.865 3.466 36.875 3.727 ;
      RECT 36.84 3.456 36.865 3.717 ;
      RECT 36.835 3.446 36.84 3.709 ;
      RECT 36.77 3.542 37.1 3.691 ;
      RECT 36.685 3.542 37.1 3.653 ;
      RECT 36.575 3.37 36.835 3.63 ;
      RECT 36.95 3.5 36.975 3.768 ;
      RECT 36.99 3.51 37 3.774 ;
      RECT 36.575 3.518 37.015 3.63 ;
      RECT 36.76 7.765 37.05 7.995 ;
      RECT 36.82 7.025 36.99 7.995 ;
      RECT 36.72 7.055 37.09 7.425 ;
      RECT 36.76 7.025 37.05 7.425 ;
      RECT 35.79 3.275 35.82 3.575 ;
      RECT 35.565 3.26 35.57 3.535 ;
      RECT 35.365 3.26 35.52 3.52 ;
      RECT 36.665 1.975 36.695 2.235 ;
      RECT 36.655 1.975 36.665 2.343 ;
      RECT 36.635 1.975 36.655 2.353 ;
      RECT 36.62 1.975 36.635 2.365 ;
      RECT 36.565 1.975 36.62 2.415 ;
      RECT 36.55 1.975 36.565 2.463 ;
      RECT 36.52 1.975 36.55 2.498 ;
      RECT 36.465 1.975 36.52 2.56 ;
      RECT 36.445 1.975 36.465 2.628 ;
      RECT 36.44 1.975 36.445 2.658 ;
      RECT 36.435 1.975 36.44 2.67 ;
      RECT 36.43 2.092 36.435 2.688 ;
      RECT 36.41 2.11 36.43 2.713 ;
      RECT 36.39 2.137 36.41 2.763 ;
      RECT 36.385 2.157 36.39 2.794 ;
      RECT 36.38 2.165 36.385 2.811 ;
      RECT 36.365 2.191 36.38 2.84 ;
      RECT 36.35 2.233 36.365 2.875 ;
      RECT 36.345 2.262 36.35 2.898 ;
      RECT 36.34 2.277 36.345 2.911 ;
      RECT 36.335 2.3 36.34 2.922 ;
      RECT 36.325 2.32 36.335 2.94 ;
      RECT 36.315 2.35 36.325 2.963 ;
      RECT 36.31 2.372 36.315 2.983 ;
      RECT 36.305 2.387 36.31 2.998 ;
      RECT 36.29 2.417 36.305 3.025 ;
      RECT 36.285 2.447 36.29 3.051 ;
      RECT 36.28 2.465 36.285 3.063 ;
      RECT 36.27 2.495 36.28 3.082 ;
      RECT 36.26 2.52 36.27 3.107 ;
      RECT 36.255 2.54 36.26 3.126 ;
      RECT 36.25 2.557 36.255 3.139 ;
      RECT 36.24 2.583 36.25 3.158 ;
      RECT 36.23 2.621 36.24 3.185 ;
      RECT 36.225 2.647 36.23 3.205 ;
      RECT 36.22 2.657 36.225 3.215 ;
      RECT 36.215 2.67 36.22 3.23 ;
      RECT 36.21 2.685 36.215 3.24 ;
      RECT 36.205 2.707 36.21 3.255 ;
      RECT 36.2 2.725 36.205 3.266 ;
      RECT 36.195 2.735 36.2 3.277 ;
      RECT 36.19 2.743 36.195 3.289 ;
      RECT 36.185 2.751 36.19 3.3 ;
      RECT 36.18 2.777 36.185 3.313 ;
      RECT 36.17 2.805 36.18 3.326 ;
      RECT 36.165 2.835 36.17 3.335 ;
      RECT 36.16 2.85 36.165 3.342 ;
      RECT 36.145 2.875 36.16 3.349 ;
      RECT 36.14 2.897 36.145 3.355 ;
      RECT 36.135 2.922 36.14 3.358 ;
      RECT 36.126 2.95 36.135 3.362 ;
      RECT 36.12 2.967 36.126 3.367 ;
      RECT 36.115 2.985 36.12 3.371 ;
      RECT 36.11 2.997 36.115 3.374 ;
      RECT 36.105 3.018 36.11 3.378 ;
      RECT 36.1 3.036 36.105 3.381 ;
      RECT 36.095 3.05 36.1 3.384 ;
      RECT 36.09 3.067 36.095 3.387 ;
      RECT 36.085 3.08 36.09 3.39 ;
      RECT 36.06 3.117 36.085 3.398 ;
      RECT 36.055 3.162 36.06 3.407 ;
      RECT 36.05 3.19 36.055 3.41 ;
      RECT 36.04 3.21 36.05 3.414 ;
      RECT 36.035 3.23 36.04 3.419 ;
      RECT 36.03 3.245 36.035 3.422 ;
      RECT 36.01 3.255 36.03 3.429 ;
      RECT 35.945 3.262 36.01 3.455 ;
      RECT 35.91 3.265 35.945 3.483 ;
      RECT 35.895 3.268 35.91 3.498 ;
      RECT 35.885 3.269 35.895 3.513 ;
      RECT 35.875 3.27 35.885 3.53 ;
      RECT 35.87 3.27 35.875 3.545 ;
      RECT 35.865 3.27 35.87 3.553 ;
      RECT 35.85 3.271 35.865 3.568 ;
      RECT 35.82 3.273 35.85 3.575 ;
      RECT 35.71 3.28 35.79 3.575 ;
      RECT 35.665 3.285 35.71 3.575 ;
      RECT 35.655 3.286 35.665 3.565 ;
      RECT 35.645 3.287 35.655 3.558 ;
      RECT 35.625 3.289 35.645 3.553 ;
      RECT 35.615 3.26 35.625 3.548 ;
      RECT 35.57 3.26 35.615 3.54 ;
      RECT 35.54 3.26 35.565 3.53 ;
      RECT 35.52 3.26 35.54 3.523 ;
      RECT 35.8 2.06 36.06 2.32 ;
      RECT 35.68 2.075 35.69 2.24 ;
      RECT 35.665 2.075 35.67 2.235 ;
      RECT 33.03 1.915 33.215 2.205 ;
      RECT 34.845 2.04 34.86 2.195 ;
      RECT 32.995 1.915 33.02 2.175 ;
      RECT 35.41 1.965 35.415 2.107 ;
      RECT 35.325 1.96 35.35 2.1 ;
      RECT 35.725 2.077 35.8 2.27 ;
      RECT 35.71 2.075 35.725 2.253 ;
      RECT 35.69 2.075 35.71 2.245 ;
      RECT 35.67 2.075 35.68 2.238 ;
      RECT 35.625 2.07 35.665 2.228 ;
      RECT 35.585 2.045 35.625 2.213 ;
      RECT 35.57 2.02 35.585 2.203 ;
      RECT 35.565 2.014 35.57 2.201 ;
      RECT 35.53 2.006 35.565 2.184 ;
      RECT 35.525 1.999 35.53 2.172 ;
      RECT 35.505 1.994 35.525 2.16 ;
      RECT 35.495 1.988 35.505 2.145 ;
      RECT 35.475 1.983 35.495 2.13 ;
      RECT 35.465 1.978 35.475 2.123 ;
      RECT 35.46 1.976 35.465 2.118 ;
      RECT 35.455 1.975 35.46 2.115 ;
      RECT 35.415 1.97 35.455 2.111 ;
      RECT 35.395 1.964 35.41 2.106 ;
      RECT 35.36 1.961 35.395 2.103 ;
      RECT 35.35 1.96 35.36 2.101 ;
      RECT 35.29 1.96 35.325 2.098 ;
      RECT 35.245 1.96 35.29 2.098 ;
      RECT 35.195 1.96 35.245 2.101 ;
      RECT 35.18 1.962 35.195 2.103 ;
      RECT 35.165 1.965 35.18 2.104 ;
      RECT 35.155 1.97 35.165 2.105 ;
      RECT 35.125 1.975 35.155 2.11 ;
      RECT 35.115 1.981 35.125 2.118 ;
      RECT 35.105 1.983 35.115 2.122 ;
      RECT 35.095 1.987 35.105 2.126 ;
      RECT 35.07 1.993 35.095 2.134 ;
      RECT 35.06 1.998 35.07 2.142 ;
      RECT 35.045 2.002 35.06 2.146 ;
      RECT 35.01 2.008 35.045 2.154 ;
      RECT 34.99 2.013 35.01 2.164 ;
      RECT 34.96 2.02 34.99 2.173 ;
      RECT 34.915 2.029 34.96 2.187 ;
      RECT 34.91 2.034 34.915 2.198 ;
      RECT 34.89 2.037 34.91 2.199 ;
      RECT 34.86 2.04 34.89 2.197 ;
      RECT 34.825 2.04 34.845 2.193 ;
      RECT 34.755 2.04 34.825 2.184 ;
      RECT 34.74 2.037 34.755 2.176 ;
      RECT 34.7 2.03 34.74 2.171 ;
      RECT 34.675 2.02 34.7 2.164 ;
      RECT 34.67 2.014 34.675 2.161 ;
      RECT 34.63 2.008 34.67 2.158 ;
      RECT 34.615 2.001 34.63 2.153 ;
      RECT 34.595 1.997 34.615 2.148 ;
      RECT 34.58 1.992 34.595 2.144 ;
      RECT 34.565 1.987 34.58 2.142 ;
      RECT 34.55 1.983 34.565 2.141 ;
      RECT 34.535 1.981 34.55 2.137 ;
      RECT 34.525 1.979 34.535 2.132 ;
      RECT 34.51 1.976 34.525 2.128 ;
      RECT 34.5 1.974 34.51 2.123 ;
      RECT 34.48 1.971 34.5 2.119 ;
      RECT 34.435 1.97 34.48 2.117 ;
      RECT 34.375 1.972 34.435 2.118 ;
      RECT 34.355 1.974 34.375 2.12 ;
      RECT 34.325 1.977 34.355 2.121 ;
      RECT 34.275 1.982 34.325 2.123 ;
      RECT 34.27 1.985 34.275 2.125 ;
      RECT 34.26 1.987 34.27 2.128 ;
      RECT 34.255 1.989 34.26 2.131 ;
      RECT 34.205 1.992 34.255 2.138 ;
      RECT 34.185 1.996 34.205 2.15 ;
      RECT 34.175 1.999 34.185 2.156 ;
      RECT 34.165 2 34.175 2.159 ;
      RECT 34.126 2.003 34.165 2.161 ;
      RECT 34.04 2.01 34.126 2.164 ;
      RECT 33.966 2.02 34.04 2.168 ;
      RECT 33.88 2.031 33.966 2.173 ;
      RECT 33.865 2.038 33.88 2.175 ;
      RECT 33.81 2.042 33.865 2.176 ;
      RECT 33.796 2.045 33.81 2.178 ;
      RECT 33.71 2.045 33.796 2.18 ;
      RECT 33.67 2.042 33.71 2.183 ;
      RECT 33.646 2.038 33.67 2.185 ;
      RECT 33.56 2.028 33.646 2.188 ;
      RECT 33.53 2.017 33.56 2.189 ;
      RECT 33.511 2.013 33.53 2.188 ;
      RECT 33.425 2.006 33.511 2.185 ;
      RECT 33.365 1.995 33.425 2.182 ;
      RECT 33.345 1.987 33.365 2.18 ;
      RECT 33.31 1.982 33.345 2.179 ;
      RECT 33.285 1.977 33.31 2.178 ;
      RECT 33.255 1.972 33.285 2.177 ;
      RECT 33.23 1.915 33.255 2.176 ;
      RECT 33.215 1.915 33.23 2.2 ;
      RECT 33.02 1.915 33.03 2.2 ;
      RECT 34.795 2.935 34.8 3.075 ;
      RECT 34.455 2.935 34.49 3.073 ;
      RECT 34.03 2.92 34.045 3.065 ;
      RECT 35.86 2.7 35.95 2.96 ;
      RECT 35.69 2.565 35.79 2.96 ;
      RECT 32.725 2.54 32.805 2.75 ;
      RECT 35.815 2.677 35.86 2.96 ;
      RECT 35.805 2.647 35.815 2.96 ;
      RECT 35.79 2.57 35.805 2.96 ;
      RECT 35.605 2.565 35.69 2.925 ;
      RECT 35.6 2.567 35.605 2.92 ;
      RECT 35.595 2.572 35.6 2.92 ;
      RECT 35.56 2.672 35.595 2.92 ;
      RECT 35.55 2.7 35.56 2.92 ;
      RECT 35.54 2.715 35.55 2.92 ;
      RECT 35.53 2.727 35.54 2.92 ;
      RECT 35.525 2.737 35.53 2.92 ;
      RECT 35.51 2.747 35.525 2.922 ;
      RECT 35.505 2.762 35.51 2.924 ;
      RECT 35.49 2.775 35.505 2.926 ;
      RECT 35.485 2.79 35.49 2.929 ;
      RECT 35.465 2.8 35.485 2.933 ;
      RECT 35.45 2.81 35.465 2.936 ;
      RECT 35.415 2.817 35.45 2.941 ;
      RECT 35.371 2.824 35.415 2.949 ;
      RECT 35.285 2.836 35.371 2.962 ;
      RECT 35.26 2.847 35.285 2.973 ;
      RECT 35.23 2.852 35.26 2.978 ;
      RECT 35.195 2.857 35.23 2.986 ;
      RECT 35.165 2.862 35.195 2.993 ;
      RECT 35.14 2.867 35.165 2.998 ;
      RECT 35.075 2.874 35.14 3.007 ;
      RECT 35.005 2.887 35.075 3.023 ;
      RECT 34.975 2.897 35.005 3.035 ;
      RECT 34.95 2.902 34.975 3.042 ;
      RECT 34.895 2.909 34.95 3.05 ;
      RECT 34.89 2.916 34.895 3.055 ;
      RECT 34.885 2.918 34.89 3.056 ;
      RECT 34.87 2.92 34.885 3.058 ;
      RECT 34.865 2.92 34.87 3.061 ;
      RECT 34.8 2.927 34.865 3.068 ;
      RECT 34.765 2.937 34.795 3.078 ;
      RECT 34.748 2.94 34.765 3.08 ;
      RECT 34.662 2.939 34.748 3.079 ;
      RECT 34.576 2.937 34.662 3.076 ;
      RECT 34.49 2.936 34.576 3.074 ;
      RECT 34.389 2.934 34.455 3.073 ;
      RECT 34.303 2.931 34.389 3.071 ;
      RECT 34.217 2.927 34.303 3.069 ;
      RECT 34.131 2.924 34.217 3.068 ;
      RECT 34.045 2.921 34.131 3.066 ;
      RECT 33.945 2.92 34.03 3.063 ;
      RECT 33.895 2.918 33.945 3.061 ;
      RECT 33.875 2.915 33.895 3.059 ;
      RECT 33.855 2.913 33.875 3.056 ;
      RECT 33.83 2.909 33.855 3.053 ;
      RECT 33.785 2.903 33.83 3.048 ;
      RECT 33.745 2.897 33.785 3.04 ;
      RECT 33.72 2.892 33.745 3.033 ;
      RECT 33.665 2.885 33.72 3.025 ;
      RECT 33.641 2.878 33.665 3.018 ;
      RECT 33.555 2.869 33.641 3.008 ;
      RECT 33.525 2.861 33.555 2.998 ;
      RECT 33.495 2.857 33.525 2.993 ;
      RECT 33.49 2.854 33.495 2.99 ;
      RECT 33.485 2.853 33.49 2.99 ;
      RECT 33.41 2.846 33.485 2.983 ;
      RECT 33.371 2.837 33.41 2.972 ;
      RECT 33.285 2.827 33.371 2.96 ;
      RECT 33.245 2.817 33.285 2.948 ;
      RECT 33.206 2.812 33.245 2.941 ;
      RECT 33.12 2.802 33.206 2.93 ;
      RECT 33.08 2.79 33.12 2.919 ;
      RECT 33.045 2.775 33.08 2.912 ;
      RECT 33.035 2.765 33.045 2.909 ;
      RECT 33.015 2.75 33.035 2.907 ;
      RECT 32.985 2.72 33.015 2.903 ;
      RECT 32.975 2.7 32.985 2.898 ;
      RECT 32.97 2.692 32.975 2.895 ;
      RECT 32.965 2.685 32.97 2.893 ;
      RECT 32.95 2.672 32.965 2.886 ;
      RECT 32.945 2.662 32.95 2.878 ;
      RECT 32.94 2.655 32.945 2.873 ;
      RECT 32.935 2.65 32.94 2.869 ;
      RECT 32.92 2.637 32.935 2.861 ;
      RECT 32.915 2.547 32.92 2.85 ;
      RECT 32.91 2.542 32.915 2.843 ;
      RECT 32.835 2.54 32.91 2.803 ;
      RECT 32.805 2.54 32.835 2.758 ;
      RECT 32.71 2.545 32.725 2.745 ;
      RECT 35.195 2.25 35.455 2.51 ;
      RECT 35.18 2.238 35.36 2.475 ;
      RECT 35.175 2.239 35.36 2.473 ;
      RECT 35.16 2.243 35.37 2.463 ;
      RECT 35.155 2.248 35.375 2.433 ;
      RECT 35.16 2.245 35.375 2.463 ;
      RECT 35.175 2.24 35.37 2.473 ;
      RECT 35.195 2.237 35.36 2.51 ;
      RECT 35.195 2.236 35.35 2.51 ;
      RECT 35.22 2.235 35.35 2.51 ;
      RECT 34.78 2.48 35.04 2.74 ;
      RECT 34.655 2.525 35.04 2.735 ;
      RECT 34.645 2.53 35.04 2.73 ;
      RECT 34.66 3.47 34.675 3.78 ;
      RECT 33.255 3.24 33.265 3.37 ;
      RECT 33.035 3.235 33.14 3.37 ;
      RECT 32.95 3.24 33 3.37 ;
      RECT 31.5 1.975 31.505 3.08 ;
      RECT 34.755 3.562 34.76 3.698 ;
      RECT 34.75 3.557 34.755 3.758 ;
      RECT 34.745 3.555 34.75 3.771 ;
      RECT 34.73 3.552 34.745 3.773 ;
      RECT 34.725 3.547 34.73 3.775 ;
      RECT 34.72 3.543 34.725 3.778 ;
      RECT 34.705 3.538 34.72 3.78 ;
      RECT 34.675 3.53 34.705 3.78 ;
      RECT 34.636 3.47 34.66 3.78 ;
      RECT 34.55 3.47 34.636 3.777 ;
      RECT 34.52 3.47 34.55 3.77 ;
      RECT 34.495 3.47 34.52 3.763 ;
      RECT 34.47 3.47 34.495 3.755 ;
      RECT 34.455 3.47 34.47 3.748 ;
      RECT 34.43 3.47 34.455 3.74 ;
      RECT 34.415 3.47 34.43 3.733 ;
      RECT 34.375 3.48 34.415 3.722 ;
      RECT 34.365 3.475 34.375 3.712 ;
      RECT 34.361 3.474 34.365 3.709 ;
      RECT 34.275 3.466 34.361 3.692 ;
      RECT 34.242 3.455 34.275 3.669 ;
      RECT 34.156 3.444 34.242 3.647 ;
      RECT 34.07 3.428 34.156 3.616 ;
      RECT 34 3.413 34.07 3.588 ;
      RECT 33.99 3.406 34 3.575 ;
      RECT 33.96 3.403 33.99 3.565 ;
      RECT 33.935 3.399 33.96 3.558 ;
      RECT 33.92 3.396 33.935 3.553 ;
      RECT 33.915 3.395 33.92 3.548 ;
      RECT 33.885 3.39 33.915 3.541 ;
      RECT 33.88 3.385 33.885 3.536 ;
      RECT 33.865 3.382 33.88 3.531 ;
      RECT 33.86 3.377 33.865 3.526 ;
      RECT 33.84 3.372 33.86 3.523 ;
      RECT 33.825 3.367 33.84 3.515 ;
      RECT 33.81 3.361 33.825 3.51 ;
      RECT 33.78 3.352 33.81 3.503 ;
      RECT 33.775 3.345 33.78 3.495 ;
      RECT 33.77 3.343 33.775 3.493 ;
      RECT 33.765 3.342 33.77 3.49 ;
      RECT 33.725 3.335 33.765 3.483 ;
      RECT 33.711 3.325 33.725 3.473 ;
      RECT 33.66 3.314 33.711 3.461 ;
      RECT 33.635 3.3 33.66 3.447 ;
      RECT 33.61 3.289 33.635 3.439 ;
      RECT 33.59 3.278 33.61 3.433 ;
      RECT 33.58 3.272 33.59 3.428 ;
      RECT 33.575 3.27 33.58 3.424 ;
      RECT 33.555 3.265 33.575 3.419 ;
      RECT 33.525 3.255 33.555 3.409 ;
      RECT 33.52 3.247 33.525 3.402 ;
      RECT 33.505 3.245 33.52 3.398 ;
      RECT 33.485 3.245 33.505 3.393 ;
      RECT 33.48 3.244 33.485 3.391 ;
      RECT 33.475 3.244 33.48 3.388 ;
      RECT 33.435 3.243 33.475 3.383 ;
      RECT 33.41 3.242 33.435 3.378 ;
      RECT 33.35 3.241 33.41 3.375 ;
      RECT 33.265 3.24 33.35 3.373 ;
      RECT 33.226 3.239 33.255 3.37 ;
      RECT 33.14 3.237 33.226 3.37 ;
      RECT 33 3.237 33.035 3.37 ;
      RECT 32.91 3.241 32.95 3.373 ;
      RECT 32.895 3.244 32.91 3.38 ;
      RECT 32.885 3.245 32.895 3.387 ;
      RECT 32.86 3.248 32.885 3.392 ;
      RECT 32.855 3.25 32.86 3.395 ;
      RECT 32.805 3.252 32.855 3.396 ;
      RECT 32.766 3.256 32.805 3.398 ;
      RECT 32.68 3.258 32.766 3.401 ;
      RECT 32.662 3.26 32.68 3.403 ;
      RECT 32.576 3.263 32.662 3.405 ;
      RECT 32.49 3.267 32.576 3.408 ;
      RECT 32.453 3.271 32.49 3.411 ;
      RECT 32.367 3.274 32.453 3.414 ;
      RECT 32.281 3.278 32.367 3.417 ;
      RECT 32.195 3.283 32.281 3.421 ;
      RECT 32.175 3.285 32.195 3.424 ;
      RECT 32.155 3.284 32.175 3.425 ;
      RECT 32.106 3.281 32.155 3.426 ;
      RECT 32.02 3.276 32.106 3.429 ;
      RECT 31.97 3.271 32.02 3.431 ;
      RECT 31.946 3.269 31.97 3.432 ;
      RECT 31.86 3.264 31.946 3.434 ;
      RECT 31.835 3.26 31.86 3.433 ;
      RECT 31.825 3.257 31.835 3.431 ;
      RECT 31.815 3.25 31.825 3.428 ;
      RECT 31.81 3.23 31.815 3.423 ;
      RECT 31.8 3.2 31.81 3.418 ;
      RECT 31.785 3.07 31.8 3.409 ;
      RECT 31.78 3.062 31.785 3.402 ;
      RECT 31.76 3.055 31.78 3.394 ;
      RECT 31.755 3.037 31.76 3.386 ;
      RECT 31.745 3.017 31.755 3.381 ;
      RECT 31.74 2.99 31.745 3.377 ;
      RECT 31.735 2.967 31.74 3.374 ;
      RECT 31.715 2.925 31.735 3.366 ;
      RECT 31.68 2.84 31.715 3.35 ;
      RECT 31.675 2.772 31.68 3.338 ;
      RECT 31.66 2.742 31.675 3.332 ;
      RECT 31.655 1.987 31.66 2.233 ;
      RECT 31.645 2.712 31.66 3.323 ;
      RECT 31.65 1.982 31.655 2.265 ;
      RECT 31.645 1.977 31.65 2.308 ;
      RECT 31.64 1.975 31.645 2.343 ;
      RECT 31.625 2.675 31.645 3.313 ;
      RECT 31.635 1.975 31.64 2.38 ;
      RECT 31.62 1.975 31.635 2.478 ;
      RECT 31.62 2.648 31.625 3.306 ;
      RECT 31.615 1.975 31.62 2.553 ;
      RECT 31.615 2.636 31.62 3.303 ;
      RECT 31.61 1.975 31.615 2.585 ;
      RECT 31.61 2.615 31.615 3.3 ;
      RECT 31.605 1.975 31.61 3.297 ;
      RECT 31.57 1.975 31.605 3.283 ;
      RECT 31.555 1.975 31.57 3.265 ;
      RECT 31.535 1.975 31.555 3.255 ;
      RECT 31.51 1.975 31.535 3.238 ;
      RECT 31.505 1.975 31.51 3.188 ;
      RECT 31.495 1.975 31.5 3.018 ;
      RECT 31.49 1.975 31.495 2.925 ;
      RECT 31.485 1.975 31.49 2.838 ;
      RECT 31.48 1.975 31.485 2.77 ;
      RECT 31.475 1.975 31.48 2.713 ;
      RECT 31.465 1.975 31.475 2.608 ;
      RECT 31.46 1.975 31.465 2.48 ;
      RECT 31.455 1.975 31.46 2.398 ;
      RECT 31.45 1.977 31.455 2.315 ;
      RECT 31.445 1.982 31.45 2.248 ;
      RECT 31.44 1.987 31.445 2.175 ;
      RECT 34.255 2.305 34.515 2.565 ;
      RECT 34.275 2.272 34.485 2.565 ;
      RECT 34.275 2.27 34.475 2.565 ;
      RECT 34.285 2.257 34.475 2.565 ;
      RECT 34.285 2.255 34.4 2.565 ;
      RECT 33.76 2.38 33.935 2.66 ;
      RECT 33.755 2.38 33.935 2.658 ;
      RECT 33.755 2.38 33.95 2.655 ;
      RECT 33.745 2.38 33.95 2.653 ;
      RECT 33.69 2.38 33.95 2.64 ;
      RECT 33.69 2.455 33.955 2.618 ;
      RECT 33.235 2.392 33.255 2.635 ;
      RECT 33.235 2.392 33.295 2.634 ;
      RECT 33.23 2.394 33.295 2.633 ;
      RECT 33.23 2.394 33.381 2.632 ;
      RECT 33.23 2.394 33.45 2.631 ;
      RECT 33.23 2.394 33.47 2.623 ;
      RECT 33.21 2.397 33.47 2.621 ;
      RECT 33.195 2.407 33.47 2.606 ;
      RECT 33.195 2.407 33.485 2.605 ;
      RECT 33.19 2.416 33.485 2.597 ;
      RECT 33.19 2.416 33.49 2.593 ;
      RECT 33.295 2.33 33.555 2.59 ;
      RECT 33.185 2.418 33.555 2.475 ;
      RECT 33.255 2.385 33.555 2.59 ;
      RECT 33.22 3.578 33.225 3.785 ;
      RECT 33.17 3.572 33.22 3.784 ;
      RECT 33.137 3.586 33.23 3.783 ;
      RECT 33.051 3.586 33.23 3.782 ;
      RECT 32.965 3.586 33.23 3.781 ;
      RECT 32.965 3.685 33.235 3.778 ;
      RECT 32.96 3.685 33.235 3.773 ;
      RECT 32.955 3.685 33.235 3.755 ;
      RECT 32.95 3.685 33.235 3.738 ;
      RECT 32.91 3.47 33.17 3.73 ;
      RECT 32.37 2.62 32.456 3.034 ;
      RECT 32.37 2.62 32.495 3.031 ;
      RECT 32.37 2.62 32.515 3.021 ;
      RECT 32.325 2.62 32.515 3.018 ;
      RECT 32.325 2.772 32.525 3.008 ;
      RECT 32.325 2.793 32.53 3.002 ;
      RECT 32.325 2.811 32.535 2.998 ;
      RECT 32.325 2.831 32.545 2.993 ;
      RECT 32.3 2.831 32.545 2.99 ;
      RECT 32.29 2.831 32.545 2.968 ;
      RECT 32.29 2.847 32.55 2.938 ;
      RECT 32.255 2.62 32.515 2.925 ;
      RECT 32.255 2.859 32.555 2.88 ;
      RECT 29.92 7.765 30.21 7.995 ;
      RECT 29.98 6.285 30.15 7.995 ;
      RECT 29.965 6.66 30.32 7.015 ;
      RECT 29.92 6.285 30.21 6.515 ;
      RECT 29.92 2.365 30.21 2.595 ;
      RECT 29.98 0.885 30.15 2.595 ;
      RECT 29.92 0.885 30.21 1.115 ;
      RECT 29.51 2.735 29.84 2.965 ;
      RECT 29.51 2.765 30.01 2.935 ;
      RECT 29.51 2.395 29.7 2.965 ;
      RECT 28.93 2.365 29.22 2.595 ;
      RECT 28.93 2.395 29.7 2.565 ;
      RECT 28.99 0.885 29.16 2.595 ;
      RECT 28.93 0.885 29.22 1.115 ;
      RECT 28.93 7.765 29.22 7.995 ;
      RECT 28.99 6.285 29.16 7.995 ;
      RECT 28.93 6.285 29.22 6.515 ;
      RECT 28.93 6.325 29.78 6.485 ;
      RECT 29.61 5.915 29.78 6.485 ;
      RECT 28.93 6.32 29.32 6.485 ;
      RECT 29.55 5.915 29.84 6.145 ;
      RECT 29.55 5.945 30.01 6.115 ;
      RECT 28.56 2.735 28.85 2.965 ;
      RECT 28.56 2.765 29.02 2.935 ;
      RECT 28.62 1.655 28.785 2.965 ;
      RECT 27.135 1.625 27.425 1.855 ;
      RECT 27.135 1.655 28.785 1.825 ;
      RECT 27.195 0.885 27.365 1.855 ;
      RECT 27.135 0.885 27.425 1.115 ;
      RECT 27.135 7.765 27.425 7.995 ;
      RECT 27.195 7.025 27.365 7.995 ;
      RECT 27.195 7.12 28.785 7.29 ;
      RECT 28.615 5.915 28.785 7.29 ;
      RECT 27.135 7.025 27.425 7.255 ;
      RECT 28.56 5.915 28.85 6.145 ;
      RECT 28.56 5.945 29.02 6.115 ;
      RECT 25.185 2.705 25.525 3.055 ;
      RECT 25.275 2.025 25.445 3.055 ;
      RECT 27.565 1.965 27.915 2.315 ;
      RECT 25.275 2.025 27.915 2.195 ;
      RECT 27.59 6.655 27.915 6.98 ;
      RECT 22.13 6.61 22.48 6.96 ;
      RECT 27.565 6.655 27.915 6.885 ;
      RECT 21.93 6.655 22.48 6.885 ;
      RECT 21.76 6.685 27.915 6.855 ;
      RECT 26.79 2.365 27.11 2.685 ;
      RECT 26.76 2.365 27.11 2.595 ;
      RECT 26.59 2.395 27.11 2.565 ;
      RECT 26.79 6.255 27.11 6.545 ;
      RECT 26.76 6.285 27.11 6.515 ;
      RECT 26.59 6.315 27.11 6.485 ;
      RECT 25.745 2.705 26.085 3.055 ;
      RECT 25.745 2.765 26.225 2.935 ;
      RECT 25.74 5.86 26.08 6.21 ;
      RECT 20.13 5.915 20.42 6.145 ;
      RECT 20.13 5.945 26.225 6.115 ;
      RECT 22.48 2.985 22.63 3.26 ;
      RECT 23.02 2.065 23.025 2.285 ;
      RECT 24.17 2.265 24.185 2.463 ;
      RECT 24.135 2.257 24.17 2.47 ;
      RECT 24.105 2.25 24.135 2.47 ;
      RECT 24.05 2.215 24.105 2.47 ;
      RECT 23.985 2.152 24.05 2.47 ;
      RECT 23.98 2.117 23.985 2.468 ;
      RECT 23.975 2.112 23.98 2.46 ;
      RECT 23.97 2.107 23.975 2.446 ;
      RECT 23.965 2.104 23.97 2.439 ;
      RECT 23.92 2.094 23.965 2.39 ;
      RECT 23.9 2.081 23.92 2.325 ;
      RECT 23.895 2.076 23.9 2.298 ;
      RECT 23.89 2.075 23.895 2.291 ;
      RECT 23.885 2.074 23.89 2.284 ;
      RECT 23.8 2.059 23.885 2.23 ;
      RECT 23.77 2.04 23.8 2.18 ;
      RECT 23.69 2.023 23.77 2.165 ;
      RECT 23.655 2.01 23.69 2.15 ;
      RECT 23.647 2.01 23.655 2.145 ;
      RECT 23.561 2.011 23.647 2.145 ;
      RECT 23.475 2.013 23.561 2.145 ;
      RECT 23.45 2.014 23.475 2.149 ;
      RECT 23.375 2.02 23.45 2.164 ;
      RECT 23.292 2.032 23.375 2.188 ;
      RECT 23.206 2.045 23.292 2.214 ;
      RECT 23.12 2.058 23.206 2.24 ;
      RECT 23.085 2.067 23.12 2.259 ;
      RECT 23.035 2.067 23.085 2.272 ;
      RECT 23.025 2.065 23.035 2.283 ;
      RECT 23.01 2.062 23.02 2.285 ;
      RECT 22.995 2.054 23.01 2.293 ;
      RECT 22.98 2.046 22.995 2.313 ;
      RECT 22.975 2.041 22.98 2.37 ;
      RECT 22.96 2.036 22.975 2.443 ;
      RECT 22.955 2.031 22.96 2.485 ;
      RECT 22.95 2.029 22.955 2.513 ;
      RECT 22.945 2.027 22.95 2.535 ;
      RECT 22.935 2.023 22.945 2.578 ;
      RECT 22.93 2.02 22.935 2.603 ;
      RECT 22.925 2.018 22.93 2.623 ;
      RECT 22.92 2.016 22.925 2.647 ;
      RECT 22.915 2.012 22.92 2.67 ;
      RECT 22.91 2.008 22.915 2.693 ;
      RECT 22.875 1.998 22.91 2.8 ;
      RECT 22.87 1.988 22.875 2.898 ;
      RECT 22.865 1.986 22.87 2.925 ;
      RECT 22.86 1.985 22.865 2.945 ;
      RECT 22.855 1.977 22.86 2.965 ;
      RECT 22.85 1.972 22.855 3 ;
      RECT 22.845 1.97 22.85 3.018 ;
      RECT 22.84 1.97 22.845 3.043 ;
      RECT 22.835 1.97 22.84 3.065 ;
      RECT 22.8 1.97 22.835 3.108 ;
      RECT 22.775 1.97 22.8 3.137 ;
      RECT 22.765 1.97 22.775 2.323 ;
      RECT 22.768 2.38 22.775 3.147 ;
      RECT 22.765 2.437 22.768 3.15 ;
      RECT 22.76 1.97 22.765 2.295 ;
      RECT 22.76 2.487 22.765 3.153 ;
      RECT 22.75 1.97 22.76 2.285 ;
      RECT 22.755 2.54 22.76 3.156 ;
      RECT 22.75 2.625 22.755 3.16 ;
      RECT 22.74 1.97 22.75 2.273 ;
      RECT 22.745 2.672 22.75 3.164 ;
      RECT 22.74 2.747 22.745 3.168 ;
      RECT 22.705 1.97 22.74 2.248 ;
      RECT 22.73 2.83 22.74 3.173 ;
      RECT 22.72 2.897 22.73 3.18 ;
      RECT 22.715 2.925 22.72 3.185 ;
      RECT 22.705 2.938 22.715 3.191 ;
      RECT 22.66 1.97 22.705 2.205 ;
      RECT 22.7 2.943 22.705 3.198 ;
      RECT 22.66 2.96 22.7 3.26 ;
      RECT 22.655 1.972 22.66 2.178 ;
      RECT 22.63 2.98 22.66 3.26 ;
      RECT 22.65 1.977 22.655 2.15 ;
      RECT 22.44 2.989 22.48 3.26 ;
      RECT 22.415 2.997 22.44 3.23 ;
      RECT 22.37 3.005 22.415 3.23 ;
      RECT 22.355 3.01 22.37 3.225 ;
      RECT 22.345 3.01 22.355 3.219 ;
      RECT 22.335 3.017 22.345 3.216 ;
      RECT 22.33 3.055 22.335 3.205 ;
      RECT 22.325 3.117 22.33 3.183 ;
      RECT 23.595 2.992 23.78 3.215 ;
      RECT 23.595 3.007 23.785 3.211 ;
      RECT 23.585 2.28 23.67 3.21 ;
      RECT 23.585 3.007 23.79 3.204 ;
      RECT 23.58 3.015 23.79 3.203 ;
      RECT 23.785 2.735 24.105 3.055 ;
      RECT 23.58 2.907 23.75 2.998 ;
      RECT 23.575 2.907 23.75 2.98 ;
      RECT 23.565 2.715 23.7 2.955 ;
      RECT 23.56 2.715 23.7 2.9 ;
      RECT 23.52 2.295 23.69 2.8 ;
      RECT 23.505 2.295 23.69 2.67 ;
      RECT 23.5 2.295 23.69 2.623 ;
      RECT 23.495 2.295 23.69 2.603 ;
      RECT 23.49 2.295 23.69 2.578 ;
      RECT 23.46 2.295 23.72 2.555 ;
      RECT 23.47 2.292 23.68 2.555 ;
      RECT 23.595 2.287 23.68 3.215 ;
      RECT 23.48 2.28 23.67 2.555 ;
      RECT 23.475 2.285 23.67 2.555 ;
      RECT 22.305 2.497 22.49 2.71 ;
      RECT 22.305 2.505 22.5 2.703 ;
      RECT 22.285 2.505 22.5 2.7 ;
      RECT 22.28 2.505 22.5 2.685 ;
      RECT 22.21 2.42 22.47 2.68 ;
      RECT 22.21 2.565 22.505 2.593 ;
      RECT 21.865 3.02 22.125 3.28 ;
      RECT 21.89 2.965 22.085 3.28 ;
      RECT 21.885 2.714 22.065 3.008 ;
      RECT 21.885 2.72 22.075 3.008 ;
      RECT 21.865 2.722 22.075 2.953 ;
      RECT 21.86 2.732 22.075 2.82 ;
      RECT 21.89 2.712 22.065 3.28 ;
      RECT 21.976 2.71 22.065 3.28 ;
      RECT 21.835 1.93 21.87 2.3 ;
      RECT 21.625 2.04 21.63 2.3 ;
      RECT 21.87 1.937 21.885 2.3 ;
      RECT 21.76 1.93 21.835 2.378 ;
      RECT 21.75 1.93 21.76 2.463 ;
      RECT 21.725 1.93 21.75 2.498 ;
      RECT 21.685 1.93 21.725 2.566 ;
      RECT 21.675 1.937 21.685 2.618 ;
      RECT 21.645 2.04 21.675 2.659 ;
      RECT 21.64 2.04 21.645 2.698 ;
      RECT 21.63 2.04 21.64 2.718 ;
      RECT 21.625 2.335 21.63 2.755 ;
      RECT 21.62 2.352 21.625 2.775 ;
      RECT 21.605 2.415 21.62 2.815 ;
      RECT 21.6 2.458 21.605 2.85 ;
      RECT 21.595 2.466 21.6 2.863 ;
      RECT 21.585 2.48 21.595 2.885 ;
      RECT 21.56 2.515 21.585 2.95 ;
      RECT 21.55 2.55 21.56 3.013 ;
      RECT 21.53 2.58 21.55 3.074 ;
      RECT 21.515 2.616 21.53 3.141 ;
      RECT 21.505 2.644 21.515 3.18 ;
      RECT 21.495 2.666 21.505 3.2 ;
      RECT 21.49 2.676 21.495 3.211 ;
      RECT 21.485 2.685 21.49 3.214 ;
      RECT 21.475 2.703 21.485 3.218 ;
      RECT 21.465 2.721 21.475 3.219 ;
      RECT 21.44 2.76 21.465 3.216 ;
      RECT 21.42 2.802 21.44 3.213 ;
      RECT 21.405 2.84 21.42 3.212 ;
      RECT 21.37 2.875 21.405 3.209 ;
      RECT 21.365 2.897 21.37 3.207 ;
      RECT 21.3 2.937 21.365 3.204 ;
      RECT 21.295 2.977 21.3 3.2 ;
      RECT 21.28 2.987 21.295 3.191 ;
      RECT 21.27 3.107 21.28 3.176 ;
      RECT 21.75 3.52 21.76 3.78 ;
      RECT 21.75 3.523 21.77 3.779 ;
      RECT 21.74 3.513 21.75 3.778 ;
      RECT 21.73 3.528 21.81 3.774 ;
      RECT 21.715 3.507 21.73 3.772 ;
      RECT 21.69 3.532 21.815 3.768 ;
      RECT 21.675 3.492 21.69 3.763 ;
      RECT 21.675 3.534 21.825 3.762 ;
      RECT 21.675 3.542 21.84 3.755 ;
      RECT 21.615 3.479 21.675 3.745 ;
      RECT 21.605 3.466 21.615 3.727 ;
      RECT 21.58 3.456 21.605 3.717 ;
      RECT 21.575 3.446 21.58 3.709 ;
      RECT 21.51 3.542 21.84 3.691 ;
      RECT 21.425 3.542 21.84 3.653 ;
      RECT 21.315 3.37 21.575 3.63 ;
      RECT 21.69 3.5 21.715 3.768 ;
      RECT 21.73 3.51 21.74 3.774 ;
      RECT 21.315 3.518 21.755 3.63 ;
      RECT 21.5 7.765 21.79 7.995 ;
      RECT 21.56 7.025 21.73 7.995 ;
      RECT 21.46 7.055 21.83 7.425 ;
      RECT 21.5 7.025 21.79 7.425 ;
      RECT 20.53 3.275 20.56 3.575 ;
      RECT 20.305 3.26 20.31 3.535 ;
      RECT 20.105 3.26 20.26 3.52 ;
      RECT 21.405 1.975 21.435 2.235 ;
      RECT 21.395 1.975 21.405 2.343 ;
      RECT 21.375 1.975 21.395 2.353 ;
      RECT 21.36 1.975 21.375 2.365 ;
      RECT 21.305 1.975 21.36 2.415 ;
      RECT 21.29 1.975 21.305 2.463 ;
      RECT 21.26 1.975 21.29 2.498 ;
      RECT 21.205 1.975 21.26 2.56 ;
      RECT 21.185 1.975 21.205 2.628 ;
      RECT 21.18 1.975 21.185 2.658 ;
      RECT 21.175 1.975 21.18 2.67 ;
      RECT 21.17 2.092 21.175 2.688 ;
      RECT 21.15 2.11 21.17 2.713 ;
      RECT 21.13 2.137 21.15 2.763 ;
      RECT 21.125 2.157 21.13 2.794 ;
      RECT 21.12 2.165 21.125 2.811 ;
      RECT 21.105 2.191 21.12 2.84 ;
      RECT 21.09 2.233 21.105 2.875 ;
      RECT 21.085 2.262 21.09 2.898 ;
      RECT 21.08 2.277 21.085 2.911 ;
      RECT 21.075 2.3 21.08 2.922 ;
      RECT 21.065 2.32 21.075 2.94 ;
      RECT 21.055 2.35 21.065 2.963 ;
      RECT 21.05 2.372 21.055 2.983 ;
      RECT 21.045 2.387 21.05 2.998 ;
      RECT 21.03 2.417 21.045 3.025 ;
      RECT 21.025 2.447 21.03 3.051 ;
      RECT 21.02 2.465 21.025 3.063 ;
      RECT 21.01 2.495 21.02 3.082 ;
      RECT 21 2.52 21.01 3.107 ;
      RECT 20.995 2.54 21 3.126 ;
      RECT 20.99 2.557 20.995 3.139 ;
      RECT 20.98 2.583 20.99 3.158 ;
      RECT 20.97 2.621 20.98 3.185 ;
      RECT 20.965 2.647 20.97 3.205 ;
      RECT 20.96 2.657 20.965 3.215 ;
      RECT 20.955 2.67 20.96 3.23 ;
      RECT 20.95 2.685 20.955 3.24 ;
      RECT 20.945 2.707 20.95 3.255 ;
      RECT 20.94 2.725 20.945 3.266 ;
      RECT 20.935 2.735 20.94 3.277 ;
      RECT 20.93 2.743 20.935 3.289 ;
      RECT 20.925 2.751 20.93 3.3 ;
      RECT 20.92 2.777 20.925 3.313 ;
      RECT 20.91 2.805 20.92 3.326 ;
      RECT 20.905 2.835 20.91 3.335 ;
      RECT 20.9 2.85 20.905 3.342 ;
      RECT 20.885 2.875 20.9 3.349 ;
      RECT 20.88 2.897 20.885 3.355 ;
      RECT 20.875 2.922 20.88 3.358 ;
      RECT 20.866 2.95 20.875 3.362 ;
      RECT 20.86 2.967 20.866 3.367 ;
      RECT 20.855 2.985 20.86 3.371 ;
      RECT 20.85 2.997 20.855 3.374 ;
      RECT 20.845 3.018 20.85 3.378 ;
      RECT 20.84 3.036 20.845 3.381 ;
      RECT 20.835 3.05 20.84 3.384 ;
      RECT 20.83 3.067 20.835 3.387 ;
      RECT 20.825 3.08 20.83 3.39 ;
      RECT 20.8 3.117 20.825 3.398 ;
      RECT 20.795 3.162 20.8 3.407 ;
      RECT 20.79 3.19 20.795 3.41 ;
      RECT 20.78 3.21 20.79 3.414 ;
      RECT 20.775 3.23 20.78 3.419 ;
      RECT 20.77 3.245 20.775 3.422 ;
      RECT 20.75 3.255 20.77 3.429 ;
      RECT 20.685 3.262 20.75 3.455 ;
      RECT 20.65 3.265 20.685 3.483 ;
      RECT 20.635 3.268 20.65 3.498 ;
      RECT 20.625 3.269 20.635 3.513 ;
      RECT 20.615 3.27 20.625 3.53 ;
      RECT 20.61 3.27 20.615 3.545 ;
      RECT 20.605 3.27 20.61 3.553 ;
      RECT 20.59 3.271 20.605 3.568 ;
      RECT 20.56 3.273 20.59 3.575 ;
      RECT 20.45 3.28 20.53 3.575 ;
      RECT 20.405 3.285 20.45 3.575 ;
      RECT 20.395 3.286 20.405 3.565 ;
      RECT 20.385 3.287 20.395 3.558 ;
      RECT 20.365 3.289 20.385 3.553 ;
      RECT 20.355 3.26 20.365 3.548 ;
      RECT 20.31 3.26 20.355 3.54 ;
      RECT 20.28 3.26 20.305 3.53 ;
      RECT 20.26 3.26 20.28 3.523 ;
      RECT 20.54 2.06 20.8 2.32 ;
      RECT 20.42 2.075 20.43 2.24 ;
      RECT 20.405 2.075 20.41 2.235 ;
      RECT 17.77 1.915 17.955 2.205 ;
      RECT 19.585 2.04 19.6 2.195 ;
      RECT 17.735 1.915 17.76 2.175 ;
      RECT 20.15 1.965 20.155 2.107 ;
      RECT 20.065 1.96 20.09 2.1 ;
      RECT 20.465 2.077 20.54 2.27 ;
      RECT 20.45 2.075 20.465 2.253 ;
      RECT 20.43 2.075 20.45 2.245 ;
      RECT 20.41 2.075 20.42 2.238 ;
      RECT 20.365 2.07 20.405 2.228 ;
      RECT 20.325 2.045 20.365 2.213 ;
      RECT 20.31 2.02 20.325 2.203 ;
      RECT 20.305 2.014 20.31 2.201 ;
      RECT 20.27 2.006 20.305 2.184 ;
      RECT 20.265 1.999 20.27 2.172 ;
      RECT 20.245 1.994 20.265 2.16 ;
      RECT 20.235 1.988 20.245 2.145 ;
      RECT 20.215 1.983 20.235 2.13 ;
      RECT 20.205 1.978 20.215 2.123 ;
      RECT 20.2 1.976 20.205 2.118 ;
      RECT 20.195 1.975 20.2 2.115 ;
      RECT 20.155 1.97 20.195 2.111 ;
      RECT 20.135 1.964 20.15 2.106 ;
      RECT 20.1 1.961 20.135 2.103 ;
      RECT 20.09 1.96 20.1 2.101 ;
      RECT 20.03 1.96 20.065 2.098 ;
      RECT 19.985 1.96 20.03 2.098 ;
      RECT 19.935 1.96 19.985 2.101 ;
      RECT 19.92 1.962 19.935 2.103 ;
      RECT 19.905 1.965 19.92 2.104 ;
      RECT 19.895 1.97 19.905 2.105 ;
      RECT 19.865 1.975 19.895 2.11 ;
      RECT 19.855 1.981 19.865 2.118 ;
      RECT 19.845 1.983 19.855 2.122 ;
      RECT 19.835 1.987 19.845 2.126 ;
      RECT 19.81 1.993 19.835 2.134 ;
      RECT 19.8 1.998 19.81 2.142 ;
      RECT 19.785 2.002 19.8 2.146 ;
      RECT 19.75 2.008 19.785 2.154 ;
      RECT 19.73 2.013 19.75 2.164 ;
      RECT 19.7 2.02 19.73 2.173 ;
      RECT 19.655 2.029 19.7 2.187 ;
      RECT 19.65 2.034 19.655 2.198 ;
      RECT 19.63 2.037 19.65 2.199 ;
      RECT 19.6 2.04 19.63 2.197 ;
      RECT 19.565 2.04 19.585 2.193 ;
      RECT 19.495 2.04 19.565 2.184 ;
      RECT 19.48 2.037 19.495 2.176 ;
      RECT 19.44 2.03 19.48 2.171 ;
      RECT 19.415 2.02 19.44 2.164 ;
      RECT 19.41 2.014 19.415 2.161 ;
      RECT 19.37 2.008 19.41 2.158 ;
      RECT 19.355 2.001 19.37 2.153 ;
      RECT 19.335 1.997 19.355 2.148 ;
      RECT 19.32 1.992 19.335 2.144 ;
      RECT 19.305 1.987 19.32 2.142 ;
      RECT 19.29 1.983 19.305 2.141 ;
      RECT 19.275 1.981 19.29 2.137 ;
      RECT 19.265 1.979 19.275 2.132 ;
      RECT 19.25 1.976 19.265 2.128 ;
      RECT 19.24 1.974 19.25 2.123 ;
      RECT 19.22 1.971 19.24 2.119 ;
      RECT 19.175 1.97 19.22 2.117 ;
      RECT 19.115 1.972 19.175 2.118 ;
      RECT 19.095 1.974 19.115 2.12 ;
      RECT 19.065 1.977 19.095 2.121 ;
      RECT 19.015 1.982 19.065 2.123 ;
      RECT 19.01 1.985 19.015 2.125 ;
      RECT 19 1.987 19.01 2.128 ;
      RECT 18.995 1.989 19 2.131 ;
      RECT 18.945 1.992 18.995 2.138 ;
      RECT 18.925 1.996 18.945 2.15 ;
      RECT 18.915 1.999 18.925 2.156 ;
      RECT 18.905 2 18.915 2.159 ;
      RECT 18.866 2.003 18.905 2.161 ;
      RECT 18.78 2.01 18.866 2.164 ;
      RECT 18.706 2.02 18.78 2.168 ;
      RECT 18.62 2.031 18.706 2.173 ;
      RECT 18.605 2.038 18.62 2.175 ;
      RECT 18.55 2.042 18.605 2.176 ;
      RECT 18.536 2.045 18.55 2.178 ;
      RECT 18.45 2.045 18.536 2.18 ;
      RECT 18.41 2.042 18.45 2.183 ;
      RECT 18.386 2.038 18.41 2.185 ;
      RECT 18.3 2.028 18.386 2.188 ;
      RECT 18.27 2.017 18.3 2.189 ;
      RECT 18.251 2.013 18.27 2.188 ;
      RECT 18.165 2.006 18.251 2.185 ;
      RECT 18.105 1.995 18.165 2.182 ;
      RECT 18.085 1.987 18.105 2.18 ;
      RECT 18.05 1.982 18.085 2.179 ;
      RECT 18.025 1.977 18.05 2.178 ;
      RECT 17.995 1.972 18.025 2.177 ;
      RECT 17.97 1.915 17.995 2.176 ;
      RECT 17.955 1.915 17.97 2.2 ;
      RECT 17.76 1.915 17.77 2.2 ;
      RECT 19.535 2.935 19.54 3.075 ;
      RECT 19.195 2.935 19.23 3.073 ;
      RECT 18.77 2.92 18.785 3.065 ;
      RECT 20.6 2.7 20.69 2.96 ;
      RECT 20.43 2.565 20.53 2.96 ;
      RECT 17.465 2.54 17.545 2.75 ;
      RECT 20.555 2.677 20.6 2.96 ;
      RECT 20.545 2.647 20.555 2.96 ;
      RECT 20.53 2.57 20.545 2.96 ;
      RECT 20.345 2.565 20.43 2.925 ;
      RECT 20.34 2.567 20.345 2.92 ;
      RECT 20.335 2.572 20.34 2.92 ;
      RECT 20.3 2.672 20.335 2.92 ;
      RECT 20.29 2.7 20.3 2.92 ;
      RECT 20.28 2.715 20.29 2.92 ;
      RECT 20.27 2.727 20.28 2.92 ;
      RECT 20.265 2.737 20.27 2.92 ;
      RECT 20.25 2.747 20.265 2.922 ;
      RECT 20.245 2.762 20.25 2.924 ;
      RECT 20.23 2.775 20.245 2.926 ;
      RECT 20.225 2.79 20.23 2.929 ;
      RECT 20.205 2.8 20.225 2.933 ;
      RECT 20.19 2.81 20.205 2.936 ;
      RECT 20.155 2.817 20.19 2.941 ;
      RECT 20.111 2.824 20.155 2.949 ;
      RECT 20.025 2.836 20.111 2.962 ;
      RECT 20 2.847 20.025 2.973 ;
      RECT 19.97 2.852 20 2.978 ;
      RECT 19.935 2.857 19.97 2.986 ;
      RECT 19.905 2.862 19.935 2.993 ;
      RECT 19.88 2.867 19.905 2.998 ;
      RECT 19.815 2.874 19.88 3.007 ;
      RECT 19.745 2.887 19.815 3.023 ;
      RECT 19.715 2.897 19.745 3.035 ;
      RECT 19.69 2.902 19.715 3.042 ;
      RECT 19.635 2.909 19.69 3.05 ;
      RECT 19.63 2.916 19.635 3.055 ;
      RECT 19.625 2.918 19.63 3.056 ;
      RECT 19.61 2.92 19.625 3.058 ;
      RECT 19.605 2.92 19.61 3.061 ;
      RECT 19.54 2.927 19.605 3.068 ;
      RECT 19.505 2.937 19.535 3.078 ;
      RECT 19.488 2.94 19.505 3.08 ;
      RECT 19.402 2.939 19.488 3.079 ;
      RECT 19.316 2.937 19.402 3.076 ;
      RECT 19.23 2.936 19.316 3.074 ;
      RECT 19.129 2.934 19.195 3.073 ;
      RECT 19.043 2.931 19.129 3.071 ;
      RECT 18.957 2.927 19.043 3.069 ;
      RECT 18.871 2.924 18.957 3.068 ;
      RECT 18.785 2.921 18.871 3.066 ;
      RECT 18.685 2.92 18.77 3.063 ;
      RECT 18.635 2.918 18.685 3.061 ;
      RECT 18.615 2.915 18.635 3.059 ;
      RECT 18.595 2.913 18.615 3.056 ;
      RECT 18.57 2.909 18.595 3.053 ;
      RECT 18.525 2.903 18.57 3.048 ;
      RECT 18.485 2.897 18.525 3.04 ;
      RECT 18.46 2.892 18.485 3.033 ;
      RECT 18.405 2.885 18.46 3.025 ;
      RECT 18.381 2.878 18.405 3.018 ;
      RECT 18.295 2.869 18.381 3.008 ;
      RECT 18.265 2.861 18.295 2.998 ;
      RECT 18.235 2.857 18.265 2.993 ;
      RECT 18.23 2.854 18.235 2.99 ;
      RECT 18.225 2.853 18.23 2.99 ;
      RECT 18.15 2.846 18.225 2.983 ;
      RECT 18.111 2.837 18.15 2.972 ;
      RECT 18.025 2.827 18.111 2.96 ;
      RECT 17.985 2.817 18.025 2.948 ;
      RECT 17.946 2.812 17.985 2.941 ;
      RECT 17.86 2.802 17.946 2.93 ;
      RECT 17.82 2.79 17.86 2.919 ;
      RECT 17.785 2.775 17.82 2.912 ;
      RECT 17.775 2.765 17.785 2.909 ;
      RECT 17.755 2.75 17.775 2.907 ;
      RECT 17.725 2.72 17.755 2.903 ;
      RECT 17.715 2.7 17.725 2.898 ;
      RECT 17.71 2.692 17.715 2.895 ;
      RECT 17.705 2.685 17.71 2.893 ;
      RECT 17.69 2.672 17.705 2.886 ;
      RECT 17.685 2.662 17.69 2.878 ;
      RECT 17.68 2.655 17.685 2.873 ;
      RECT 17.675 2.65 17.68 2.869 ;
      RECT 17.66 2.637 17.675 2.861 ;
      RECT 17.655 2.547 17.66 2.85 ;
      RECT 17.65 2.542 17.655 2.843 ;
      RECT 17.575 2.54 17.65 2.803 ;
      RECT 17.545 2.54 17.575 2.758 ;
      RECT 17.45 2.545 17.465 2.745 ;
      RECT 19.935 2.25 20.195 2.51 ;
      RECT 19.92 2.238 20.1 2.475 ;
      RECT 19.915 2.239 20.1 2.473 ;
      RECT 19.9 2.243 20.11 2.463 ;
      RECT 19.895 2.248 20.115 2.433 ;
      RECT 19.9 2.245 20.115 2.463 ;
      RECT 19.915 2.24 20.11 2.473 ;
      RECT 19.935 2.237 20.1 2.51 ;
      RECT 19.935 2.236 20.09 2.51 ;
      RECT 19.96 2.235 20.09 2.51 ;
      RECT 19.52 2.48 19.78 2.74 ;
      RECT 19.395 2.525 19.78 2.735 ;
      RECT 19.385 2.53 19.78 2.73 ;
      RECT 19.4 3.47 19.415 3.78 ;
      RECT 17.995 3.24 18.005 3.37 ;
      RECT 17.775 3.235 17.88 3.37 ;
      RECT 17.69 3.24 17.74 3.37 ;
      RECT 16.24 1.975 16.245 3.08 ;
      RECT 19.495 3.562 19.5 3.698 ;
      RECT 19.49 3.557 19.495 3.758 ;
      RECT 19.485 3.555 19.49 3.771 ;
      RECT 19.47 3.552 19.485 3.773 ;
      RECT 19.465 3.547 19.47 3.775 ;
      RECT 19.46 3.543 19.465 3.778 ;
      RECT 19.445 3.538 19.46 3.78 ;
      RECT 19.415 3.53 19.445 3.78 ;
      RECT 19.376 3.47 19.4 3.78 ;
      RECT 19.29 3.47 19.376 3.777 ;
      RECT 19.26 3.47 19.29 3.77 ;
      RECT 19.235 3.47 19.26 3.763 ;
      RECT 19.21 3.47 19.235 3.755 ;
      RECT 19.195 3.47 19.21 3.748 ;
      RECT 19.17 3.47 19.195 3.74 ;
      RECT 19.155 3.47 19.17 3.733 ;
      RECT 19.115 3.48 19.155 3.722 ;
      RECT 19.105 3.475 19.115 3.712 ;
      RECT 19.101 3.474 19.105 3.709 ;
      RECT 19.015 3.466 19.101 3.692 ;
      RECT 18.982 3.455 19.015 3.669 ;
      RECT 18.896 3.444 18.982 3.647 ;
      RECT 18.81 3.428 18.896 3.616 ;
      RECT 18.74 3.413 18.81 3.588 ;
      RECT 18.73 3.406 18.74 3.575 ;
      RECT 18.7 3.403 18.73 3.565 ;
      RECT 18.675 3.399 18.7 3.558 ;
      RECT 18.66 3.396 18.675 3.553 ;
      RECT 18.655 3.395 18.66 3.548 ;
      RECT 18.625 3.39 18.655 3.541 ;
      RECT 18.62 3.385 18.625 3.536 ;
      RECT 18.605 3.382 18.62 3.531 ;
      RECT 18.6 3.377 18.605 3.526 ;
      RECT 18.58 3.372 18.6 3.523 ;
      RECT 18.565 3.367 18.58 3.515 ;
      RECT 18.55 3.361 18.565 3.51 ;
      RECT 18.52 3.352 18.55 3.503 ;
      RECT 18.515 3.345 18.52 3.495 ;
      RECT 18.51 3.343 18.515 3.493 ;
      RECT 18.505 3.342 18.51 3.49 ;
      RECT 18.465 3.335 18.505 3.483 ;
      RECT 18.451 3.325 18.465 3.473 ;
      RECT 18.4 3.314 18.451 3.461 ;
      RECT 18.375 3.3 18.4 3.447 ;
      RECT 18.35 3.289 18.375 3.439 ;
      RECT 18.33 3.278 18.35 3.433 ;
      RECT 18.32 3.272 18.33 3.428 ;
      RECT 18.315 3.27 18.32 3.424 ;
      RECT 18.295 3.265 18.315 3.419 ;
      RECT 18.265 3.255 18.295 3.409 ;
      RECT 18.26 3.247 18.265 3.402 ;
      RECT 18.245 3.245 18.26 3.398 ;
      RECT 18.225 3.245 18.245 3.393 ;
      RECT 18.22 3.244 18.225 3.391 ;
      RECT 18.215 3.244 18.22 3.388 ;
      RECT 18.175 3.243 18.215 3.383 ;
      RECT 18.15 3.242 18.175 3.378 ;
      RECT 18.09 3.241 18.15 3.375 ;
      RECT 18.005 3.24 18.09 3.373 ;
      RECT 17.966 3.239 17.995 3.37 ;
      RECT 17.88 3.237 17.966 3.37 ;
      RECT 17.74 3.237 17.775 3.37 ;
      RECT 17.65 3.241 17.69 3.373 ;
      RECT 17.635 3.244 17.65 3.38 ;
      RECT 17.625 3.245 17.635 3.387 ;
      RECT 17.6 3.248 17.625 3.392 ;
      RECT 17.595 3.25 17.6 3.395 ;
      RECT 17.545 3.252 17.595 3.396 ;
      RECT 17.506 3.256 17.545 3.398 ;
      RECT 17.42 3.258 17.506 3.401 ;
      RECT 17.402 3.26 17.42 3.403 ;
      RECT 17.316 3.263 17.402 3.405 ;
      RECT 17.23 3.267 17.316 3.408 ;
      RECT 17.193 3.271 17.23 3.411 ;
      RECT 17.107 3.274 17.193 3.414 ;
      RECT 17.021 3.278 17.107 3.417 ;
      RECT 16.935 3.283 17.021 3.421 ;
      RECT 16.915 3.285 16.935 3.424 ;
      RECT 16.895 3.284 16.915 3.425 ;
      RECT 16.846 3.281 16.895 3.426 ;
      RECT 16.76 3.276 16.846 3.429 ;
      RECT 16.71 3.271 16.76 3.431 ;
      RECT 16.686 3.269 16.71 3.432 ;
      RECT 16.6 3.264 16.686 3.434 ;
      RECT 16.575 3.26 16.6 3.433 ;
      RECT 16.565 3.257 16.575 3.431 ;
      RECT 16.555 3.25 16.565 3.428 ;
      RECT 16.55 3.23 16.555 3.423 ;
      RECT 16.54 3.2 16.55 3.418 ;
      RECT 16.525 3.07 16.54 3.409 ;
      RECT 16.52 3.062 16.525 3.402 ;
      RECT 16.5 3.055 16.52 3.394 ;
      RECT 16.495 3.037 16.5 3.386 ;
      RECT 16.485 3.017 16.495 3.381 ;
      RECT 16.48 2.99 16.485 3.377 ;
      RECT 16.475 2.967 16.48 3.374 ;
      RECT 16.455 2.925 16.475 3.366 ;
      RECT 16.42 2.84 16.455 3.35 ;
      RECT 16.415 2.772 16.42 3.338 ;
      RECT 16.4 2.742 16.415 3.332 ;
      RECT 16.395 1.987 16.4 2.233 ;
      RECT 16.385 2.712 16.4 3.323 ;
      RECT 16.39 1.982 16.395 2.265 ;
      RECT 16.385 1.977 16.39 2.308 ;
      RECT 16.38 1.975 16.385 2.343 ;
      RECT 16.365 2.675 16.385 3.313 ;
      RECT 16.375 1.975 16.38 2.38 ;
      RECT 16.36 1.975 16.375 2.478 ;
      RECT 16.36 2.648 16.365 3.306 ;
      RECT 16.355 1.975 16.36 2.553 ;
      RECT 16.355 2.636 16.36 3.303 ;
      RECT 16.35 1.975 16.355 2.585 ;
      RECT 16.35 2.615 16.355 3.3 ;
      RECT 16.345 1.975 16.35 3.297 ;
      RECT 16.31 1.975 16.345 3.283 ;
      RECT 16.295 1.975 16.31 3.265 ;
      RECT 16.275 1.975 16.295 3.255 ;
      RECT 16.25 1.975 16.275 3.238 ;
      RECT 16.245 1.975 16.25 3.188 ;
      RECT 16.235 1.975 16.24 3.018 ;
      RECT 16.23 1.975 16.235 2.925 ;
      RECT 16.225 1.975 16.23 2.838 ;
      RECT 16.22 1.975 16.225 2.77 ;
      RECT 16.215 1.975 16.22 2.713 ;
      RECT 16.205 1.975 16.215 2.608 ;
      RECT 16.2 1.975 16.205 2.48 ;
      RECT 16.195 1.975 16.2 2.398 ;
      RECT 16.19 1.977 16.195 2.315 ;
      RECT 16.185 1.982 16.19 2.248 ;
      RECT 16.18 1.987 16.185 2.175 ;
      RECT 18.995 2.305 19.255 2.565 ;
      RECT 19.015 2.272 19.225 2.565 ;
      RECT 19.015 2.27 19.215 2.565 ;
      RECT 19.025 2.257 19.215 2.565 ;
      RECT 19.025 2.255 19.14 2.565 ;
      RECT 18.5 2.38 18.675 2.66 ;
      RECT 18.495 2.38 18.675 2.658 ;
      RECT 18.495 2.38 18.69 2.655 ;
      RECT 18.485 2.38 18.69 2.653 ;
      RECT 18.43 2.38 18.69 2.64 ;
      RECT 18.43 2.455 18.695 2.618 ;
      RECT 17.975 2.392 17.995 2.635 ;
      RECT 17.975 2.392 18.035 2.634 ;
      RECT 17.97 2.394 18.035 2.633 ;
      RECT 17.97 2.394 18.121 2.632 ;
      RECT 17.97 2.394 18.19 2.631 ;
      RECT 17.97 2.394 18.21 2.623 ;
      RECT 17.95 2.397 18.21 2.621 ;
      RECT 17.935 2.407 18.21 2.606 ;
      RECT 17.935 2.407 18.225 2.605 ;
      RECT 17.93 2.416 18.225 2.597 ;
      RECT 17.93 2.416 18.23 2.593 ;
      RECT 18.035 2.33 18.295 2.59 ;
      RECT 17.925 2.418 18.295 2.475 ;
      RECT 17.995 2.385 18.295 2.59 ;
      RECT 17.96 3.578 17.965 3.785 ;
      RECT 17.91 3.572 17.96 3.784 ;
      RECT 17.877 3.586 17.97 3.783 ;
      RECT 17.791 3.586 17.97 3.782 ;
      RECT 17.705 3.586 17.97 3.781 ;
      RECT 17.705 3.685 17.975 3.778 ;
      RECT 17.7 3.685 17.975 3.773 ;
      RECT 17.695 3.685 17.975 3.755 ;
      RECT 17.69 3.685 17.975 3.738 ;
      RECT 17.65 3.47 17.91 3.73 ;
      RECT 17.11 2.62 17.196 3.034 ;
      RECT 17.11 2.62 17.235 3.031 ;
      RECT 17.11 2.62 17.255 3.021 ;
      RECT 17.065 2.62 17.255 3.018 ;
      RECT 17.065 2.772 17.265 3.008 ;
      RECT 17.065 2.793 17.27 3.002 ;
      RECT 17.065 2.811 17.275 2.998 ;
      RECT 17.065 2.831 17.285 2.993 ;
      RECT 17.04 2.831 17.285 2.99 ;
      RECT 17.03 2.831 17.285 2.968 ;
      RECT 17.03 2.847 17.29 2.938 ;
      RECT 16.995 2.62 17.255 2.925 ;
      RECT 16.995 2.859 17.295 2.88 ;
      RECT 14.66 7.765 14.95 7.995 ;
      RECT 14.72 6.285 14.89 7.995 ;
      RECT 14.71 6.655 15.06 7.005 ;
      RECT 14.66 6.285 14.95 6.515 ;
      RECT 14.66 2.365 14.95 2.595 ;
      RECT 14.72 0.885 14.89 2.595 ;
      RECT 14.66 0.885 14.95 1.115 ;
      RECT 14.25 2.735 14.58 2.965 ;
      RECT 14.25 2.765 14.75 2.935 ;
      RECT 14.25 2.395 14.44 2.965 ;
      RECT 13.67 2.365 13.96 2.595 ;
      RECT 13.67 2.395 14.44 2.565 ;
      RECT 13.73 0.885 13.9 2.595 ;
      RECT 13.67 0.885 13.96 1.115 ;
      RECT 13.67 7.765 13.96 7.995 ;
      RECT 13.73 6.285 13.9 7.995 ;
      RECT 13.67 6.285 13.96 6.515 ;
      RECT 13.67 6.325 14.52 6.485 ;
      RECT 14.35 5.915 14.52 6.485 ;
      RECT 13.67 6.32 14.06 6.485 ;
      RECT 14.29 5.915 14.58 6.145 ;
      RECT 14.29 5.945 14.75 6.115 ;
      RECT 13.3 2.735 13.59 2.965 ;
      RECT 13.3 2.765 13.76 2.935 ;
      RECT 13.36 1.655 13.525 2.965 ;
      RECT 11.875 1.625 12.165 1.855 ;
      RECT 11.875 1.655 13.525 1.825 ;
      RECT 11.935 0.885 12.105 1.855 ;
      RECT 11.875 0.885 12.165 1.115 ;
      RECT 11.875 7.765 12.165 7.995 ;
      RECT 11.935 7.025 12.105 7.995 ;
      RECT 11.935 7.12 13.525 7.29 ;
      RECT 13.355 5.915 13.525 7.29 ;
      RECT 11.875 7.025 12.165 7.255 ;
      RECT 13.3 5.915 13.59 6.145 ;
      RECT 13.3 5.945 13.76 6.115 ;
      RECT 9.925 2.705 10.265 3.055 ;
      RECT 10.015 2.025 10.185 3.055 ;
      RECT 12.305 1.965 12.655 2.315 ;
      RECT 10.015 2.025 12.655 2.195 ;
      RECT 12.33 6.655 12.655 6.98 ;
      RECT 6.87 6.605 7.22 6.955 ;
      RECT 12.305 6.655 12.655 6.885 ;
      RECT 6.67 6.655 7.22 6.885 ;
      RECT 6.5 6.685 12.655 6.855 ;
      RECT 11.53 2.365 11.85 2.685 ;
      RECT 11.5 2.365 11.85 2.595 ;
      RECT 11.33 2.395 11.85 2.565 ;
      RECT 11.53 6.255 11.85 6.545 ;
      RECT 11.5 6.285 11.85 6.515 ;
      RECT 11.33 6.315 11.85 6.485 ;
      RECT 10.485 2.705 10.825 3.055 ;
      RECT 10.485 2.765 10.965 2.935 ;
      RECT 10.48 5.86 10.82 6.21 ;
      RECT 4.87 5.915 5.16 6.145 ;
      RECT 4.87 5.945 10.965 6.115 ;
      RECT 7.22 2.985 7.37 3.26 ;
      RECT 7.76 2.065 7.765 2.285 ;
      RECT 8.91 2.265 8.925 2.463 ;
      RECT 8.875 2.257 8.91 2.47 ;
      RECT 8.845 2.25 8.875 2.47 ;
      RECT 8.79 2.215 8.845 2.47 ;
      RECT 8.725 2.152 8.79 2.47 ;
      RECT 8.72 2.117 8.725 2.468 ;
      RECT 8.715 2.112 8.72 2.46 ;
      RECT 8.71 2.107 8.715 2.446 ;
      RECT 8.705 2.104 8.71 2.439 ;
      RECT 8.66 2.094 8.705 2.39 ;
      RECT 8.64 2.081 8.66 2.325 ;
      RECT 8.635 2.076 8.64 2.298 ;
      RECT 8.63 2.075 8.635 2.291 ;
      RECT 8.625 2.074 8.63 2.284 ;
      RECT 8.54 2.059 8.625 2.23 ;
      RECT 8.51 2.04 8.54 2.18 ;
      RECT 8.43 2.023 8.51 2.165 ;
      RECT 8.395 2.01 8.43 2.15 ;
      RECT 8.387 2.01 8.395 2.145 ;
      RECT 8.301 2.011 8.387 2.145 ;
      RECT 8.215 2.013 8.301 2.145 ;
      RECT 8.19 2.014 8.215 2.149 ;
      RECT 8.115 2.02 8.19 2.164 ;
      RECT 8.032 2.032 8.115 2.188 ;
      RECT 7.946 2.045 8.032 2.214 ;
      RECT 7.86 2.058 7.946 2.24 ;
      RECT 7.825 2.067 7.86 2.259 ;
      RECT 7.775 2.067 7.825 2.272 ;
      RECT 7.765 2.065 7.775 2.283 ;
      RECT 7.75 2.062 7.76 2.285 ;
      RECT 7.735 2.054 7.75 2.293 ;
      RECT 7.72 2.046 7.735 2.313 ;
      RECT 7.715 2.041 7.72 2.37 ;
      RECT 7.7 2.036 7.715 2.443 ;
      RECT 7.695 2.031 7.7 2.485 ;
      RECT 7.69 2.029 7.695 2.513 ;
      RECT 7.685 2.027 7.69 2.535 ;
      RECT 7.675 2.023 7.685 2.578 ;
      RECT 7.67 2.02 7.675 2.603 ;
      RECT 7.665 2.018 7.67 2.623 ;
      RECT 7.66 2.016 7.665 2.647 ;
      RECT 7.655 2.012 7.66 2.67 ;
      RECT 7.65 2.008 7.655 2.693 ;
      RECT 7.615 1.998 7.65 2.8 ;
      RECT 7.61 1.988 7.615 2.898 ;
      RECT 7.605 1.986 7.61 2.925 ;
      RECT 7.6 1.985 7.605 2.945 ;
      RECT 7.595 1.977 7.6 2.965 ;
      RECT 7.59 1.972 7.595 3 ;
      RECT 7.585 1.97 7.59 3.018 ;
      RECT 7.58 1.97 7.585 3.043 ;
      RECT 7.575 1.97 7.58 3.065 ;
      RECT 7.54 1.97 7.575 3.108 ;
      RECT 7.515 1.97 7.54 3.137 ;
      RECT 7.505 1.97 7.515 2.323 ;
      RECT 7.508 2.38 7.515 3.147 ;
      RECT 7.505 2.437 7.508 3.15 ;
      RECT 7.5 1.97 7.505 2.295 ;
      RECT 7.5 2.487 7.505 3.153 ;
      RECT 7.49 1.97 7.5 2.285 ;
      RECT 7.495 2.54 7.5 3.156 ;
      RECT 7.49 2.625 7.495 3.16 ;
      RECT 7.48 1.97 7.49 2.273 ;
      RECT 7.485 2.672 7.49 3.164 ;
      RECT 7.48 2.747 7.485 3.168 ;
      RECT 7.445 1.97 7.48 2.248 ;
      RECT 7.47 2.83 7.48 3.173 ;
      RECT 7.46 2.897 7.47 3.18 ;
      RECT 7.455 2.925 7.46 3.185 ;
      RECT 7.445 2.938 7.455 3.191 ;
      RECT 7.4 1.97 7.445 2.205 ;
      RECT 7.44 2.943 7.445 3.198 ;
      RECT 7.4 2.96 7.44 3.26 ;
      RECT 7.395 1.972 7.4 2.178 ;
      RECT 7.37 2.98 7.4 3.26 ;
      RECT 7.39 1.977 7.395 2.15 ;
      RECT 7.18 2.989 7.22 3.26 ;
      RECT 7.155 2.997 7.18 3.23 ;
      RECT 7.11 3.005 7.155 3.23 ;
      RECT 7.095 3.01 7.11 3.225 ;
      RECT 7.085 3.01 7.095 3.219 ;
      RECT 7.075 3.017 7.085 3.216 ;
      RECT 7.07 3.055 7.075 3.205 ;
      RECT 7.065 3.117 7.07 3.183 ;
      RECT 8.335 2.992 8.52 3.215 ;
      RECT 8.335 3.007 8.525 3.211 ;
      RECT 8.325 2.28 8.41 3.21 ;
      RECT 8.325 3.007 8.53 3.204 ;
      RECT 8.32 3.015 8.53 3.203 ;
      RECT 8.525 2.735 8.845 3.055 ;
      RECT 8.32 2.907 8.49 2.998 ;
      RECT 8.315 2.907 8.49 2.98 ;
      RECT 8.305 2.715 8.44 2.955 ;
      RECT 8.3 2.715 8.44 2.9 ;
      RECT 8.26 2.295 8.43 2.8 ;
      RECT 8.245 2.295 8.43 2.67 ;
      RECT 8.24 2.295 8.43 2.623 ;
      RECT 8.235 2.295 8.43 2.603 ;
      RECT 8.23 2.295 8.43 2.578 ;
      RECT 8.2 2.295 8.46 2.555 ;
      RECT 8.21 2.292 8.42 2.555 ;
      RECT 8.335 2.287 8.42 3.215 ;
      RECT 8.22 2.28 8.41 2.555 ;
      RECT 8.215 2.285 8.41 2.555 ;
      RECT 7.045 2.497 7.23 2.71 ;
      RECT 7.045 2.505 7.24 2.703 ;
      RECT 7.025 2.505 7.24 2.7 ;
      RECT 7.02 2.505 7.24 2.685 ;
      RECT 6.95 2.42 7.21 2.68 ;
      RECT 6.95 2.565 7.245 2.593 ;
      RECT 6.605 3.02 6.865 3.28 ;
      RECT 6.63 2.965 6.825 3.28 ;
      RECT 6.625 2.714 6.805 3.008 ;
      RECT 6.625 2.72 6.815 3.008 ;
      RECT 6.605 2.722 6.815 2.953 ;
      RECT 6.6 2.732 6.815 2.82 ;
      RECT 6.63 2.712 6.805 3.28 ;
      RECT 6.716 2.71 6.805 3.28 ;
      RECT 6.575 1.93 6.61 2.3 ;
      RECT 6.365 2.04 6.37 2.3 ;
      RECT 6.61 1.937 6.625 2.3 ;
      RECT 6.5 1.93 6.575 2.378 ;
      RECT 6.49 1.93 6.5 2.463 ;
      RECT 6.465 1.93 6.49 2.498 ;
      RECT 6.425 1.93 6.465 2.566 ;
      RECT 6.415 1.937 6.425 2.618 ;
      RECT 6.385 2.04 6.415 2.659 ;
      RECT 6.38 2.04 6.385 2.698 ;
      RECT 6.37 2.04 6.38 2.718 ;
      RECT 6.365 2.335 6.37 2.755 ;
      RECT 6.36 2.352 6.365 2.775 ;
      RECT 6.345 2.415 6.36 2.815 ;
      RECT 6.34 2.458 6.345 2.85 ;
      RECT 6.335 2.466 6.34 2.863 ;
      RECT 6.325 2.48 6.335 2.885 ;
      RECT 6.3 2.515 6.325 2.95 ;
      RECT 6.29 2.55 6.3 3.013 ;
      RECT 6.27 2.58 6.29 3.074 ;
      RECT 6.255 2.616 6.27 3.141 ;
      RECT 6.245 2.644 6.255 3.18 ;
      RECT 6.235 2.666 6.245 3.2 ;
      RECT 6.23 2.676 6.235 3.211 ;
      RECT 6.225 2.685 6.23 3.214 ;
      RECT 6.215 2.703 6.225 3.218 ;
      RECT 6.205 2.721 6.215 3.219 ;
      RECT 6.18 2.76 6.205 3.216 ;
      RECT 6.16 2.802 6.18 3.213 ;
      RECT 6.145 2.84 6.16 3.212 ;
      RECT 6.11 2.875 6.145 3.209 ;
      RECT 6.105 2.897 6.11 3.207 ;
      RECT 6.04 2.937 6.105 3.204 ;
      RECT 6.035 2.977 6.04 3.2 ;
      RECT 6.02 2.987 6.035 3.191 ;
      RECT 6.01 3.107 6.02 3.176 ;
      RECT 6.49 3.52 6.5 3.78 ;
      RECT 6.49 3.523 6.51 3.779 ;
      RECT 6.48 3.513 6.49 3.778 ;
      RECT 6.47 3.528 6.55 3.774 ;
      RECT 6.455 3.507 6.47 3.772 ;
      RECT 6.43 3.532 6.555 3.768 ;
      RECT 6.415 3.492 6.43 3.763 ;
      RECT 6.415 3.534 6.565 3.762 ;
      RECT 6.415 3.542 6.58 3.755 ;
      RECT 6.355 3.479 6.415 3.745 ;
      RECT 6.345 3.466 6.355 3.727 ;
      RECT 6.32 3.456 6.345 3.717 ;
      RECT 6.315 3.446 6.32 3.709 ;
      RECT 6.25 3.542 6.58 3.691 ;
      RECT 6.165 3.542 6.58 3.653 ;
      RECT 6.055 3.37 6.315 3.63 ;
      RECT 6.43 3.5 6.455 3.768 ;
      RECT 6.47 3.51 6.48 3.774 ;
      RECT 6.055 3.518 6.495 3.63 ;
      RECT 6.24 7.765 6.53 7.995 ;
      RECT 6.3 7.025 6.47 7.995 ;
      RECT 6.2 7.055 6.57 7.425 ;
      RECT 6.24 7.025 6.53 7.425 ;
      RECT 5.27 3.275 5.3 3.575 ;
      RECT 5.045 3.26 5.05 3.535 ;
      RECT 4.845 3.26 5 3.52 ;
      RECT 6.145 1.975 6.175 2.235 ;
      RECT 6.135 1.975 6.145 2.343 ;
      RECT 6.115 1.975 6.135 2.353 ;
      RECT 6.1 1.975 6.115 2.365 ;
      RECT 6.045 1.975 6.1 2.415 ;
      RECT 6.03 1.975 6.045 2.463 ;
      RECT 6 1.975 6.03 2.498 ;
      RECT 5.945 1.975 6 2.56 ;
      RECT 5.925 1.975 5.945 2.628 ;
      RECT 5.92 1.975 5.925 2.658 ;
      RECT 5.915 1.975 5.92 2.67 ;
      RECT 5.91 2.092 5.915 2.688 ;
      RECT 5.89 2.11 5.91 2.713 ;
      RECT 5.87 2.137 5.89 2.763 ;
      RECT 5.865 2.157 5.87 2.794 ;
      RECT 5.86 2.165 5.865 2.811 ;
      RECT 5.845 2.191 5.86 2.84 ;
      RECT 5.83 2.233 5.845 2.875 ;
      RECT 5.825 2.262 5.83 2.898 ;
      RECT 5.82 2.277 5.825 2.911 ;
      RECT 5.815 2.3 5.82 2.922 ;
      RECT 5.805 2.32 5.815 2.94 ;
      RECT 5.795 2.35 5.805 2.963 ;
      RECT 5.79 2.372 5.795 2.983 ;
      RECT 5.785 2.387 5.79 2.998 ;
      RECT 5.77 2.417 5.785 3.025 ;
      RECT 5.765 2.447 5.77 3.051 ;
      RECT 5.76 2.465 5.765 3.063 ;
      RECT 5.75 2.495 5.76 3.082 ;
      RECT 5.74 2.52 5.75 3.107 ;
      RECT 5.735 2.54 5.74 3.126 ;
      RECT 5.73 2.557 5.735 3.139 ;
      RECT 5.72 2.583 5.73 3.158 ;
      RECT 5.71 2.621 5.72 3.185 ;
      RECT 5.705 2.647 5.71 3.205 ;
      RECT 5.7 2.657 5.705 3.215 ;
      RECT 5.695 2.67 5.7 3.23 ;
      RECT 5.69 2.685 5.695 3.24 ;
      RECT 5.685 2.707 5.69 3.255 ;
      RECT 5.68 2.725 5.685 3.266 ;
      RECT 5.675 2.735 5.68 3.277 ;
      RECT 5.67 2.743 5.675 3.289 ;
      RECT 5.665 2.751 5.67 3.3 ;
      RECT 5.66 2.777 5.665 3.313 ;
      RECT 5.65 2.805 5.66 3.326 ;
      RECT 5.645 2.835 5.65 3.335 ;
      RECT 5.64 2.85 5.645 3.342 ;
      RECT 5.625 2.875 5.64 3.349 ;
      RECT 5.62 2.897 5.625 3.355 ;
      RECT 5.615 2.922 5.62 3.358 ;
      RECT 5.606 2.95 5.615 3.362 ;
      RECT 5.6 2.967 5.606 3.367 ;
      RECT 5.595 2.985 5.6 3.371 ;
      RECT 5.59 2.997 5.595 3.374 ;
      RECT 5.585 3.018 5.59 3.378 ;
      RECT 5.58 3.036 5.585 3.381 ;
      RECT 5.575 3.05 5.58 3.384 ;
      RECT 5.57 3.067 5.575 3.387 ;
      RECT 5.565 3.08 5.57 3.39 ;
      RECT 5.54 3.117 5.565 3.398 ;
      RECT 5.535 3.162 5.54 3.407 ;
      RECT 5.53 3.19 5.535 3.41 ;
      RECT 5.52 3.21 5.53 3.414 ;
      RECT 5.515 3.23 5.52 3.419 ;
      RECT 5.51 3.245 5.515 3.422 ;
      RECT 5.49 3.255 5.51 3.429 ;
      RECT 5.425 3.262 5.49 3.455 ;
      RECT 5.39 3.265 5.425 3.483 ;
      RECT 5.375 3.268 5.39 3.498 ;
      RECT 5.365 3.269 5.375 3.513 ;
      RECT 5.355 3.27 5.365 3.53 ;
      RECT 5.35 3.27 5.355 3.545 ;
      RECT 5.345 3.27 5.35 3.553 ;
      RECT 5.33 3.271 5.345 3.568 ;
      RECT 5.3 3.273 5.33 3.575 ;
      RECT 5.19 3.28 5.27 3.575 ;
      RECT 5.145 3.285 5.19 3.575 ;
      RECT 5.135 3.286 5.145 3.565 ;
      RECT 5.125 3.287 5.135 3.558 ;
      RECT 5.105 3.289 5.125 3.553 ;
      RECT 5.095 3.26 5.105 3.548 ;
      RECT 5.05 3.26 5.095 3.54 ;
      RECT 5.02 3.26 5.045 3.53 ;
      RECT 5 3.26 5.02 3.523 ;
      RECT 5.28 2.06 5.54 2.32 ;
      RECT 5.16 2.075 5.17 2.24 ;
      RECT 5.145 2.075 5.15 2.235 ;
      RECT 2.51 1.915 2.695 2.205 ;
      RECT 4.325 2.04 4.34 2.195 ;
      RECT 2.475 1.915 2.5 2.175 ;
      RECT 4.89 1.965 4.895 2.107 ;
      RECT 4.805 1.96 4.83 2.1 ;
      RECT 5.205 2.077 5.28 2.27 ;
      RECT 5.19 2.075 5.205 2.253 ;
      RECT 5.17 2.075 5.19 2.245 ;
      RECT 5.15 2.075 5.16 2.238 ;
      RECT 5.105 2.07 5.145 2.228 ;
      RECT 5.065 2.045 5.105 2.213 ;
      RECT 5.05 2.02 5.065 2.203 ;
      RECT 5.045 2.014 5.05 2.201 ;
      RECT 5.01 2.006 5.045 2.184 ;
      RECT 5.005 1.999 5.01 2.172 ;
      RECT 4.985 1.994 5.005 2.16 ;
      RECT 4.975 1.988 4.985 2.145 ;
      RECT 4.955 1.983 4.975 2.13 ;
      RECT 4.945 1.978 4.955 2.123 ;
      RECT 4.94 1.976 4.945 2.118 ;
      RECT 4.935 1.975 4.94 2.115 ;
      RECT 4.895 1.97 4.935 2.111 ;
      RECT 4.875 1.964 4.89 2.106 ;
      RECT 4.84 1.961 4.875 2.103 ;
      RECT 4.83 1.96 4.84 2.101 ;
      RECT 4.77 1.96 4.805 2.098 ;
      RECT 4.725 1.96 4.77 2.098 ;
      RECT 4.675 1.96 4.725 2.101 ;
      RECT 4.66 1.962 4.675 2.103 ;
      RECT 4.645 1.965 4.66 2.104 ;
      RECT 4.635 1.97 4.645 2.105 ;
      RECT 4.605 1.975 4.635 2.11 ;
      RECT 4.595 1.981 4.605 2.118 ;
      RECT 4.585 1.983 4.595 2.122 ;
      RECT 4.575 1.987 4.585 2.126 ;
      RECT 4.55 1.993 4.575 2.134 ;
      RECT 4.54 1.998 4.55 2.142 ;
      RECT 4.525 2.002 4.54 2.146 ;
      RECT 4.49 2.008 4.525 2.154 ;
      RECT 4.47 2.013 4.49 2.164 ;
      RECT 4.44 2.02 4.47 2.173 ;
      RECT 4.395 2.029 4.44 2.187 ;
      RECT 4.39 2.034 4.395 2.198 ;
      RECT 4.37 2.037 4.39 2.199 ;
      RECT 4.34 2.04 4.37 2.197 ;
      RECT 4.305 2.04 4.325 2.193 ;
      RECT 4.235 2.04 4.305 2.184 ;
      RECT 4.22 2.037 4.235 2.176 ;
      RECT 4.18 2.03 4.22 2.171 ;
      RECT 4.155 2.02 4.18 2.164 ;
      RECT 4.15 2.014 4.155 2.161 ;
      RECT 4.11 2.008 4.15 2.158 ;
      RECT 4.095 2.001 4.11 2.153 ;
      RECT 4.075 1.997 4.095 2.148 ;
      RECT 4.06 1.992 4.075 2.144 ;
      RECT 4.045 1.987 4.06 2.142 ;
      RECT 4.03 1.983 4.045 2.141 ;
      RECT 4.015 1.981 4.03 2.137 ;
      RECT 4.005 1.979 4.015 2.132 ;
      RECT 3.99 1.976 4.005 2.128 ;
      RECT 3.98 1.974 3.99 2.123 ;
      RECT 3.96 1.971 3.98 2.119 ;
      RECT 3.915 1.97 3.96 2.117 ;
      RECT 3.855 1.972 3.915 2.118 ;
      RECT 3.835 1.974 3.855 2.12 ;
      RECT 3.805 1.977 3.835 2.121 ;
      RECT 3.755 1.982 3.805 2.123 ;
      RECT 3.75 1.985 3.755 2.125 ;
      RECT 3.74 1.987 3.75 2.128 ;
      RECT 3.735 1.989 3.74 2.131 ;
      RECT 3.685 1.992 3.735 2.138 ;
      RECT 3.665 1.996 3.685 2.15 ;
      RECT 3.655 1.999 3.665 2.156 ;
      RECT 3.645 2 3.655 2.159 ;
      RECT 3.606 2.003 3.645 2.161 ;
      RECT 3.52 2.01 3.606 2.164 ;
      RECT 3.446 2.02 3.52 2.168 ;
      RECT 3.36 2.031 3.446 2.173 ;
      RECT 3.345 2.038 3.36 2.175 ;
      RECT 3.29 2.042 3.345 2.176 ;
      RECT 3.276 2.045 3.29 2.178 ;
      RECT 3.19 2.045 3.276 2.18 ;
      RECT 3.15 2.042 3.19 2.183 ;
      RECT 3.126 2.038 3.15 2.185 ;
      RECT 3.04 2.028 3.126 2.188 ;
      RECT 3.01 2.017 3.04 2.189 ;
      RECT 2.991 2.013 3.01 2.188 ;
      RECT 2.905 2.006 2.991 2.185 ;
      RECT 2.845 1.995 2.905 2.182 ;
      RECT 2.825 1.987 2.845 2.18 ;
      RECT 2.79 1.982 2.825 2.179 ;
      RECT 2.765 1.977 2.79 2.178 ;
      RECT 2.735 1.972 2.765 2.177 ;
      RECT 2.71 1.915 2.735 2.176 ;
      RECT 2.695 1.915 2.71 2.2 ;
      RECT 2.5 1.915 2.51 2.2 ;
      RECT 4.275 2.935 4.28 3.075 ;
      RECT 3.935 2.935 3.97 3.073 ;
      RECT 3.51 2.92 3.525 3.065 ;
      RECT 5.34 2.7 5.43 2.96 ;
      RECT 5.17 2.565 5.27 2.96 ;
      RECT 2.205 2.54 2.285 2.75 ;
      RECT 5.295 2.677 5.34 2.96 ;
      RECT 5.285 2.647 5.295 2.96 ;
      RECT 5.27 2.57 5.285 2.96 ;
      RECT 5.085 2.565 5.17 2.925 ;
      RECT 5.08 2.567 5.085 2.92 ;
      RECT 5.075 2.572 5.08 2.92 ;
      RECT 5.04 2.672 5.075 2.92 ;
      RECT 5.03 2.7 5.04 2.92 ;
      RECT 5.02 2.715 5.03 2.92 ;
      RECT 5.01 2.727 5.02 2.92 ;
      RECT 5.005 2.737 5.01 2.92 ;
      RECT 4.99 2.747 5.005 2.922 ;
      RECT 4.985 2.762 4.99 2.924 ;
      RECT 4.97 2.775 4.985 2.926 ;
      RECT 4.965 2.79 4.97 2.929 ;
      RECT 4.945 2.8 4.965 2.933 ;
      RECT 4.93 2.81 4.945 2.936 ;
      RECT 4.895 2.817 4.93 2.941 ;
      RECT 4.851 2.824 4.895 2.949 ;
      RECT 4.765 2.836 4.851 2.962 ;
      RECT 4.74 2.847 4.765 2.973 ;
      RECT 4.71 2.852 4.74 2.978 ;
      RECT 4.675 2.857 4.71 2.986 ;
      RECT 4.645 2.862 4.675 2.993 ;
      RECT 4.62 2.867 4.645 2.998 ;
      RECT 4.555 2.874 4.62 3.007 ;
      RECT 4.485 2.887 4.555 3.023 ;
      RECT 4.455 2.897 4.485 3.035 ;
      RECT 4.43 2.902 4.455 3.042 ;
      RECT 4.375 2.909 4.43 3.05 ;
      RECT 4.37 2.916 4.375 3.055 ;
      RECT 4.365 2.918 4.37 3.056 ;
      RECT 4.35 2.92 4.365 3.058 ;
      RECT 4.345 2.92 4.35 3.061 ;
      RECT 4.28 2.927 4.345 3.068 ;
      RECT 4.245 2.937 4.275 3.078 ;
      RECT 4.228 2.94 4.245 3.08 ;
      RECT 4.142 2.939 4.228 3.079 ;
      RECT 4.056 2.937 4.142 3.076 ;
      RECT 3.97 2.936 4.056 3.074 ;
      RECT 3.869 2.934 3.935 3.073 ;
      RECT 3.783 2.931 3.869 3.071 ;
      RECT 3.697 2.927 3.783 3.069 ;
      RECT 3.611 2.924 3.697 3.068 ;
      RECT 3.525 2.921 3.611 3.066 ;
      RECT 3.425 2.92 3.51 3.063 ;
      RECT 3.375 2.918 3.425 3.061 ;
      RECT 3.355 2.915 3.375 3.059 ;
      RECT 3.335 2.913 3.355 3.056 ;
      RECT 3.31 2.909 3.335 3.053 ;
      RECT 3.265 2.903 3.31 3.048 ;
      RECT 3.225 2.897 3.265 3.04 ;
      RECT 3.2 2.892 3.225 3.033 ;
      RECT 3.145 2.885 3.2 3.025 ;
      RECT 3.121 2.878 3.145 3.018 ;
      RECT 3.035 2.869 3.121 3.008 ;
      RECT 3.005 2.861 3.035 2.998 ;
      RECT 2.975 2.857 3.005 2.993 ;
      RECT 2.97 2.854 2.975 2.99 ;
      RECT 2.965 2.853 2.97 2.99 ;
      RECT 2.89 2.846 2.965 2.983 ;
      RECT 2.851 2.837 2.89 2.972 ;
      RECT 2.765 2.827 2.851 2.96 ;
      RECT 2.725 2.817 2.765 2.948 ;
      RECT 2.686 2.812 2.725 2.941 ;
      RECT 2.6 2.802 2.686 2.93 ;
      RECT 2.56 2.79 2.6 2.919 ;
      RECT 2.525 2.775 2.56 2.912 ;
      RECT 2.515 2.765 2.525 2.909 ;
      RECT 2.495 2.75 2.515 2.907 ;
      RECT 2.465 2.72 2.495 2.903 ;
      RECT 2.455 2.7 2.465 2.898 ;
      RECT 2.45 2.692 2.455 2.895 ;
      RECT 2.445 2.685 2.45 2.893 ;
      RECT 2.43 2.672 2.445 2.886 ;
      RECT 2.425 2.662 2.43 2.878 ;
      RECT 2.42 2.655 2.425 2.873 ;
      RECT 2.415 2.65 2.42 2.869 ;
      RECT 2.4 2.637 2.415 2.861 ;
      RECT 2.395 2.547 2.4 2.85 ;
      RECT 2.39 2.542 2.395 2.843 ;
      RECT 2.315 2.54 2.39 2.803 ;
      RECT 2.285 2.54 2.315 2.758 ;
      RECT 2.19 2.545 2.205 2.745 ;
      RECT 4.675 2.25 4.935 2.51 ;
      RECT 4.66 2.238 4.84 2.475 ;
      RECT 4.655 2.239 4.84 2.473 ;
      RECT 4.64 2.243 4.85 2.463 ;
      RECT 4.635 2.248 4.855 2.433 ;
      RECT 4.64 2.245 4.855 2.463 ;
      RECT 4.655 2.24 4.85 2.473 ;
      RECT 4.675 2.237 4.84 2.51 ;
      RECT 4.675 2.236 4.83 2.51 ;
      RECT 4.7 2.235 4.83 2.51 ;
      RECT 4.26 2.48 4.52 2.74 ;
      RECT 4.135 2.525 4.52 2.735 ;
      RECT 4.125 2.53 4.52 2.73 ;
      RECT 4.14 3.47 4.155 3.78 ;
      RECT 2.735 3.24 2.745 3.37 ;
      RECT 2.515 3.235 2.62 3.37 ;
      RECT 2.43 3.24 2.48 3.37 ;
      RECT 0.98 1.975 0.985 3.08 ;
      RECT 4.235 3.562 4.24 3.698 ;
      RECT 4.23 3.557 4.235 3.758 ;
      RECT 4.225 3.555 4.23 3.771 ;
      RECT 4.21 3.552 4.225 3.773 ;
      RECT 4.205 3.547 4.21 3.775 ;
      RECT 4.2 3.543 4.205 3.778 ;
      RECT 4.185 3.538 4.2 3.78 ;
      RECT 4.155 3.53 4.185 3.78 ;
      RECT 4.116 3.47 4.14 3.78 ;
      RECT 4.03 3.47 4.116 3.777 ;
      RECT 4 3.47 4.03 3.77 ;
      RECT 3.975 3.47 4 3.763 ;
      RECT 3.95 3.47 3.975 3.755 ;
      RECT 3.935 3.47 3.95 3.748 ;
      RECT 3.91 3.47 3.935 3.74 ;
      RECT 3.895 3.47 3.91 3.733 ;
      RECT 3.855 3.48 3.895 3.722 ;
      RECT 3.845 3.475 3.855 3.712 ;
      RECT 3.841 3.474 3.845 3.709 ;
      RECT 3.755 3.466 3.841 3.692 ;
      RECT 3.722 3.455 3.755 3.669 ;
      RECT 3.636 3.444 3.722 3.647 ;
      RECT 3.55 3.428 3.636 3.616 ;
      RECT 3.48 3.413 3.55 3.588 ;
      RECT 3.47 3.406 3.48 3.575 ;
      RECT 3.44 3.403 3.47 3.565 ;
      RECT 3.415 3.399 3.44 3.558 ;
      RECT 3.4 3.396 3.415 3.553 ;
      RECT 3.395 3.395 3.4 3.548 ;
      RECT 3.365 3.39 3.395 3.541 ;
      RECT 3.36 3.385 3.365 3.536 ;
      RECT 3.345 3.382 3.36 3.531 ;
      RECT 3.34 3.377 3.345 3.526 ;
      RECT 3.32 3.372 3.34 3.523 ;
      RECT 3.305 3.367 3.32 3.515 ;
      RECT 3.29 3.361 3.305 3.51 ;
      RECT 3.26 3.352 3.29 3.503 ;
      RECT 3.255 3.345 3.26 3.495 ;
      RECT 3.25 3.343 3.255 3.493 ;
      RECT 3.245 3.342 3.25 3.49 ;
      RECT 3.205 3.335 3.245 3.483 ;
      RECT 3.191 3.325 3.205 3.473 ;
      RECT 3.14 3.314 3.191 3.461 ;
      RECT 3.115 3.3 3.14 3.447 ;
      RECT 3.09 3.289 3.115 3.439 ;
      RECT 3.07 3.278 3.09 3.433 ;
      RECT 3.06 3.272 3.07 3.428 ;
      RECT 3.055 3.27 3.06 3.424 ;
      RECT 3.035 3.265 3.055 3.419 ;
      RECT 3.005 3.255 3.035 3.409 ;
      RECT 3 3.247 3.005 3.402 ;
      RECT 2.985 3.245 3 3.398 ;
      RECT 2.965 3.245 2.985 3.393 ;
      RECT 2.96 3.244 2.965 3.391 ;
      RECT 2.955 3.244 2.96 3.388 ;
      RECT 2.915 3.243 2.955 3.383 ;
      RECT 2.89 3.242 2.915 3.378 ;
      RECT 2.83 3.241 2.89 3.375 ;
      RECT 2.745 3.24 2.83 3.373 ;
      RECT 2.706 3.239 2.735 3.37 ;
      RECT 2.62 3.237 2.706 3.37 ;
      RECT 2.48 3.237 2.515 3.37 ;
      RECT 2.39 3.241 2.43 3.373 ;
      RECT 2.375 3.244 2.39 3.38 ;
      RECT 2.365 3.245 2.375 3.387 ;
      RECT 2.34 3.248 2.365 3.392 ;
      RECT 2.335 3.25 2.34 3.395 ;
      RECT 2.285 3.252 2.335 3.396 ;
      RECT 2.246 3.256 2.285 3.398 ;
      RECT 2.16 3.258 2.246 3.401 ;
      RECT 2.142 3.26 2.16 3.403 ;
      RECT 2.056 3.263 2.142 3.405 ;
      RECT 1.97 3.267 2.056 3.408 ;
      RECT 1.933 3.271 1.97 3.411 ;
      RECT 1.847 3.274 1.933 3.414 ;
      RECT 1.761 3.278 1.847 3.417 ;
      RECT 1.675 3.283 1.761 3.421 ;
      RECT 1.655 3.285 1.675 3.424 ;
      RECT 1.635 3.284 1.655 3.425 ;
      RECT 1.586 3.281 1.635 3.426 ;
      RECT 1.5 3.276 1.586 3.429 ;
      RECT 1.45 3.271 1.5 3.431 ;
      RECT 1.426 3.269 1.45 3.432 ;
      RECT 1.34 3.264 1.426 3.434 ;
      RECT 1.315 3.26 1.34 3.433 ;
      RECT 1.305 3.257 1.315 3.431 ;
      RECT 1.295 3.25 1.305 3.428 ;
      RECT 1.29 3.23 1.295 3.423 ;
      RECT 1.28 3.2 1.29 3.418 ;
      RECT 1.265 3.07 1.28 3.409 ;
      RECT 1.26 3.062 1.265 3.402 ;
      RECT 1.24 3.055 1.26 3.394 ;
      RECT 1.235 3.037 1.24 3.386 ;
      RECT 1.225 3.017 1.235 3.381 ;
      RECT 1.22 2.99 1.225 3.377 ;
      RECT 1.215 2.967 1.22 3.374 ;
      RECT 1.195 2.925 1.215 3.366 ;
      RECT 1.16 2.84 1.195 3.35 ;
      RECT 1.155 2.772 1.16 3.338 ;
      RECT 1.14 2.742 1.155 3.332 ;
      RECT 1.135 1.987 1.14 2.233 ;
      RECT 1.125 2.712 1.14 3.323 ;
      RECT 1.13 1.982 1.135 2.265 ;
      RECT 1.125 1.977 1.13 2.308 ;
      RECT 1.12 1.975 1.125 2.343 ;
      RECT 1.105 2.675 1.125 3.313 ;
      RECT 1.115 1.975 1.12 2.38 ;
      RECT 1.1 1.975 1.115 2.478 ;
      RECT 1.1 2.648 1.105 3.306 ;
      RECT 1.095 1.975 1.1 2.553 ;
      RECT 1.095 2.636 1.1 3.303 ;
      RECT 1.09 1.975 1.095 2.585 ;
      RECT 1.09 2.615 1.095 3.3 ;
      RECT 1.085 1.975 1.09 3.297 ;
      RECT 1.05 1.975 1.085 3.283 ;
      RECT 1.035 1.975 1.05 3.265 ;
      RECT 1.015 1.975 1.035 3.255 ;
      RECT 0.99 1.975 1.015 3.238 ;
      RECT 0.985 1.975 0.99 3.188 ;
      RECT 0.975 1.975 0.98 3.018 ;
      RECT 0.97 1.975 0.975 2.925 ;
      RECT 0.965 1.975 0.97 2.838 ;
      RECT 0.96 1.975 0.965 2.77 ;
      RECT 0.955 1.975 0.96 2.713 ;
      RECT 0.945 1.975 0.955 2.608 ;
      RECT 0.94 1.975 0.945 2.48 ;
      RECT 0.935 1.975 0.94 2.398 ;
      RECT 0.93 1.977 0.935 2.315 ;
      RECT 0.925 1.982 0.93 2.248 ;
      RECT 0.92 1.987 0.925 2.175 ;
      RECT 3.735 2.305 3.995 2.565 ;
      RECT 3.755 2.272 3.965 2.565 ;
      RECT 3.755 2.27 3.955 2.565 ;
      RECT 3.765 2.257 3.955 2.565 ;
      RECT 3.765 2.255 3.88 2.565 ;
      RECT 3.24 2.38 3.415 2.66 ;
      RECT 3.235 2.38 3.415 2.658 ;
      RECT 3.235 2.38 3.43 2.655 ;
      RECT 3.225 2.38 3.43 2.653 ;
      RECT 3.17 2.38 3.43 2.64 ;
      RECT 3.17 2.455 3.435 2.618 ;
      RECT 2.715 2.392 2.735 2.635 ;
      RECT 2.715 2.392 2.775 2.634 ;
      RECT 2.71 2.394 2.775 2.633 ;
      RECT 2.71 2.394 2.861 2.632 ;
      RECT 2.71 2.394 2.93 2.631 ;
      RECT 2.71 2.394 2.95 2.623 ;
      RECT 2.69 2.397 2.95 2.621 ;
      RECT 2.675 2.407 2.95 2.606 ;
      RECT 2.675 2.407 2.965 2.605 ;
      RECT 2.67 2.416 2.965 2.597 ;
      RECT 2.67 2.416 2.97 2.593 ;
      RECT 2.775 2.33 3.035 2.59 ;
      RECT 2.665 2.418 3.035 2.475 ;
      RECT 2.735 2.385 3.035 2.59 ;
      RECT 2.7 3.578 2.705 3.785 ;
      RECT 2.65 3.572 2.7 3.784 ;
      RECT 2.617 3.586 2.71 3.783 ;
      RECT 2.531 3.586 2.71 3.782 ;
      RECT 2.445 3.586 2.71 3.781 ;
      RECT 2.445 3.685 2.715 3.778 ;
      RECT 2.44 3.685 2.715 3.773 ;
      RECT 2.435 3.685 2.715 3.755 ;
      RECT 2.43 3.685 2.715 3.738 ;
      RECT 2.39 3.47 2.65 3.73 ;
      RECT 1.85 2.62 1.936 3.034 ;
      RECT 1.85 2.62 1.975 3.031 ;
      RECT 1.85 2.62 1.995 3.021 ;
      RECT 1.805 2.62 1.995 3.018 ;
      RECT 1.805 2.772 2.005 3.008 ;
      RECT 1.805 2.793 2.01 3.002 ;
      RECT 1.805 2.811 2.015 2.998 ;
      RECT 1.805 2.831 2.025 2.993 ;
      RECT 1.78 2.831 2.025 2.99 ;
      RECT 1.77 2.831 2.025 2.968 ;
      RECT 1.77 2.847 2.03 2.938 ;
      RECT 1.735 2.62 1.995 2.925 ;
      RECT 1.735 2.859 2.035 2.88 ;
      RECT -0.825 6.655 -0.535 6.885 ;
      RECT -0.995 6.685 -0.535 6.855 ;
      RECT -1.255 7.765 -0.965 7.995 ;
      RECT -1.195 7.025 -1.025 7.995 ;
      RECT -1.285 7.025 -0.935 7.315 ;
      RECT -1.66 6.285 -1.31 6.575 ;
      RECT -1.8 6.315 -1.31 6.485 ;
      RECT -2.625 5.915 -2.335 6.145 ;
      RECT -2.625 5.945 -2.165 6.115 ;
      RECT 65.36 3.265 65.62 3.525 ;
      RECT 50.1 3.265 50.36 3.525 ;
      RECT 34.84 3.265 35.1 3.525 ;
      RECT 19.58 3.265 19.84 3.525 ;
      RECT 4.32 3.265 4.58 3.525 ;
    LAYER mcon ;
      RECT 75.76 0.915 75.93 1.085 ;
      RECT 75.76 2.395 75.93 2.565 ;
      RECT 75.76 6.315 75.93 6.485 ;
      RECT 75.76 7.795 75.93 7.965 ;
      RECT 75.41 0.105 75.58 0.275 ;
      RECT 75.41 4.165 75.58 4.335 ;
      RECT 75.41 4.545 75.58 4.715 ;
      RECT 75.41 8.605 75.58 8.775 ;
      RECT 75.39 2.765 75.56 2.935 ;
      RECT 75.39 5.945 75.56 6.115 ;
      RECT 74.77 0.915 74.94 1.085 ;
      RECT 74.77 2.395 74.94 2.565 ;
      RECT 74.77 6.315 74.94 6.485 ;
      RECT 74.77 7.795 74.94 7.965 ;
      RECT 74.42 0.105 74.59 0.275 ;
      RECT 74.42 4.165 74.59 4.335 ;
      RECT 74.42 4.545 74.59 4.715 ;
      RECT 74.42 8.605 74.59 8.775 ;
      RECT 74.4 2.765 74.57 2.935 ;
      RECT 74.4 5.945 74.57 6.115 ;
      RECT 73.715 0.105 73.885 0.275 ;
      RECT 73.715 4.165 73.885 4.335 ;
      RECT 73.715 4.545 73.885 4.715 ;
      RECT 73.715 8.605 73.885 8.775 ;
      RECT 73.405 2.025 73.575 2.195 ;
      RECT 73.405 6.685 73.575 6.855 ;
      RECT 73.035 0.105 73.205 0.275 ;
      RECT 73.035 8.605 73.205 8.775 ;
      RECT 72.975 0.915 73.145 1.085 ;
      RECT 72.975 1.655 73.145 1.825 ;
      RECT 72.975 7.055 73.145 7.225 ;
      RECT 72.975 7.795 73.145 7.965 ;
      RECT 72.6 2.395 72.77 2.565 ;
      RECT 72.6 6.315 72.77 6.485 ;
      RECT 72.355 0.105 72.525 0.275 ;
      RECT 72.355 8.605 72.525 8.775 ;
      RECT 71.675 0.105 71.845 0.275 ;
      RECT 71.675 8.605 71.845 8.775 ;
      RECT 71.605 2.765 71.775 2.935 ;
      RECT 71.605 5.945 71.775 6.115 ;
      RECT 70.215 1.415 70.385 1.585 ;
      RECT 70.215 4.135 70.385 4.305 ;
      RECT 69.775 2.28 69.945 2.45 ;
      RECT 69.755 1.415 69.925 1.585 ;
      RECT 69.755 4.135 69.925 4.305 ;
      RECT 69.38 3.025 69.55 3.195 ;
      RECT 69.295 1.415 69.465 1.585 ;
      RECT 69.295 4.135 69.465 4.305 ;
      RECT 69.27 2.3 69.44 2.47 ;
      RECT 68.835 1.415 69.005 1.585 ;
      RECT 68.835 4.135 69.005 4.305 ;
      RECT 68.45 1.99 68.62 2.16 ;
      RECT 68.375 1.415 68.545 1.585 ;
      RECT 68.375 4.135 68.545 4.305 ;
      RECT 68.135 3.03 68.305 3.2 ;
      RECT 68.09 2.52 68.26 2.69 ;
      RECT 68.08 4.545 68.25 4.715 ;
      RECT 68.08 8.605 68.25 8.775 ;
      RECT 67.915 1.415 68.085 1.585 ;
      RECT 67.915 4.135 68.085 4.305 ;
      RECT 67.77 6.685 67.94 6.855 ;
      RECT 67.665 2.73 67.835 2.9 ;
      RECT 67.475 1.95 67.645 2.12 ;
      RECT 67.455 1.415 67.625 1.585 ;
      RECT 67.455 4.135 67.625 4.305 ;
      RECT 67.425 3.56 67.595 3.73 ;
      RECT 67.4 8.605 67.57 8.775 ;
      RECT 67.34 7.055 67.51 7.225 ;
      RECT 67.34 7.795 67.51 7.965 ;
      RECT 67.09 3 67.26 3.17 ;
      RECT 66.995 1.415 67.165 1.585 ;
      RECT 66.995 2.16 67.165 2.33 ;
      RECT 66.995 4.135 67.165 4.305 ;
      RECT 66.965 6.315 67.135 6.485 ;
      RECT 66.72 8.605 66.89 8.775 ;
      RECT 66.535 1.415 66.705 1.585 ;
      RECT 66.535 4.135 66.705 4.305 ;
      RECT 66.195 3.385 66.365 3.555 ;
      RECT 66.135 2.585 66.305 2.755 ;
      RECT 66.075 1.415 66.245 1.585 ;
      RECT 66.075 4.135 66.245 4.305 ;
      RECT 66.04 8.605 66.21 8.775 ;
      RECT 65.97 5.945 66.14 6.115 ;
      RECT 65.695 2.255 65.865 2.425 ;
      RECT 65.615 1.415 65.785 1.585 ;
      RECT 65.615 4.135 65.785 4.305 ;
      RECT 65.43 3.305 65.6 3.475 ;
      RECT 65.185 2.545 65.355 2.715 ;
      RECT 65.155 1.415 65.325 1.585 ;
      RECT 65.155 4.135 65.325 4.305 ;
      RECT 65.09 3.575 65.26 3.745 ;
      RECT 64.815 2.27 64.985 2.44 ;
      RECT 64.695 1.415 64.865 1.585 ;
      RECT 64.695 4.135 64.865 4.305 ;
      RECT 64.285 2.47 64.455 2.64 ;
      RECT 64.235 1.415 64.405 1.585 ;
      RECT 64.235 4.135 64.405 4.305 ;
      RECT 63.775 1.415 63.945 1.585 ;
      RECT 63.775 4.135 63.945 4.305 ;
      RECT 63.765 2.415 63.935 2.585 ;
      RECT 63.56 2.015 63.73 2.185 ;
      RECT 63.56 3.595 63.73 3.765 ;
      RECT 63.315 1.415 63.485 1.585 ;
      RECT 63.315 4.135 63.485 4.305 ;
      RECT 63.25 2.56 63.42 2.73 ;
      RECT 62.855 1.415 63.025 1.585 ;
      RECT 62.855 4.135 63.025 4.305 ;
      RECT 62.84 2.785 63.01 2.955 ;
      RECT 62.395 1.415 62.565 1.585 ;
      RECT 62.395 4.135 62.565 4.305 ;
      RECT 62.13 3.085 62.3 3.255 ;
      RECT 61.985 1.995 62.155 2.165 ;
      RECT 61.935 1.415 62.105 1.585 ;
      RECT 61.935 4.135 62.105 4.305 ;
      RECT 60.5 0.915 60.67 1.085 ;
      RECT 60.5 2.395 60.67 2.565 ;
      RECT 60.5 6.315 60.67 6.485 ;
      RECT 60.5 7.795 60.67 7.965 ;
      RECT 60.15 0.105 60.32 0.275 ;
      RECT 60.15 4.165 60.32 4.335 ;
      RECT 60.15 4.545 60.32 4.715 ;
      RECT 60.15 8.605 60.32 8.775 ;
      RECT 60.13 2.765 60.3 2.935 ;
      RECT 60.13 5.945 60.3 6.115 ;
      RECT 59.51 0.915 59.68 1.085 ;
      RECT 59.51 2.395 59.68 2.565 ;
      RECT 59.51 6.315 59.68 6.485 ;
      RECT 59.51 7.795 59.68 7.965 ;
      RECT 59.16 0.105 59.33 0.275 ;
      RECT 59.16 4.165 59.33 4.335 ;
      RECT 59.16 4.545 59.33 4.715 ;
      RECT 59.16 8.605 59.33 8.775 ;
      RECT 59.14 2.765 59.31 2.935 ;
      RECT 59.14 5.945 59.31 6.115 ;
      RECT 58.455 0.105 58.625 0.275 ;
      RECT 58.455 4.165 58.625 4.335 ;
      RECT 58.455 4.545 58.625 4.715 ;
      RECT 58.455 8.605 58.625 8.775 ;
      RECT 58.145 2.025 58.315 2.195 ;
      RECT 58.145 6.685 58.315 6.855 ;
      RECT 57.775 0.105 57.945 0.275 ;
      RECT 57.775 8.605 57.945 8.775 ;
      RECT 57.715 0.915 57.885 1.085 ;
      RECT 57.715 1.655 57.885 1.825 ;
      RECT 57.715 7.055 57.885 7.225 ;
      RECT 57.715 7.795 57.885 7.965 ;
      RECT 57.34 2.395 57.51 2.565 ;
      RECT 57.34 6.315 57.51 6.485 ;
      RECT 57.095 0.105 57.265 0.275 ;
      RECT 57.095 8.605 57.265 8.775 ;
      RECT 56.415 0.105 56.585 0.275 ;
      RECT 56.415 8.605 56.585 8.775 ;
      RECT 56.345 2.765 56.515 2.935 ;
      RECT 56.345 5.945 56.515 6.115 ;
      RECT 54.955 1.415 55.125 1.585 ;
      RECT 54.955 4.135 55.125 4.305 ;
      RECT 54.515 2.28 54.685 2.45 ;
      RECT 54.495 1.415 54.665 1.585 ;
      RECT 54.495 4.135 54.665 4.305 ;
      RECT 54.12 3.025 54.29 3.195 ;
      RECT 54.035 1.415 54.205 1.585 ;
      RECT 54.035 4.135 54.205 4.305 ;
      RECT 54.01 2.3 54.18 2.47 ;
      RECT 53.575 1.415 53.745 1.585 ;
      RECT 53.575 4.135 53.745 4.305 ;
      RECT 53.19 1.99 53.36 2.16 ;
      RECT 53.115 1.415 53.285 1.585 ;
      RECT 53.115 4.135 53.285 4.305 ;
      RECT 52.875 3.03 53.045 3.2 ;
      RECT 52.83 2.52 53 2.69 ;
      RECT 52.82 4.545 52.99 4.715 ;
      RECT 52.82 8.605 52.99 8.775 ;
      RECT 52.655 1.415 52.825 1.585 ;
      RECT 52.655 4.135 52.825 4.305 ;
      RECT 52.51 6.685 52.68 6.855 ;
      RECT 52.405 2.73 52.575 2.9 ;
      RECT 52.215 1.95 52.385 2.12 ;
      RECT 52.195 1.415 52.365 1.585 ;
      RECT 52.195 4.135 52.365 4.305 ;
      RECT 52.165 3.56 52.335 3.73 ;
      RECT 52.14 8.605 52.31 8.775 ;
      RECT 52.08 7.055 52.25 7.225 ;
      RECT 52.08 7.795 52.25 7.965 ;
      RECT 51.83 3 52 3.17 ;
      RECT 51.735 1.415 51.905 1.585 ;
      RECT 51.735 2.16 51.905 2.33 ;
      RECT 51.735 4.135 51.905 4.305 ;
      RECT 51.705 6.315 51.875 6.485 ;
      RECT 51.46 8.605 51.63 8.775 ;
      RECT 51.275 1.415 51.445 1.585 ;
      RECT 51.275 4.135 51.445 4.305 ;
      RECT 50.935 3.385 51.105 3.555 ;
      RECT 50.875 2.585 51.045 2.755 ;
      RECT 50.815 1.415 50.985 1.585 ;
      RECT 50.815 4.135 50.985 4.305 ;
      RECT 50.78 8.605 50.95 8.775 ;
      RECT 50.71 5.945 50.88 6.115 ;
      RECT 50.435 2.255 50.605 2.425 ;
      RECT 50.355 1.415 50.525 1.585 ;
      RECT 50.355 4.135 50.525 4.305 ;
      RECT 50.17 3.305 50.34 3.475 ;
      RECT 49.925 2.545 50.095 2.715 ;
      RECT 49.895 1.415 50.065 1.585 ;
      RECT 49.895 4.135 50.065 4.305 ;
      RECT 49.83 3.575 50 3.745 ;
      RECT 49.555 2.27 49.725 2.44 ;
      RECT 49.435 1.415 49.605 1.585 ;
      RECT 49.435 4.135 49.605 4.305 ;
      RECT 49.025 2.47 49.195 2.64 ;
      RECT 48.975 1.415 49.145 1.585 ;
      RECT 48.975 4.135 49.145 4.305 ;
      RECT 48.515 1.415 48.685 1.585 ;
      RECT 48.515 4.135 48.685 4.305 ;
      RECT 48.505 2.415 48.675 2.585 ;
      RECT 48.3 2.015 48.47 2.185 ;
      RECT 48.3 3.595 48.47 3.765 ;
      RECT 48.055 1.415 48.225 1.585 ;
      RECT 48.055 4.135 48.225 4.305 ;
      RECT 47.99 2.56 48.16 2.73 ;
      RECT 47.595 1.415 47.765 1.585 ;
      RECT 47.595 4.135 47.765 4.305 ;
      RECT 47.58 2.785 47.75 2.955 ;
      RECT 47.135 1.415 47.305 1.585 ;
      RECT 47.135 4.135 47.305 4.305 ;
      RECT 46.87 3.085 47.04 3.255 ;
      RECT 46.725 1.995 46.895 2.165 ;
      RECT 46.675 1.415 46.845 1.585 ;
      RECT 46.675 4.135 46.845 4.305 ;
      RECT 45.24 0.915 45.41 1.085 ;
      RECT 45.24 2.395 45.41 2.565 ;
      RECT 45.24 6.315 45.41 6.485 ;
      RECT 45.24 7.795 45.41 7.965 ;
      RECT 44.89 0.105 45.06 0.275 ;
      RECT 44.89 4.165 45.06 4.335 ;
      RECT 44.89 4.545 45.06 4.715 ;
      RECT 44.89 8.605 45.06 8.775 ;
      RECT 44.87 2.765 45.04 2.935 ;
      RECT 44.87 5.945 45.04 6.115 ;
      RECT 44.25 0.915 44.42 1.085 ;
      RECT 44.25 2.395 44.42 2.565 ;
      RECT 44.25 6.315 44.42 6.485 ;
      RECT 44.25 7.795 44.42 7.965 ;
      RECT 43.9 0.105 44.07 0.275 ;
      RECT 43.9 4.165 44.07 4.335 ;
      RECT 43.9 4.545 44.07 4.715 ;
      RECT 43.9 8.605 44.07 8.775 ;
      RECT 43.88 2.765 44.05 2.935 ;
      RECT 43.88 5.945 44.05 6.115 ;
      RECT 43.195 0.105 43.365 0.275 ;
      RECT 43.195 4.165 43.365 4.335 ;
      RECT 43.195 4.545 43.365 4.715 ;
      RECT 43.195 8.605 43.365 8.775 ;
      RECT 42.885 2.025 43.055 2.195 ;
      RECT 42.885 6.685 43.055 6.855 ;
      RECT 42.515 0.105 42.685 0.275 ;
      RECT 42.515 8.605 42.685 8.775 ;
      RECT 42.455 0.915 42.625 1.085 ;
      RECT 42.455 1.655 42.625 1.825 ;
      RECT 42.455 7.055 42.625 7.225 ;
      RECT 42.455 7.795 42.625 7.965 ;
      RECT 42.08 2.395 42.25 2.565 ;
      RECT 42.08 6.315 42.25 6.485 ;
      RECT 41.835 0.105 42.005 0.275 ;
      RECT 41.835 8.605 42.005 8.775 ;
      RECT 41.155 0.105 41.325 0.275 ;
      RECT 41.155 8.605 41.325 8.775 ;
      RECT 41.085 2.765 41.255 2.935 ;
      RECT 41.085 5.945 41.255 6.115 ;
      RECT 39.695 1.415 39.865 1.585 ;
      RECT 39.695 4.135 39.865 4.305 ;
      RECT 39.255 2.28 39.425 2.45 ;
      RECT 39.235 1.415 39.405 1.585 ;
      RECT 39.235 4.135 39.405 4.305 ;
      RECT 38.86 3.025 39.03 3.195 ;
      RECT 38.775 1.415 38.945 1.585 ;
      RECT 38.775 4.135 38.945 4.305 ;
      RECT 38.75 2.3 38.92 2.47 ;
      RECT 38.315 1.415 38.485 1.585 ;
      RECT 38.315 4.135 38.485 4.305 ;
      RECT 37.93 1.99 38.1 2.16 ;
      RECT 37.855 1.415 38.025 1.585 ;
      RECT 37.855 4.135 38.025 4.305 ;
      RECT 37.615 3.03 37.785 3.2 ;
      RECT 37.57 2.52 37.74 2.69 ;
      RECT 37.56 4.545 37.73 4.715 ;
      RECT 37.56 8.605 37.73 8.775 ;
      RECT 37.395 1.415 37.565 1.585 ;
      RECT 37.395 4.135 37.565 4.305 ;
      RECT 37.25 6.685 37.42 6.855 ;
      RECT 37.145 2.73 37.315 2.9 ;
      RECT 36.955 1.95 37.125 2.12 ;
      RECT 36.935 1.415 37.105 1.585 ;
      RECT 36.935 4.135 37.105 4.305 ;
      RECT 36.905 3.56 37.075 3.73 ;
      RECT 36.88 8.605 37.05 8.775 ;
      RECT 36.82 7.055 36.99 7.225 ;
      RECT 36.82 7.795 36.99 7.965 ;
      RECT 36.57 3 36.74 3.17 ;
      RECT 36.475 1.415 36.645 1.585 ;
      RECT 36.475 2.16 36.645 2.33 ;
      RECT 36.475 4.135 36.645 4.305 ;
      RECT 36.445 6.315 36.615 6.485 ;
      RECT 36.2 8.605 36.37 8.775 ;
      RECT 36.015 1.415 36.185 1.585 ;
      RECT 36.015 4.135 36.185 4.305 ;
      RECT 35.675 3.385 35.845 3.555 ;
      RECT 35.615 2.585 35.785 2.755 ;
      RECT 35.555 1.415 35.725 1.585 ;
      RECT 35.555 4.135 35.725 4.305 ;
      RECT 35.52 8.605 35.69 8.775 ;
      RECT 35.45 5.945 35.62 6.115 ;
      RECT 35.175 2.255 35.345 2.425 ;
      RECT 35.095 1.415 35.265 1.585 ;
      RECT 35.095 4.135 35.265 4.305 ;
      RECT 34.91 3.305 35.08 3.475 ;
      RECT 34.665 2.545 34.835 2.715 ;
      RECT 34.635 1.415 34.805 1.585 ;
      RECT 34.635 4.135 34.805 4.305 ;
      RECT 34.57 3.575 34.74 3.745 ;
      RECT 34.295 2.27 34.465 2.44 ;
      RECT 34.175 1.415 34.345 1.585 ;
      RECT 34.175 4.135 34.345 4.305 ;
      RECT 33.765 2.47 33.935 2.64 ;
      RECT 33.715 1.415 33.885 1.585 ;
      RECT 33.715 4.135 33.885 4.305 ;
      RECT 33.255 1.415 33.425 1.585 ;
      RECT 33.255 4.135 33.425 4.305 ;
      RECT 33.245 2.415 33.415 2.585 ;
      RECT 33.04 2.015 33.21 2.185 ;
      RECT 33.04 3.595 33.21 3.765 ;
      RECT 32.795 1.415 32.965 1.585 ;
      RECT 32.795 4.135 32.965 4.305 ;
      RECT 32.73 2.56 32.9 2.73 ;
      RECT 32.335 1.415 32.505 1.585 ;
      RECT 32.335 4.135 32.505 4.305 ;
      RECT 32.32 2.785 32.49 2.955 ;
      RECT 31.875 1.415 32.045 1.585 ;
      RECT 31.875 4.135 32.045 4.305 ;
      RECT 31.61 3.085 31.78 3.255 ;
      RECT 31.465 1.995 31.635 2.165 ;
      RECT 31.415 1.415 31.585 1.585 ;
      RECT 31.415 4.135 31.585 4.305 ;
      RECT 29.98 0.915 30.15 1.085 ;
      RECT 29.98 2.395 30.15 2.565 ;
      RECT 29.98 6.315 30.15 6.485 ;
      RECT 29.98 7.795 30.15 7.965 ;
      RECT 29.63 0.105 29.8 0.275 ;
      RECT 29.63 4.165 29.8 4.335 ;
      RECT 29.63 4.545 29.8 4.715 ;
      RECT 29.63 8.605 29.8 8.775 ;
      RECT 29.61 2.765 29.78 2.935 ;
      RECT 29.61 5.945 29.78 6.115 ;
      RECT 28.99 0.915 29.16 1.085 ;
      RECT 28.99 2.395 29.16 2.565 ;
      RECT 28.99 6.315 29.16 6.485 ;
      RECT 28.99 7.795 29.16 7.965 ;
      RECT 28.64 0.105 28.81 0.275 ;
      RECT 28.64 4.165 28.81 4.335 ;
      RECT 28.64 4.545 28.81 4.715 ;
      RECT 28.64 8.605 28.81 8.775 ;
      RECT 28.62 2.765 28.79 2.935 ;
      RECT 28.62 5.945 28.79 6.115 ;
      RECT 27.935 0.105 28.105 0.275 ;
      RECT 27.935 4.165 28.105 4.335 ;
      RECT 27.935 4.545 28.105 4.715 ;
      RECT 27.935 8.605 28.105 8.775 ;
      RECT 27.625 2.025 27.795 2.195 ;
      RECT 27.625 6.685 27.795 6.855 ;
      RECT 27.255 0.105 27.425 0.275 ;
      RECT 27.255 8.605 27.425 8.775 ;
      RECT 27.195 0.915 27.365 1.085 ;
      RECT 27.195 1.655 27.365 1.825 ;
      RECT 27.195 7.055 27.365 7.225 ;
      RECT 27.195 7.795 27.365 7.965 ;
      RECT 26.82 2.395 26.99 2.565 ;
      RECT 26.82 6.315 26.99 6.485 ;
      RECT 26.575 0.105 26.745 0.275 ;
      RECT 26.575 8.605 26.745 8.775 ;
      RECT 25.895 0.105 26.065 0.275 ;
      RECT 25.895 8.605 26.065 8.775 ;
      RECT 25.825 2.765 25.995 2.935 ;
      RECT 25.825 5.945 25.995 6.115 ;
      RECT 24.435 1.415 24.605 1.585 ;
      RECT 24.435 4.135 24.605 4.305 ;
      RECT 23.995 2.28 24.165 2.45 ;
      RECT 23.975 1.415 24.145 1.585 ;
      RECT 23.975 4.135 24.145 4.305 ;
      RECT 23.6 3.025 23.77 3.195 ;
      RECT 23.515 1.415 23.685 1.585 ;
      RECT 23.515 4.135 23.685 4.305 ;
      RECT 23.49 2.3 23.66 2.47 ;
      RECT 23.055 1.415 23.225 1.585 ;
      RECT 23.055 4.135 23.225 4.305 ;
      RECT 22.67 1.99 22.84 2.16 ;
      RECT 22.595 1.415 22.765 1.585 ;
      RECT 22.595 4.135 22.765 4.305 ;
      RECT 22.355 3.03 22.525 3.2 ;
      RECT 22.31 2.52 22.48 2.69 ;
      RECT 22.3 4.545 22.47 4.715 ;
      RECT 22.3 8.605 22.47 8.775 ;
      RECT 22.135 1.415 22.305 1.585 ;
      RECT 22.135 4.135 22.305 4.305 ;
      RECT 21.99 6.685 22.16 6.855 ;
      RECT 21.885 2.73 22.055 2.9 ;
      RECT 21.695 1.95 21.865 2.12 ;
      RECT 21.675 1.415 21.845 1.585 ;
      RECT 21.675 4.135 21.845 4.305 ;
      RECT 21.645 3.56 21.815 3.73 ;
      RECT 21.62 8.605 21.79 8.775 ;
      RECT 21.56 7.055 21.73 7.225 ;
      RECT 21.56 7.795 21.73 7.965 ;
      RECT 21.31 3 21.48 3.17 ;
      RECT 21.215 1.415 21.385 1.585 ;
      RECT 21.215 2.16 21.385 2.33 ;
      RECT 21.215 4.135 21.385 4.305 ;
      RECT 21.185 6.315 21.355 6.485 ;
      RECT 20.94 8.605 21.11 8.775 ;
      RECT 20.755 1.415 20.925 1.585 ;
      RECT 20.755 4.135 20.925 4.305 ;
      RECT 20.415 3.385 20.585 3.555 ;
      RECT 20.355 2.585 20.525 2.755 ;
      RECT 20.295 1.415 20.465 1.585 ;
      RECT 20.295 4.135 20.465 4.305 ;
      RECT 20.26 8.605 20.43 8.775 ;
      RECT 20.19 5.945 20.36 6.115 ;
      RECT 19.915 2.255 20.085 2.425 ;
      RECT 19.835 1.415 20.005 1.585 ;
      RECT 19.835 4.135 20.005 4.305 ;
      RECT 19.65 3.305 19.82 3.475 ;
      RECT 19.405 2.545 19.575 2.715 ;
      RECT 19.375 1.415 19.545 1.585 ;
      RECT 19.375 4.135 19.545 4.305 ;
      RECT 19.31 3.575 19.48 3.745 ;
      RECT 19.035 2.27 19.205 2.44 ;
      RECT 18.915 1.415 19.085 1.585 ;
      RECT 18.915 4.135 19.085 4.305 ;
      RECT 18.505 2.47 18.675 2.64 ;
      RECT 18.455 1.415 18.625 1.585 ;
      RECT 18.455 4.135 18.625 4.305 ;
      RECT 17.995 1.415 18.165 1.585 ;
      RECT 17.995 4.135 18.165 4.305 ;
      RECT 17.985 2.415 18.155 2.585 ;
      RECT 17.78 2.015 17.95 2.185 ;
      RECT 17.78 3.595 17.95 3.765 ;
      RECT 17.535 1.415 17.705 1.585 ;
      RECT 17.535 4.135 17.705 4.305 ;
      RECT 17.47 2.56 17.64 2.73 ;
      RECT 17.075 1.415 17.245 1.585 ;
      RECT 17.075 4.135 17.245 4.305 ;
      RECT 17.06 2.785 17.23 2.955 ;
      RECT 16.615 1.415 16.785 1.585 ;
      RECT 16.615 4.135 16.785 4.305 ;
      RECT 16.35 3.085 16.52 3.255 ;
      RECT 16.205 1.995 16.375 2.165 ;
      RECT 16.155 1.415 16.325 1.585 ;
      RECT 16.155 4.135 16.325 4.305 ;
      RECT 14.72 0.915 14.89 1.085 ;
      RECT 14.72 2.395 14.89 2.565 ;
      RECT 14.72 6.315 14.89 6.485 ;
      RECT 14.72 7.795 14.89 7.965 ;
      RECT 14.37 0.105 14.54 0.275 ;
      RECT 14.37 4.165 14.54 4.335 ;
      RECT 14.37 4.545 14.54 4.715 ;
      RECT 14.37 8.605 14.54 8.775 ;
      RECT 14.35 2.765 14.52 2.935 ;
      RECT 14.35 5.945 14.52 6.115 ;
      RECT 13.73 0.915 13.9 1.085 ;
      RECT 13.73 2.395 13.9 2.565 ;
      RECT 13.73 6.315 13.9 6.485 ;
      RECT 13.73 7.795 13.9 7.965 ;
      RECT 13.38 0.105 13.55 0.275 ;
      RECT 13.38 4.165 13.55 4.335 ;
      RECT 13.38 4.545 13.55 4.715 ;
      RECT 13.38 8.605 13.55 8.775 ;
      RECT 13.36 2.765 13.53 2.935 ;
      RECT 13.36 5.945 13.53 6.115 ;
      RECT 12.675 0.105 12.845 0.275 ;
      RECT 12.675 4.165 12.845 4.335 ;
      RECT 12.675 4.545 12.845 4.715 ;
      RECT 12.675 8.605 12.845 8.775 ;
      RECT 12.365 2.025 12.535 2.195 ;
      RECT 12.365 6.685 12.535 6.855 ;
      RECT 11.995 0.105 12.165 0.275 ;
      RECT 11.995 8.605 12.165 8.775 ;
      RECT 11.935 0.915 12.105 1.085 ;
      RECT 11.935 1.655 12.105 1.825 ;
      RECT 11.935 7.055 12.105 7.225 ;
      RECT 11.935 7.795 12.105 7.965 ;
      RECT 11.56 2.395 11.73 2.565 ;
      RECT 11.56 6.315 11.73 6.485 ;
      RECT 11.315 0.105 11.485 0.275 ;
      RECT 11.315 8.605 11.485 8.775 ;
      RECT 10.635 0.105 10.805 0.275 ;
      RECT 10.635 8.605 10.805 8.775 ;
      RECT 10.565 2.765 10.735 2.935 ;
      RECT 10.565 5.945 10.735 6.115 ;
      RECT 9.175 1.415 9.345 1.585 ;
      RECT 9.175 4.135 9.345 4.305 ;
      RECT 8.735 2.28 8.905 2.45 ;
      RECT 8.715 1.415 8.885 1.585 ;
      RECT 8.715 4.135 8.885 4.305 ;
      RECT 8.34 3.025 8.51 3.195 ;
      RECT 8.255 1.415 8.425 1.585 ;
      RECT 8.255 4.135 8.425 4.305 ;
      RECT 8.23 2.3 8.4 2.47 ;
      RECT 7.795 1.415 7.965 1.585 ;
      RECT 7.795 4.135 7.965 4.305 ;
      RECT 7.41 1.99 7.58 2.16 ;
      RECT 7.335 1.415 7.505 1.585 ;
      RECT 7.335 4.135 7.505 4.305 ;
      RECT 7.095 3.03 7.265 3.2 ;
      RECT 7.05 2.52 7.22 2.69 ;
      RECT 7.04 4.545 7.21 4.715 ;
      RECT 7.04 8.605 7.21 8.775 ;
      RECT 6.875 1.415 7.045 1.585 ;
      RECT 6.875 4.135 7.045 4.305 ;
      RECT 6.73 6.685 6.9 6.855 ;
      RECT 6.625 2.73 6.795 2.9 ;
      RECT 6.435 1.95 6.605 2.12 ;
      RECT 6.415 1.415 6.585 1.585 ;
      RECT 6.415 4.135 6.585 4.305 ;
      RECT 6.385 3.56 6.555 3.73 ;
      RECT 6.36 8.605 6.53 8.775 ;
      RECT 6.3 7.055 6.47 7.225 ;
      RECT 6.3 7.795 6.47 7.965 ;
      RECT 6.05 3 6.22 3.17 ;
      RECT 5.955 1.415 6.125 1.585 ;
      RECT 5.955 2.16 6.125 2.33 ;
      RECT 5.955 4.135 6.125 4.305 ;
      RECT 5.925 6.315 6.095 6.485 ;
      RECT 5.68 8.605 5.85 8.775 ;
      RECT 5.495 1.415 5.665 1.585 ;
      RECT 5.495 4.135 5.665 4.305 ;
      RECT 5.155 3.385 5.325 3.555 ;
      RECT 5.095 2.585 5.265 2.755 ;
      RECT 5.035 1.415 5.205 1.585 ;
      RECT 5.035 4.135 5.205 4.305 ;
      RECT 5 8.605 5.17 8.775 ;
      RECT 4.93 5.945 5.1 6.115 ;
      RECT 4.655 2.255 4.825 2.425 ;
      RECT 4.575 1.415 4.745 1.585 ;
      RECT 4.575 4.135 4.745 4.305 ;
      RECT 4.39 3.305 4.56 3.475 ;
      RECT 4.145 2.545 4.315 2.715 ;
      RECT 4.115 1.415 4.285 1.585 ;
      RECT 4.115 4.135 4.285 4.305 ;
      RECT 4.05 3.575 4.22 3.745 ;
      RECT 3.775 2.27 3.945 2.44 ;
      RECT 3.655 1.415 3.825 1.585 ;
      RECT 3.655 4.135 3.825 4.305 ;
      RECT 3.245 2.47 3.415 2.64 ;
      RECT 3.195 1.415 3.365 1.585 ;
      RECT 3.195 4.135 3.365 4.305 ;
      RECT 2.735 1.415 2.905 1.585 ;
      RECT 2.735 4.135 2.905 4.305 ;
      RECT 2.725 2.415 2.895 2.585 ;
      RECT 2.52 2.015 2.69 2.185 ;
      RECT 2.52 3.595 2.69 3.765 ;
      RECT 2.275 1.415 2.445 1.585 ;
      RECT 2.275 4.135 2.445 4.305 ;
      RECT 2.21 2.56 2.38 2.73 ;
      RECT 1.815 1.415 1.985 1.585 ;
      RECT 1.815 4.135 1.985 4.305 ;
      RECT 1.8 2.785 1.97 2.955 ;
      RECT 1.355 1.415 1.525 1.585 ;
      RECT 1.355 4.135 1.525 4.305 ;
      RECT 1.09 3.085 1.26 3.255 ;
      RECT 0.945 1.995 1.115 2.165 ;
      RECT 0.895 1.415 1.065 1.585 ;
      RECT 0.895 4.135 1.065 4.305 ;
      RECT -0.455 4.545 -0.285 4.715 ;
      RECT -0.455 8.605 -0.285 8.775 ;
      RECT -0.765 6.685 -0.595 6.855 ;
      RECT -1.135 8.605 -0.965 8.775 ;
      RECT -1.195 7.055 -1.025 7.225 ;
      RECT -1.195 7.795 -1.025 7.965 ;
      RECT -1.57 6.315 -1.4 6.485 ;
      RECT -1.815 8.605 -1.645 8.775 ;
      RECT -2.495 8.605 -2.325 8.775 ;
      RECT -2.565 5.945 -2.395 6.115 ;
    LAYER li ;
      RECT 69.76 0 69.93 2.085 ;
      RECT 68.82 0 68.99 2.085 ;
      RECT 67.86 0 68.03 2.085 ;
      RECT 65.94 0 66.11 2.085 ;
      RECT 64.98 0 65.15 2.085 ;
      RECT 63.06 0 63.23 2.085 ;
      RECT 54.5 0 54.67 2.085 ;
      RECT 53.56 0 53.73 2.085 ;
      RECT 52.6 0 52.77 2.085 ;
      RECT 50.68 0 50.85 2.085 ;
      RECT 49.72 0 49.89 2.085 ;
      RECT 47.8 0 47.97 2.085 ;
      RECT 39.24 0 39.41 2.085 ;
      RECT 38.3 0 38.47 2.085 ;
      RECT 37.34 0 37.51 2.085 ;
      RECT 35.42 0 35.59 2.085 ;
      RECT 34.46 0 34.63 2.085 ;
      RECT 32.54 0 32.71 2.085 ;
      RECT 23.98 0 24.15 2.085 ;
      RECT 23.04 0 23.21 2.085 ;
      RECT 22.08 0 22.25 2.085 ;
      RECT 20.16 0 20.33 2.085 ;
      RECT 19.2 0 19.37 2.085 ;
      RECT 17.28 0 17.45 2.085 ;
      RECT 8.72 0 8.89 2.085 ;
      RECT 7.78 0 7.95 2.085 ;
      RECT 6.82 0 6.99 2.085 ;
      RECT 4.9 0 5.07 2.085 ;
      RECT 3.94 0 4.11 2.085 ;
      RECT 2.02 0 2.19 2.085 ;
      RECT 66.815 0 67.01 1.595 ;
      RECT 63.06 0 63.335 1.595 ;
      RECT 51.555 0 51.75 1.595 ;
      RECT 47.8 0 48.075 1.595 ;
      RECT 36.295 0 36.49 1.595 ;
      RECT 32.54 0 32.815 1.595 ;
      RECT 21.035 0 21.23 1.595 ;
      RECT 17.28 0 17.555 1.595 ;
      RECT 5.775 0 5.97 1.595 ;
      RECT 2.02 0 2.295 1.595 ;
      RECT 61.79 0 70.53 1.585 ;
      RECT 46.53 0 55.27 1.585 ;
      RECT 31.27 0 40.01 1.585 ;
      RECT 16.01 0 24.75 1.585 ;
      RECT 0.75 0 9.49 1.585 ;
      RECT 75.33 0 75.5 0.935 ;
      RECT 74.34 0 74.51 0.935 ;
      RECT 71.595 0 71.765 0.935 ;
      RECT 60.07 0 60.24 0.935 ;
      RECT 59.08 0 59.25 0.935 ;
      RECT 56.335 0 56.505 0.935 ;
      RECT 44.81 0 44.98 0.935 ;
      RECT 43.82 0 43.99 0.935 ;
      RECT 41.075 0 41.245 0.935 ;
      RECT 29.55 0 29.72 0.935 ;
      RECT 28.56 0 28.73 0.935 ;
      RECT 25.815 0 25.985 0.935 ;
      RECT 14.29 0 14.46 0.935 ;
      RECT 13.3 0 13.47 0.935 ;
      RECT 10.555 0 10.725 0.935 ;
      RECT -2.75 0 76.3 0.305 ;
      RECT -0.765 4.14 -0.595 8.305 ;
      RECT 75.33 3.405 75.5 5.475 ;
      RECT 74.34 3.405 74.51 5.475 ;
      RECT 71.595 3.405 71.765 5.475 ;
      RECT 65.96 3.635 66.13 5.475 ;
      RECT 60.07 3.405 60.24 5.475 ;
      RECT 59.08 3.405 59.25 5.475 ;
      RECT 56.335 3.405 56.505 5.475 ;
      RECT 50.7 3.635 50.87 5.475 ;
      RECT 44.81 3.405 44.98 5.475 ;
      RECT 43.82 3.405 43.99 5.475 ;
      RECT 41.075 3.405 41.245 5.475 ;
      RECT 35.44 3.635 35.61 5.475 ;
      RECT 29.55 3.405 29.72 5.475 ;
      RECT 28.56 3.405 28.73 5.475 ;
      RECT 25.815 3.405 25.985 5.475 ;
      RECT 20.18 3.635 20.35 5.475 ;
      RECT 14.29 3.405 14.46 5.475 ;
      RECT 13.3 3.405 13.47 5.475 ;
      RECT 10.555 3.405 10.725 5.475 ;
      RECT 4.92 3.635 5.09 5.475 ;
      RECT -2.575 4.14 -2.405 5.475 ;
      RECT -2.75 4.14 76.3 4.745 ;
      RECT 61.79 4.135 76.3 4.745 ;
      RECT 46.53 4.135 61.04 4.745 ;
      RECT 31.27 4.135 45.78 4.745 ;
      RECT 16.01 4.135 30.52 4.745 ;
      RECT 0.75 4.135 15.26 4.745 ;
      RECT 68.82 3.635 68.99 4.745 ;
      RECT 66.9 3.635 67.07 4.745 ;
      RECT 64.5 3.635 64.67 4.745 ;
      RECT 62.58 3.635 62.75 4.745 ;
      RECT 53.56 3.635 53.73 4.745 ;
      RECT 51.64 3.635 51.81 4.745 ;
      RECT 49.24 3.635 49.41 4.745 ;
      RECT 47.32 3.635 47.49 4.745 ;
      RECT 38.3 3.635 38.47 4.745 ;
      RECT 36.38 3.635 36.55 4.745 ;
      RECT 33.98 3.635 34.15 4.745 ;
      RECT 32.06 3.635 32.23 4.745 ;
      RECT 23.04 3.635 23.21 4.745 ;
      RECT 21.12 3.635 21.29 4.745 ;
      RECT 18.72 3.635 18.89 4.745 ;
      RECT 16.8 3.635 16.97 4.745 ;
      RECT 7.78 3.635 7.95 4.745 ;
      RECT 5.86 3.635 6.03 4.745 ;
      RECT 3.46 3.635 3.63 4.745 ;
      RECT 1.54 3.635 1.71 4.745 ;
      RECT -2.75 8.575 76.3 8.88 ;
      RECT 75.33 7.945 75.5 8.88 ;
      RECT 74.34 7.945 74.51 8.88 ;
      RECT 71.595 7.945 71.765 8.88 ;
      RECT 65.96 7.945 66.13 8.88 ;
      RECT 60.07 7.945 60.24 8.88 ;
      RECT 59.08 7.945 59.25 8.88 ;
      RECT 56.335 7.945 56.505 8.88 ;
      RECT 50.7 7.945 50.87 8.88 ;
      RECT 44.81 7.945 44.98 8.88 ;
      RECT 43.82 7.945 43.99 8.88 ;
      RECT 41.075 7.945 41.245 8.88 ;
      RECT 35.44 7.945 35.61 8.88 ;
      RECT 29.55 7.945 29.72 8.88 ;
      RECT 28.56 7.945 28.73 8.88 ;
      RECT 25.815 7.945 25.985 8.88 ;
      RECT 20.18 7.945 20.35 8.88 ;
      RECT 14.29 7.945 14.46 8.88 ;
      RECT 13.3 7.945 13.47 8.88 ;
      RECT 10.555 7.945 10.725 8.88 ;
      RECT 4.92 7.945 5.09 8.88 ;
      RECT -2.575 7.945 -2.405 8.88 ;
      RECT 75.39 1.74 75.56 2.935 ;
      RECT 75.39 1.74 75.855 1.91 ;
      RECT 75.39 6.97 75.855 7.14 ;
      RECT 75.39 5.945 75.56 7.14 ;
      RECT 74.4 1.74 74.57 2.935 ;
      RECT 74.4 1.74 74.865 1.91 ;
      RECT 74.4 6.97 74.865 7.14 ;
      RECT 74.4 5.945 74.57 7.14 ;
      RECT 72.545 2.635 72.715 3.865 ;
      RECT 72.6 0.855 72.77 2.805 ;
      RECT 72.545 0.575 72.715 1.025 ;
      RECT 72.545 7.855 72.715 8.305 ;
      RECT 72.6 6.075 72.77 8.025 ;
      RECT 72.545 5.015 72.715 6.245 ;
      RECT 72.025 0.575 72.195 3.865 ;
      RECT 72.025 2.075 72.43 2.405 ;
      RECT 72.025 1.235 72.43 1.565 ;
      RECT 72.025 5.015 72.195 8.305 ;
      RECT 72.025 7.315 72.43 7.645 ;
      RECT 72.025 6.475 72.43 6.805 ;
      RECT 69.95 3.126 69.955 3.298 ;
      RECT 69.945 3.119 69.95 3.388 ;
      RECT 69.94 3.113 69.945 3.407 ;
      RECT 69.92 3.107 69.94 3.417 ;
      RECT 69.905 3.102 69.92 3.425 ;
      RECT 69.868 3.096 69.905 3.423 ;
      RECT 69.782 3.082 69.868 3.419 ;
      RECT 69.696 3.064 69.782 3.414 ;
      RECT 69.61 3.045 69.696 3.408 ;
      RECT 69.58 3.033 69.61 3.404 ;
      RECT 69.56 3.027 69.58 3.403 ;
      RECT 69.495 3.025 69.56 3.401 ;
      RECT 69.48 3.025 69.495 3.393 ;
      RECT 69.465 3.025 69.48 3.38 ;
      RECT 69.46 3.025 69.465 3.37 ;
      RECT 69.445 3.025 69.46 3.348 ;
      RECT 69.43 3.025 69.445 3.315 ;
      RECT 69.425 3.025 69.43 3.293 ;
      RECT 69.415 3.025 69.425 3.275 ;
      RECT 69.4 3.025 69.415 3.253 ;
      RECT 69.38 3.025 69.4 3.215 ;
      RECT 69.73 2.31 69.765 2.749 ;
      RECT 69.73 2.31 69.77 2.748 ;
      RECT 69.675 2.37 69.77 2.747 ;
      RECT 69.54 2.542 69.77 2.746 ;
      RECT 69.65 2.42 69.77 2.746 ;
      RECT 69.54 2.542 69.795 2.736 ;
      RECT 69.595 2.487 69.875 2.653 ;
      RECT 69.77 2.281 69.775 2.744 ;
      RECT 69.625 2.457 69.915 2.53 ;
      RECT 69.64 2.44 69.77 2.746 ;
      RECT 69.775 2.28 69.945 2.468 ;
      RECT 69.765 2.283 69.945 2.468 ;
      RECT 69.27 2.16 69.44 2.47 ;
      RECT 69.27 2.16 69.445 2.443 ;
      RECT 69.27 2.16 69.45 2.42 ;
      RECT 69.27 2.16 69.46 2.37 ;
      RECT 69.265 2.265 69.46 2.34 ;
      RECT 69.3 1.835 69.47 2.313 ;
      RECT 69.3 1.835 69.485 2.234 ;
      RECT 69.29 2.045 69.485 2.234 ;
      RECT 69.3 1.845 69.495 2.149 ;
      RECT 69.23 2.587 69.235 2.79 ;
      RECT 69.22 2.575 69.23 2.9 ;
      RECT 69.195 2.575 69.22 2.94 ;
      RECT 69.115 2.575 69.195 3.025 ;
      RECT 69.105 2.575 69.115 3.095 ;
      RECT 69.08 2.575 69.105 3.118 ;
      RECT 69.06 2.575 69.08 3.153 ;
      RECT 69.015 2.585 69.06 3.196 ;
      RECT 69.005 2.597 69.015 3.233 ;
      RECT 68.985 2.611 69.005 3.253 ;
      RECT 68.975 2.629 68.985 3.269 ;
      RECT 68.96 2.655 68.975 3.279 ;
      RECT 68.945 2.696 68.96 3.293 ;
      RECT 68.935 2.731 68.945 3.303 ;
      RECT 68.93 2.747 68.935 3.308 ;
      RECT 68.92 2.762 68.93 3.313 ;
      RECT 68.9 2.805 68.92 3.323 ;
      RECT 68.88 2.842 68.9 3.336 ;
      RECT 68.845 2.865 68.88 3.354 ;
      RECT 68.835 2.879 68.845 3.37 ;
      RECT 68.815 2.889 68.835 3.38 ;
      RECT 68.81 2.898 68.815 3.388 ;
      RECT 68.8 2.905 68.81 3.395 ;
      RECT 68.79 2.912 68.8 3.403 ;
      RECT 68.775 2.922 68.79 3.411 ;
      RECT 68.765 2.936 68.775 3.421 ;
      RECT 68.755 2.948 68.765 3.433 ;
      RECT 68.74 2.97 68.755 3.446 ;
      RECT 68.73 2.992 68.74 3.457 ;
      RECT 68.72 3.012 68.73 3.466 ;
      RECT 68.715 3.027 68.72 3.473 ;
      RECT 68.685 3.06 68.715 3.487 ;
      RECT 68.675 3.095 68.685 3.502 ;
      RECT 68.67 3.102 68.675 3.508 ;
      RECT 68.65 3.117 68.67 3.515 ;
      RECT 68.645 3.132 68.65 3.523 ;
      RECT 68.64 3.141 68.645 3.528 ;
      RECT 68.625 3.147 68.64 3.535 ;
      RECT 68.62 3.153 68.625 3.543 ;
      RECT 68.615 3.157 68.62 3.55 ;
      RECT 68.61 3.161 68.615 3.56 ;
      RECT 68.6 3.166 68.61 3.57 ;
      RECT 68.58 3.177 68.6 3.598 ;
      RECT 68.565 3.189 68.58 3.625 ;
      RECT 68.545 3.202 68.565 3.65 ;
      RECT 68.525 3.217 68.545 3.674 ;
      RECT 68.51 3.232 68.525 3.689 ;
      RECT 68.505 3.243 68.51 3.698 ;
      RECT 68.44 3.288 68.505 3.708 ;
      RECT 68.405 3.347 68.44 3.721 ;
      RECT 68.4 3.37 68.405 3.727 ;
      RECT 68.395 3.377 68.4 3.729 ;
      RECT 68.38 3.387 68.395 3.732 ;
      RECT 68.35 3.412 68.38 3.736 ;
      RECT 68.345 3.43 68.35 3.74 ;
      RECT 68.34 3.437 68.345 3.741 ;
      RECT 68.32 3.445 68.34 3.745 ;
      RECT 68.31 3.452 68.32 3.749 ;
      RECT 68.266 3.463 68.31 3.756 ;
      RECT 68.18 3.491 68.266 3.772 ;
      RECT 68.12 3.515 68.18 3.79 ;
      RECT 68.075 3.525 68.12 3.804 ;
      RECT 68.016 3.533 68.075 3.818 ;
      RECT 67.93 3.54 68.016 3.837 ;
      RECT 67.905 3.545 67.93 3.852 ;
      RECT 67.825 3.548 67.905 3.855 ;
      RECT 67.745 3.552 67.825 3.842 ;
      RECT 67.736 3.555 67.745 3.827 ;
      RECT 67.65 3.555 67.736 3.812 ;
      RECT 67.59 3.557 67.65 3.789 ;
      RECT 67.586 3.56 67.59 3.779 ;
      RECT 67.5 3.56 67.586 3.764 ;
      RECT 67.425 3.56 67.5 3.74 ;
      RECT 68.74 2.569 68.75 2.745 ;
      RECT 68.695 2.536 68.74 2.745 ;
      RECT 68.65 2.487 68.695 2.745 ;
      RECT 68.62 2.457 68.65 2.746 ;
      RECT 68.615 2.44 68.62 2.747 ;
      RECT 68.59 2.42 68.615 2.748 ;
      RECT 68.575 2.395 68.59 2.749 ;
      RECT 68.57 2.382 68.575 2.75 ;
      RECT 68.565 2.376 68.57 2.748 ;
      RECT 68.56 2.368 68.565 2.742 ;
      RECT 68.535 2.36 68.56 2.722 ;
      RECT 68.515 2.349 68.535 2.693 ;
      RECT 68.485 2.334 68.515 2.664 ;
      RECT 68.465 2.32 68.485 2.636 ;
      RECT 68.455 2.314 68.465 2.615 ;
      RECT 68.45 2.311 68.455 2.598 ;
      RECT 68.445 2.308 68.45 2.583 ;
      RECT 68.43 2.303 68.445 2.548 ;
      RECT 68.425 2.299 68.43 2.515 ;
      RECT 68.405 2.294 68.425 2.491 ;
      RECT 68.375 2.286 68.405 2.456 ;
      RECT 68.36 2.28 68.375 2.433 ;
      RECT 68.32 2.273 68.36 2.418 ;
      RECT 68.295 2.265 68.32 2.398 ;
      RECT 68.275 2.26 68.295 2.388 ;
      RECT 68.24 2.254 68.275 2.383 ;
      RECT 68.195 2.245 68.24 2.382 ;
      RECT 68.165 2.241 68.195 2.384 ;
      RECT 68.08 2.249 68.165 2.388 ;
      RECT 68.01 2.26 68.08 2.41 ;
      RECT 67.997 2.266 68.01 2.433 ;
      RECT 67.911 2.273 67.997 2.455 ;
      RECT 67.825 2.285 67.911 2.492 ;
      RECT 67.825 2.662 67.835 2.9 ;
      RECT 67.82 2.291 67.825 2.515 ;
      RECT 67.815 2.547 67.825 2.9 ;
      RECT 67.815 2.292 67.82 2.52 ;
      RECT 67.81 2.293 67.815 2.9 ;
      RECT 67.786 2.295 67.81 2.901 ;
      RECT 67.7 2.303 67.786 2.903 ;
      RECT 67.68 2.317 67.7 2.906 ;
      RECT 67.675 2.345 67.68 2.907 ;
      RECT 67.67 2.357 67.675 2.908 ;
      RECT 67.665 2.372 67.67 2.909 ;
      RECT 67.655 2.402 67.665 2.91 ;
      RECT 67.65 2.44 67.655 2.908 ;
      RECT 67.645 2.46 67.65 2.903 ;
      RECT 67.63 2.495 67.645 2.888 ;
      RECT 67.62 2.547 67.63 2.868 ;
      RECT 67.615 2.577 67.62 2.856 ;
      RECT 67.6 2.59 67.615 2.839 ;
      RECT 67.575 2.594 67.6 2.806 ;
      RECT 67.56 2.592 67.575 2.783 ;
      RECT 67.545 2.591 67.56 2.78 ;
      RECT 67.485 2.589 67.545 2.778 ;
      RECT 67.475 2.587 67.485 2.773 ;
      RECT 67.435 2.586 67.475 2.77 ;
      RECT 67.365 2.583 67.435 2.768 ;
      RECT 67.31 2.581 67.365 2.763 ;
      RECT 67.24 2.575 67.31 2.758 ;
      RECT 67.231 2.575 67.24 2.755 ;
      RECT 67.145 2.575 67.231 2.75 ;
      RECT 67.14 2.575 67.145 2.745 ;
      RECT 68.445 1.81 68.62 2.16 ;
      RECT 68.445 1.825 68.63 2.158 ;
      RECT 68.42 1.775 68.565 2.155 ;
      RECT 68.4 1.776 68.565 2.148 ;
      RECT 68.39 1.777 68.575 2.143 ;
      RECT 68.36 1.778 68.575 2.13 ;
      RECT 68.31 1.779 68.575 2.106 ;
      RECT 68.305 1.781 68.575 2.091 ;
      RECT 68.305 1.847 68.635 2.085 ;
      RECT 68.285 1.788 68.59 2.065 ;
      RECT 68.275 1.797 68.6 1.92 ;
      RECT 68.285 1.792 68.6 2.065 ;
      RECT 68.305 1.782 68.59 2.091 ;
      RECT 67.89 3.107 68.06 3.395 ;
      RECT 67.885 3.125 68.07 3.39 ;
      RECT 67.85 3.133 68.135 3.31 ;
      RECT 67.85 3.133 68.221 3.3 ;
      RECT 67.85 3.133 68.275 3.246 ;
      RECT 68.135 3.03 68.305 3.214 ;
      RECT 67.85 3.185 68.31 3.202 ;
      RECT 67.835 3.155 68.305 3.198 ;
      RECT 68.095 3.037 68.135 3.349 ;
      RECT 67.975 3.074 68.305 3.214 ;
      RECT 68.07 3.049 68.095 3.375 ;
      RECT 68.06 3.056 68.305 3.214 ;
      RECT 68.191 2.52 68.26 2.779 ;
      RECT 68.191 2.575 68.265 2.778 ;
      RECT 68.105 2.575 68.265 2.777 ;
      RECT 68.1 2.575 68.27 2.77 ;
      RECT 68.09 2.52 68.26 2.765 ;
      RECT 67.47 1.819 67.645 2.12 ;
      RECT 67.455 1.807 67.47 2.105 ;
      RECT 67.425 1.806 67.455 2.058 ;
      RECT 67.425 1.824 67.65 2.053 ;
      RECT 67.41 1.808 67.47 2.018 ;
      RECT 67.405 1.83 67.66 1.918 ;
      RECT 67.405 1.813 67.556 1.918 ;
      RECT 67.405 1.815 67.56 1.918 ;
      RECT 67.41 1.811 67.556 2.018 ;
      RECT 67.515 3.047 67.52 3.395 ;
      RECT 67.505 3.037 67.515 3.401 ;
      RECT 67.47 3.027 67.505 3.403 ;
      RECT 67.432 3.022 67.47 3.407 ;
      RECT 67.346 3.015 67.432 3.414 ;
      RECT 67.26 3.005 67.346 3.424 ;
      RECT 67.215 3 67.26 3.432 ;
      RECT 67.211 3 67.215 3.436 ;
      RECT 67.125 3 67.211 3.443 ;
      RECT 67.11 3 67.125 3.443 ;
      RECT 67.1 2.998 67.11 3.415 ;
      RECT 67.09 2.994 67.1 3.358 ;
      RECT 67.07 2.988 67.09 3.29 ;
      RECT 67.065 2.984 67.07 3.238 ;
      RECT 67.055 2.983 67.065 3.205 ;
      RECT 67.005 2.981 67.055 3.19 ;
      RECT 66.98 2.979 67.005 3.185 ;
      RECT 66.937 2.977 66.98 3.181 ;
      RECT 66.851 2.973 66.937 3.169 ;
      RECT 66.765 2.968 66.851 3.153 ;
      RECT 66.735 2.965 66.765 3.14 ;
      RECT 66.71 2.964 66.735 3.128 ;
      RECT 66.705 2.964 66.71 3.118 ;
      RECT 66.665 2.963 66.705 3.11 ;
      RECT 66.65 2.962 66.665 3.103 ;
      RECT 66.6 2.961 66.65 3.095 ;
      RECT 66.598 2.96 66.6 3.09 ;
      RECT 66.512 2.958 66.598 3.09 ;
      RECT 66.426 2.953 66.512 3.09 ;
      RECT 66.34 2.949 66.426 3.09 ;
      RECT 66.291 2.945 66.34 3.088 ;
      RECT 66.205 2.942 66.291 3.083 ;
      RECT 66.182 2.939 66.205 3.079 ;
      RECT 66.096 2.936 66.182 3.074 ;
      RECT 66.01 2.932 66.096 3.065 ;
      RECT 65.985 2.925 66.01 3.06 ;
      RECT 65.925 2.89 65.985 3.057 ;
      RECT 65.905 2.815 65.925 3.054 ;
      RECT 65.9 2.757 65.905 3.053 ;
      RECT 65.875 2.697 65.9 3.052 ;
      RECT 65.8 2.575 65.875 3.048 ;
      RECT 65.79 2.575 65.8 3.04 ;
      RECT 65.775 2.575 65.79 3.03 ;
      RECT 65.76 2.575 65.775 3 ;
      RECT 65.745 2.575 65.76 2.945 ;
      RECT 65.73 2.575 65.745 2.883 ;
      RECT 65.705 2.575 65.73 2.808 ;
      RECT 65.7 2.575 65.705 2.758 ;
      RECT 67.045 2.12 67.065 2.429 ;
      RECT 67.031 2.122 67.08 2.426 ;
      RECT 67.031 2.127 67.1 2.417 ;
      RECT 66.945 2.125 67.08 2.411 ;
      RECT 66.945 2.133 67.135 2.394 ;
      RECT 66.91 2.135 67.135 2.393 ;
      RECT 66.88 2.143 67.135 2.384 ;
      RECT 66.87 2.148 67.155 2.37 ;
      RECT 66.91 2.138 67.155 2.37 ;
      RECT 66.91 2.141 67.165 2.358 ;
      RECT 66.88 2.143 67.175 2.345 ;
      RECT 66.88 2.147 67.185 2.288 ;
      RECT 66.87 2.152 67.19 2.203 ;
      RECT 67.031 2.12 67.065 2.426 ;
      RECT 66.91 7.855 67.08 8.305 ;
      RECT 66.965 6.075 67.135 8.025 ;
      RECT 66.91 5.015 67.08 6.245 ;
      RECT 66.47 2.223 66.475 2.435 ;
      RECT 66.345 2.22 66.36 2.435 ;
      RECT 65.81 2.25 65.88 2.435 ;
      RECT 65.695 2.25 65.73 2.43 ;
      RECT 66.816 2.552 66.835 2.746 ;
      RECT 66.73 2.507 66.816 2.747 ;
      RECT 66.72 2.46 66.73 2.749 ;
      RECT 66.715 2.44 66.72 2.75 ;
      RECT 66.695 2.405 66.715 2.751 ;
      RECT 66.68 2.355 66.695 2.752 ;
      RECT 66.66 2.292 66.68 2.753 ;
      RECT 66.65 2.255 66.66 2.754 ;
      RECT 66.635 2.244 66.65 2.755 ;
      RECT 66.63 2.236 66.635 2.753 ;
      RECT 66.62 2.235 66.63 2.745 ;
      RECT 66.59 2.232 66.62 2.724 ;
      RECT 66.515 2.227 66.59 2.669 ;
      RECT 66.5 2.223 66.515 2.615 ;
      RECT 66.49 2.223 66.5 2.51 ;
      RECT 66.475 2.223 66.49 2.443 ;
      RECT 66.46 2.223 66.47 2.433 ;
      RECT 66.405 2.222 66.46 2.43 ;
      RECT 66.36 2.22 66.405 2.433 ;
      RECT 66.332 2.22 66.345 2.436 ;
      RECT 66.246 2.224 66.332 2.438 ;
      RECT 66.16 2.23 66.246 2.443 ;
      RECT 66.14 2.234 66.16 2.445 ;
      RECT 66.138 2.235 66.14 2.444 ;
      RECT 66.052 2.237 66.138 2.443 ;
      RECT 65.966 2.242 66.052 2.44 ;
      RECT 65.88 2.247 65.966 2.437 ;
      RECT 65.73 2.25 65.81 2.433 ;
      RECT 66.39 5.015 66.56 8.305 ;
      RECT 66.39 7.315 66.795 7.645 ;
      RECT 66.39 6.475 66.795 6.805 ;
      RECT 66.506 3.225 66.555 3.559 ;
      RECT 66.506 3.225 66.56 3.558 ;
      RECT 66.42 3.225 66.56 3.557 ;
      RECT 66.195 3.333 66.565 3.555 ;
      RECT 66.42 3.225 66.59 3.548 ;
      RECT 66.39 3.237 66.595 3.539 ;
      RECT 66.375 3.255 66.6 3.536 ;
      RECT 66.19 3.339 66.6 3.463 ;
      RECT 66.185 3.346 66.6 3.423 ;
      RECT 66.2 3.312 66.6 3.536 ;
      RECT 66.361 3.258 66.565 3.555 ;
      RECT 66.275 3.278 66.6 3.536 ;
      RECT 66.375 3.252 66.595 3.539 ;
      RECT 66.145 2.576 66.335 2.77 ;
      RECT 66.14 2.578 66.335 2.769 ;
      RECT 66.135 2.582 66.35 2.766 ;
      RECT 66.15 2.575 66.35 2.766 ;
      RECT 66.135 2.685 66.355 2.761 ;
      RECT 65.43 3.185 65.521 3.483 ;
      RECT 65.425 3.187 65.6 3.478 ;
      RECT 65.43 3.185 65.6 3.478 ;
      RECT 65.425 3.191 65.62 3.476 ;
      RECT 65.425 3.246 65.66 3.475 ;
      RECT 65.425 3.281 65.675 3.469 ;
      RECT 65.425 3.315 65.685 3.459 ;
      RECT 65.415 3.195 65.62 3.31 ;
      RECT 65.415 3.215 65.635 3.31 ;
      RECT 65.415 3.198 65.625 3.31 ;
      RECT 65.64 1.966 65.645 2.028 ;
      RECT 65.635 1.888 65.64 2.051 ;
      RECT 65.63 1.845 65.635 2.062 ;
      RECT 65.625 1.835 65.63 2.074 ;
      RECT 65.62 1.835 65.625 2.083 ;
      RECT 65.595 1.835 65.62 2.115 ;
      RECT 65.59 1.835 65.595 2.148 ;
      RECT 65.575 1.835 65.59 2.173 ;
      RECT 65.565 1.835 65.575 2.2 ;
      RECT 65.56 1.835 65.565 2.213 ;
      RECT 65.555 1.835 65.56 2.228 ;
      RECT 65.545 1.835 65.555 2.243 ;
      RECT 65.54 1.835 65.545 2.263 ;
      RECT 65.515 1.835 65.54 2.298 ;
      RECT 65.47 1.835 65.515 2.343 ;
      RECT 65.46 1.835 65.47 2.356 ;
      RECT 65.375 1.92 65.46 2.363 ;
      RECT 65.34 2.042 65.375 2.372 ;
      RECT 65.335 2.082 65.34 2.376 ;
      RECT 65.315 2.105 65.335 2.378 ;
      RECT 65.31 2.135 65.315 2.381 ;
      RECT 65.3 2.147 65.31 2.382 ;
      RECT 65.255 2.17 65.3 2.387 ;
      RECT 65.215 2.2 65.255 2.395 ;
      RECT 65.18 2.212 65.215 2.401 ;
      RECT 65.175 2.217 65.18 2.405 ;
      RECT 65.105 2.227 65.175 2.412 ;
      RECT 65.065 2.237 65.105 2.422 ;
      RECT 65.045 2.242 65.065 2.428 ;
      RECT 65.035 2.246 65.045 2.433 ;
      RECT 65.03 2.249 65.035 2.436 ;
      RECT 65.02 2.25 65.03 2.437 ;
      RECT 64.995 2.252 65.02 2.441 ;
      RECT 64.985 2.257 64.995 2.444 ;
      RECT 64.94 2.265 64.985 2.445 ;
      RECT 64.815 2.27 64.94 2.445 ;
      RECT 65.37 2.567 65.39 2.749 ;
      RECT 65.321 2.552 65.37 2.748 ;
      RECT 65.235 2.567 65.39 2.746 ;
      RECT 65.22 2.567 65.39 2.745 ;
      RECT 65.185 2.545 65.355 2.73 ;
      RECT 65.255 3.565 65.27 3.774 ;
      RECT 65.255 3.573 65.275 3.773 ;
      RECT 65.2 3.573 65.275 3.772 ;
      RECT 65.18 3.577 65.28 3.77 ;
      RECT 65.16 3.527 65.2 3.769 ;
      RECT 65.105 3.585 65.285 3.767 ;
      RECT 65.07 3.542 65.2 3.765 ;
      RECT 65.066 3.545 65.255 3.764 ;
      RECT 64.98 3.553 65.255 3.762 ;
      RECT 64.98 3.597 65.29 3.755 ;
      RECT 64.97 3.69 65.29 3.753 ;
      RECT 64.98 3.609 65.295 3.738 ;
      RECT 64.98 3.63 65.31 3.708 ;
      RECT 64.98 3.657 65.315 3.678 ;
      RECT 65.105 3.535 65.2 3.767 ;
      RECT 64.735 2.58 64.74 3.118 ;
      RECT 64.54 2.91 64.545 3.105 ;
      RECT 62.84 2.575 62.855 2.955 ;
      RECT 64.905 2.575 64.91 2.745 ;
      RECT 64.9 2.575 64.905 2.755 ;
      RECT 64.895 2.575 64.9 2.768 ;
      RECT 64.87 2.575 64.895 2.81 ;
      RECT 64.845 2.575 64.87 2.883 ;
      RECT 64.83 2.575 64.845 2.935 ;
      RECT 64.825 2.575 64.83 2.965 ;
      RECT 64.8 2.575 64.825 3.005 ;
      RECT 64.785 2.575 64.8 3.06 ;
      RECT 64.78 2.575 64.785 3.093 ;
      RECT 64.755 2.575 64.78 3.113 ;
      RECT 64.74 2.575 64.755 3.119 ;
      RECT 64.67 2.61 64.735 3.115 ;
      RECT 64.62 2.665 64.67 3.11 ;
      RECT 64.61 2.697 64.62 3.108 ;
      RECT 64.605 2.722 64.61 3.108 ;
      RECT 64.585 2.795 64.605 3.108 ;
      RECT 64.575 2.875 64.585 3.107 ;
      RECT 64.56 2.905 64.575 3.107 ;
      RECT 64.545 2.91 64.56 3.106 ;
      RECT 64.485 2.912 64.54 3.103 ;
      RECT 64.455 2.917 64.485 3.099 ;
      RECT 64.453 2.92 64.455 3.098 ;
      RECT 64.367 2.922 64.453 3.095 ;
      RECT 64.281 2.928 64.367 3.089 ;
      RECT 64.195 2.933 64.281 3.083 ;
      RECT 64.122 2.938 64.195 3.084 ;
      RECT 64.036 2.944 64.122 3.092 ;
      RECT 63.95 2.95 64.036 3.101 ;
      RECT 63.93 2.954 63.95 3.106 ;
      RECT 63.883 2.956 63.93 3.109 ;
      RECT 63.797 2.961 63.883 3.115 ;
      RECT 63.711 2.966 63.797 3.124 ;
      RECT 63.625 2.972 63.711 3.132 ;
      RECT 63.54 2.97 63.625 3.141 ;
      RECT 63.536 2.965 63.54 3.145 ;
      RECT 63.45 2.96 63.536 3.137 ;
      RECT 63.386 2.951 63.45 3.125 ;
      RECT 63.3 2.942 63.386 3.112 ;
      RECT 63.276 2.935 63.3 3.103 ;
      RECT 63.19 2.929 63.276 3.09 ;
      RECT 63.15 2.922 63.19 3.076 ;
      RECT 63.145 2.912 63.15 3.072 ;
      RECT 63.135 2.9 63.145 3.071 ;
      RECT 63.115 2.87 63.135 3.068 ;
      RECT 63.06 2.79 63.115 3.062 ;
      RECT 63.04 2.709 63.06 3.057 ;
      RECT 63.02 2.667 63.04 3.053 ;
      RECT 62.995 2.62 63.02 3.047 ;
      RECT 62.99 2.595 62.995 3.044 ;
      RECT 62.955 2.575 62.99 3.039 ;
      RECT 62.946 2.575 62.955 3.032 ;
      RECT 62.86 2.575 62.946 3.002 ;
      RECT 62.855 2.575 62.86 2.965 ;
      RECT 62.82 2.575 62.84 2.887 ;
      RECT 62.815 2.617 62.82 2.852 ;
      RECT 62.81 2.692 62.815 2.808 ;
      RECT 64.26 2.497 64.435 2.745 ;
      RECT 64.26 2.497 64.44 2.743 ;
      RECT 64.255 2.529 64.44 2.703 ;
      RECT 64.285 2.47 64.455 2.69 ;
      RECT 64.25 2.547 64.455 2.623 ;
      RECT 63.56 2.01 63.73 2.185 ;
      RECT 63.56 2.01 63.902 2.177 ;
      RECT 63.56 2.01 63.985 2.171 ;
      RECT 63.56 2.01 64.02 2.167 ;
      RECT 63.56 2.01 64.04 2.166 ;
      RECT 63.56 2.01 64.126 2.162 ;
      RECT 64.02 1.835 64.19 2.157 ;
      RECT 63.595 1.942 64.22 2.155 ;
      RECT 63.585 1.997 64.225 2.153 ;
      RECT 63.56 2.033 64.235 2.148 ;
      RECT 63.56 2.06 64.24 2.078 ;
      RECT 63.625 1.885 64.2 2.155 ;
      RECT 63.816 1.87 64.2 2.155 ;
      RECT 63.65 1.873 64.2 2.155 ;
      RECT 63.73 1.871 63.816 2.182 ;
      RECT 63.816 1.868 64.195 2.155 ;
      RECT 64 1.845 64.195 2.155 ;
      RECT 63.902 1.866 64.195 2.155 ;
      RECT 63.985 1.86 64 2.168 ;
      RECT 64.135 3.225 64.14 3.425 ;
      RECT 63.6 3.29 63.645 3.425 ;
      RECT 64.17 3.225 64.19 3.398 ;
      RECT 64.14 3.225 64.17 3.413 ;
      RECT 64.075 3.225 64.135 3.45 ;
      RECT 64.06 3.225 64.075 3.48 ;
      RECT 64.045 3.225 64.06 3.493 ;
      RECT 64.025 3.225 64.045 3.508 ;
      RECT 64.02 3.225 64.025 3.517 ;
      RECT 64.01 3.229 64.02 3.522 ;
      RECT 63.995 3.239 64.01 3.533 ;
      RECT 63.97 3.255 63.995 3.543 ;
      RECT 63.96 3.269 63.97 3.545 ;
      RECT 63.94 3.281 63.96 3.542 ;
      RECT 63.91 3.302 63.94 3.536 ;
      RECT 63.9 3.314 63.91 3.531 ;
      RECT 63.89 3.312 63.9 3.528 ;
      RECT 63.875 3.311 63.89 3.523 ;
      RECT 63.87 3.31 63.875 3.518 ;
      RECT 63.835 3.308 63.87 3.508 ;
      RECT 63.815 3.305 63.835 3.49 ;
      RECT 63.805 3.303 63.815 3.485 ;
      RECT 63.795 3.302 63.805 3.48 ;
      RECT 63.76 3.3 63.795 3.468 ;
      RECT 63.705 3.296 63.76 3.448 ;
      RECT 63.695 3.294 63.705 3.433 ;
      RECT 63.69 3.294 63.695 3.428 ;
      RECT 63.645 3.292 63.69 3.425 ;
      RECT 63.55 3.29 63.6 3.429 ;
      RECT 63.54 3.291 63.55 3.434 ;
      RECT 63.48 3.298 63.54 3.448 ;
      RECT 63.455 3.306 63.48 3.468 ;
      RECT 63.445 3.31 63.455 3.48 ;
      RECT 63.44 3.311 63.445 3.485 ;
      RECT 63.425 3.313 63.44 3.488 ;
      RECT 63.41 3.315 63.425 3.493 ;
      RECT 63.405 3.315 63.41 3.496 ;
      RECT 63.36 3.32 63.405 3.507 ;
      RECT 63.355 3.324 63.36 3.519 ;
      RECT 63.33 3.32 63.355 3.523 ;
      RECT 63.32 3.316 63.33 3.527 ;
      RECT 63.31 3.315 63.32 3.531 ;
      RECT 63.295 3.305 63.31 3.537 ;
      RECT 63.29 3.293 63.295 3.541 ;
      RECT 63.285 3.29 63.29 3.542 ;
      RECT 63.28 3.287 63.285 3.544 ;
      RECT 63.265 3.275 63.28 3.543 ;
      RECT 63.25 3.257 63.265 3.54 ;
      RECT 63.23 3.236 63.25 3.533 ;
      RECT 63.165 3.225 63.23 3.505 ;
      RECT 63.161 3.225 63.165 3.484 ;
      RECT 63.075 3.225 63.161 3.454 ;
      RECT 63.06 3.225 63.075 3.41 ;
      RECT 63.635 2.325 63.64 2.56 ;
      RECT 62.765 2.241 62.77 2.445 ;
      RECT 63.345 2.27 63.35 2.425 ;
      RECT 63.265 2.25 63.27 2.425 ;
      RECT 63.935 2.392 63.95 2.745 ;
      RECT 63.861 2.377 63.935 2.745 ;
      RECT 63.775 2.36 63.861 2.745 ;
      RECT 63.765 2.35 63.775 2.743 ;
      RECT 63.76 2.348 63.765 2.738 ;
      RECT 63.745 2.346 63.76 2.724 ;
      RECT 63.675 2.338 63.745 2.664 ;
      RECT 63.655 2.329 63.675 2.598 ;
      RECT 63.65 2.326 63.655 2.578 ;
      RECT 63.64 2.325 63.65 2.568 ;
      RECT 63.63 2.325 63.635 2.552 ;
      RECT 63.62 2.324 63.63 2.542 ;
      RECT 63.61 2.322 63.62 2.53 ;
      RECT 63.595 2.319 63.61 2.51 ;
      RECT 63.585 2.317 63.595 2.495 ;
      RECT 63.565 2.314 63.585 2.483 ;
      RECT 63.56 2.312 63.565 2.473 ;
      RECT 63.535 2.31 63.56 2.46 ;
      RECT 63.505 2.305 63.535 2.445 ;
      RECT 63.425 2.296 63.505 2.436 ;
      RECT 63.38 2.285 63.425 2.429 ;
      RECT 63.36 2.276 63.38 2.426 ;
      RECT 63.35 2.271 63.36 2.425 ;
      RECT 63.305 2.265 63.345 2.425 ;
      RECT 63.29 2.257 63.305 2.425 ;
      RECT 63.27 2.252 63.29 2.425 ;
      RECT 63.25 2.249 63.265 2.425 ;
      RECT 63.167 2.248 63.25 2.424 ;
      RECT 63.081 2.247 63.167 2.42 ;
      RECT 62.995 2.245 63.081 2.417 ;
      RECT 62.942 2.244 62.995 2.419 ;
      RECT 62.856 2.243 62.942 2.428 ;
      RECT 62.77 2.242 62.856 2.44 ;
      RECT 62.75 2.241 62.765 2.448 ;
      RECT 62.67 2.24 62.75 2.46 ;
      RECT 62.645 2.24 62.67 2.473 ;
      RECT 62.62 2.24 62.645 2.488 ;
      RECT 62.615 2.24 62.62 2.51 ;
      RECT 62.61 2.24 62.615 2.528 ;
      RECT 62.605 2.24 62.61 2.545 ;
      RECT 62.6 2.24 62.605 2.558 ;
      RECT 62.595 2.24 62.6 2.568 ;
      RECT 62.555 2.24 62.595 2.653 ;
      RECT 62.54 2.24 62.555 2.738 ;
      RECT 62.53 2.241 62.54 2.75 ;
      RECT 62.495 2.246 62.53 2.755 ;
      RECT 62.455 2.255 62.495 2.755 ;
      RECT 62.44 2.265 62.455 2.755 ;
      RECT 62.435 2.275 62.44 2.755 ;
      RECT 62.415 2.302 62.435 2.755 ;
      RECT 62.365 2.385 62.415 2.755 ;
      RECT 62.36 2.447 62.365 2.755 ;
      RECT 62.35 2.46 62.36 2.755 ;
      RECT 62.34 2.482 62.35 2.755 ;
      RECT 62.33 2.507 62.34 2.75 ;
      RECT 62.325 2.545 62.33 2.743 ;
      RECT 62.315 2.655 62.325 2.738 ;
      RECT 63.71 3.576 63.725 3.835 ;
      RECT 63.71 3.591 63.73 3.834 ;
      RECT 63.626 3.591 63.73 3.832 ;
      RECT 63.626 3.605 63.735 3.831 ;
      RECT 63.54 3.647 63.74 3.828 ;
      RECT 63.535 3.59 63.725 3.823 ;
      RECT 63.535 3.661 63.745 3.82 ;
      RECT 63.53 3.692 63.745 3.818 ;
      RECT 63.535 3.689 63.76 3.808 ;
      RECT 63.53 3.735 63.775 3.793 ;
      RECT 63.53 3.763 63.78 3.778 ;
      RECT 63.54 3.565 63.71 3.828 ;
      RECT 63.3 2.575 63.47 2.745 ;
      RECT 63.265 2.575 63.47 2.74 ;
      RECT 63.255 2.575 63.47 2.733 ;
      RECT 63.25 2.56 63.42 2.73 ;
      RECT 62.08 3.097 62.345 3.54 ;
      RECT 62.075 3.068 62.29 3.538 ;
      RECT 62.07 3.222 62.35 3.533 ;
      RECT 62.075 3.117 62.35 3.533 ;
      RECT 62.075 3.128 62.36 3.52 ;
      RECT 62.075 3.075 62.32 3.538 ;
      RECT 62.08 3.062 62.29 3.54 ;
      RECT 62.08 3.06 62.24 3.54 ;
      RECT 62.181 3.052 62.24 3.54 ;
      RECT 62.095 3.053 62.24 3.54 ;
      RECT 62.181 3.051 62.23 3.54 ;
      RECT 61.985 1.866 62.16 2.165 ;
      RECT 62.035 1.828 62.16 2.165 ;
      RECT 62.02 1.83 62.246 2.157 ;
      RECT 62.02 1.833 62.285 2.144 ;
      RECT 62.02 1.834 62.295 2.13 ;
      RECT 61.975 1.885 62.295 2.12 ;
      RECT 62.02 1.835 62.3 2.115 ;
      RECT 61.975 2.045 62.305 2.105 ;
      RECT 61.96 1.905 62.3 2.045 ;
      RECT 61.955 1.921 62.3 1.985 ;
      RECT 62 1.845 62.3 2.115 ;
      RECT 62.035 1.826 62.121 2.165 ;
      RECT 60.13 1.74 60.3 2.935 ;
      RECT 60.13 1.74 60.595 1.91 ;
      RECT 60.13 6.97 60.595 7.14 ;
      RECT 60.13 5.945 60.3 7.14 ;
      RECT 59.14 1.74 59.31 2.935 ;
      RECT 59.14 1.74 59.605 1.91 ;
      RECT 59.14 6.97 59.605 7.14 ;
      RECT 59.14 5.945 59.31 7.14 ;
      RECT 57.285 2.635 57.455 3.865 ;
      RECT 57.34 0.855 57.51 2.805 ;
      RECT 57.285 0.575 57.455 1.025 ;
      RECT 57.285 7.855 57.455 8.305 ;
      RECT 57.34 6.075 57.51 8.025 ;
      RECT 57.285 5.015 57.455 6.245 ;
      RECT 56.765 0.575 56.935 3.865 ;
      RECT 56.765 2.075 57.17 2.405 ;
      RECT 56.765 1.235 57.17 1.565 ;
      RECT 56.765 5.015 56.935 8.305 ;
      RECT 56.765 7.315 57.17 7.645 ;
      RECT 56.765 6.475 57.17 6.805 ;
      RECT 54.69 3.126 54.695 3.298 ;
      RECT 54.685 3.119 54.69 3.388 ;
      RECT 54.68 3.113 54.685 3.407 ;
      RECT 54.66 3.107 54.68 3.417 ;
      RECT 54.645 3.102 54.66 3.425 ;
      RECT 54.608 3.096 54.645 3.423 ;
      RECT 54.522 3.082 54.608 3.419 ;
      RECT 54.436 3.064 54.522 3.414 ;
      RECT 54.35 3.045 54.436 3.408 ;
      RECT 54.32 3.033 54.35 3.404 ;
      RECT 54.3 3.027 54.32 3.403 ;
      RECT 54.235 3.025 54.3 3.401 ;
      RECT 54.22 3.025 54.235 3.393 ;
      RECT 54.205 3.025 54.22 3.38 ;
      RECT 54.2 3.025 54.205 3.37 ;
      RECT 54.185 3.025 54.2 3.348 ;
      RECT 54.17 3.025 54.185 3.315 ;
      RECT 54.165 3.025 54.17 3.293 ;
      RECT 54.155 3.025 54.165 3.275 ;
      RECT 54.14 3.025 54.155 3.253 ;
      RECT 54.12 3.025 54.14 3.215 ;
      RECT 54.47 2.31 54.505 2.749 ;
      RECT 54.47 2.31 54.51 2.748 ;
      RECT 54.415 2.37 54.51 2.747 ;
      RECT 54.28 2.542 54.51 2.746 ;
      RECT 54.39 2.42 54.51 2.746 ;
      RECT 54.28 2.542 54.535 2.736 ;
      RECT 54.335 2.487 54.615 2.653 ;
      RECT 54.51 2.281 54.515 2.744 ;
      RECT 54.365 2.457 54.655 2.53 ;
      RECT 54.38 2.44 54.51 2.746 ;
      RECT 54.515 2.28 54.685 2.468 ;
      RECT 54.505 2.283 54.685 2.468 ;
      RECT 54.01 2.16 54.18 2.47 ;
      RECT 54.01 2.16 54.185 2.443 ;
      RECT 54.01 2.16 54.19 2.42 ;
      RECT 54.01 2.16 54.2 2.37 ;
      RECT 54.005 2.265 54.2 2.34 ;
      RECT 54.04 1.835 54.21 2.313 ;
      RECT 54.04 1.835 54.225 2.234 ;
      RECT 54.03 2.045 54.225 2.234 ;
      RECT 54.04 1.845 54.235 2.149 ;
      RECT 53.97 2.587 53.975 2.79 ;
      RECT 53.96 2.575 53.97 2.9 ;
      RECT 53.935 2.575 53.96 2.94 ;
      RECT 53.855 2.575 53.935 3.025 ;
      RECT 53.845 2.575 53.855 3.095 ;
      RECT 53.82 2.575 53.845 3.118 ;
      RECT 53.8 2.575 53.82 3.153 ;
      RECT 53.755 2.585 53.8 3.196 ;
      RECT 53.745 2.597 53.755 3.233 ;
      RECT 53.725 2.611 53.745 3.253 ;
      RECT 53.715 2.629 53.725 3.269 ;
      RECT 53.7 2.655 53.715 3.279 ;
      RECT 53.685 2.696 53.7 3.293 ;
      RECT 53.675 2.731 53.685 3.303 ;
      RECT 53.67 2.747 53.675 3.308 ;
      RECT 53.66 2.762 53.67 3.313 ;
      RECT 53.64 2.805 53.66 3.323 ;
      RECT 53.62 2.842 53.64 3.336 ;
      RECT 53.585 2.865 53.62 3.354 ;
      RECT 53.575 2.879 53.585 3.37 ;
      RECT 53.555 2.889 53.575 3.38 ;
      RECT 53.55 2.898 53.555 3.388 ;
      RECT 53.54 2.905 53.55 3.395 ;
      RECT 53.53 2.912 53.54 3.403 ;
      RECT 53.515 2.922 53.53 3.411 ;
      RECT 53.505 2.936 53.515 3.421 ;
      RECT 53.495 2.948 53.505 3.433 ;
      RECT 53.48 2.97 53.495 3.446 ;
      RECT 53.47 2.992 53.48 3.457 ;
      RECT 53.46 3.012 53.47 3.466 ;
      RECT 53.455 3.027 53.46 3.473 ;
      RECT 53.425 3.06 53.455 3.487 ;
      RECT 53.415 3.095 53.425 3.502 ;
      RECT 53.41 3.102 53.415 3.508 ;
      RECT 53.39 3.117 53.41 3.515 ;
      RECT 53.385 3.132 53.39 3.523 ;
      RECT 53.38 3.141 53.385 3.528 ;
      RECT 53.365 3.147 53.38 3.535 ;
      RECT 53.36 3.153 53.365 3.543 ;
      RECT 53.355 3.157 53.36 3.55 ;
      RECT 53.35 3.161 53.355 3.56 ;
      RECT 53.34 3.166 53.35 3.57 ;
      RECT 53.32 3.177 53.34 3.598 ;
      RECT 53.305 3.189 53.32 3.625 ;
      RECT 53.285 3.202 53.305 3.65 ;
      RECT 53.265 3.217 53.285 3.674 ;
      RECT 53.25 3.232 53.265 3.689 ;
      RECT 53.245 3.243 53.25 3.698 ;
      RECT 53.18 3.288 53.245 3.708 ;
      RECT 53.145 3.347 53.18 3.721 ;
      RECT 53.14 3.37 53.145 3.727 ;
      RECT 53.135 3.377 53.14 3.729 ;
      RECT 53.12 3.387 53.135 3.732 ;
      RECT 53.09 3.412 53.12 3.736 ;
      RECT 53.085 3.43 53.09 3.74 ;
      RECT 53.08 3.437 53.085 3.741 ;
      RECT 53.06 3.445 53.08 3.745 ;
      RECT 53.05 3.452 53.06 3.749 ;
      RECT 53.006 3.463 53.05 3.756 ;
      RECT 52.92 3.491 53.006 3.772 ;
      RECT 52.86 3.515 52.92 3.79 ;
      RECT 52.815 3.525 52.86 3.804 ;
      RECT 52.756 3.533 52.815 3.818 ;
      RECT 52.67 3.54 52.756 3.837 ;
      RECT 52.645 3.545 52.67 3.852 ;
      RECT 52.565 3.548 52.645 3.855 ;
      RECT 52.485 3.552 52.565 3.842 ;
      RECT 52.476 3.555 52.485 3.827 ;
      RECT 52.39 3.555 52.476 3.812 ;
      RECT 52.33 3.557 52.39 3.789 ;
      RECT 52.326 3.56 52.33 3.779 ;
      RECT 52.24 3.56 52.326 3.764 ;
      RECT 52.165 3.56 52.24 3.74 ;
      RECT 53.48 2.569 53.49 2.745 ;
      RECT 53.435 2.536 53.48 2.745 ;
      RECT 53.39 2.487 53.435 2.745 ;
      RECT 53.36 2.457 53.39 2.746 ;
      RECT 53.355 2.44 53.36 2.747 ;
      RECT 53.33 2.42 53.355 2.748 ;
      RECT 53.315 2.395 53.33 2.749 ;
      RECT 53.31 2.382 53.315 2.75 ;
      RECT 53.305 2.376 53.31 2.748 ;
      RECT 53.3 2.368 53.305 2.742 ;
      RECT 53.275 2.36 53.3 2.722 ;
      RECT 53.255 2.349 53.275 2.693 ;
      RECT 53.225 2.334 53.255 2.664 ;
      RECT 53.205 2.32 53.225 2.636 ;
      RECT 53.195 2.314 53.205 2.615 ;
      RECT 53.19 2.311 53.195 2.598 ;
      RECT 53.185 2.308 53.19 2.583 ;
      RECT 53.17 2.303 53.185 2.548 ;
      RECT 53.165 2.299 53.17 2.515 ;
      RECT 53.145 2.294 53.165 2.491 ;
      RECT 53.115 2.286 53.145 2.456 ;
      RECT 53.1 2.28 53.115 2.433 ;
      RECT 53.06 2.273 53.1 2.418 ;
      RECT 53.035 2.265 53.06 2.398 ;
      RECT 53.015 2.26 53.035 2.388 ;
      RECT 52.98 2.254 53.015 2.383 ;
      RECT 52.935 2.245 52.98 2.382 ;
      RECT 52.905 2.241 52.935 2.384 ;
      RECT 52.82 2.249 52.905 2.388 ;
      RECT 52.75 2.26 52.82 2.41 ;
      RECT 52.737 2.266 52.75 2.433 ;
      RECT 52.651 2.273 52.737 2.455 ;
      RECT 52.565 2.285 52.651 2.492 ;
      RECT 52.565 2.662 52.575 2.9 ;
      RECT 52.56 2.291 52.565 2.515 ;
      RECT 52.555 2.547 52.565 2.9 ;
      RECT 52.555 2.292 52.56 2.52 ;
      RECT 52.55 2.293 52.555 2.9 ;
      RECT 52.526 2.295 52.55 2.901 ;
      RECT 52.44 2.303 52.526 2.903 ;
      RECT 52.42 2.317 52.44 2.906 ;
      RECT 52.415 2.345 52.42 2.907 ;
      RECT 52.41 2.357 52.415 2.908 ;
      RECT 52.405 2.372 52.41 2.909 ;
      RECT 52.395 2.402 52.405 2.91 ;
      RECT 52.39 2.44 52.395 2.908 ;
      RECT 52.385 2.46 52.39 2.903 ;
      RECT 52.37 2.495 52.385 2.888 ;
      RECT 52.36 2.547 52.37 2.868 ;
      RECT 52.355 2.577 52.36 2.856 ;
      RECT 52.34 2.59 52.355 2.839 ;
      RECT 52.315 2.594 52.34 2.806 ;
      RECT 52.3 2.592 52.315 2.783 ;
      RECT 52.285 2.591 52.3 2.78 ;
      RECT 52.225 2.589 52.285 2.778 ;
      RECT 52.215 2.587 52.225 2.773 ;
      RECT 52.175 2.586 52.215 2.77 ;
      RECT 52.105 2.583 52.175 2.768 ;
      RECT 52.05 2.581 52.105 2.763 ;
      RECT 51.98 2.575 52.05 2.758 ;
      RECT 51.971 2.575 51.98 2.755 ;
      RECT 51.885 2.575 51.971 2.75 ;
      RECT 51.88 2.575 51.885 2.745 ;
      RECT 53.185 1.81 53.36 2.16 ;
      RECT 53.185 1.825 53.37 2.158 ;
      RECT 53.16 1.775 53.305 2.155 ;
      RECT 53.14 1.776 53.305 2.148 ;
      RECT 53.13 1.777 53.315 2.143 ;
      RECT 53.1 1.778 53.315 2.13 ;
      RECT 53.05 1.779 53.315 2.106 ;
      RECT 53.045 1.781 53.315 2.091 ;
      RECT 53.045 1.847 53.375 2.085 ;
      RECT 53.025 1.788 53.33 2.065 ;
      RECT 53.015 1.797 53.34 1.92 ;
      RECT 53.025 1.792 53.34 2.065 ;
      RECT 53.045 1.782 53.33 2.091 ;
      RECT 52.63 3.107 52.8 3.395 ;
      RECT 52.625 3.125 52.81 3.39 ;
      RECT 52.59 3.133 52.875 3.31 ;
      RECT 52.59 3.133 52.961 3.3 ;
      RECT 52.59 3.133 53.015 3.246 ;
      RECT 52.875 3.03 53.045 3.214 ;
      RECT 52.59 3.185 53.05 3.202 ;
      RECT 52.575 3.155 53.045 3.198 ;
      RECT 52.835 3.037 52.875 3.349 ;
      RECT 52.715 3.074 53.045 3.214 ;
      RECT 52.81 3.049 52.835 3.375 ;
      RECT 52.8 3.056 53.045 3.214 ;
      RECT 52.931 2.52 53 2.779 ;
      RECT 52.931 2.575 53.005 2.778 ;
      RECT 52.845 2.575 53.005 2.777 ;
      RECT 52.84 2.575 53.01 2.77 ;
      RECT 52.83 2.52 53 2.765 ;
      RECT 52.21 1.819 52.385 2.12 ;
      RECT 52.195 1.807 52.21 2.105 ;
      RECT 52.165 1.806 52.195 2.058 ;
      RECT 52.165 1.824 52.39 2.053 ;
      RECT 52.15 1.808 52.21 2.018 ;
      RECT 52.145 1.83 52.4 1.918 ;
      RECT 52.145 1.813 52.296 1.918 ;
      RECT 52.145 1.815 52.3 1.918 ;
      RECT 52.15 1.811 52.296 2.018 ;
      RECT 52.255 3.047 52.26 3.395 ;
      RECT 52.245 3.037 52.255 3.401 ;
      RECT 52.21 3.027 52.245 3.403 ;
      RECT 52.172 3.022 52.21 3.407 ;
      RECT 52.086 3.015 52.172 3.414 ;
      RECT 52 3.005 52.086 3.424 ;
      RECT 51.955 3 52 3.432 ;
      RECT 51.951 3 51.955 3.436 ;
      RECT 51.865 3 51.951 3.443 ;
      RECT 51.85 3 51.865 3.443 ;
      RECT 51.84 2.998 51.85 3.415 ;
      RECT 51.83 2.994 51.84 3.358 ;
      RECT 51.81 2.988 51.83 3.29 ;
      RECT 51.805 2.984 51.81 3.238 ;
      RECT 51.795 2.983 51.805 3.205 ;
      RECT 51.745 2.981 51.795 3.19 ;
      RECT 51.72 2.979 51.745 3.185 ;
      RECT 51.677 2.977 51.72 3.181 ;
      RECT 51.591 2.973 51.677 3.169 ;
      RECT 51.505 2.968 51.591 3.153 ;
      RECT 51.475 2.965 51.505 3.14 ;
      RECT 51.45 2.964 51.475 3.128 ;
      RECT 51.445 2.964 51.45 3.118 ;
      RECT 51.405 2.963 51.445 3.11 ;
      RECT 51.39 2.962 51.405 3.103 ;
      RECT 51.34 2.961 51.39 3.095 ;
      RECT 51.338 2.96 51.34 3.09 ;
      RECT 51.252 2.958 51.338 3.09 ;
      RECT 51.166 2.953 51.252 3.09 ;
      RECT 51.08 2.949 51.166 3.09 ;
      RECT 51.031 2.945 51.08 3.088 ;
      RECT 50.945 2.942 51.031 3.083 ;
      RECT 50.922 2.939 50.945 3.079 ;
      RECT 50.836 2.936 50.922 3.074 ;
      RECT 50.75 2.932 50.836 3.065 ;
      RECT 50.725 2.925 50.75 3.06 ;
      RECT 50.665 2.89 50.725 3.057 ;
      RECT 50.645 2.815 50.665 3.054 ;
      RECT 50.64 2.757 50.645 3.053 ;
      RECT 50.615 2.697 50.64 3.052 ;
      RECT 50.54 2.575 50.615 3.048 ;
      RECT 50.53 2.575 50.54 3.04 ;
      RECT 50.515 2.575 50.53 3.03 ;
      RECT 50.5 2.575 50.515 3 ;
      RECT 50.485 2.575 50.5 2.945 ;
      RECT 50.47 2.575 50.485 2.883 ;
      RECT 50.445 2.575 50.47 2.808 ;
      RECT 50.44 2.575 50.445 2.758 ;
      RECT 51.785 2.12 51.805 2.429 ;
      RECT 51.771 2.122 51.82 2.426 ;
      RECT 51.771 2.127 51.84 2.417 ;
      RECT 51.685 2.125 51.82 2.411 ;
      RECT 51.685 2.133 51.875 2.394 ;
      RECT 51.65 2.135 51.875 2.393 ;
      RECT 51.62 2.143 51.875 2.384 ;
      RECT 51.61 2.148 51.895 2.37 ;
      RECT 51.65 2.138 51.895 2.37 ;
      RECT 51.65 2.141 51.905 2.358 ;
      RECT 51.62 2.143 51.915 2.345 ;
      RECT 51.62 2.147 51.925 2.288 ;
      RECT 51.61 2.152 51.93 2.203 ;
      RECT 51.771 2.12 51.805 2.426 ;
      RECT 51.65 7.855 51.82 8.305 ;
      RECT 51.705 6.075 51.875 8.025 ;
      RECT 51.65 5.015 51.82 6.245 ;
      RECT 51.21 2.223 51.215 2.435 ;
      RECT 51.085 2.22 51.1 2.435 ;
      RECT 50.55 2.25 50.62 2.435 ;
      RECT 50.435 2.25 50.47 2.43 ;
      RECT 51.556 2.552 51.575 2.746 ;
      RECT 51.47 2.507 51.556 2.747 ;
      RECT 51.46 2.46 51.47 2.749 ;
      RECT 51.455 2.44 51.46 2.75 ;
      RECT 51.435 2.405 51.455 2.751 ;
      RECT 51.42 2.355 51.435 2.752 ;
      RECT 51.4 2.292 51.42 2.753 ;
      RECT 51.39 2.255 51.4 2.754 ;
      RECT 51.375 2.244 51.39 2.755 ;
      RECT 51.37 2.236 51.375 2.753 ;
      RECT 51.36 2.235 51.37 2.745 ;
      RECT 51.33 2.232 51.36 2.724 ;
      RECT 51.255 2.227 51.33 2.669 ;
      RECT 51.24 2.223 51.255 2.615 ;
      RECT 51.23 2.223 51.24 2.51 ;
      RECT 51.215 2.223 51.23 2.443 ;
      RECT 51.2 2.223 51.21 2.433 ;
      RECT 51.145 2.222 51.2 2.43 ;
      RECT 51.1 2.22 51.145 2.433 ;
      RECT 51.072 2.22 51.085 2.436 ;
      RECT 50.986 2.224 51.072 2.438 ;
      RECT 50.9 2.23 50.986 2.443 ;
      RECT 50.88 2.234 50.9 2.445 ;
      RECT 50.878 2.235 50.88 2.444 ;
      RECT 50.792 2.237 50.878 2.443 ;
      RECT 50.706 2.242 50.792 2.44 ;
      RECT 50.62 2.247 50.706 2.437 ;
      RECT 50.47 2.25 50.55 2.433 ;
      RECT 51.13 5.015 51.3 8.305 ;
      RECT 51.13 7.315 51.535 7.645 ;
      RECT 51.13 6.475 51.535 6.805 ;
      RECT 51.246 3.225 51.295 3.559 ;
      RECT 51.246 3.225 51.3 3.558 ;
      RECT 51.16 3.225 51.3 3.557 ;
      RECT 50.935 3.333 51.305 3.555 ;
      RECT 51.16 3.225 51.33 3.548 ;
      RECT 51.13 3.237 51.335 3.539 ;
      RECT 51.115 3.255 51.34 3.536 ;
      RECT 50.93 3.339 51.34 3.463 ;
      RECT 50.925 3.346 51.34 3.423 ;
      RECT 50.94 3.312 51.34 3.536 ;
      RECT 51.101 3.258 51.305 3.555 ;
      RECT 51.015 3.278 51.34 3.536 ;
      RECT 51.115 3.252 51.335 3.539 ;
      RECT 50.885 2.576 51.075 2.77 ;
      RECT 50.88 2.578 51.075 2.769 ;
      RECT 50.875 2.582 51.09 2.766 ;
      RECT 50.89 2.575 51.09 2.766 ;
      RECT 50.875 2.685 51.095 2.761 ;
      RECT 50.17 3.185 50.261 3.483 ;
      RECT 50.165 3.187 50.34 3.478 ;
      RECT 50.17 3.185 50.34 3.478 ;
      RECT 50.165 3.191 50.36 3.476 ;
      RECT 50.165 3.246 50.4 3.475 ;
      RECT 50.165 3.281 50.415 3.469 ;
      RECT 50.165 3.315 50.425 3.459 ;
      RECT 50.155 3.195 50.36 3.31 ;
      RECT 50.155 3.215 50.375 3.31 ;
      RECT 50.155 3.198 50.365 3.31 ;
      RECT 50.38 1.966 50.385 2.028 ;
      RECT 50.375 1.888 50.38 2.051 ;
      RECT 50.37 1.845 50.375 2.062 ;
      RECT 50.365 1.835 50.37 2.074 ;
      RECT 50.36 1.835 50.365 2.083 ;
      RECT 50.335 1.835 50.36 2.115 ;
      RECT 50.33 1.835 50.335 2.148 ;
      RECT 50.315 1.835 50.33 2.173 ;
      RECT 50.305 1.835 50.315 2.2 ;
      RECT 50.3 1.835 50.305 2.213 ;
      RECT 50.295 1.835 50.3 2.228 ;
      RECT 50.285 1.835 50.295 2.243 ;
      RECT 50.28 1.835 50.285 2.263 ;
      RECT 50.255 1.835 50.28 2.298 ;
      RECT 50.21 1.835 50.255 2.343 ;
      RECT 50.2 1.835 50.21 2.356 ;
      RECT 50.115 1.92 50.2 2.363 ;
      RECT 50.08 2.042 50.115 2.372 ;
      RECT 50.075 2.082 50.08 2.376 ;
      RECT 50.055 2.105 50.075 2.378 ;
      RECT 50.05 2.135 50.055 2.381 ;
      RECT 50.04 2.147 50.05 2.382 ;
      RECT 49.995 2.17 50.04 2.387 ;
      RECT 49.955 2.2 49.995 2.395 ;
      RECT 49.92 2.212 49.955 2.401 ;
      RECT 49.915 2.217 49.92 2.405 ;
      RECT 49.845 2.227 49.915 2.412 ;
      RECT 49.805 2.237 49.845 2.422 ;
      RECT 49.785 2.242 49.805 2.428 ;
      RECT 49.775 2.246 49.785 2.433 ;
      RECT 49.77 2.249 49.775 2.436 ;
      RECT 49.76 2.25 49.77 2.437 ;
      RECT 49.735 2.252 49.76 2.441 ;
      RECT 49.725 2.257 49.735 2.444 ;
      RECT 49.68 2.265 49.725 2.445 ;
      RECT 49.555 2.27 49.68 2.445 ;
      RECT 50.11 2.567 50.13 2.749 ;
      RECT 50.061 2.552 50.11 2.748 ;
      RECT 49.975 2.567 50.13 2.746 ;
      RECT 49.96 2.567 50.13 2.745 ;
      RECT 49.925 2.545 50.095 2.73 ;
      RECT 49.995 3.565 50.01 3.774 ;
      RECT 49.995 3.573 50.015 3.773 ;
      RECT 49.94 3.573 50.015 3.772 ;
      RECT 49.92 3.577 50.02 3.77 ;
      RECT 49.9 3.527 49.94 3.769 ;
      RECT 49.845 3.585 50.025 3.767 ;
      RECT 49.81 3.542 49.94 3.765 ;
      RECT 49.806 3.545 49.995 3.764 ;
      RECT 49.72 3.553 49.995 3.762 ;
      RECT 49.72 3.597 50.03 3.755 ;
      RECT 49.71 3.69 50.03 3.753 ;
      RECT 49.72 3.609 50.035 3.738 ;
      RECT 49.72 3.63 50.05 3.708 ;
      RECT 49.72 3.657 50.055 3.678 ;
      RECT 49.845 3.535 49.94 3.767 ;
      RECT 49.475 2.58 49.48 3.118 ;
      RECT 49.28 2.91 49.285 3.105 ;
      RECT 47.58 2.575 47.595 2.955 ;
      RECT 49.645 2.575 49.65 2.745 ;
      RECT 49.64 2.575 49.645 2.755 ;
      RECT 49.635 2.575 49.64 2.768 ;
      RECT 49.61 2.575 49.635 2.81 ;
      RECT 49.585 2.575 49.61 2.883 ;
      RECT 49.57 2.575 49.585 2.935 ;
      RECT 49.565 2.575 49.57 2.965 ;
      RECT 49.54 2.575 49.565 3.005 ;
      RECT 49.525 2.575 49.54 3.06 ;
      RECT 49.52 2.575 49.525 3.093 ;
      RECT 49.495 2.575 49.52 3.113 ;
      RECT 49.48 2.575 49.495 3.119 ;
      RECT 49.41 2.61 49.475 3.115 ;
      RECT 49.36 2.665 49.41 3.11 ;
      RECT 49.35 2.697 49.36 3.108 ;
      RECT 49.345 2.722 49.35 3.108 ;
      RECT 49.325 2.795 49.345 3.108 ;
      RECT 49.315 2.875 49.325 3.107 ;
      RECT 49.3 2.905 49.315 3.107 ;
      RECT 49.285 2.91 49.3 3.106 ;
      RECT 49.225 2.912 49.28 3.103 ;
      RECT 49.195 2.917 49.225 3.099 ;
      RECT 49.193 2.92 49.195 3.098 ;
      RECT 49.107 2.922 49.193 3.095 ;
      RECT 49.021 2.928 49.107 3.089 ;
      RECT 48.935 2.933 49.021 3.083 ;
      RECT 48.862 2.938 48.935 3.084 ;
      RECT 48.776 2.944 48.862 3.092 ;
      RECT 48.69 2.95 48.776 3.101 ;
      RECT 48.67 2.954 48.69 3.106 ;
      RECT 48.623 2.956 48.67 3.109 ;
      RECT 48.537 2.961 48.623 3.115 ;
      RECT 48.451 2.966 48.537 3.124 ;
      RECT 48.365 2.972 48.451 3.132 ;
      RECT 48.28 2.97 48.365 3.141 ;
      RECT 48.276 2.965 48.28 3.145 ;
      RECT 48.19 2.96 48.276 3.137 ;
      RECT 48.126 2.951 48.19 3.125 ;
      RECT 48.04 2.942 48.126 3.112 ;
      RECT 48.016 2.935 48.04 3.103 ;
      RECT 47.93 2.929 48.016 3.09 ;
      RECT 47.89 2.922 47.93 3.076 ;
      RECT 47.885 2.912 47.89 3.072 ;
      RECT 47.875 2.9 47.885 3.071 ;
      RECT 47.855 2.87 47.875 3.068 ;
      RECT 47.8 2.79 47.855 3.062 ;
      RECT 47.78 2.709 47.8 3.057 ;
      RECT 47.76 2.667 47.78 3.053 ;
      RECT 47.735 2.62 47.76 3.047 ;
      RECT 47.73 2.595 47.735 3.044 ;
      RECT 47.695 2.575 47.73 3.039 ;
      RECT 47.686 2.575 47.695 3.032 ;
      RECT 47.6 2.575 47.686 3.002 ;
      RECT 47.595 2.575 47.6 2.965 ;
      RECT 47.56 2.575 47.58 2.887 ;
      RECT 47.555 2.617 47.56 2.852 ;
      RECT 47.55 2.692 47.555 2.808 ;
      RECT 49 2.497 49.175 2.745 ;
      RECT 49 2.497 49.18 2.743 ;
      RECT 48.995 2.529 49.18 2.703 ;
      RECT 49.025 2.47 49.195 2.69 ;
      RECT 48.99 2.547 49.195 2.623 ;
      RECT 48.3 2.01 48.47 2.185 ;
      RECT 48.3 2.01 48.642 2.177 ;
      RECT 48.3 2.01 48.725 2.171 ;
      RECT 48.3 2.01 48.76 2.167 ;
      RECT 48.3 2.01 48.78 2.166 ;
      RECT 48.3 2.01 48.866 2.162 ;
      RECT 48.76 1.835 48.93 2.157 ;
      RECT 48.335 1.942 48.96 2.155 ;
      RECT 48.325 1.997 48.965 2.153 ;
      RECT 48.3 2.033 48.975 2.148 ;
      RECT 48.3 2.06 48.98 2.078 ;
      RECT 48.365 1.885 48.94 2.155 ;
      RECT 48.556 1.87 48.94 2.155 ;
      RECT 48.39 1.873 48.94 2.155 ;
      RECT 48.47 1.871 48.556 2.182 ;
      RECT 48.556 1.868 48.935 2.155 ;
      RECT 48.74 1.845 48.935 2.155 ;
      RECT 48.642 1.866 48.935 2.155 ;
      RECT 48.725 1.86 48.74 2.168 ;
      RECT 48.875 3.225 48.88 3.425 ;
      RECT 48.34 3.29 48.385 3.425 ;
      RECT 48.91 3.225 48.93 3.398 ;
      RECT 48.88 3.225 48.91 3.413 ;
      RECT 48.815 3.225 48.875 3.45 ;
      RECT 48.8 3.225 48.815 3.48 ;
      RECT 48.785 3.225 48.8 3.493 ;
      RECT 48.765 3.225 48.785 3.508 ;
      RECT 48.76 3.225 48.765 3.517 ;
      RECT 48.75 3.229 48.76 3.522 ;
      RECT 48.735 3.239 48.75 3.533 ;
      RECT 48.71 3.255 48.735 3.543 ;
      RECT 48.7 3.269 48.71 3.545 ;
      RECT 48.68 3.281 48.7 3.542 ;
      RECT 48.65 3.302 48.68 3.536 ;
      RECT 48.64 3.314 48.65 3.531 ;
      RECT 48.63 3.312 48.64 3.528 ;
      RECT 48.615 3.311 48.63 3.523 ;
      RECT 48.61 3.31 48.615 3.518 ;
      RECT 48.575 3.308 48.61 3.508 ;
      RECT 48.555 3.305 48.575 3.49 ;
      RECT 48.545 3.303 48.555 3.485 ;
      RECT 48.535 3.302 48.545 3.48 ;
      RECT 48.5 3.3 48.535 3.468 ;
      RECT 48.445 3.296 48.5 3.448 ;
      RECT 48.435 3.294 48.445 3.433 ;
      RECT 48.43 3.294 48.435 3.428 ;
      RECT 48.385 3.292 48.43 3.425 ;
      RECT 48.29 3.29 48.34 3.429 ;
      RECT 48.28 3.291 48.29 3.434 ;
      RECT 48.22 3.298 48.28 3.448 ;
      RECT 48.195 3.306 48.22 3.468 ;
      RECT 48.185 3.31 48.195 3.48 ;
      RECT 48.18 3.311 48.185 3.485 ;
      RECT 48.165 3.313 48.18 3.488 ;
      RECT 48.15 3.315 48.165 3.493 ;
      RECT 48.145 3.315 48.15 3.496 ;
      RECT 48.1 3.32 48.145 3.507 ;
      RECT 48.095 3.324 48.1 3.519 ;
      RECT 48.07 3.32 48.095 3.523 ;
      RECT 48.06 3.316 48.07 3.527 ;
      RECT 48.05 3.315 48.06 3.531 ;
      RECT 48.035 3.305 48.05 3.537 ;
      RECT 48.03 3.293 48.035 3.541 ;
      RECT 48.025 3.29 48.03 3.542 ;
      RECT 48.02 3.287 48.025 3.544 ;
      RECT 48.005 3.275 48.02 3.543 ;
      RECT 47.99 3.257 48.005 3.54 ;
      RECT 47.97 3.236 47.99 3.533 ;
      RECT 47.905 3.225 47.97 3.505 ;
      RECT 47.901 3.225 47.905 3.484 ;
      RECT 47.815 3.225 47.901 3.454 ;
      RECT 47.8 3.225 47.815 3.41 ;
      RECT 48.375 2.325 48.38 2.56 ;
      RECT 47.505 2.241 47.51 2.445 ;
      RECT 48.085 2.27 48.09 2.425 ;
      RECT 48.005 2.25 48.01 2.425 ;
      RECT 48.675 2.392 48.69 2.745 ;
      RECT 48.601 2.377 48.675 2.745 ;
      RECT 48.515 2.36 48.601 2.745 ;
      RECT 48.505 2.35 48.515 2.743 ;
      RECT 48.5 2.348 48.505 2.738 ;
      RECT 48.485 2.346 48.5 2.724 ;
      RECT 48.415 2.338 48.485 2.664 ;
      RECT 48.395 2.329 48.415 2.598 ;
      RECT 48.39 2.326 48.395 2.578 ;
      RECT 48.38 2.325 48.39 2.568 ;
      RECT 48.37 2.325 48.375 2.552 ;
      RECT 48.36 2.324 48.37 2.542 ;
      RECT 48.35 2.322 48.36 2.53 ;
      RECT 48.335 2.319 48.35 2.51 ;
      RECT 48.325 2.317 48.335 2.495 ;
      RECT 48.305 2.314 48.325 2.483 ;
      RECT 48.3 2.312 48.305 2.473 ;
      RECT 48.275 2.31 48.3 2.46 ;
      RECT 48.245 2.305 48.275 2.445 ;
      RECT 48.165 2.296 48.245 2.436 ;
      RECT 48.12 2.285 48.165 2.429 ;
      RECT 48.1 2.276 48.12 2.426 ;
      RECT 48.09 2.271 48.1 2.425 ;
      RECT 48.045 2.265 48.085 2.425 ;
      RECT 48.03 2.257 48.045 2.425 ;
      RECT 48.01 2.252 48.03 2.425 ;
      RECT 47.99 2.249 48.005 2.425 ;
      RECT 47.907 2.248 47.99 2.424 ;
      RECT 47.821 2.247 47.907 2.42 ;
      RECT 47.735 2.245 47.821 2.417 ;
      RECT 47.682 2.244 47.735 2.419 ;
      RECT 47.596 2.243 47.682 2.428 ;
      RECT 47.51 2.242 47.596 2.44 ;
      RECT 47.49 2.241 47.505 2.448 ;
      RECT 47.41 2.24 47.49 2.46 ;
      RECT 47.385 2.24 47.41 2.473 ;
      RECT 47.36 2.24 47.385 2.488 ;
      RECT 47.355 2.24 47.36 2.51 ;
      RECT 47.35 2.24 47.355 2.528 ;
      RECT 47.345 2.24 47.35 2.545 ;
      RECT 47.34 2.24 47.345 2.558 ;
      RECT 47.335 2.24 47.34 2.568 ;
      RECT 47.295 2.24 47.335 2.653 ;
      RECT 47.28 2.24 47.295 2.738 ;
      RECT 47.27 2.241 47.28 2.75 ;
      RECT 47.235 2.246 47.27 2.755 ;
      RECT 47.195 2.255 47.235 2.755 ;
      RECT 47.18 2.265 47.195 2.755 ;
      RECT 47.175 2.275 47.18 2.755 ;
      RECT 47.155 2.302 47.175 2.755 ;
      RECT 47.105 2.385 47.155 2.755 ;
      RECT 47.1 2.447 47.105 2.755 ;
      RECT 47.09 2.46 47.1 2.755 ;
      RECT 47.08 2.482 47.09 2.755 ;
      RECT 47.07 2.507 47.08 2.75 ;
      RECT 47.065 2.545 47.07 2.743 ;
      RECT 47.055 2.655 47.065 2.738 ;
      RECT 48.45 3.576 48.465 3.835 ;
      RECT 48.45 3.591 48.47 3.834 ;
      RECT 48.366 3.591 48.47 3.832 ;
      RECT 48.366 3.605 48.475 3.831 ;
      RECT 48.28 3.647 48.48 3.828 ;
      RECT 48.275 3.59 48.465 3.823 ;
      RECT 48.275 3.661 48.485 3.82 ;
      RECT 48.27 3.692 48.485 3.818 ;
      RECT 48.275 3.689 48.5 3.808 ;
      RECT 48.27 3.735 48.515 3.793 ;
      RECT 48.27 3.763 48.52 3.778 ;
      RECT 48.28 3.565 48.45 3.828 ;
      RECT 48.04 2.575 48.21 2.745 ;
      RECT 48.005 2.575 48.21 2.74 ;
      RECT 47.995 2.575 48.21 2.733 ;
      RECT 47.99 2.56 48.16 2.73 ;
      RECT 46.82 3.097 47.085 3.54 ;
      RECT 46.815 3.068 47.03 3.538 ;
      RECT 46.81 3.222 47.09 3.533 ;
      RECT 46.815 3.117 47.09 3.533 ;
      RECT 46.815 3.128 47.1 3.52 ;
      RECT 46.815 3.075 47.06 3.538 ;
      RECT 46.82 3.062 47.03 3.54 ;
      RECT 46.82 3.06 46.98 3.54 ;
      RECT 46.921 3.052 46.98 3.54 ;
      RECT 46.835 3.053 46.98 3.54 ;
      RECT 46.921 3.051 46.97 3.54 ;
      RECT 46.725 1.866 46.9 2.165 ;
      RECT 46.775 1.828 46.9 2.165 ;
      RECT 46.76 1.83 46.986 2.157 ;
      RECT 46.76 1.833 47.025 2.144 ;
      RECT 46.76 1.834 47.035 2.13 ;
      RECT 46.715 1.885 47.035 2.12 ;
      RECT 46.76 1.835 47.04 2.115 ;
      RECT 46.715 2.045 47.045 2.105 ;
      RECT 46.7 1.905 47.04 2.045 ;
      RECT 46.695 1.921 47.04 1.985 ;
      RECT 46.74 1.845 47.04 2.115 ;
      RECT 46.775 1.826 46.861 2.165 ;
      RECT 44.87 1.74 45.04 2.935 ;
      RECT 44.87 1.74 45.335 1.91 ;
      RECT 44.87 6.97 45.335 7.14 ;
      RECT 44.87 5.945 45.04 7.14 ;
      RECT 43.88 1.74 44.05 2.935 ;
      RECT 43.88 1.74 44.345 1.91 ;
      RECT 43.88 6.97 44.345 7.14 ;
      RECT 43.88 5.945 44.05 7.14 ;
      RECT 42.025 2.635 42.195 3.865 ;
      RECT 42.08 0.855 42.25 2.805 ;
      RECT 42.025 0.575 42.195 1.025 ;
      RECT 42.025 7.855 42.195 8.305 ;
      RECT 42.08 6.075 42.25 8.025 ;
      RECT 42.025 5.015 42.195 6.245 ;
      RECT 41.505 0.575 41.675 3.865 ;
      RECT 41.505 2.075 41.91 2.405 ;
      RECT 41.505 1.235 41.91 1.565 ;
      RECT 41.505 5.015 41.675 8.305 ;
      RECT 41.505 7.315 41.91 7.645 ;
      RECT 41.505 6.475 41.91 6.805 ;
      RECT 39.43 3.126 39.435 3.298 ;
      RECT 39.425 3.119 39.43 3.388 ;
      RECT 39.42 3.113 39.425 3.407 ;
      RECT 39.4 3.107 39.42 3.417 ;
      RECT 39.385 3.102 39.4 3.425 ;
      RECT 39.348 3.096 39.385 3.423 ;
      RECT 39.262 3.082 39.348 3.419 ;
      RECT 39.176 3.064 39.262 3.414 ;
      RECT 39.09 3.045 39.176 3.408 ;
      RECT 39.06 3.033 39.09 3.404 ;
      RECT 39.04 3.027 39.06 3.403 ;
      RECT 38.975 3.025 39.04 3.401 ;
      RECT 38.96 3.025 38.975 3.393 ;
      RECT 38.945 3.025 38.96 3.38 ;
      RECT 38.94 3.025 38.945 3.37 ;
      RECT 38.925 3.025 38.94 3.348 ;
      RECT 38.91 3.025 38.925 3.315 ;
      RECT 38.905 3.025 38.91 3.293 ;
      RECT 38.895 3.025 38.905 3.275 ;
      RECT 38.88 3.025 38.895 3.253 ;
      RECT 38.86 3.025 38.88 3.215 ;
      RECT 39.21 2.31 39.245 2.749 ;
      RECT 39.21 2.31 39.25 2.748 ;
      RECT 39.155 2.37 39.25 2.747 ;
      RECT 39.02 2.542 39.25 2.746 ;
      RECT 39.13 2.42 39.25 2.746 ;
      RECT 39.02 2.542 39.275 2.736 ;
      RECT 39.075 2.487 39.355 2.653 ;
      RECT 39.25 2.281 39.255 2.744 ;
      RECT 39.105 2.457 39.395 2.53 ;
      RECT 39.12 2.44 39.25 2.746 ;
      RECT 39.255 2.28 39.425 2.468 ;
      RECT 39.245 2.283 39.425 2.468 ;
      RECT 38.75 2.16 38.92 2.47 ;
      RECT 38.75 2.16 38.925 2.443 ;
      RECT 38.75 2.16 38.93 2.42 ;
      RECT 38.75 2.16 38.94 2.37 ;
      RECT 38.745 2.265 38.94 2.34 ;
      RECT 38.78 1.835 38.95 2.313 ;
      RECT 38.78 1.835 38.965 2.234 ;
      RECT 38.77 2.045 38.965 2.234 ;
      RECT 38.78 1.845 38.975 2.149 ;
      RECT 38.71 2.587 38.715 2.79 ;
      RECT 38.7 2.575 38.71 2.9 ;
      RECT 38.675 2.575 38.7 2.94 ;
      RECT 38.595 2.575 38.675 3.025 ;
      RECT 38.585 2.575 38.595 3.095 ;
      RECT 38.56 2.575 38.585 3.118 ;
      RECT 38.54 2.575 38.56 3.153 ;
      RECT 38.495 2.585 38.54 3.196 ;
      RECT 38.485 2.597 38.495 3.233 ;
      RECT 38.465 2.611 38.485 3.253 ;
      RECT 38.455 2.629 38.465 3.269 ;
      RECT 38.44 2.655 38.455 3.279 ;
      RECT 38.425 2.696 38.44 3.293 ;
      RECT 38.415 2.731 38.425 3.303 ;
      RECT 38.41 2.747 38.415 3.308 ;
      RECT 38.4 2.762 38.41 3.313 ;
      RECT 38.38 2.805 38.4 3.323 ;
      RECT 38.36 2.842 38.38 3.336 ;
      RECT 38.325 2.865 38.36 3.354 ;
      RECT 38.315 2.879 38.325 3.37 ;
      RECT 38.295 2.889 38.315 3.38 ;
      RECT 38.29 2.898 38.295 3.388 ;
      RECT 38.28 2.905 38.29 3.395 ;
      RECT 38.27 2.912 38.28 3.403 ;
      RECT 38.255 2.922 38.27 3.411 ;
      RECT 38.245 2.936 38.255 3.421 ;
      RECT 38.235 2.948 38.245 3.433 ;
      RECT 38.22 2.97 38.235 3.446 ;
      RECT 38.21 2.992 38.22 3.457 ;
      RECT 38.2 3.012 38.21 3.466 ;
      RECT 38.195 3.027 38.2 3.473 ;
      RECT 38.165 3.06 38.195 3.487 ;
      RECT 38.155 3.095 38.165 3.502 ;
      RECT 38.15 3.102 38.155 3.508 ;
      RECT 38.13 3.117 38.15 3.515 ;
      RECT 38.125 3.132 38.13 3.523 ;
      RECT 38.12 3.141 38.125 3.528 ;
      RECT 38.105 3.147 38.12 3.535 ;
      RECT 38.1 3.153 38.105 3.543 ;
      RECT 38.095 3.157 38.1 3.55 ;
      RECT 38.09 3.161 38.095 3.56 ;
      RECT 38.08 3.166 38.09 3.57 ;
      RECT 38.06 3.177 38.08 3.598 ;
      RECT 38.045 3.189 38.06 3.625 ;
      RECT 38.025 3.202 38.045 3.65 ;
      RECT 38.005 3.217 38.025 3.674 ;
      RECT 37.99 3.232 38.005 3.689 ;
      RECT 37.985 3.243 37.99 3.698 ;
      RECT 37.92 3.288 37.985 3.708 ;
      RECT 37.885 3.347 37.92 3.721 ;
      RECT 37.88 3.37 37.885 3.727 ;
      RECT 37.875 3.377 37.88 3.729 ;
      RECT 37.86 3.387 37.875 3.732 ;
      RECT 37.83 3.412 37.86 3.736 ;
      RECT 37.825 3.43 37.83 3.74 ;
      RECT 37.82 3.437 37.825 3.741 ;
      RECT 37.8 3.445 37.82 3.745 ;
      RECT 37.79 3.452 37.8 3.749 ;
      RECT 37.746 3.463 37.79 3.756 ;
      RECT 37.66 3.491 37.746 3.772 ;
      RECT 37.6 3.515 37.66 3.79 ;
      RECT 37.555 3.525 37.6 3.804 ;
      RECT 37.496 3.533 37.555 3.818 ;
      RECT 37.41 3.54 37.496 3.837 ;
      RECT 37.385 3.545 37.41 3.852 ;
      RECT 37.305 3.548 37.385 3.855 ;
      RECT 37.225 3.552 37.305 3.842 ;
      RECT 37.216 3.555 37.225 3.827 ;
      RECT 37.13 3.555 37.216 3.812 ;
      RECT 37.07 3.557 37.13 3.789 ;
      RECT 37.066 3.56 37.07 3.779 ;
      RECT 36.98 3.56 37.066 3.764 ;
      RECT 36.905 3.56 36.98 3.74 ;
      RECT 38.22 2.569 38.23 2.745 ;
      RECT 38.175 2.536 38.22 2.745 ;
      RECT 38.13 2.487 38.175 2.745 ;
      RECT 38.1 2.457 38.13 2.746 ;
      RECT 38.095 2.44 38.1 2.747 ;
      RECT 38.07 2.42 38.095 2.748 ;
      RECT 38.055 2.395 38.07 2.749 ;
      RECT 38.05 2.382 38.055 2.75 ;
      RECT 38.045 2.376 38.05 2.748 ;
      RECT 38.04 2.368 38.045 2.742 ;
      RECT 38.015 2.36 38.04 2.722 ;
      RECT 37.995 2.349 38.015 2.693 ;
      RECT 37.965 2.334 37.995 2.664 ;
      RECT 37.945 2.32 37.965 2.636 ;
      RECT 37.935 2.314 37.945 2.615 ;
      RECT 37.93 2.311 37.935 2.598 ;
      RECT 37.925 2.308 37.93 2.583 ;
      RECT 37.91 2.303 37.925 2.548 ;
      RECT 37.905 2.299 37.91 2.515 ;
      RECT 37.885 2.294 37.905 2.491 ;
      RECT 37.855 2.286 37.885 2.456 ;
      RECT 37.84 2.28 37.855 2.433 ;
      RECT 37.8 2.273 37.84 2.418 ;
      RECT 37.775 2.265 37.8 2.398 ;
      RECT 37.755 2.26 37.775 2.388 ;
      RECT 37.72 2.254 37.755 2.383 ;
      RECT 37.675 2.245 37.72 2.382 ;
      RECT 37.645 2.241 37.675 2.384 ;
      RECT 37.56 2.249 37.645 2.388 ;
      RECT 37.49 2.26 37.56 2.41 ;
      RECT 37.477 2.266 37.49 2.433 ;
      RECT 37.391 2.273 37.477 2.455 ;
      RECT 37.305 2.285 37.391 2.492 ;
      RECT 37.305 2.662 37.315 2.9 ;
      RECT 37.3 2.291 37.305 2.515 ;
      RECT 37.295 2.547 37.305 2.9 ;
      RECT 37.295 2.292 37.3 2.52 ;
      RECT 37.29 2.293 37.295 2.9 ;
      RECT 37.266 2.295 37.29 2.901 ;
      RECT 37.18 2.303 37.266 2.903 ;
      RECT 37.16 2.317 37.18 2.906 ;
      RECT 37.155 2.345 37.16 2.907 ;
      RECT 37.15 2.357 37.155 2.908 ;
      RECT 37.145 2.372 37.15 2.909 ;
      RECT 37.135 2.402 37.145 2.91 ;
      RECT 37.13 2.44 37.135 2.908 ;
      RECT 37.125 2.46 37.13 2.903 ;
      RECT 37.11 2.495 37.125 2.888 ;
      RECT 37.1 2.547 37.11 2.868 ;
      RECT 37.095 2.577 37.1 2.856 ;
      RECT 37.08 2.59 37.095 2.839 ;
      RECT 37.055 2.594 37.08 2.806 ;
      RECT 37.04 2.592 37.055 2.783 ;
      RECT 37.025 2.591 37.04 2.78 ;
      RECT 36.965 2.589 37.025 2.778 ;
      RECT 36.955 2.587 36.965 2.773 ;
      RECT 36.915 2.586 36.955 2.77 ;
      RECT 36.845 2.583 36.915 2.768 ;
      RECT 36.79 2.581 36.845 2.763 ;
      RECT 36.72 2.575 36.79 2.758 ;
      RECT 36.711 2.575 36.72 2.755 ;
      RECT 36.625 2.575 36.711 2.75 ;
      RECT 36.62 2.575 36.625 2.745 ;
      RECT 37.925 1.81 38.1 2.16 ;
      RECT 37.925 1.825 38.11 2.158 ;
      RECT 37.9 1.775 38.045 2.155 ;
      RECT 37.88 1.776 38.045 2.148 ;
      RECT 37.87 1.777 38.055 2.143 ;
      RECT 37.84 1.778 38.055 2.13 ;
      RECT 37.79 1.779 38.055 2.106 ;
      RECT 37.785 1.781 38.055 2.091 ;
      RECT 37.785 1.847 38.115 2.085 ;
      RECT 37.765 1.788 38.07 2.065 ;
      RECT 37.755 1.797 38.08 1.92 ;
      RECT 37.765 1.792 38.08 2.065 ;
      RECT 37.785 1.782 38.07 2.091 ;
      RECT 37.37 3.107 37.54 3.395 ;
      RECT 37.365 3.125 37.55 3.39 ;
      RECT 37.33 3.133 37.615 3.31 ;
      RECT 37.33 3.133 37.701 3.3 ;
      RECT 37.33 3.133 37.755 3.246 ;
      RECT 37.615 3.03 37.785 3.214 ;
      RECT 37.33 3.185 37.79 3.202 ;
      RECT 37.315 3.155 37.785 3.198 ;
      RECT 37.575 3.037 37.615 3.349 ;
      RECT 37.455 3.074 37.785 3.214 ;
      RECT 37.55 3.049 37.575 3.375 ;
      RECT 37.54 3.056 37.785 3.214 ;
      RECT 37.671 2.52 37.74 2.779 ;
      RECT 37.671 2.575 37.745 2.778 ;
      RECT 37.585 2.575 37.745 2.777 ;
      RECT 37.58 2.575 37.75 2.77 ;
      RECT 37.57 2.52 37.74 2.765 ;
      RECT 36.95 1.819 37.125 2.12 ;
      RECT 36.935 1.807 36.95 2.105 ;
      RECT 36.905 1.806 36.935 2.058 ;
      RECT 36.905 1.824 37.13 2.053 ;
      RECT 36.89 1.808 36.95 2.018 ;
      RECT 36.885 1.83 37.14 1.918 ;
      RECT 36.885 1.813 37.036 1.918 ;
      RECT 36.885 1.815 37.04 1.918 ;
      RECT 36.89 1.811 37.036 2.018 ;
      RECT 36.995 3.047 37 3.395 ;
      RECT 36.985 3.037 36.995 3.401 ;
      RECT 36.95 3.027 36.985 3.403 ;
      RECT 36.912 3.022 36.95 3.407 ;
      RECT 36.826 3.015 36.912 3.414 ;
      RECT 36.74 3.005 36.826 3.424 ;
      RECT 36.695 3 36.74 3.432 ;
      RECT 36.691 3 36.695 3.436 ;
      RECT 36.605 3 36.691 3.443 ;
      RECT 36.59 3 36.605 3.443 ;
      RECT 36.58 2.998 36.59 3.415 ;
      RECT 36.57 2.994 36.58 3.358 ;
      RECT 36.55 2.988 36.57 3.29 ;
      RECT 36.545 2.984 36.55 3.238 ;
      RECT 36.535 2.983 36.545 3.205 ;
      RECT 36.485 2.981 36.535 3.19 ;
      RECT 36.46 2.979 36.485 3.185 ;
      RECT 36.417 2.977 36.46 3.181 ;
      RECT 36.331 2.973 36.417 3.169 ;
      RECT 36.245 2.968 36.331 3.153 ;
      RECT 36.215 2.965 36.245 3.14 ;
      RECT 36.19 2.964 36.215 3.128 ;
      RECT 36.185 2.964 36.19 3.118 ;
      RECT 36.145 2.963 36.185 3.11 ;
      RECT 36.13 2.962 36.145 3.103 ;
      RECT 36.08 2.961 36.13 3.095 ;
      RECT 36.078 2.96 36.08 3.09 ;
      RECT 35.992 2.958 36.078 3.09 ;
      RECT 35.906 2.953 35.992 3.09 ;
      RECT 35.82 2.949 35.906 3.09 ;
      RECT 35.771 2.945 35.82 3.088 ;
      RECT 35.685 2.942 35.771 3.083 ;
      RECT 35.662 2.939 35.685 3.079 ;
      RECT 35.576 2.936 35.662 3.074 ;
      RECT 35.49 2.932 35.576 3.065 ;
      RECT 35.465 2.925 35.49 3.06 ;
      RECT 35.405 2.89 35.465 3.057 ;
      RECT 35.385 2.815 35.405 3.054 ;
      RECT 35.38 2.757 35.385 3.053 ;
      RECT 35.355 2.697 35.38 3.052 ;
      RECT 35.28 2.575 35.355 3.048 ;
      RECT 35.27 2.575 35.28 3.04 ;
      RECT 35.255 2.575 35.27 3.03 ;
      RECT 35.24 2.575 35.255 3 ;
      RECT 35.225 2.575 35.24 2.945 ;
      RECT 35.21 2.575 35.225 2.883 ;
      RECT 35.185 2.575 35.21 2.808 ;
      RECT 35.18 2.575 35.185 2.758 ;
      RECT 36.525 2.12 36.545 2.429 ;
      RECT 36.511 2.122 36.56 2.426 ;
      RECT 36.511 2.127 36.58 2.417 ;
      RECT 36.425 2.125 36.56 2.411 ;
      RECT 36.425 2.133 36.615 2.394 ;
      RECT 36.39 2.135 36.615 2.393 ;
      RECT 36.36 2.143 36.615 2.384 ;
      RECT 36.35 2.148 36.635 2.37 ;
      RECT 36.39 2.138 36.635 2.37 ;
      RECT 36.39 2.141 36.645 2.358 ;
      RECT 36.36 2.143 36.655 2.345 ;
      RECT 36.36 2.147 36.665 2.288 ;
      RECT 36.35 2.152 36.67 2.203 ;
      RECT 36.511 2.12 36.545 2.426 ;
      RECT 36.39 7.855 36.56 8.305 ;
      RECT 36.445 6.075 36.615 8.025 ;
      RECT 36.39 5.015 36.56 6.245 ;
      RECT 35.95 2.223 35.955 2.435 ;
      RECT 35.825 2.22 35.84 2.435 ;
      RECT 35.29 2.25 35.36 2.435 ;
      RECT 35.175 2.25 35.21 2.43 ;
      RECT 36.296 2.552 36.315 2.746 ;
      RECT 36.21 2.507 36.296 2.747 ;
      RECT 36.2 2.46 36.21 2.749 ;
      RECT 36.195 2.44 36.2 2.75 ;
      RECT 36.175 2.405 36.195 2.751 ;
      RECT 36.16 2.355 36.175 2.752 ;
      RECT 36.14 2.292 36.16 2.753 ;
      RECT 36.13 2.255 36.14 2.754 ;
      RECT 36.115 2.244 36.13 2.755 ;
      RECT 36.11 2.236 36.115 2.753 ;
      RECT 36.1 2.235 36.11 2.745 ;
      RECT 36.07 2.232 36.1 2.724 ;
      RECT 35.995 2.227 36.07 2.669 ;
      RECT 35.98 2.223 35.995 2.615 ;
      RECT 35.97 2.223 35.98 2.51 ;
      RECT 35.955 2.223 35.97 2.443 ;
      RECT 35.94 2.223 35.95 2.433 ;
      RECT 35.885 2.222 35.94 2.43 ;
      RECT 35.84 2.22 35.885 2.433 ;
      RECT 35.812 2.22 35.825 2.436 ;
      RECT 35.726 2.224 35.812 2.438 ;
      RECT 35.64 2.23 35.726 2.443 ;
      RECT 35.62 2.234 35.64 2.445 ;
      RECT 35.618 2.235 35.62 2.444 ;
      RECT 35.532 2.237 35.618 2.443 ;
      RECT 35.446 2.242 35.532 2.44 ;
      RECT 35.36 2.247 35.446 2.437 ;
      RECT 35.21 2.25 35.29 2.433 ;
      RECT 35.87 5.015 36.04 8.305 ;
      RECT 35.87 7.315 36.275 7.645 ;
      RECT 35.87 6.475 36.275 6.805 ;
      RECT 35.986 3.225 36.035 3.559 ;
      RECT 35.986 3.225 36.04 3.558 ;
      RECT 35.9 3.225 36.04 3.557 ;
      RECT 35.675 3.333 36.045 3.555 ;
      RECT 35.9 3.225 36.07 3.548 ;
      RECT 35.87 3.237 36.075 3.539 ;
      RECT 35.855 3.255 36.08 3.536 ;
      RECT 35.67 3.339 36.08 3.463 ;
      RECT 35.665 3.346 36.08 3.423 ;
      RECT 35.68 3.312 36.08 3.536 ;
      RECT 35.841 3.258 36.045 3.555 ;
      RECT 35.755 3.278 36.08 3.536 ;
      RECT 35.855 3.252 36.075 3.539 ;
      RECT 35.625 2.576 35.815 2.77 ;
      RECT 35.62 2.578 35.815 2.769 ;
      RECT 35.615 2.582 35.83 2.766 ;
      RECT 35.63 2.575 35.83 2.766 ;
      RECT 35.615 2.685 35.835 2.761 ;
      RECT 34.91 3.185 35.001 3.483 ;
      RECT 34.905 3.187 35.08 3.478 ;
      RECT 34.91 3.185 35.08 3.478 ;
      RECT 34.905 3.191 35.1 3.476 ;
      RECT 34.905 3.246 35.14 3.475 ;
      RECT 34.905 3.281 35.155 3.469 ;
      RECT 34.905 3.315 35.165 3.459 ;
      RECT 34.895 3.195 35.1 3.31 ;
      RECT 34.895 3.215 35.115 3.31 ;
      RECT 34.895 3.198 35.105 3.31 ;
      RECT 35.12 1.966 35.125 2.028 ;
      RECT 35.115 1.888 35.12 2.051 ;
      RECT 35.11 1.845 35.115 2.062 ;
      RECT 35.105 1.835 35.11 2.074 ;
      RECT 35.1 1.835 35.105 2.083 ;
      RECT 35.075 1.835 35.1 2.115 ;
      RECT 35.07 1.835 35.075 2.148 ;
      RECT 35.055 1.835 35.07 2.173 ;
      RECT 35.045 1.835 35.055 2.2 ;
      RECT 35.04 1.835 35.045 2.213 ;
      RECT 35.035 1.835 35.04 2.228 ;
      RECT 35.025 1.835 35.035 2.243 ;
      RECT 35.02 1.835 35.025 2.263 ;
      RECT 34.995 1.835 35.02 2.298 ;
      RECT 34.95 1.835 34.995 2.343 ;
      RECT 34.94 1.835 34.95 2.356 ;
      RECT 34.855 1.92 34.94 2.363 ;
      RECT 34.82 2.042 34.855 2.372 ;
      RECT 34.815 2.082 34.82 2.376 ;
      RECT 34.795 2.105 34.815 2.378 ;
      RECT 34.79 2.135 34.795 2.381 ;
      RECT 34.78 2.147 34.79 2.382 ;
      RECT 34.735 2.17 34.78 2.387 ;
      RECT 34.695 2.2 34.735 2.395 ;
      RECT 34.66 2.212 34.695 2.401 ;
      RECT 34.655 2.217 34.66 2.405 ;
      RECT 34.585 2.227 34.655 2.412 ;
      RECT 34.545 2.237 34.585 2.422 ;
      RECT 34.525 2.242 34.545 2.428 ;
      RECT 34.515 2.246 34.525 2.433 ;
      RECT 34.51 2.249 34.515 2.436 ;
      RECT 34.5 2.25 34.51 2.437 ;
      RECT 34.475 2.252 34.5 2.441 ;
      RECT 34.465 2.257 34.475 2.444 ;
      RECT 34.42 2.265 34.465 2.445 ;
      RECT 34.295 2.27 34.42 2.445 ;
      RECT 34.85 2.567 34.87 2.749 ;
      RECT 34.801 2.552 34.85 2.748 ;
      RECT 34.715 2.567 34.87 2.746 ;
      RECT 34.7 2.567 34.87 2.745 ;
      RECT 34.665 2.545 34.835 2.73 ;
      RECT 34.735 3.565 34.75 3.774 ;
      RECT 34.735 3.573 34.755 3.773 ;
      RECT 34.68 3.573 34.755 3.772 ;
      RECT 34.66 3.577 34.76 3.77 ;
      RECT 34.64 3.527 34.68 3.769 ;
      RECT 34.585 3.585 34.765 3.767 ;
      RECT 34.55 3.542 34.68 3.765 ;
      RECT 34.546 3.545 34.735 3.764 ;
      RECT 34.46 3.553 34.735 3.762 ;
      RECT 34.46 3.597 34.77 3.755 ;
      RECT 34.45 3.69 34.77 3.753 ;
      RECT 34.46 3.609 34.775 3.738 ;
      RECT 34.46 3.63 34.79 3.708 ;
      RECT 34.46 3.657 34.795 3.678 ;
      RECT 34.585 3.535 34.68 3.767 ;
      RECT 34.215 2.58 34.22 3.118 ;
      RECT 34.02 2.91 34.025 3.105 ;
      RECT 32.32 2.575 32.335 2.955 ;
      RECT 34.385 2.575 34.39 2.745 ;
      RECT 34.38 2.575 34.385 2.755 ;
      RECT 34.375 2.575 34.38 2.768 ;
      RECT 34.35 2.575 34.375 2.81 ;
      RECT 34.325 2.575 34.35 2.883 ;
      RECT 34.31 2.575 34.325 2.935 ;
      RECT 34.305 2.575 34.31 2.965 ;
      RECT 34.28 2.575 34.305 3.005 ;
      RECT 34.265 2.575 34.28 3.06 ;
      RECT 34.26 2.575 34.265 3.093 ;
      RECT 34.235 2.575 34.26 3.113 ;
      RECT 34.22 2.575 34.235 3.119 ;
      RECT 34.15 2.61 34.215 3.115 ;
      RECT 34.1 2.665 34.15 3.11 ;
      RECT 34.09 2.697 34.1 3.108 ;
      RECT 34.085 2.722 34.09 3.108 ;
      RECT 34.065 2.795 34.085 3.108 ;
      RECT 34.055 2.875 34.065 3.107 ;
      RECT 34.04 2.905 34.055 3.107 ;
      RECT 34.025 2.91 34.04 3.106 ;
      RECT 33.965 2.912 34.02 3.103 ;
      RECT 33.935 2.917 33.965 3.099 ;
      RECT 33.933 2.92 33.935 3.098 ;
      RECT 33.847 2.922 33.933 3.095 ;
      RECT 33.761 2.928 33.847 3.089 ;
      RECT 33.675 2.933 33.761 3.083 ;
      RECT 33.602 2.938 33.675 3.084 ;
      RECT 33.516 2.944 33.602 3.092 ;
      RECT 33.43 2.95 33.516 3.101 ;
      RECT 33.41 2.954 33.43 3.106 ;
      RECT 33.363 2.956 33.41 3.109 ;
      RECT 33.277 2.961 33.363 3.115 ;
      RECT 33.191 2.966 33.277 3.124 ;
      RECT 33.105 2.972 33.191 3.132 ;
      RECT 33.02 2.97 33.105 3.141 ;
      RECT 33.016 2.965 33.02 3.145 ;
      RECT 32.93 2.96 33.016 3.137 ;
      RECT 32.866 2.951 32.93 3.125 ;
      RECT 32.78 2.942 32.866 3.112 ;
      RECT 32.756 2.935 32.78 3.103 ;
      RECT 32.67 2.929 32.756 3.09 ;
      RECT 32.63 2.922 32.67 3.076 ;
      RECT 32.625 2.912 32.63 3.072 ;
      RECT 32.615 2.9 32.625 3.071 ;
      RECT 32.595 2.87 32.615 3.068 ;
      RECT 32.54 2.79 32.595 3.062 ;
      RECT 32.52 2.709 32.54 3.057 ;
      RECT 32.5 2.667 32.52 3.053 ;
      RECT 32.475 2.62 32.5 3.047 ;
      RECT 32.47 2.595 32.475 3.044 ;
      RECT 32.435 2.575 32.47 3.039 ;
      RECT 32.426 2.575 32.435 3.032 ;
      RECT 32.34 2.575 32.426 3.002 ;
      RECT 32.335 2.575 32.34 2.965 ;
      RECT 32.3 2.575 32.32 2.887 ;
      RECT 32.295 2.617 32.3 2.852 ;
      RECT 32.29 2.692 32.295 2.808 ;
      RECT 33.74 2.497 33.915 2.745 ;
      RECT 33.74 2.497 33.92 2.743 ;
      RECT 33.735 2.529 33.92 2.703 ;
      RECT 33.765 2.47 33.935 2.69 ;
      RECT 33.73 2.547 33.935 2.623 ;
      RECT 33.04 2.01 33.21 2.185 ;
      RECT 33.04 2.01 33.382 2.177 ;
      RECT 33.04 2.01 33.465 2.171 ;
      RECT 33.04 2.01 33.5 2.167 ;
      RECT 33.04 2.01 33.52 2.166 ;
      RECT 33.04 2.01 33.606 2.162 ;
      RECT 33.5 1.835 33.67 2.157 ;
      RECT 33.075 1.942 33.7 2.155 ;
      RECT 33.065 1.997 33.705 2.153 ;
      RECT 33.04 2.033 33.715 2.148 ;
      RECT 33.04 2.06 33.72 2.078 ;
      RECT 33.105 1.885 33.68 2.155 ;
      RECT 33.296 1.87 33.68 2.155 ;
      RECT 33.13 1.873 33.68 2.155 ;
      RECT 33.21 1.871 33.296 2.182 ;
      RECT 33.296 1.868 33.675 2.155 ;
      RECT 33.48 1.845 33.675 2.155 ;
      RECT 33.382 1.866 33.675 2.155 ;
      RECT 33.465 1.86 33.48 2.168 ;
      RECT 33.615 3.225 33.62 3.425 ;
      RECT 33.08 3.29 33.125 3.425 ;
      RECT 33.65 3.225 33.67 3.398 ;
      RECT 33.62 3.225 33.65 3.413 ;
      RECT 33.555 3.225 33.615 3.45 ;
      RECT 33.54 3.225 33.555 3.48 ;
      RECT 33.525 3.225 33.54 3.493 ;
      RECT 33.505 3.225 33.525 3.508 ;
      RECT 33.5 3.225 33.505 3.517 ;
      RECT 33.49 3.229 33.5 3.522 ;
      RECT 33.475 3.239 33.49 3.533 ;
      RECT 33.45 3.255 33.475 3.543 ;
      RECT 33.44 3.269 33.45 3.545 ;
      RECT 33.42 3.281 33.44 3.542 ;
      RECT 33.39 3.302 33.42 3.536 ;
      RECT 33.38 3.314 33.39 3.531 ;
      RECT 33.37 3.312 33.38 3.528 ;
      RECT 33.355 3.311 33.37 3.523 ;
      RECT 33.35 3.31 33.355 3.518 ;
      RECT 33.315 3.308 33.35 3.508 ;
      RECT 33.295 3.305 33.315 3.49 ;
      RECT 33.285 3.303 33.295 3.485 ;
      RECT 33.275 3.302 33.285 3.48 ;
      RECT 33.24 3.3 33.275 3.468 ;
      RECT 33.185 3.296 33.24 3.448 ;
      RECT 33.175 3.294 33.185 3.433 ;
      RECT 33.17 3.294 33.175 3.428 ;
      RECT 33.125 3.292 33.17 3.425 ;
      RECT 33.03 3.29 33.08 3.429 ;
      RECT 33.02 3.291 33.03 3.434 ;
      RECT 32.96 3.298 33.02 3.448 ;
      RECT 32.935 3.306 32.96 3.468 ;
      RECT 32.925 3.31 32.935 3.48 ;
      RECT 32.92 3.311 32.925 3.485 ;
      RECT 32.905 3.313 32.92 3.488 ;
      RECT 32.89 3.315 32.905 3.493 ;
      RECT 32.885 3.315 32.89 3.496 ;
      RECT 32.84 3.32 32.885 3.507 ;
      RECT 32.835 3.324 32.84 3.519 ;
      RECT 32.81 3.32 32.835 3.523 ;
      RECT 32.8 3.316 32.81 3.527 ;
      RECT 32.79 3.315 32.8 3.531 ;
      RECT 32.775 3.305 32.79 3.537 ;
      RECT 32.77 3.293 32.775 3.541 ;
      RECT 32.765 3.29 32.77 3.542 ;
      RECT 32.76 3.287 32.765 3.544 ;
      RECT 32.745 3.275 32.76 3.543 ;
      RECT 32.73 3.257 32.745 3.54 ;
      RECT 32.71 3.236 32.73 3.533 ;
      RECT 32.645 3.225 32.71 3.505 ;
      RECT 32.641 3.225 32.645 3.484 ;
      RECT 32.555 3.225 32.641 3.454 ;
      RECT 32.54 3.225 32.555 3.41 ;
      RECT 33.115 2.325 33.12 2.56 ;
      RECT 32.245 2.241 32.25 2.445 ;
      RECT 32.825 2.27 32.83 2.425 ;
      RECT 32.745 2.25 32.75 2.425 ;
      RECT 33.415 2.392 33.43 2.745 ;
      RECT 33.341 2.377 33.415 2.745 ;
      RECT 33.255 2.36 33.341 2.745 ;
      RECT 33.245 2.35 33.255 2.743 ;
      RECT 33.24 2.348 33.245 2.738 ;
      RECT 33.225 2.346 33.24 2.724 ;
      RECT 33.155 2.338 33.225 2.664 ;
      RECT 33.135 2.329 33.155 2.598 ;
      RECT 33.13 2.326 33.135 2.578 ;
      RECT 33.12 2.325 33.13 2.568 ;
      RECT 33.11 2.325 33.115 2.552 ;
      RECT 33.1 2.324 33.11 2.542 ;
      RECT 33.09 2.322 33.1 2.53 ;
      RECT 33.075 2.319 33.09 2.51 ;
      RECT 33.065 2.317 33.075 2.495 ;
      RECT 33.045 2.314 33.065 2.483 ;
      RECT 33.04 2.312 33.045 2.473 ;
      RECT 33.015 2.31 33.04 2.46 ;
      RECT 32.985 2.305 33.015 2.445 ;
      RECT 32.905 2.296 32.985 2.436 ;
      RECT 32.86 2.285 32.905 2.429 ;
      RECT 32.84 2.276 32.86 2.426 ;
      RECT 32.83 2.271 32.84 2.425 ;
      RECT 32.785 2.265 32.825 2.425 ;
      RECT 32.77 2.257 32.785 2.425 ;
      RECT 32.75 2.252 32.77 2.425 ;
      RECT 32.73 2.249 32.745 2.425 ;
      RECT 32.647 2.248 32.73 2.424 ;
      RECT 32.561 2.247 32.647 2.42 ;
      RECT 32.475 2.245 32.561 2.417 ;
      RECT 32.422 2.244 32.475 2.419 ;
      RECT 32.336 2.243 32.422 2.428 ;
      RECT 32.25 2.242 32.336 2.44 ;
      RECT 32.23 2.241 32.245 2.448 ;
      RECT 32.15 2.24 32.23 2.46 ;
      RECT 32.125 2.24 32.15 2.473 ;
      RECT 32.1 2.24 32.125 2.488 ;
      RECT 32.095 2.24 32.1 2.51 ;
      RECT 32.09 2.24 32.095 2.528 ;
      RECT 32.085 2.24 32.09 2.545 ;
      RECT 32.08 2.24 32.085 2.558 ;
      RECT 32.075 2.24 32.08 2.568 ;
      RECT 32.035 2.24 32.075 2.653 ;
      RECT 32.02 2.24 32.035 2.738 ;
      RECT 32.01 2.241 32.02 2.75 ;
      RECT 31.975 2.246 32.01 2.755 ;
      RECT 31.935 2.255 31.975 2.755 ;
      RECT 31.92 2.265 31.935 2.755 ;
      RECT 31.915 2.275 31.92 2.755 ;
      RECT 31.895 2.302 31.915 2.755 ;
      RECT 31.845 2.385 31.895 2.755 ;
      RECT 31.84 2.447 31.845 2.755 ;
      RECT 31.83 2.46 31.84 2.755 ;
      RECT 31.82 2.482 31.83 2.755 ;
      RECT 31.81 2.507 31.82 2.75 ;
      RECT 31.805 2.545 31.81 2.743 ;
      RECT 31.795 2.655 31.805 2.738 ;
      RECT 33.19 3.576 33.205 3.835 ;
      RECT 33.19 3.591 33.21 3.834 ;
      RECT 33.106 3.591 33.21 3.832 ;
      RECT 33.106 3.605 33.215 3.831 ;
      RECT 33.02 3.647 33.22 3.828 ;
      RECT 33.015 3.59 33.205 3.823 ;
      RECT 33.015 3.661 33.225 3.82 ;
      RECT 33.01 3.692 33.225 3.818 ;
      RECT 33.015 3.689 33.24 3.808 ;
      RECT 33.01 3.735 33.255 3.793 ;
      RECT 33.01 3.763 33.26 3.778 ;
      RECT 33.02 3.565 33.19 3.828 ;
      RECT 32.78 2.575 32.95 2.745 ;
      RECT 32.745 2.575 32.95 2.74 ;
      RECT 32.735 2.575 32.95 2.733 ;
      RECT 32.73 2.56 32.9 2.73 ;
      RECT 31.56 3.097 31.825 3.54 ;
      RECT 31.555 3.068 31.77 3.538 ;
      RECT 31.55 3.222 31.83 3.533 ;
      RECT 31.555 3.117 31.83 3.533 ;
      RECT 31.555 3.128 31.84 3.52 ;
      RECT 31.555 3.075 31.8 3.538 ;
      RECT 31.56 3.062 31.77 3.54 ;
      RECT 31.56 3.06 31.72 3.54 ;
      RECT 31.661 3.052 31.72 3.54 ;
      RECT 31.575 3.053 31.72 3.54 ;
      RECT 31.661 3.051 31.71 3.54 ;
      RECT 31.465 1.866 31.64 2.165 ;
      RECT 31.515 1.828 31.64 2.165 ;
      RECT 31.5 1.83 31.726 2.157 ;
      RECT 31.5 1.833 31.765 2.144 ;
      RECT 31.5 1.834 31.775 2.13 ;
      RECT 31.455 1.885 31.775 2.12 ;
      RECT 31.5 1.835 31.78 2.115 ;
      RECT 31.455 2.045 31.785 2.105 ;
      RECT 31.44 1.905 31.78 2.045 ;
      RECT 31.435 1.921 31.78 1.985 ;
      RECT 31.48 1.845 31.78 2.115 ;
      RECT 31.515 1.826 31.601 2.165 ;
      RECT 29.61 1.74 29.78 2.935 ;
      RECT 29.61 1.74 30.075 1.91 ;
      RECT 29.61 6.97 30.075 7.14 ;
      RECT 29.61 5.945 29.78 7.14 ;
      RECT 28.62 1.74 28.79 2.935 ;
      RECT 28.62 1.74 29.085 1.91 ;
      RECT 28.62 6.97 29.085 7.14 ;
      RECT 28.62 5.945 28.79 7.14 ;
      RECT 26.765 2.635 26.935 3.865 ;
      RECT 26.82 0.855 26.99 2.805 ;
      RECT 26.765 0.575 26.935 1.025 ;
      RECT 26.765 7.855 26.935 8.305 ;
      RECT 26.82 6.075 26.99 8.025 ;
      RECT 26.765 5.015 26.935 6.245 ;
      RECT 26.245 0.575 26.415 3.865 ;
      RECT 26.245 2.075 26.65 2.405 ;
      RECT 26.245 1.235 26.65 1.565 ;
      RECT 26.245 5.015 26.415 8.305 ;
      RECT 26.245 7.315 26.65 7.645 ;
      RECT 26.245 6.475 26.65 6.805 ;
      RECT 24.17 3.126 24.175 3.298 ;
      RECT 24.165 3.119 24.17 3.388 ;
      RECT 24.16 3.113 24.165 3.407 ;
      RECT 24.14 3.107 24.16 3.417 ;
      RECT 24.125 3.102 24.14 3.425 ;
      RECT 24.088 3.096 24.125 3.423 ;
      RECT 24.002 3.082 24.088 3.419 ;
      RECT 23.916 3.064 24.002 3.414 ;
      RECT 23.83 3.045 23.916 3.408 ;
      RECT 23.8 3.033 23.83 3.404 ;
      RECT 23.78 3.027 23.8 3.403 ;
      RECT 23.715 3.025 23.78 3.401 ;
      RECT 23.7 3.025 23.715 3.393 ;
      RECT 23.685 3.025 23.7 3.38 ;
      RECT 23.68 3.025 23.685 3.37 ;
      RECT 23.665 3.025 23.68 3.348 ;
      RECT 23.65 3.025 23.665 3.315 ;
      RECT 23.645 3.025 23.65 3.293 ;
      RECT 23.635 3.025 23.645 3.275 ;
      RECT 23.62 3.025 23.635 3.253 ;
      RECT 23.6 3.025 23.62 3.215 ;
      RECT 23.95 2.31 23.985 2.749 ;
      RECT 23.95 2.31 23.99 2.748 ;
      RECT 23.895 2.37 23.99 2.747 ;
      RECT 23.76 2.542 23.99 2.746 ;
      RECT 23.87 2.42 23.99 2.746 ;
      RECT 23.76 2.542 24.015 2.736 ;
      RECT 23.815 2.487 24.095 2.653 ;
      RECT 23.99 2.281 23.995 2.744 ;
      RECT 23.845 2.457 24.135 2.53 ;
      RECT 23.86 2.44 23.99 2.746 ;
      RECT 23.995 2.28 24.165 2.468 ;
      RECT 23.985 2.283 24.165 2.468 ;
      RECT 23.49 2.16 23.66 2.47 ;
      RECT 23.49 2.16 23.665 2.443 ;
      RECT 23.49 2.16 23.67 2.42 ;
      RECT 23.49 2.16 23.68 2.37 ;
      RECT 23.485 2.265 23.68 2.34 ;
      RECT 23.52 1.835 23.69 2.313 ;
      RECT 23.52 1.835 23.705 2.234 ;
      RECT 23.51 2.045 23.705 2.234 ;
      RECT 23.52 1.845 23.715 2.149 ;
      RECT 23.45 2.587 23.455 2.79 ;
      RECT 23.44 2.575 23.45 2.9 ;
      RECT 23.415 2.575 23.44 2.94 ;
      RECT 23.335 2.575 23.415 3.025 ;
      RECT 23.325 2.575 23.335 3.095 ;
      RECT 23.3 2.575 23.325 3.118 ;
      RECT 23.28 2.575 23.3 3.153 ;
      RECT 23.235 2.585 23.28 3.196 ;
      RECT 23.225 2.597 23.235 3.233 ;
      RECT 23.205 2.611 23.225 3.253 ;
      RECT 23.195 2.629 23.205 3.269 ;
      RECT 23.18 2.655 23.195 3.279 ;
      RECT 23.165 2.696 23.18 3.293 ;
      RECT 23.155 2.731 23.165 3.303 ;
      RECT 23.15 2.747 23.155 3.308 ;
      RECT 23.14 2.762 23.15 3.313 ;
      RECT 23.12 2.805 23.14 3.323 ;
      RECT 23.1 2.842 23.12 3.336 ;
      RECT 23.065 2.865 23.1 3.354 ;
      RECT 23.055 2.879 23.065 3.37 ;
      RECT 23.035 2.889 23.055 3.38 ;
      RECT 23.03 2.898 23.035 3.388 ;
      RECT 23.02 2.905 23.03 3.395 ;
      RECT 23.01 2.912 23.02 3.403 ;
      RECT 22.995 2.922 23.01 3.411 ;
      RECT 22.985 2.936 22.995 3.421 ;
      RECT 22.975 2.948 22.985 3.433 ;
      RECT 22.96 2.97 22.975 3.446 ;
      RECT 22.95 2.992 22.96 3.457 ;
      RECT 22.94 3.012 22.95 3.466 ;
      RECT 22.935 3.027 22.94 3.473 ;
      RECT 22.905 3.06 22.935 3.487 ;
      RECT 22.895 3.095 22.905 3.502 ;
      RECT 22.89 3.102 22.895 3.508 ;
      RECT 22.87 3.117 22.89 3.515 ;
      RECT 22.865 3.132 22.87 3.523 ;
      RECT 22.86 3.141 22.865 3.528 ;
      RECT 22.845 3.147 22.86 3.535 ;
      RECT 22.84 3.153 22.845 3.543 ;
      RECT 22.835 3.157 22.84 3.55 ;
      RECT 22.83 3.161 22.835 3.56 ;
      RECT 22.82 3.166 22.83 3.57 ;
      RECT 22.8 3.177 22.82 3.598 ;
      RECT 22.785 3.189 22.8 3.625 ;
      RECT 22.765 3.202 22.785 3.65 ;
      RECT 22.745 3.217 22.765 3.674 ;
      RECT 22.73 3.232 22.745 3.689 ;
      RECT 22.725 3.243 22.73 3.698 ;
      RECT 22.66 3.288 22.725 3.708 ;
      RECT 22.625 3.347 22.66 3.721 ;
      RECT 22.62 3.37 22.625 3.727 ;
      RECT 22.615 3.377 22.62 3.729 ;
      RECT 22.6 3.387 22.615 3.732 ;
      RECT 22.57 3.412 22.6 3.736 ;
      RECT 22.565 3.43 22.57 3.74 ;
      RECT 22.56 3.437 22.565 3.741 ;
      RECT 22.54 3.445 22.56 3.745 ;
      RECT 22.53 3.452 22.54 3.749 ;
      RECT 22.486 3.463 22.53 3.756 ;
      RECT 22.4 3.491 22.486 3.772 ;
      RECT 22.34 3.515 22.4 3.79 ;
      RECT 22.295 3.525 22.34 3.804 ;
      RECT 22.236 3.533 22.295 3.818 ;
      RECT 22.15 3.54 22.236 3.837 ;
      RECT 22.125 3.545 22.15 3.852 ;
      RECT 22.045 3.548 22.125 3.855 ;
      RECT 21.965 3.552 22.045 3.842 ;
      RECT 21.956 3.555 21.965 3.827 ;
      RECT 21.87 3.555 21.956 3.812 ;
      RECT 21.81 3.557 21.87 3.789 ;
      RECT 21.806 3.56 21.81 3.779 ;
      RECT 21.72 3.56 21.806 3.764 ;
      RECT 21.645 3.56 21.72 3.74 ;
      RECT 22.96 2.569 22.97 2.745 ;
      RECT 22.915 2.536 22.96 2.745 ;
      RECT 22.87 2.487 22.915 2.745 ;
      RECT 22.84 2.457 22.87 2.746 ;
      RECT 22.835 2.44 22.84 2.747 ;
      RECT 22.81 2.42 22.835 2.748 ;
      RECT 22.795 2.395 22.81 2.749 ;
      RECT 22.79 2.382 22.795 2.75 ;
      RECT 22.785 2.376 22.79 2.748 ;
      RECT 22.78 2.368 22.785 2.742 ;
      RECT 22.755 2.36 22.78 2.722 ;
      RECT 22.735 2.349 22.755 2.693 ;
      RECT 22.705 2.334 22.735 2.664 ;
      RECT 22.685 2.32 22.705 2.636 ;
      RECT 22.675 2.314 22.685 2.615 ;
      RECT 22.67 2.311 22.675 2.598 ;
      RECT 22.665 2.308 22.67 2.583 ;
      RECT 22.65 2.303 22.665 2.548 ;
      RECT 22.645 2.299 22.65 2.515 ;
      RECT 22.625 2.294 22.645 2.491 ;
      RECT 22.595 2.286 22.625 2.456 ;
      RECT 22.58 2.28 22.595 2.433 ;
      RECT 22.54 2.273 22.58 2.418 ;
      RECT 22.515 2.265 22.54 2.398 ;
      RECT 22.495 2.26 22.515 2.388 ;
      RECT 22.46 2.254 22.495 2.383 ;
      RECT 22.415 2.245 22.46 2.382 ;
      RECT 22.385 2.241 22.415 2.384 ;
      RECT 22.3 2.249 22.385 2.388 ;
      RECT 22.23 2.26 22.3 2.41 ;
      RECT 22.217 2.266 22.23 2.433 ;
      RECT 22.131 2.273 22.217 2.455 ;
      RECT 22.045 2.285 22.131 2.492 ;
      RECT 22.045 2.662 22.055 2.9 ;
      RECT 22.04 2.291 22.045 2.515 ;
      RECT 22.035 2.547 22.045 2.9 ;
      RECT 22.035 2.292 22.04 2.52 ;
      RECT 22.03 2.293 22.035 2.9 ;
      RECT 22.006 2.295 22.03 2.901 ;
      RECT 21.92 2.303 22.006 2.903 ;
      RECT 21.9 2.317 21.92 2.906 ;
      RECT 21.895 2.345 21.9 2.907 ;
      RECT 21.89 2.357 21.895 2.908 ;
      RECT 21.885 2.372 21.89 2.909 ;
      RECT 21.875 2.402 21.885 2.91 ;
      RECT 21.87 2.44 21.875 2.908 ;
      RECT 21.865 2.46 21.87 2.903 ;
      RECT 21.85 2.495 21.865 2.888 ;
      RECT 21.84 2.547 21.85 2.868 ;
      RECT 21.835 2.577 21.84 2.856 ;
      RECT 21.82 2.59 21.835 2.839 ;
      RECT 21.795 2.594 21.82 2.806 ;
      RECT 21.78 2.592 21.795 2.783 ;
      RECT 21.765 2.591 21.78 2.78 ;
      RECT 21.705 2.589 21.765 2.778 ;
      RECT 21.695 2.587 21.705 2.773 ;
      RECT 21.655 2.586 21.695 2.77 ;
      RECT 21.585 2.583 21.655 2.768 ;
      RECT 21.53 2.581 21.585 2.763 ;
      RECT 21.46 2.575 21.53 2.758 ;
      RECT 21.451 2.575 21.46 2.755 ;
      RECT 21.365 2.575 21.451 2.75 ;
      RECT 21.36 2.575 21.365 2.745 ;
      RECT 22.665 1.81 22.84 2.16 ;
      RECT 22.665 1.825 22.85 2.158 ;
      RECT 22.64 1.775 22.785 2.155 ;
      RECT 22.62 1.776 22.785 2.148 ;
      RECT 22.61 1.777 22.795 2.143 ;
      RECT 22.58 1.778 22.795 2.13 ;
      RECT 22.53 1.779 22.795 2.106 ;
      RECT 22.525 1.781 22.795 2.091 ;
      RECT 22.525 1.847 22.855 2.085 ;
      RECT 22.505 1.788 22.81 2.065 ;
      RECT 22.495 1.797 22.82 1.92 ;
      RECT 22.505 1.792 22.82 2.065 ;
      RECT 22.525 1.782 22.81 2.091 ;
      RECT 22.11 3.107 22.28 3.395 ;
      RECT 22.105 3.125 22.29 3.39 ;
      RECT 22.07 3.133 22.355 3.31 ;
      RECT 22.07 3.133 22.441 3.3 ;
      RECT 22.07 3.133 22.495 3.246 ;
      RECT 22.355 3.03 22.525 3.214 ;
      RECT 22.07 3.185 22.53 3.202 ;
      RECT 22.055 3.155 22.525 3.198 ;
      RECT 22.315 3.037 22.355 3.349 ;
      RECT 22.195 3.074 22.525 3.214 ;
      RECT 22.29 3.049 22.315 3.375 ;
      RECT 22.28 3.056 22.525 3.214 ;
      RECT 22.411 2.52 22.48 2.779 ;
      RECT 22.411 2.575 22.485 2.778 ;
      RECT 22.325 2.575 22.485 2.777 ;
      RECT 22.32 2.575 22.49 2.77 ;
      RECT 22.31 2.52 22.48 2.765 ;
      RECT 21.69 1.819 21.865 2.12 ;
      RECT 21.675 1.807 21.69 2.105 ;
      RECT 21.645 1.806 21.675 2.058 ;
      RECT 21.645 1.824 21.87 2.053 ;
      RECT 21.63 1.808 21.69 2.018 ;
      RECT 21.625 1.83 21.88 1.918 ;
      RECT 21.625 1.813 21.776 1.918 ;
      RECT 21.625 1.815 21.78 1.918 ;
      RECT 21.63 1.811 21.776 2.018 ;
      RECT 21.735 3.047 21.74 3.395 ;
      RECT 21.725 3.037 21.735 3.401 ;
      RECT 21.69 3.027 21.725 3.403 ;
      RECT 21.652 3.022 21.69 3.407 ;
      RECT 21.566 3.015 21.652 3.414 ;
      RECT 21.48 3.005 21.566 3.424 ;
      RECT 21.435 3 21.48 3.432 ;
      RECT 21.431 3 21.435 3.436 ;
      RECT 21.345 3 21.431 3.443 ;
      RECT 21.33 3 21.345 3.443 ;
      RECT 21.32 2.998 21.33 3.415 ;
      RECT 21.31 2.994 21.32 3.358 ;
      RECT 21.29 2.988 21.31 3.29 ;
      RECT 21.285 2.984 21.29 3.238 ;
      RECT 21.275 2.983 21.285 3.205 ;
      RECT 21.225 2.981 21.275 3.19 ;
      RECT 21.2 2.979 21.225 3.185 ;
      RECT 21.157 2.977 21.2 3.181 ;
      RECT 21.071 2.973 21.157 3.169 ;
      RECT 20.985 2.968 21.071 3.153 ;
      RECT 20.955 2.965 20.985 3.14 ;
      RECT 20.93 2.964 20.955 3.128 ;
      RECT 20.925 2.964 20.93 3.118 ;
      RECT 20.885 2.963 20.925 3.11 ;
      RECT 20.87 2.962 20.885 3.103 ;
      RECT 20.82 2.961 20.87 3.095 ;
      RECT 20.818 2.96 20.82 3.09 ;
      RECT 20.732 2.958 20.818 3.09 ;
      RECT 20.646 2.953 20.732 3.09 ;
      RECT 20.56 2.949 20.646 3.09 ;
      RECT 20.511 2.945 20.56 3.088 ;
      RECT 20.425 2.942 20.511 3.083 ;
      RECT 20.402 2.939 20.425 3.079 ;
      RECT 20.316 2.936 20.402 3.074 ;
      RECT 20.23 2.932 20.316 3.065 ;
      RECT 20.205 2.925 20.23 3.06 ;
      RECT 20.145 2.89 20.205 3.057 ;
      RECT 20.125 2.815 20.145 3.054 ;
      RECT 20.12 2.757 20.125 3.053 ;
      RECT 20.095 2.697 20.12 3.052 ;
      RECT 20.02 2.575 20.095 3.048 ;
      RECT 20.01 2.575 20.02 3.04 ;
      RECT 19.995 2.575 20.01 3.03 ;
      RECT 19.98 2.575 19.995 3 ;
      RECT 19.965 2.575 19.98 2.945 ;
      RECT 19.95 2.575 19.965 2.883 ;
      RECT 19.925 2.575 19.95 2.808 ;
      RECT 19.92 2.575 19.925 2.758 ;
      RECT 21.265 2.12 21.285 2.429 ;
      RECT 21.251 2.122 21.3 2.426 ;
      RECT 21.251 2.127 21.32 2.417 ;
      RECT 21.165 2.125 21.3 2.411 ;
      RECT 21.165 2.133 21.355 2.394 ;
      RECT 21.13 2.135 21.355 2.393 ;
      RECT 21.1 2.143 21.355 2.384 ;
      RECT 21.09 2.148 21.375 2.37 ;
      RECT 21.13 2.138 21.375 2.37 ;
      RECT 21.13 2.141 21.385 2.358 ;
      RECT 21.1 2.143 21.395 2.345 ;
      RECT 21.1 2.147 21.405 2.288 ;
      RECT 21.09 2.152 21.41 2.203 ;
      RECT 21.251 2.12 21.285 2.426 ;
      RECT 21.13 7.855 21.3 8.305 ;
      RECT 21.185 6.075 21.355 8.025 ;
      RECT 21.13 5.015 21.3 6.245 ;
      RECT 20.69 2.223 20.695 2.435 ;
      RECT 20.565 2.22 20.58 2.435 ;
      RECT 20.03 2.25 20.1 2.435 ;
      RECT 19.915 2.25 19.95 2.43 ;
      RECT 21.036 2.552 21.055 2.746 ;
      RECT 20.95 2.507 21.036 2.747 ;
      RECT 20.94 2.46 20.95 2.749 ;
      RECT 20.935 2.44 20.94 2.75 ;
      RECT 20.915 2.405 20.935 2.751 ;
      RECT 20.9 2.355 20.915 2.752 ;
      RECT 20.88 2.292 20.9 2.753 ;
      RECT 20.87 2.255 20.88 2.754 ;
      RECT 20.855 2.244 20.87 2.755 ;
      RECT 20.85 2.236 20.855 2.753 ;
      RECT 20.84 2.235 20.85 2.745 ;
      RECT 20.81 2.232 20.84 2.724 ;
      RECT 20.735 2.227 20.81 2.669 ;
      RECT 20.72 2.223 20.735 2.615 ;
      RECT 20.71 2.223 20.72 2.51 ;
      RECT 20.695 2.223 20.71 2.443 ;
      RECT 20.68 2.223 20.69 2.433 ;
      RECT 20.625 2.222 20.68 2.43 ;
      RECT 20.58 2.22 20.625 2.433 ;
      RECT 20.552 2.22 20.565 2.436 ;
      RECT 20.466 2.224 20.552 2.438 ;
      RECT 20.38 2.23 20.466 2.443 ;
      RECT 20.36 2.234 20.38 2.445 ;
      RECT 20.358 2.235 20.36 2.444 ;
      RECT 20.272 2.237 20.358 2.443 ;
      RECT 20.186 2.242 20.272 2.44 ;
      RECT 20.1 2.247 20.186 2.437 ;
      RECT 19.95 2.25 20.03 2.433 ;
      RECT 20.61 5.015 20.78 8.305 ;
      RECT 20.61 7.315 21.015 7.645 ;
      RECT 20.61 6.475 21.015 6.805 ;
      RECT 20.726 3.225 20.775 3.559 ;
      RECT 20.726 3.225 20.78 3.558 ;
      RECT 20.64 3.225 20.78 3.557 ;
      RECT 20.415 3.333 20.785 3.555 ;
      RECT 20.64 3.225 20.81 3.548 ;
      RECT 20.61 3.237 20.815 3.539 ;
      RECT 20.595 3.255 20.82 3.536 ;
      RECT 20.41 3.339 20.82 3.463 ;
      RECT 20.405 3.346 20.82 3.423 ;
      RECT 20.42 3.312 20.82 3.536 ;
      RECT 20.581 3.258 20.785 3.555 ;
      RECT 20.495 3.278 20.82 3.536 ;
      RECT 20.595 3.252 20.815 3.539 ;
      RECT 20.365 2.576 20.555 2.77 ;
      RECT 20.36 2.578 20.555 2.769 ;
      RECT 20.355 2.582 20.57 2.766 ;
      RECT 20.37 2.575 20.57 2.766 ;
      RECT 20.355 2.685 20.575 2.761 ;
      RECT 19.65 3.185 19.741 3.483 ;
      RECT 19.645 3.187 19.82 3.478 ;
      RECT 19.65 3.185 19.82 3.478 ;
      RECT 19.645 3.191 19.84 3.476 ;
      RECT 19.645 3.246 19.88 3.475 ;
      RECT 19.645 3.281 19.895 3.469 ;
      RECT 19.645 3.315 19.905 3.459 ;
      RECT 19.635 3.195 19.84 3.31 ;
      RECT 19.635 3.215 19.855 3.31 ;
      RECT 19.635 3.198 19.845 3.31 ;
      RECT 19.86 1.966 19.865 2.028 ;
      RECT 19.855 1.888 19.86 2.051 ;
      RECT 19.85 1.845 19.855 2.062 ;
      RECT 19.845 1.835 19.85 2.074 ;
      RECT 19.84 1.835 19.845 2.083 ;
      RECT 19.815 1.835 19.84 2.115 ;
      RECT 19.81 1.835 19.815 2.148 ;
      RECT 19.795 1.835 19.81 2.173 ;
      RECT 19.785 1.835 19.795 2.2 ;
      RECT 19.78 1.835 19.785 2.213 ;
      RECT 19.775 1.835 19.78 2.228 ;
      RECT 19.765 1.835 19.775 2.243 ;
      RECT 19.76 1.835 19.765 2.263 ;
      RECT 19.735 1.835 19.76 2.298 ;
      RECT 19.69 1.835 19.735 2.343 ;
      RECT 19.68 1.835 19.69 2.356 ;
      RECT 19.595 1.92 19.68 2.363 ;
      RECT 19.56 2.042 19.595 2.372 ;
      RECT 19.555 2.082 19.56 2.376 ;
      RECT 19.535 2.105 19.555 2.378 ;
      RECT 19.53 2.135 19.535 2.381 ;
      RECT 19.52 2.147 19.53 2.382 ;
      RECT 19.475 2.17 19.52 2.387 ;
      RECT 19.435 2.2 19.475 2.395 ;
      RECT 19.4 2.212 19.435 2.401 ;
      RECT 19.395 2.217 19.4 2.405 ;
      RECT 19.325 2.227 19.395 2.412 ;
      RECT 19.285 2.237 19.325 2.422 ;
      RECT 19.265 2.242 19.285 2.428 ;
      RECT 19.255 2.246 19.265 2.433 ;
      RECT 19.25 2.249 19.255 2.436 ;
      RECT 19.24 2.25 19.25 2.437 ;
      RECT 19.215 2.252 19.24 2.441 ;
      RECT 19.205 2.257 19.215 2.444 ;
      RECT 19.16 2.265 19.205 2.445 ;
      RECT 19.035 2.27 19.16 2.445 ;
      RECT 19.59 2.567 19.61 2.749 ;
      RECT 19.541 2.552 19.59 2.748 ;
      RECT 19.455 2.567 19.61 2.746 ;
      RECT 19.44 2.567 19.61 2.745 ;
      RECT 19.405 2.545 19.575 2.73 ;
      RECT 19.475 3.565 19.49 3.774 ;
      RECT 19.475 3.573 19.495 3.773 ;
      RECT 19.42 3.573 19.495 3.772 ;
      RECT 19.4 3.577 19.5 3.77 ;
      RECT 19.38 3.527 19.42 3.769 ;
      RECT 19.325 3.585 19.505 3.767 ;
      RECT 19.29 3.542 19.42 3.765 ;
      RECT 19.286 3.545 19.475 3.764 ;
      RECT 19.2 3.553 19.475 3.762 ;
      RECT 19.2 3.597 19.51 3.755 ;
      RECT 19.19 3.69 19.51 3.753 ;
      RECT 19.2 3.609 19.515 3.738 ;
      RECT 19.2 3.63 19.53 3.708 ;
      RECT 19.2 3.657 19.535 3.678 ;
      RECT 19.325 3.535 19.42 3.767 ;
      RECT 18.955 2.58 18.96 3.118 ;
      RECT 18.76 2.91 18.765 3.105 ;
      RECT 17.06 2.575 17.075 2.955 ;
      RECT 19.125 2.575 19.13 2.745 ;
      RECT 19.12 2.575 19.125 2.755 ;
      RECT 19.115 2.575 19.12 2.768 ;
      RECT 19.09 2.575 19.115 2.81 ;
      RECT 19.065 2.575 19.09 2.883 ;
      RECT 19.05 2.575 19.065 2.935 ;
      RECT 19.045 2.575 19.05 2.965 ;
      RECT 19.02 2.575 19.045 3.005 ;
      RECT 19.005 2.575 19.02 3.06 ;
      RECT 19 2.575 19.005 3.093 ;
      RECT 18.975 2.575 19 3.113 ;
      RECT 18.96 2.575 18.975 3.119 ;
      RECT 18.89 2.61 18.955 3.115 ;
      RECT 18.84 2.665 18.89 3.11 ;
      RECT 18.83 2.697 18.84 3.108 ;
      RECT 18.825 2.722 18.83 3.108 ;
      RECT 18.805 2.795 18.825 3.108 ;
      RECT 18.795 2.875 18.805 3.107 ;
      RECT 18.78 2.905 18.795 3.107 ;
      RECT 18.765 2.91 18.78 3.106 ;
      RECT 18.705 2.912 18.76 3.103 ;
      RECT 18.675 2.917 18.705 3.099 ;
      RECT 18.673 2.92 18.675 3.098 ;
      RECT 18.587 2.922 18.673 3.095 ;
      RECT 18.501 2.928 18.587 3.089 ;
      RECT 18.415 2.933 18.501 3.083 ;
      RECT 18.342 2.938 18.415 3.084 ;
      RECT 18.256 2.944 18.342 3.092 ;
      RECT 18.17 2.95 18.256 3.101 ;
      RECT 18.15 2.954 18.17 3.106 ;
      RECT 18.103 2.956 18.15 3.109 ;
      RECT 18.017 2.961 18.103 3.115 ;
      RECT 17.931 2.966 18.017 3.124 ;
      RECT 17.845 2.972 17.931 3.132 ;
      RECT 17.76 2.97 17.845 3.141 ;
      RECT 17.756 2.965 17.76 3.145 ;
      RECT 17.67 2.96 17.756 3.137 ;
      RECT 17.606 2.951 17.67 3.125 ;
      RECT 17.52 2.942 17.606 3.112 ;
      RECT 17.496 2.935 17.52 3.103 ;
      RECT 17.41 2.929 17.496 3.09 ;
      RECT 17.37 2.922 17.41 3.076 ;
      RECT 17.365 2.912 17.37 3.072 ;
      RECT 17.355 2.9 17.365 3.071 ;
      RECT 17.335 2.87 17.355 3.068 ;
      RECT 17.28 2.79 17.335 3.062 ;
      RECT 17.26 2.709 17.28 3.057 ;
      RECT 17.24 2.667 17.26 3.053 ;
      RECT 17.215 2.62 17.24 3.047 ;
      RECT 17.21 2.595 17.215 3.044 ;
      RECT 17.175 2.575 17.21 3.039 ;
      RECT 17.166 2.575 17.175 3.032 ;
      RECT 17.08 2.575 17.166 3.002 ;
      RECT 17.075 2.575 17.08 2.965 ;
      RECT 17.04 2.575 17.06 2.887 ;
      RECT 17.035 2.617 17.04 2.852 ;
      RECT 17.03 2.692 17.035 2.808 ;
      RECT 18.48 2.497 18.655 2.745 ;
      RECT 18.48 2.497 18.66 2.743 ;
      RECT 18.475 2.529 18.66 2.703 ;
      RECT 18.505 2.47 18.675 2.69 ;
      RECT 18.47 2.547 18.675 2.623 ;
      RECT 17.78 2.01 17.95 2.185 ;
      RECT 17.78 2.01 18.122 2.177 ;
      RECT 17.78 2.01 18.205 2.171 ;
      RECT 17.78 2.01 18.24 2.167 ;
      RECT 17.78 2.01 18.26 2.166 ;
      RECT 17.78 2.01 18.346 2.162 ;
      RECT 18.24 1.835 18.41 2.157 ;
      RECT 17.815 1.942 18.44 2.155 ;
      RECT 17.805 1.997 18.445 2.153 ;
      RECT 17.78 2.033 18.455 2.148 ;
      RECT 17.78 2.06 18.46 2.078 ;
      RECT 17.845 1.885 18.42 2.155 ;
      RECT 18.036 1.87 18.42 2.155 ;
      RECT 17.87 1.873 18.42 2.155 ;
      RECT 17.95 1.871 18.036 2.182 ;
      RECT 18.036 1.868 18.415 2.155 ;
      RECT 18.22 1.845 18.415 2.155 ;
      RECT 18.122 1.866 18.415 2.155 ;
      RECT 18.205 1.86 18.22 2.168 ;
      RECT 18.355 3.225 18.36 3.425 ;
      RECT 17.82 3.29 17.865 3.425 ;
      RECT 18.39 3.225 18.41 3.398 ;
      RECT 18.36 3.225 18.39 3.413 ;
      RECT 18.295 3.225 18.355 3.45 ;
      RECT 18.28 3.225 18.295 3.48 ;
      RECT 18.265 3.225 18.28 3.493 ;
      RECT 18.245 3.225 18.265 3.508 ;
      RECT 18.24 3.225 18.245 3.517 ;
      RECT 18.23 3.229 18.24 3.522 ;
      RECT 18.215 3.239 18.23 3.533 ;
      RECT 18.19 3.255 18.215 3.543 ;
      RECT 18.18 3.269 18.19 3.545 ;
      RECT 18.16 3.281 18.18 3.542 ;
      RECT 18.13 3.302 18.16 3.536 ;
      RECT 18.12 3.314 18.13 3.531 ;
      RECT 18.11 3.312 18.12 3.528 ;
      RECT 18.095 3.311 18.11 3.523 ;
      RECT 18.09 3.31 18.095 3.518 ;
      RECT 18.055 3.308 18.09 3.508 ;
      RECT 18.035 3.305 18.055 3.49 ;
      RECT 18.025 3.303 18.035 3.485 ;
      RECT 18.015 3.302 18.025 3.48 ;
      RECT 17.98 3.3 18.015 3.468 ;
      RECT 17.925 3.296 17.98 3.448 ;
      RECT 17.915 3.294 17.925 3.433 ;
      RECT 17.91 3.294 17.915 3.428 ;
      RECT 17.865 3.292 17.91 3.425 ;
      RECT 17.77 3.29 17.82 3.429 ;
      RECT 17.76 3.291 17.77 3.434 ;
      RECT 17.7 3.298 17.76 3.448 ;
      RECT 17.675 3.306 17.7 3.468 ;
      RECT 17.665 3.31 17.675 3.48 ;
      RECT 17.66 3.311 17.665 3.485 ;
      RECT 17.645 3.313 17.66 3.488 ;
      RECT 17.63 3.315 17.645 3.493 ;
      RECT 17.625 3.315 17.63 3.496 ;
      RECT 17.58 3.32 17.625 3.507 ;
      RECT 17.575 3.324 17.58 3.519 ;
      RECT 17.55 3.32 17.575 3.523 ;
      RECT 17.54 3.316 17.55 3.527 ;
      RECT 17.53 3.315 17.54 3.531 ;
      RECT 17.515 3.305 17.53 3.537 ;
      RECT 17.51 3.293 17.515 3.541 ;
      RECT 17.505 3.29 17.51 3.542 ;
      RECT 17.5 3.287 17.505 3.544 ;
      RECT 17.485 3.275 17.5 3.543 ;
      RECT 17.47 3.257 17.485 3.54 ;
      RECT 17.45 3.236 17.47 3.533 ;
      RECT 17.385 3.225 17.45 3.505 ;
      RECT 17.381 3.225 17.385 3.484 ;
      RECT 17.295 3.225 17.381 3.454 ;
      RECT 17.28 3.225 17.295 3.41 ;
      RECT 17.855 2.325 17.86 2.56 ;
      RECT 16.985 2.241 16.99 2.445 ;
      RECT 17.565 2.27 17.57 2.425 ;
      RECT 17.485 2.25 17.49 2.425 ;
      RECT 18.155 2.392 18.17 2.745 ;
      RECT 18.081 2.377 18.155 2.745 ;
      RECT 17.995 2.36 18.081 2.745 ;
      RECT 17.985 2.35 17.995 2.743 ;
      RECT 17.98 2.348 17.985 2.738 ;
      RECT 17.965 2.346 17.98 2.724 ;
      RECT 17.895 2.338 17.965 2.664 ;
      RECT 17.875 2.329 17.895 2.598 ;
      RECT 17.87 2.326 17.875 2.578 ;
      RECT 17.86 2.325 17.87 2.568 ;
      RECT 17.85 2.325 17.855 2.552 ;
      RECT 17.84 2.324 17.85 2.542 ;
      RECT 17.83 2.322 17.84 2.53 ;
      RECT 17.815 2.319 17.83 2.51 ;
      RECT 17.805 2.317 17.815 2.495 ;
      RECT 17.785 2.314 17.805 2.483 ;
      RECT 17.78 2.312 17.785 2.473 ;
      RECT 17.755 2.31 17.78 2.46 ;
      RECT 17.725 2.305 17.755 2.445 ;
      RECT 17.645 2.296 17.725 2.436 ;
      RECT 17.6 2.285 17.645 2.429 ;
      RECT 17.58 2.276 17.6 2.426 ;
      RECT 17.57 2.271 17.58 2.425 ;
      RECT 17.525 2.265 17.565 2.425 ;
      RECT 17.51 2.257 17.525 2.425 ;
      RECT 17.49 2.252 17.51 2.425 ;
      RECT 17.47 2.249 17.485 2.425 ;
      RECT 17.387 2.248 17.47 2.424 ;
      RECT 17.301 2.247 17.387 2.42 ;
      RECT 17.215 2.245 17.301 2.417 ;
      RECT 17.162 2.244 17.215 2.419 ;
      RECT 17.076 2.243 17.162 2.428 ;
      RECT 16.99 2.242 17.076 2.44 ;
      RECT 16.97 2.241 16.985 2.448 ;
      RECT 16.89 2.24 16.97 2.46 ;
      RECT 16.865 2.24 16.89 2.473 ;
      RECT 16.84 2.24 16.865 2.488 ;
      RECT 16.835 2.24 16.84 2.51 ;
      RECT 16.83 2.24 16.835 2.528 ;
      RECT 16.825 2.24 16.83 2.545 ;
      RECT 16.82 2.24 16.825 2.558 ;
      RECT 16.815 2.24 16.82 2.568 ;
      RECT 16.775 2.24 16.815 2.653 ;
      RECT 16.76 2.24 16.775 2.738 ;
      RECT 16.75 2.241 16.76 2.75 ;
      RECT 16.715 2.246 16.75 2.755 ;
      RECT 16.675 2.255 16.715 2.755 ;
      RECT 16.66 2.265 16.675 2.755 ;
      RECT 16.655 2.275 16.66 2.755 ;
      RECT 16.635 2.302 16.655 2.755 ;
      RECT 16.585 2.385 16.635 2.755 ;
      RECT 16.58 2.447 16.585 2.755 ;
      RECT 16.57 2.46 16.58 2.755 ;
      RECT 16.56 2.482 16.57 2.755 ;
      RECT 16.55 2.507 16.56 2.75 ;
      RECT 16.545 2.545 16.55 2.743 ;
      RECT 16.535 2.655 16.545 2.738 ;
      RECT 17.93 3.576 17.945 3.835 ;
      RECT 17.93 3.591 17.95 3.834 ;
      RECT 17.846 3.591 17.95 3.832 ;
      RECT 17.846 3.605 17.955 3.831 ;
      RECT 17.76 3.647 17.96 3.828 ;
      RECT 17.755 3.59 17.945 3.823 ;
      RECT 17.755 3.661 17.965 3.82 ;
      RECT 17.75 3.692 17.965 3.818 ;
      RECT 17.755 3.689 17.98 3.808 ;
      RECT 17.75 3.735 17.995 3.793 ;
      RECT 17.75 3.763 18 3.778 ;
      RECT 17.76 3.565 17.93 3.828 ;
      RECT 17.52 2.575 17.69 2.745 ;
      RECT 17.485 2.575 17.69 2.74 ;
      RECT 17.475 2.575 17.69 2.733 ;
      RECT 17.47 2.56 17.64 2.73 ;
      RECT 16.3 3.097 16.565 3.54 ;
      RECT 16.295 3.068 16.51 3.538 ;
      RECT 16.29 3.222 16.57 3.533 ;
      RECT 16.295 3.117 16.57 3.533 ;
      RECT 16.295 3.128 16.58 3.52 ;
      RECT 16.295 3.075 16.54 3.538 ;
      RECT 16.3 3.062 16.51 3.54 ;
      RECT 16.3 3.06 16.46 3.54 ;
      RECT 16.401 3.052 16.46 3.54 ;
      RECT 16.315 3.053 16.46 3.54 ;
      RECT 16.401 3.051 16.45 3.54 ;
      RECT 16.205 1.866 16.38 2.165 ;
      RECT 16.255 1.828 16.38 2.165 ;
      RECT 16.24 1.83 16.466 2.157 ;
      RECT 16.24 1.833 16.505 2.144 ;
      RECT 16.24 1.834 16.515 2.13 ;
      RECT 16.195 1.885 16.515 2.12 ;
      RECT 16.24 1.835 16.52 2.115 ;
      RECT 16.195 2.045 16.525 2.105 ;
      RECT 16.18 1.905 16.52 2.045 ;
      RECT 16.175 1.921 16.52 1.985 ;
      RECT 16.22 1.845 16.52 2.115 ;
      RECT 16.255 1.826 16.341 2.165 ;
      RECT 14.35 1.74 14.52 2.935 ;
      RECT 14.35 1.74 14.815 1.91 ;
      RECT 14.35 6.97 14.815 7.14 ;
      RECT 14.35 5.945 14.52 7.14 ;
      RECT 13.36 1.74 13.53 2.935 ;
      RECT 13.36 1.74 13.825 1.91 ;
      RECT 13.36 6.97 13.825 7.14 ;
      RECT 13.36 5.945 13.53 7.14 ;
      RECT 11.505 2.635 11.675 3.865 ;
      RECT 11.56 0.855 11.73 2.805 ;
      RECT 11.505 0.575 11.675 1.025 ;
      RECT 11.505 7.855 11.675 8.305 ;
      RECT 11.56 6.075 11.73 8.025 ;
      RECT 11.505 5.015 11.675 6.245 ;
      RECT 10.985 0.575 11.155 3.865 ;
      RECT 10.985 2.075 11.39 2.405 ;
      RECT 10.985 1.235 11.39 1.565 ;
      RECT 10.985 5.015 11.155 8.305 ;
      RECT 10.985 7.315 11.39 7.645 ;
      RECT 10.985 6.475 11.39 6.805 ;
      RECT 8.91 3.126 8.915 3.298 ;
      RECT 8.905 3.119 8.91 3.388 ;
      RECT 8.9 3.113 8.905 3.407 ;
      RECT 8.88 3.107 8.9 3.417 ;
      RECT 8.865 3.102 8.88 3.425 ;
      RECT 8.828 3.096 8.865 3.423 ;
      RECT 8.742 3.082 8.828 3.419 ;
      RECT 8.656 3.064 8.742 3.414 ;
      RECT 8.57 3.045 8.656 3.408 ;
      RECT 8.54 3.033 8.57 3.404 ;
      RECT 8.52 3.027 8.54 3.403 ;
      RECT 8.455 3.025 8.52 3.401 ;
      RECT 8.44 3.025 8.455 3.393 ;
      RECT 8.425 3.025 8.44 3.38 ;
      RECT 8.42 3.025 8.425 3.37 ;
      RECT 8.405 3.025 8.42 3.348 ;
      RECT 8.39 3.025 8.405 3.315 ;
      RECT 8.385 3.025 8.39 3.293 ;
      RECT 8.375 3.025 8.385 3.275 ;
      RECT 8.36 3.025 8.375 3.253 ;
      RECT 8.34 3.025 8.36 3.215 ;
      RECT 8.69 2.31 8.725 2.749 ;
      RECT 8.69 2.31 8.73 2.748 ;
      RECT 8.635 2.37 8.73 2.747 ;
      RECT 8.5 2.542 8.73 2.746 ;
      RECT 8.61 2.42 8.73 2.746 ;
      RECT 8.5 2.542 8.755 2.736 ;
      RECT 8.555 2.487 8.835 2.653 ;
      RECT 8.73 2.281 8.735 2.744 ;
      RECT 8.585 2.457 8.875 2.53 ;
      RECT 8.6 2.44 8.73 2.746 ;
      RECT 8.735 2.28 8.905 2.468 ;
      RECT 8.725 2.283 8.905 2.468 ;
      RECT 8.23 2.16 8.4 2.47 ;
      RECT 8.23 2.16 8.405 2.443 ;
      RECT 8.23 2.16 8.41 2.42 ;
      RECT 8.23 2.16 8.42 2.37 ;
      RECT 8.225 2.265 8.42 2.34 ;
      RECT 8.26 1.835 8.43 2.313 ;
      RECT 8.26 1.835 8.445 2.234 ;
      RECT 8.25 2.045 8.445 2.234 ;
      RECT 8.26 1.845 8.455 2.149 ;
      RECT 8.19 2.587 8.195 2.79 ;
      RECT 8.18 2.575 8.19 2.9 ;
      RECT 8.155 2.575 8.18 2.94 ;
      RECT 8.075 2.575 8.155 3.025 ;
      RECT 8.065 2.575 8.075 3.095 ;
      RECT 8.04 2.575 8.065 3.118 ;
      RECT 8.02 2.575 8.04 3.153 ;
      RECT 7.975 2.585 8.02 3.196 ;
      RECT 7.965 2.597 7.975 3.233 ;
      RECT 7.945 2.611 7.965 3.253 ;
      RECT 7.935 2.629 7.945 3.269 ;
      RECT 7.92 2.655 7.935 3.279 ;
      RECT 7.905 2.696 7.92 3.293 ;
      RECT 7.895 2.731 7.905 3.303 ;
      RECT 7.89 2.747 7.895 3.308 ;
      RECT 7.88 2.762 7.89 3.313 ;
      RECT 7.86 2.805 7.88 3.323 ;
      RECT 7.84 2.842 7.86 3.336 ;
      RECT 7.805 2.865 7.84 3.354 ;
      RECT 7.795 2.879 7.805 3.37 ;
      RECT 7.775 2.889 7.795 3.38 ;
      RECT 7.77 2.898 7.775 3.388 ;
      RECT 7.76 2.905 7.77 3.395 ;
      RECT 7.75 2.912 7.76 3.403 ;
      RECT 7.735 2.922 7.75 3.411 ;
      RECT 7.725 2.936 7.735 3.421 ;
      RECT 7.715 2.948 7.725 3.433 ;
      RECT 7.7 2.97 7.715 3.446 ;
      RECT 7.69 2.992 7.7 3.457 ;
      RECT 7.68 3.012 7.69 3.466 ;
      RECT 7.675 3.027 7.68 3.473 ;
      RECT 7.645 3.06 7.675 3.487 ;
      RECT 7.635 3.095 7.645 3.502 ;
      RECT 7.63 3.102 7.635 3.508 ;
      RECT 7.61 3.117 7.63 3.515 ;
      RECT 7.605 3.132 7.61 3.523 ;
      RECT 7.6 3.141 7.605 3.528 ;
      RECT 7.585 3.147 7.6 3.535 ;
      RECT 7.58 3.153 7.585 3.543 ;
      RECT 7.575 3.157 7.58 3.55 ;
      RECT 7.57 3.161 7.575 3.56 ;
      RECT 7.56 3.166 7.57 3.57 ;
      RECT 7.54 3.177 7.56 3.598 ;
      RECT 7.525 3.189 7.54 3.625 ;
      RECT 7.505 3.202 7.525 3.65 ;
      RECT 7.485 3.217 7.505 3.674 ;
      RECT 7.47 3.232 7.485 3.689 ;
      RECT 7.465 3.243 7.47 3.698 ;
      RECT 7.4 3.288 7.465 3.708 ;
      RECT 7.365 3.347 7.4 3.721 ;
      RECT 7.36 3.37 7.365 3.727 ;
      RECT 7.355 3.377 7.36 3.729 ;
      RECT 7.34 3.387 7.355 3.732 ;
      RECT 7.31 3.412 7.34 3.736 ;
      RECT 7.305 3.43 7.31 3.74 ;
      RECT 7.3 3.437 7.305 3.741 ;
      RECT 7.28 3.445 7.3 3.745 ;
      RECT 7.27 3.452 7.28 3.749 ;
      RECT 7.226 3.463 7.27 3.756 ;
      RECT 7.14 3.491 7.226 3.772 ;
      RECT 7.08 3.515 7.14 3.79 ;
      RECT 7.035 3.525 7.08 3.804 ;
      RECT 6.976 3.533 7.035 3.818 ;
      RECT 6.89 3.54 6.976 3.837 ;
      RECT 6.865 3.545 6.89 3.852 ;
      RECT 6.785 3.548 6.865 3.855 ;
      RECT 6.705 3.552 6.785 3.842 ;
      RECT 6.696 3.555 6.705 3.827 ;
      RECT 6.61 3.555 6.696 3.812 ;
      RECT 6.55 3.557 6.61 3.789 ;
      RECT 6.546 3.56 6.55 3.779 ;
      RECT 6.46 3.56 6.546 3.764 ;
      RECT 6.385 3.56 6.46 3.74 ;
      RECT 7.7 2.569 7.71 2.745 ;
      RECT 7.655 2.536 7.7 2.745 ;
      RECT 7.61 2.487 7.655 2.745 ;
      RECT 7.58 2.457 7.61 2.746 ;
      RECT 7.575 2.44 7.58 2.747 ;
      RECT 7.55 2.42 7.575 2.748 ;
      RECT 7.535 2.395 7.55 2.749 ;
      RECT 7.53 2.382 7.535 2.75 ;
      RECT 7.525 2.376 7.53 2.748 ;
      RECT 7.52 2.368 7.525 2.742 ;
      RECT 7.495 2.36 7.52 2.722 ;
      RECT 7.475 2.349 7.495 2.693 ;
      RECT 7.445 2.334 7.475 2.664 ;
      RECT 7.425 2.32 7.445 2.636 ;
      RECT 7.415 2.314 7.425 2.615 ;
      RECT 7.41 2.311 7.415 2.598 ;
      RECT 7.405 2.308 7.41 2.583 ;
      RECT 7.39 2.303 7.405 2.548 ;
      RECT 7.385 2.299 7.39 2.515 ;
      RECT 7.365 2.294 7.385 2.491 ;
      RECT 7.335 2.286 7.365 2.456 ;
      RECT 7.32 2.28 7.335 2.433 ;
      RECT 7.28 2.273 7.32 2.418 ;
      RECT 7.255 2.265 7.28 2.398 ;
      RECT 7.235 2.26 7.255 2.388 ;
      RECT 7.2 2.254 7.235 2.383 ;
      RECT 7.155 2.245 7.2 2.382 ;
      RECT 7.125 2.241 7.155 2.384 ;
      RECT 7.04 2.249 7.125 2.388 ;
      RECT 6.97 2.26 7.04 2.41 ;
      RECT 6.957 2.266 6.97 2.433 ;
      RECT 6.871 2.273 6.957 2.455 ;
      RECT 6.785 2.285 6.871 2.492 ;
      RECT 6.785 2.662 6.795 2.9 ;
      RECT 6.78 2.291 6.785 2.515 ;
      RECT 6.775 2.547 6.785 2.9 ;
      RECT 6.775 2.292 6.78 2.52 ;
      RECT 6.77 2.293 6.775 2.9 ;
      RECT 6.746 2.295 6.77 2.901 ;
      RECT 6.66 2.303 6.746 2.903 ;
      RECT 6.64 2.317 6.66 2.906 ;
      RECT 6.635 2.345 6.64 2.907 ;
      RECT 6.63 2.357 6.635 2.908 ;
      RECT 6.625 2.372 6.63 2.909 ;
      RECT 6.615 2.402 6.625 2.91 ;
      RECT 6.61 2.44 6.615 2.908 ;
      RECT 6.605 2.46 6.61 2.903 ;
      RECT 6.59 2.495 6.605 2.888 ;
      RECT 6.58 2.547 6.59 2.868 ;
      RECT 6.575 2.577 6.58 2.856 ;
      RECT 6.56 2.59 6.575 2.839 ;
      RECT 6.535 2.594 6.56 2.806 ;
      RECT 6.52 2.592 6.535 2.783 ;
      RECT 6.505 2.591 6.52 2.78 ;
      RECT 6.445 2.589 6.505 2.778 ;
      RECT 6.435 2.587 6.445 2.773 ;
      RECT 6.395 2.586 6.435 2.77 ;
      RECT 6.325 2.583 6.395 2.768 ;
      RECT 6.27 2.581 6.325 2.763 ;
      RECT 6.2 2.575 6.27 2.758 ;
      RECT 6.191 2.575 6.2 2.755 ;
      RECT 6.105 2.575 6.191 2.75 ;
      RECT 6.1 2.575 6.105 2.745 ;
      RECT 7.405 1.81 7.58 2.16 ;
      RECT 7.405 1.825 7.59 2.158 ;
      RECT 7.38 1.775 7.525 2.155 ;
      RECT 7.36 1.776 7.525 2.148 ;
      RECT 7.35 1.777 7.535 2.143 ;
      RECT 7.32 1.778 7.535 2.13 ;
      RECT 7.27 1.779 7.535 2.106 ;
      RECT 7.265 1.781 7.535 2.091 ;
      RECT 7.265 1.847 7.595 2.085 ;
      RECT 7.245 1.788 7.55 2.065 ;
      RECT 7.235 1.797 7.56 1.92 ;
      RECT 7.245 1.792 7.56 2.065 ;
      RECT 7.265 1.782 7.55 2.091 ;
      RECT 6.85 3.107 7.02 3.395 ;
      RECT 6.845 3.125 7.03 3.39 ;
      RECT 6.81 3.133 7.095 3.31 ;
      RECT 6.81 3.133 7.181 3.3 ;
      RECT 6.81 3.133 7.235 3.246 ;
      RECT 7.095 3.03 7.265 3.214 ;
      RECT 6.81 3.185 7.27 3.202 ;
      RECT 6.795 3.155 7.265 3.198 ;
      RECT 7.055 3.037 7.095 3.349 ;
      RECT 6.935 3.074 7.265 3.214 ;
      RECT 7.03 3.049 7.055 3.375 ;
      RECT 7.02 3.056 7.265 3.214 ;
      RECT 7.151 2.52 7.22 2.779 ;
      RECT 7.151 2.575 7.225 2.778 ;
      RECT 7.065 2.575 7.225 2.777 ;
      RECT 7.06 2.575 7.23 2.77 ;
      RECT 7.05 2.52 7.22 2.765 ;
      RECT 6.43 1.819 6.605 2.12 ;
      RECT 6.415 1.807 6.43 2.105 ;
      RECT 6.385 1.806 6.415 2.058 ;
      RECT 6.385 1.824 6.61 2.053 ;
      RECT 6.37 1.808 6.43 2.018 ;
      RECT 6.365 1.83 6.62 1.918 ;
      RECT 6.365 1.813 6.516 1.918 ;
      RECT 6.365 1.815 6.52 1.918 ;
      RECT 6.37 1.811 6.516 2.018 ;
      RECT 6.475 3.047 6.48 3.395 ;
      RECT 6.465 3.037 6.475 3.401 ;
      RECT 6.43 3.027 6.465 3.403 ;
      RECT 6.392 3.022 6.43 3.407 ;
      RECT 6.306 3.015 6.392 3.414 ;
      RECT 6.22 3.005 6.306 3.424 ;
      RECT 6.175 3 6.22 3.432 ;
      RECT 6.171 3 6.175 3.436 ;
      RECT 6.085 3 6.171 3.443 ;
      RECT 6.07 3 6.085 3.443 ;
      RECT 6.06 2.998 6.07 3.415 ;
      RECT 6.05 2.994 6.06 3.358 ;
      RECT 6.03 2.988 6.05 3.29 ;
      RECT 6.025 2.984 6.03 3.238 ;
      RECT 6.015 2.983 6.025 3.205 ;
      RECT 5.965 2.981 6.015 3.19 ;
      RECT 5.94 2.979 5.965 3.185 ;
      RECT 5.897 2.977 5.94 3.181 ;
      RECT 5.811 2.973 5.897 3.169 ;
      RECT 5.725 2.968 5.811 3.153 ;
      RECT 5.695 2.965 5.725 3.14 ;
      RECT 5.67 2.964 5.695 3.128 ;
      RECT 5.665 2.964 5.67 3.118 ;
      RECT 5.625 2.963 5.665 3.11 ;
      RECT 5.61 2.962 5.625 3.103 ;
      RECT 5.56 2.961 5.61 3.095 ;
      RECT 5.558 2.96 5.56 3.09 ;
      RECT 5.472 2.958 5.558 3.09 ;
      RECT 5.386 2.953 5.472 3.09 ;
      RECT 5.3 2.949 5.386 3.09 ;
      RECT 5.251 2.945 5.3 3.088 ;
      RECT 5.165 2.942 5.251 3.083 ;
      RECT 5.142 2.939 5.165 3.079 ;
      RECT 5.056 2.936 5.142 3.074 ;
      RECT 4.97 2.932 5.056 3.065 ;
      RECT 4.945 2.925 4.97 3.06 ;
      RECT 4.885 2.89 4.945 3.057 ;
      RECT 4.865 2.815 4.885 3.054 ;
      RECT 4.86 2.757 4.865 3.053 ;
      RECT 4.835 2.697 4.86 3.052 ;
      RECT 4.76 2.575 4.835 3.048 ;
      RECT 4.75 2.575 4.76 3.04 ;
      RECT 4.735 2.575 4.75 3.03 ;
      RECT 4.72 2.575 4.735 3 ;
      RECT 4.705 2.575 4.72 2.945 ;
      RECT 4.69 2.575 4.705 2.883 ;
      RECT 4.665 2.575 4.69 2.808 ;
      RECT 4.66 2.575 4.665 2.758 ;
      RECT 6.005 2.12 6.025 2.429 ;
      RECT 5.991 2.122 6.04 2.426 ;
      RECT 5.991 2.127 6.06 2.417 ;
      RECT 5.905 2.125 6.04 2.411 ;
      RECT 5.905 2.133 6.095 2.394 ;
      RECT 5.87 2.135 6.095 2.393 ;
      RECT 5.84 2.143 6.095 2.384 ;
      RECT 5.83 2.148 6.115 2.37 ;
      RECT 5.87 2.138 6.115 2.37 ;
      RECT 5.87 2.141 6.125 2.358 ;
      RECT 5.84 2.143 6.135 2.345 ;
      RECT 5.84 2.147 6.145 2.288 ;
      RECT 5.83 2.152 6.15 2.203 ;
      RECT 5.991 2.12 6.025 2.426 ;
      RECT 5.87 7.855 6.04 8.305 ;
      RECT 5.925 6.075 6.095 8.025 ;
      RECT 5.87 5.015 6.04 6.245 ;
      RECT 5.43 2.223 5.435 2.435 ;
      RECT 5.305 2.22 5.32 2.435 ;
      RECT 4.77 2.25 4.84 2.435 ;
      RECT 4.655 2.25 4.69 2.43 ;
      RECT 5.776 2.552 5.795 2.746 ;
      RECT 5.69 2.507 5.776 2.747 ;
      RECT 5.68 2.46 5.69 2.749 ;
      RECT 5.675 2.44 5.68 2.75 ;
      RECT 5.655 2.405 5.675 2.751 ;
      RECT 5.64 2.355 5.655 2.752 ;
      RECT 5.62 2.292 5.64 2.753 ;
      RECT 5.61 2.255 5.62 2.754 ;
      RECT 5.595 2.244 5.61 2.755 ;
      RECT 5.59 2.236 5.595 2.753 ;
      RECT 5.58 2.235 5.59 2.745 ;
      RECT 5.55 2.232 5.58 2.724 ;
      RECT 5.475 2.227 5.55 2.669 ;
      RECT 5.46 2.223 5.475 2.615 ;
      RECT 5.45 2.223 5.46 2.51 ;
      RECT 5.435 2.223 5.45 2.443 ;
      RECT 5.42 2.223 5.43 2.433 ;
      RECT 5.365 2.222 5.42 2.43 ;
      RECT 5.32 2.22 5.365 2.433 ;
      RECT 5.292 2.22 5.305 2.436 ;
      RECT 5.206 2.224 5.292 2.438 ;
      RECT 5.12 2.23 5.206 2.443 ;
      RECT 5.1 2.234 5.12 2.445 ;
      RECT 5.098 2.235 5.1 2.444 ;
      RECT 5.012 2.237 5.098 2.443 ;
      RECT 4.926 2.242 5.012 2.44 ;
      RECT 4.84 2.247 4.926 2.437 ;
      RECT 4.69 2.25 4.77 2.433 ;
      RECT 5.35 5.015 5.52 8.305 ;
      RECT 5.35 7.315 5.755 7.645 ;
      RECT 5.35 6.475 5.755 6.805 ;
      RECT 5.466 3.225 5.515 3.559 ;
      RECT 5.466 3.225 5.52 3.558 ;
      RECT 5.38 3.225 5.52 3.557 ;
      RECT 5.155 3.333 5.525 3.555 ;
      RECT 5.38 3.225 5.55 3.548 ;
      RECT 5.35 3.237 5.555 3.539 ;
      RECT 5.335 3.255 5.56 3.536 ;
      RECT 5.15 3.339 5.56 3.463 ;
      RECT 5.145 3.346 5.56 3.423 ;
      RECT 5.16 3.312 5.56 3.536 ;
      RECT 5.321 3.258 5.525 3.555 ;
      RECT 5.235 3.278 5.56 3.536 ;
      RECT 5.335 3.252 5.555 3.539 ;
      RECT 5.105 2.576 5.295 2.77 ;
      RECT 5.1 2.578 5.295 2.769 ;
      RECT 5.095 2.582 5.31 2.766 ;
      RECT 5.11 2.575 5.31 2.766 ;
      RECT 5.095 2.685 5.315 2.761 ;
      RECT 4.39 3.185 4.481 3.483 ;
      RECT 4.385 3.187 4.56 3.478 ;
      RECT 4.39 3.185 4.56 3.478 ;
      RECT 4.385 3.191 4.58 3.476 ;
      RECT 4.385 3.246 4.62 3.475 ;
      RECT 4.385 3.281 4.635 3.469 ;
      RECT 4.385 3.315 4.645 3.459 ;
      RECT 4.375 3.195 4.58 3.31 ;
      RECT 4.375 3.215 4.595 3.31 ;
      RECT 4.375 3.198 4.585 3.31 ;
      RECT 4.6 1.966 4.605 2.028 ;
      RECT 4.595 1.888 4.6 2.051 ;
      RECT 4.59 1.845 4.595 2.062 ;
      RECT 4.585 1.835 4.59 2.074 ;
      RECT 4.58 1.835 4.585 2.083 ;
      RECT 4.555 1.835 4.58 2.115 ;
      RECT 4.55 1.835 4.555 2.148 ;
      RECT 4.535 1.835 4.55 2.173 ;
      RECT 4.525 1.835 4.535 2.2 ;
      RECT 4.52 1.835 4.525 2.213 ;
      RECT 4.515 1.835 4.52 2.228 ;
      RECT 4.505 1.835 4.515 2.243 ;
      RECT 4.5 1.835 4.505 2.263 ;
      RECT 4.475 1.835 4.5 2.298 ;
      RECT 4.43 1.835 4.475 2.343 ;
      RECT 4.42 1.835 4.43 2.356 ;
      RECT 4.335 1.92 4.42 2.363 ;
      RECT 4.3 2.042 4.335 2.372 ;
      RECT 4.295 2.082 4.3 2.376 ;
      RECT 4.275 2.105 4.295 2.378 ;
      RECT 4.27 2.135 4.275 2.381 ;
      RECT 4.26 2.147 4.27 2.382 ;
      RECT 4.215 2.17 4.26 2.387 ;
      RECT 4.175 2.2 4.215 2.395 ;
      RECT 4.14 2.212 4.175 2.401 ;
      RECT 4.135 2.217 4.14 2.405 ;
      RECT 4.065 2.227 4.135 2.412 ;
      RECT 4.025 2.237 4.065 2.422 ;
      RECT 4.005 2.242 4.025 2.428 ;
      RECT 3.995 2.246 4.005 2.433 ;
      RECT 3.99 2.249 3.995 2.436 ;
      RECT 3.98 2.25 3.99 2.437 ;
      RECT 3.955 2.252 3.98 2.441 ;
      RECT 3.945 2.257 3.955 2.444 ;
      RECT 3.9 2.265 3.945 2.445 ;
      RECT 3.775 2.27 3.9 2.445 ;
      RECT 4.33 2.567 4.35 2.749 ;
      RECT 4.281 2.552 4.33 2.748 ;
      RECT 4.195 2.567 4.35 2.746 ;
      RECT 4.18 2.567 4.35 2.745 ;
      RECT 4.145 2.545 4.315 2.73 ;
      RECT 4.215 3.565 4.23 3.774 ;
      RECT 4.215 3.573 4.235 3.773 ;
      RECT 4.16 3.573 4.235 3.772 ;
      RECT 4.14 3.577 4.24 3.77 ;
      RECT 4.12 3.527 4.16 3.769 ;
      RECT 4.065 3.585 4.245 3.767 ;
      RECT 4.03 3.542 4.16 3.765 ;
      RECT 4.026 3.545 4.215 3.764 ;
      RECT 3.94 3.553 4.215 3.762 ;
      RECT 3.94 3.597 4.25 3.755 ;
      RECT 3.93 3.69 4.25 3.753 ;
      RECT 3.94 3.609 4.255 3.738 ;
      RECT 3.94 3.63 4.27 3.708 ;
      RECT 3.94 3.657 4.275 3.678 ;
      RECT 4.065 3.535 4.16 3.767 ;
      RECT 3.695 2.58 3.7 3.118 ;
      RECT 3.5 2.91 3.505 3.105 ;
      RECT 1.8 2.575 1.815 2.955 ;
      RECT 3.865 2.575 3.87 2.745 ;
      RECT 3.86 2.575 3.865 2.755 ;
      RECT 3.855 2.575 3.86 2.768 ;
      RECT 3.83 2.575 3.855 2.81 ;
      RECT 3.805 2.575 3.83 2.883 ;
      RECT 3.79 2.575 3.805 2.935 ;
      RECT 3.785 2.575 3.79 2.965 ;
      RECT 3.76 2.575 3.785 3.005 ;
      RECT 3.745 2.575 3.76 3.06 ;
      RECT 3.74 2.575 3.745 3.093 ;
      RECT 3.715 2.575 3.74 3.113 ;
      RECT 3.7 2.575 3.715 3.119 ;
      RECT 3.63 2.61 3.695 3.115 ;
      RECT 3.58 2.665 3.63 3.11 ;
      RECT 3.57 2.697 3.58 3.108 ;
      RECT 3.565 2.722 3.57 3.108 ;
      RECT 3.545 2.795 3.565 3.108 ;
      RECT 3.535 2.875 3.545 3.107 ;
      RECT 3.52 2.905 3.535 3.107 ;
      RECT 3.505 2.91 3.52 3.106 ;
      RECT 3.445 2.912 3.5 3.103 ;
      RECT 3.415 2.917 3.445 3.099 ;
      RECT 3.413 2.92 3.415 3.098 ;
      RECT 3.327 2.922 3.413 3.095 ;
      RECT 3.241 2.928 3.327 3.089 ;
      RECT 3.155 2.933 3.241 3.083 ;
      RECT 3.082 2.938 3.155 3.084 ;
      RECT 2.996 2.944 3.082 3.092 ;
      RECT 2.91 2.95 2.996 3.101 ;
      RECT 2.89 2.954 2.91 3.106 ;
      RECT 2.843 2.956 2.89 3.109 ;
      RECT 2.757 2.961 2.843 3.115 ;
      RECT 2.671 2.966 2.757 3.124 ;
      RECT 2.585 2.972 2.671 3.132 ;
      RECT 2.5 2.97 2.585 3.141 ;
      RECT 2.496 2.965 2.5 3.145 ;
      RECT 2.41 2.96 2.496 3.137 ;
      RECT 2.346 2.951 2.41 3.125 ;
      RECT 2.26 2.942 2.346 3.112 ;
      RECT 2.236 2.935 2.26 3.103 ;
      RECT 2.15 2.929 2.236 3.09 ;
      RECT 2.11 2.922 2.15 3.076 ;
      RECT 2.105 2.912 2.11 3.072 ;
      RECT 2.095 2.9 2.105 3.071 ;
      RECT 2.075 2.87 2.095 3.068 ;
      RECT 2.02 2.79 2.075 3.062 ;
      RECT 2 2.709 2.02 3.057 ;
      RECT 1.98 2.667 2 3.053 ;
      RECT 1.955 2.62 1.98 3.047 ;
      RECT 1.95 2.595 1.955 3.044 ;
      RECT 1.915 2.575 1.95 3.039 ;
      RECT 1.906 2.575 1.915 3.032 ;
      RECT 1.82 2.575 1.906 3.002 ;
      RECT 1.815 2.575 1.82 2.965 ;
      RECT 1.78 2.575 1.8 2.887 ;
      RECT 1.775 2.617 1.78 2.852 ;
      RECT 1.77 2.692 1.775 2.808 ;
      RECT 3.22 2.497 3.395 2.745 ;
      RECT 3.22 2.497 3.4 2.743 ;
      RECT 3.215 2.529 3.4 2.703 ;
      RECT 3.245 2.47 3.415 2.69 ;
      RECT 3.21 2.547 3.415 2.623 ;
      RECT 2.52 2.01 2.69 2.185 ;
      RECT 2.52 2.01 2.862 2.177 ;
      RECT 2.52 2.01 2.945 2.171 ;
      RECT 2.52 2.01 2.98 2.167 ;
      RECT 2.52 2.01 3 2.166 ;
      RECT 2.52 2.01 3.086 2.162 ;
      RECT 2.98 1.835 3.15 2.157 ;
      RECT 2.555 1.942 3.18 2.155 ;
      RECT 2.545 1.997 3.185 2.153 ;
      RECT 2.52 2.033 3.195 2.148 ;
      RECT 2.52 2.06 3.2 2.078 ;
      RECT 2.585 1.885 3.16 2.155 ;
      RECT 2.776 1.87 3.16 2.155 ;
      RECT 2.61 1.873 3.16 2.155 ;
      RECT 2.69 1.871 2.776 2.182 ;
      RECT 2.776 1.868 3.155 2.155 ;
      RECT 2.96 1.845 3.155 2.155 ;
      RECT 2.862 1.866 3.155 2.155 ;
      RECT 2.945 1.86 2.96 2.168 ;
      RECT 3.095 3.225 3.1 3.425 ;
      RECT 2.56 3.29 2.605 3.425 ;
      RECT 3.13 3.225 3.15 3.398 ;
      RECT 3.1 3.225 3.13 3.413 ;
      RECT 3.035 3.225 3.095 3.45 ;
      RECT 3.02 3.225 3.035 3.48 ;
      RECT 3.005 3.225 3.02 3.493 ;
      RECT 2.985 3.225 3.005 3.508 ;
      RECT 2.98 3.225 2.985 3.517 ;
      RECT 2.97 3.229 2.98 3.522 ;
      RECT 2.955 3.239 2.97 3.533 ;
      RECT 2.93 3.255 2.955 3.543 ;
      RECT 2.92 3.269 2.93 3.545 ;
      RECT 2.9 3.281 2.92 3.542 ;
      RECT 2.87 3.302 2.9 3.536 ;
      RECT 2.86 3.314 2.87 3.531 ;
      RECT 2.85 3.312 2.86 3.528 ;
      RECT 2.835 3.311 2.85 3.523 ;
      RECT 2.83 3.31 2.835 3.518 ;
      RECT 2.795 3.308 2.83 3.508 ;
      RECT 2.775 3.305 2.795 3.49 ;
      RECT 2.765 3.303 2.775 3.485 ;
      RECT 2.755 3.302 2.765 3.48 ;
      RECT 2.72 3.3 2.755 3.468 ;
      RECT 2.665 3.296 2.72 3.448 ;
      RECT 2.655 3.294 2.665 3.433 ;
      RECT 2.65 3.294 2.655 3.428 ;
      RECT 2.605 3.292 2.65 3.425 ;
      RECT 2.51 3.29 2.56 3.429 ;
      RECT 2.5 3.291 2.51 3.434 ;
      RECT 2.44 3.298 2.5 3.448 ;
      RECT 2.415 3.306 2.44 3.468 ;
      RECT 2.405 3.31 2.415 3.48 ;
      RECT 2.4 3.311 2.405 3.485 ;
      RECT 2.385 3.313 2.4 3.488 ;
      RECT 2.37 3.315 2.385 3.493 ;
      RECT 2.365 3.315 2.37 3.496 ;
      RECT 2.32 3.32 2.365 3.507 ;
      RECT 2.315 3.324 2.32 3.519 ;
      RECT 2.29 3.32 2.315 3.523 ;
      RECT 2.28 3.316 2.29 3.527 ;
      RECT 2.27 3.315 2.28 3.531 ;
      RECT 2.255 3.305 2.27 3.537 ;
      RECT 2.25 3.293 2.255 3.541 ;
      RECT 2.245 3.29 2.25 3.542 ;
      RECT 2.24 3.287 2.245 3.544 ;
      RECT 2.225 3.275 2.24 3.543 ;
      RECT 2.21 3.257 2.225 3.54 ;
      RECT 2.19 3.236 2.21 3.533 ;
      RECT 2.125 3.225 2.19 3.505 ;
      RECT 2.121 3.225 2.125 3.484 ;
      RECT 2.035 3.225 2.121 3.454 ;
      RECT 2.02 3.225 2.035 3.41 ;
      RECT 2.595 2.325 2.6 2.56 ;
      RECT 1.725 2.241 1.73 2.445 ;
      RECT 2.305 2.27 2.31 2.425 ;
      RECT 2.225 2.25 2.23 2.425 ;
      RECT 2.895 2.392 2.91 2.745 ;
      RECT 2.821 2.377 2.895 2.745 ;
      RECT 2.735 2.36 2.821 2.745 ;
      RECT 2.725 2.35 2.735 2.743 ;
      RECT 2.72 2.348 2.725 2.738 ;
      RECT 2.705 2.346 2.72 2.724 ;
      RECT 2.635 2.338 2.705 2.664 ;
      RECT 2.615 2.329 2.635 2.598 ;
      RECT 2.61 2.326 2.615 2.578 ;
      RECT 2.6 2.325 2.61 2.568 ;
      RECT 2.59 2.325 2.595 2.552 ;
      RECT 2.58 2.324 2.59 2.542 ;
      RECT 2.57 2.322 2.58 2.53 ;
      RECT 2.555 2.319 2.57 2.51 ;
      RECT 2.545 2.317 2.555 2.495 ;
      RECT 2.525 2.314 2.545 2.483 ;
      RECT 2.52 2.312 2.525 2.473 ;
      RECT 2.495 2.31 2.52 2.46 ;
      RECT 2.465 2.305 2.495 2.445 ;
      RECT 2.385 2.296 2.465 2.436 ;
      RECT 2.34 2.285 2.385 2.429 ;
      RECT 2.32 2.276 2.34 2.426 ;
      RECT 2.31 2.271 2.32 2.425 ;
      RECT 2.265 2.265 2.305 2.425 ;
      RECT 2.25 2.257 2.265 2.425 ;
      RECT 2.23 2.252 2.25 2.425 ;
      RECT 2.21 2.249 2.225 2.425 ;
      RECT 2.127 2.248 2.21 2.424 ;
      RECT 2.041 2.247 2.127 2.42 ;
      RECT 1.955 2.245 2.041 2.417 ;
      RECT 1.902 2.244 1.955 2.419 ;
      RECT 1.816 2.243 1.902 2.428 ;
      RECT 1.73 2.242 1.816 2.44 ;
      RECT 1.71 2.241 1.725 2.448 ;
      RECT 1.63 2.24 1.71 2.46 ;
      RECT 1.605 2.24 1.63 2.473 ;
      RECT 1.58 2.24 1.605 2.488 ;
      RECT 1.575 2.24 1.58 2.51 ;
      RECT 1.57 2.24 1.575 2.528 ;
      RECT 1.565 2.24 1.57 2.545 ;
      RECT 1.56 2.24 1.565 2.558 ;
      RECT 1.555 2.24 1.56 2.568 ;
      RECT 1.515 2.24 1.555 2.653 ;
      RECT 1.5 2.24 1.515 2.738 ;
      RECT 1.49 2.241 1.5 2.75 ;
      RECT 1.455 2.246 1.49 2.755 ;
      RECT 1.415 2.255 1.455 2.755 ;
      RECT 1.4 2.265 1.415 2.755 ;
      RECT 1.395 2.275 1.4 2.755 ;
      RECT 1.375 2.302 1.395 2.755 ;
      RECT 1.325 2.385 1.375 2.755 ;
      RECT 1.32 2.447 1.325 2.755 ;
      RECT 1.31 2.46 1.32 2.755 ;
      RECT 1.3 2.482 1.31 2.755 ;
      RECT 1.29 2.507 1.3 2.75 ;
      RECT 1.285 2.545 1.29 2.743 ;
      RECT 1.275 2.655 1.285 2.738 ;
      RECT 2.67 3.576 2.685 3.835 ;
      RECT 2.67 3.591 2.69 3.834 ;
      RECT 2.586 3.591 2.69 3.832 ;
      RECT 2.586 3.605 2.695 3.831 ;
      RECT 2.5 3.647 2.7 3.828 ;
      RECT 2.495 3.59 2.685 3.823 ;
      RECT 2.495 3.661 2.705 3.82 ;
      RECT 2.49 3.692 2.705 3.818 ;
      RECT 2.495 3.689 2.72 3.808 ;
      RECT 2.49 3.735 2.735 3.793 ;
      RECT 2.49 3.763 2.74 3.778 ;
      RECT 2.5 3.565 2.67 3.828 ;
      RECT 2.26 2.575 2.43 2.745 ;
      RECT 2.225 2.575 2.43 2.74 ;
      RECT 2.215 2.575 2.43 2.733 ;
      RECT 2.21 2.56 2.38 2.73 ;
      RECT 1.04 3.097 1.305 3.54 ;
      RECT 1.035 3.068 1.25 3.538 ;
      RECT 1.03 3.222 1.31 3.533 ;
      RECT 1.035 3.117 1.31 3.533 ;
      RECT 1.035 3.128 1.32 3.52 ;
      RECT 1.035 3.075 1.28 3.538 ;
      RECT 1.04 3.062 1.25 3.54 ;
      RECT 1.04 3.06 1.2 3.54 ;
      RECT 1.141 3.052 1.2 3.54 ;
      RECT 1.055 3.053 1.2 3.54 ;
      RECT 1.141 3.051 1.19 3.54 ;
      RECT 0.945 1.866 1.12 2.165 ;
      RECT 0.995 1.828 1.12 2.165 ;
      RECT 0.98 1.83 1.206 2.157 ;
      RECT 0.98 1.833 1.245 2.144 ;
      RECT 0.98 1.834 1.255 2.13 ;
      RECT 0.935 1.885 1.255 2.12 ;
      RECT 0.98 1.835 1.26 2.115 ;
      RECT 0.935 2.045 1.265 2.105 ;
      RECT 0.92 1.905 1.26 2.045 ;
      RECT 0.915 1.921 1.26 1.985 ;
      RECT 0.96 1.845 1.26 2.115 ;
      RECT 0.995 1.826 1.081 2.165 ;
      RECT -1.625 7.855 -1.455 8.305 ;
      RECT -1.57 6.075 -1.4 8.025 ;
      RECT -1.625 5.015 -1.455 6.245 ;
      RECT -2.145 5.015 -1.975 8.305 ;
      RECT -2.145 7.315 -1.74 7.645 ;
      RECT -2.145 6.475 -1.74 6.805 ;
      RECT 75.76 0.575 75.93 1.085 ;
      RECT 75.76 2.395 75.93 3.865 ;
      RECT 75.76 5.015 75.93 6.485 ;
      RECT 75.76 7.795 75.93 8.305 ;
      RECT 74.77 0.575 74.94 1.085 ;
      RECT 74.77 2.395 74.94 3.865 ;
      RECT 74.77 5.015 74.94 6.485 ;
      RECT 74.77 7.795 74.94 8.305 ;
      RECT 73.405 0.575 73.575 3.865 ;
      RECT 73.405 5.015 73.575 8.305 ;
      RECT 72.975 0.575 73.145 1.085 ;
      RECT 72.975 1.655 73.145 3.865 ;
      RECT 72.975 5.015 73.145 7.225 ;
      RECT 72.975 7.795 73.145 8.305 ;
      RECT 71.605 1.66 71.775 2.935 ;
      RECT 71.605 5.945 71.775 7.22 ;
      RECT 67.77 5.015 67.94 8.305 ;
      RECT 67.34 5.015 67.51 7.225 ;
      RECT 67.34 7.795 67.51 8.305 ;
      RECT 65.97 5.945 66.14 7.22 ;
      RECT 60.5 0.575 60.67 1.085 ;
      RECT 60.5 2.395 60.67 3.865 ;
      RECT 60.5 5.015 60.67 6.485 ;
      RECT 60.5 7.795 60.67 8.305 ;
      RECT 59.51 0.575 59.68 1.085 ;
      RECT 59.51 2.395 59.68 3.865 ;
      RECT 59.51 5.015 59.68 6.485 ;
      RECT 59.51 7.795 59.68 8.305 ;
      RECT 58.145 0.575 58.315 3.865 ;
      RECT 58.145 5.015 58.315 8.305 ;
      RECT 57.715 0.575 57.885 1.085 ;
      RECT 57.715 1.655 57.885 3.865 ;
      RECT 57.715 5.015 57.885 7.225 ;
      RECT 57.715 7.795 57.885 8.305 ;
      RECT 56.345 1.66 56.515 2.935 ;
      RECT 56.345 5.945 56.515 7.22 ;
      RECT 52.51 5.015 52.68 8.305 ;
      RECT 52.08 5.015 52.25 7.225 ;
      RECT 52.08 7.795 52.25 8.305 ;
      RECT 50.71 5.945 50.88 7.22 ;
      RECT 45.24 0.575 45.41 1.085 ;
      RECT 45.24 2.395 45.41 3.865 ;
      RECT 45.24 5.015 45.41 6.485 ;
      RECT 45.24 7.795 45.41 8.305 ;
      RECT 44.25 0.575 44.42 1.085 ;
      RECT 44.25 2.395 44.42 3.865 ;
      RECT 44.25 5.015 44.42 6.485 ;
      RECT 44.25 7.795 44.42 8.305 ;
      RECT 42.885 0.575 43.055 3.865 ;
      RECT 42.885 5.015 43.055 8.305 ;
      RECT 42.455 0.575 42.625 1.085 ;
      RECT 42.455 1.655 42.625 3.865 ;
      RECT 42.455 5.015 42.625 7.225 ;
      RECT 42.455 7.795 42.625 8.305 ;
      RECT 41.085 1.66 41.255 2.935 ;
      RECT 41.085 5.945 41.255 7.22 ;
      RECT 37.25 5.015 37.42 8.305 ;
      RECT 36.82 5.015 36.99 7.225 ;
      RECT 36.82 7.795 36.99 8.305 ;
      RECT 35.45 5.945 35.62 7.22 ;
      RECT 29.98 0.575 30.15 1.085 ;
      RECT 29.98 2.395 30.15 3.865 ;
      RECT 29.98 5.015 30.15 6.485 ;
      RECT 29.98 7.795 30.15 8.305 ;
      RECT 28.99 0.575 29.16 1.085 ;
      RECT 28.99 2.395 29.16 3.865 ;
      RECT 28.99 5.015 29.16 6.485 ;
      RECT 28.99 7.795 29.16 8.305 ;
      RECT 27.625 0.575 27.795 3.865 ;
      RECT 27.625 5.015 27.795 8.305 ;
      RECT 27.195 0.575 27.365 1.085 ;
      RECT 27.195 1.655 27.365 3.865 ;
      RECT 27.195 5.015 27.365 7.225 ;
      RECT 27.195 7.795 27.365 8.305 ;
      RECT 25.825 1.66 25.995 2.935 ;
      RECT 25.825 5.945 25.995 7.22 ;
      RECT 21.99 5.015 22.16 8.305 ;
      RECT 21.56 5.015 21.73 7.225 ;
      RECT 21.56 7.795 21.73 8.305 ;
      RECT 20.19 5.945 20.36 7.22 ;
      RECT 14.72 0.575 14.89 1.085 ;
      RECT 14.72 2.395 14.89 3.865 ;
      RECT 14.72 5.015 14.89 6.485 ;
      RECT 14.72 7.795 14.89 8.305 ;
      RECT 13.73 0.575 13.9 1.085 ;
      RECT 13.73 2.395 13.9 3.865 ;
      RECT 13.73 5.015 13.9 6.485 ;
      RECT 13.73 7.795 13.9 8.305 ;
      RECT 12.365 0.575 12.535 3.865 ;
      RECT 12.365 5.015 12.535 8.305 ;
      RECT 11.935 0.575 12.105 1.085 ;
      RECT 11.935 1.655 12.105 3.865 ;
      RECT 11.935 5.015 12.105 7.225 ;
      RECT 11.935 7.795 12.105 8.305 ;
      RECT 10.565 1.66 10.735 2.935 ;
      RECT 10.565 5.945 10.735 7.22 ;
      RECT 6.73 5.015 6.9 8.305 ;
      RECT 6.3 5.015 6.47 7.225 ;
      RECT 6.3 7.795 6.47 8.305 ;
      RECT 4.93 5.945 5.1 7.22 ;
      RECT -1.195 5.015 -1.025 7.225 ;
      RECT -1.195 7.795 -1.025 8.305 ;
      RECT -2.565 5.945 -2.395 7.22 ;
  END
END sky130_osu_ring_oscillator_mpr2ya_8_b0r2

END LIBRARY
