magic
tech sky130A
magscale 1 2
timestamp 1715040497
<< nwell >>
rect 252441 702384 252880 702819
rect 324443 702424 324882 702859
rect 360475 701955 360914 702390
rect 432435 701818 432874 702253
rect 504430 701572 504869 702007
rect 576278 697362 576717 697797
rect 576278 644186 576717 644621
rect 576278 591146 576717 591581
rect 504184 554054 504623 554489
rect 576278 537970 576717 538405
rect 576278 484794 576717 485229
rect 576278 431754 576717 432189
rect 576278 378578 576717 379013
rect 576278 325402 576717 325837
rect 576278 272362 576717 272797
rect 576278 232515 576717 232950
<< nsubdiff >>
rect 324481 702558 324505 702592
rect 324539 702558 324565 702592
rect 252479 702518 252503 702552
rect 252537 702518 252563 702552
rect 360513 702089 360537 702123
rect 360571 702089 360597 702123
rect 432473 701952 432497 701986
rect 432531 701952 432557 701986
rect 504468 701706 504492 701740
rect 504526 701706 504552 701740
rect 576316 697629 576340 697663
rect 576374 697629 576400 697663
rect 576316 644453 576340 644487
rect 576374 644453 576400 644487
rect 576316 591413 576340 591447
rect 576374 591413 576400 591447
rect 504222 554321 504246 554355
rect 504280 554321 504306 554355
rect 576316 538237 576340 538271
rect 576374 538237 576400 538271
rect 576316 485061 576340 485095
rect 576374 485061 576400 485095
rect 576316 432021 576340 432055
rect 576374 432021 576400 432055
rect 576316 378845 576340 378879
rect 576374 378845 576400 378879
rect 576316 325669 576340 325703
rect 576374 325669 576400 325703
rect 576316 272629 576340 272663
rect 576374 272629 576400 272663
rect 576316 232782 576340 232816
rect 576374 232782 576400 232816
<< nsubdiffcont >>
rect 324505 702558 324539 702592
rect 252503 702518 252537 702552
rect 360537 702089 360571 702123
rect 432497 701952 432531 701986
rect 504492 701706 504526 701740
rect 576340 697629 576374 697663
rect 576340 644453 576374 644487
rect 576340 591413 576374 591447
rect 504246 554321 504280 554355
rect 576340 538237 576374 538271
rect 576340 485061 576374 485095
rect 576340 432021 576374 432055
rect 576340 378845 576374 378879
rect 576340 325669 576374 325703
rect 576340 272629 576374 272663
rect 576340 232782 576374 232816
<< poly >>
rect 324733 702703 324783 702710
rect 252734 702663 252784 702673
rect 252734 702611 252785 702663
rect 324733 702651 324784 702703
rect 324733 702645 324783 702651
rect 252734 702604 252784 702611
rect 360760 702234 360810 702243
rect 360760 702182 360811 702234
rect 360760 702174 360810 702182
rect 432730 702097 432780 702105
rect 432730 702045 432781 702097
rect 432730 702036 432780 702045
rect 504726 701851 504776 701862
rect 504726 701799 504777 701851
rect 504726 701792 504776 701799
<< locali >>
rect 324729 702703 324783 702710
rect 324729 702692 324784 702703
rect 252730 702663 252784 702673
rect 252730 702652 252785 702663
rect 252730 702618 252742 702652
rect 252776 702618 252785 702652
rect 324729 702658 324741 702692
rect 324775 702658 324784 702692
rect 324729 702651 324784 702658
rect 324729 702645 324783 702651
rect 252730 702611 252785 702618
rect 252730 702604 252784 702611
rect 324481 702558 324505 702592
rect 324539 702558 324565 702592
rect 252479 702518 252503 702552
rect 252537 702518 252563 702552
rect 360756 702234 360810 702243
rect 360756 702223 360811 702234
rect 360756 702189 360768 702223
rect 360802 702189 360811 702223
rect 360756 702182 360811 702189
rect 360756 702174 360810 702182
rect 360513 702089 360537 702123
rect 360571 702089 360597 702123
rect 432726 702097 432780 702105
rect 432726 702086 432781 702097
rect 432726 702052 432738 702086
rect 432772 702052 432781 702086
rect 432726 702045 432781 702052
rect 432726 702036 432780 702045
rect 432473 701952 432497 701986
rect 432531 701952 432557 701986
rect 504722 701851 504776 701862
rect 504722 701840 504777 701851
rect 504722 701806 504734 701840
rect 504768 701806 504777 701840
rect 504722 701799 504777 701806
rect 504722 701792 504776 701799
rect 504468 701706 504492 701740
rect 504526 701706 504552 701740
rect 576316 697629 576340 697663
rect 576374 697629 576400 697663
rect 576316 644453 576340 644487
rect 576374 644453 576400 644487
rect 576316 591413 576340 591447
rect 576374 591413 576400 591447
rect 504222 554321 504246 554355
rect 504280 554321 504306 554355
rect 576316 538237 576340 538271
rect 576374 538237 576400 538271
rect 576316 485061 576340 485095
rect 576374 485061 576400 485095
rect 576316 432021 576340 432055
rect 576374 432021 576400 432055
rect 576316 378845 576340 378879
rect 576374 378845 576400 378879
rect 576316 325669 576340 325703
rect 576374 325669 576400 325703
rect 576316 272629 576340 272663
rect 576374 272629 576400 272663
rect 576316 232782 576340 232816
rect 576374 232782 576400 232816
<< viali >>
rect 252742 702618 252776 702652
rect 324741 702658 324775 702692
rect 360768 702189 360802 702223
rect 432738 702052 432772 702086
rect 504734 701806 504768 701840
rect 576613 697187 576647 697221
rect 576613 644011 576647 644045
rect 576613 590971 576647 591005
rect 504519 554015 504553 554049
rect 576613 537795 576647 537829
rect 576613 484619 576647 484653
rect 576613 431579 576647 431613
rect 478943 431411 478977 431445
rect 485831 431411 485865 431445
rect 478581 410399 478615 410433
rect 485111 410399 485145 410433
rect 479474 389455 479508 389489
rect 490610 389455 490644 389489
rect 576613 378403 576647 378437
rect 477091 356815 477125 356849
rect 480143 356815 480177 356849
rect 482075 340835 482109 340869
rect 475442 340359 475476 340393
rect 478759 340359 478793 340393
rect 576613 325227 576647 325261
rect 478939 320367 478973 320401
rect 485827 320367 485861 320401
rect 478580 305407 478614 305441
rect 485110 305407 485144 305441
rect 490610 285959 490644 285993
rect 479474 285823 479508 285857
rect 576613 272187 576647 272221
rect 477101 265831 477135 265865
rect 576613 232340 576647 232374
<< metal1 >>
rect 326234 703378 326854 703384
rect 254234 703338 254854 703344
rect 254234 703286 254262 703338
rect 254314 703286 254326 703338
rect 254378 703286 254390 703338
rect 254442 703286 254454 703338
rect 254506 703286 254518 703338
rect 254570 703286 254582 703338
rect 254634 703286 254646 703338
rect 254698 703286 254710 703338
rect 254762 703286 254774 703338
rect 254826 703286 254854 703338
rect 254234 703274 254854 703286
rect 254234 703222 254262 703274
rect 254314 703222 254326 703274
rect 254378 703222 254390 703274
rect 254442 703222 254454 703274
rect 254506 703222 254518 703274
rect 254570 703222 254582 703274
rect 254634 703222 254646 703274
rect 254698 703222 254710 703274
rect 254762 703222 254774 703274
rect 254826 703222 254854 703274
rect 254234 703210 254854 703222
rect 254234 703158 254262 703210
rect 254314 703158 254326 703210
rect 254378 703158 254390 703210
rect 254442 703158 254454 703210
rect 254506 703158 254518 703210
rect 254570 703158 254582 703210
rect 254634 703158 254646 703210
rect 254698 703158 254710 703210
rect 254762 703158 254774 703210
rect 254826 703158 254854 703210
rect 326234 703326 326262 703378
rect 326314 703326 326326 703378
rect 326378 703326 326390 703378
rect 326442 703326 326454 703378
rect 326506 703326 326518 703378
rect 326570 703326 326582 703378
rect 326634 703326 326646 703378
rect 326698 703326 326710 703378
rect 326762 703326 326774 703378
rect 326826 703326 326854 703378
rect 326234 703314 326854 703326
rect 326234 703262 326262 703314
rect 326314 703262 326326 703314
rect 326378 703262 326390 703314
rect 326442 703262 326454 703314
rect 326506 703262 326518 703314
rect 326570 703262 326582 703314
rect 326634 703262 326646 703314
rect 326698 703262 326710 703314
rect 326762 703262 326774 703314
rect 326826 703262 326854 703314
rect 326234 703250 326854 703262
rect 326234 703198 326262 703250
rect 326314 703198 326326 703250
rect 326378 703198 326390 703250
rect 326442 703198 326454 703250
rect 326506 703198 326518 703250
rect 326570 703198 326582 703250
rect 326634 703198 326646 703250
rect 326698 703198 326710 703250
rect 326762 703198 326774 703250
rect 326826 703198 326854 703250
rect 326234 703186 326854 703198
rect 326234 703160 326262 703186
rect 254234 703146 254854 703158
rect 254234 703120 254262 703146
rect 252794 703094 254262 703120
rect 254314 703094 254326 703146
rect 254378 703094 254390 703146
rect 254442 703094 254454 703146
rect 254506 703094 254518 703146
rect 254570 703094 254582 703146
rect 254634 703094 254646 703146
rect 254698 703094 254710 703146
rect 254762 703094 254774 703146
rect 254826 703120 254854 703146
rect 324796 703134 326262 703160
rect 326314 703134 326326 703186
rect 326378 703134 326390 703186
rect 326442 703134 326454 703186
rect 326506 703134 326518 703186
rect 326570 703134 326582 703186
rect 326634 703134 326646 703186
rect 326698 703134 326710 703186
rect 326762 703134 326774 703186
rect 326826 703160 326854 703186
rect 326826 703134 326870 703160
rect 324796 703122 326870 703134
rect 254826 703094 254870 703120
rect 252794 703082 254870 703094
rect 252794 703030 254262 703082
rect 254314 703030 254326 703082
rect 254378 703030 254390 703082
rect 254442 703030 254454 703082
rect 254506 703030 254518 703082
rect 254570 703030 254582 703082
rect 254634 703030 254646 703082
rect 254698 703030 254710 703082
rect 254762 703030 254774 703082
rect 254826 703030 254870 703082
rect 324796 703070 326262 703122
rect 326314 703070 326326 703122
rect 326378 703070 326390 703122
rect 326442 703070 326454 703122
rect 326506 703070 326518 703122
rect 326570 703070 326582 703122
rect 326634 703070 326646 703122
rect 326698 703070 326710 703122
rect 326762 703070 326774 703122
rect 326826 703070 326870 703122
rect 324796 703064 326870 703070
rect 252794 703024 254870 703030
rect 362234 702909 362854 702915
rect 362234 702857 362262 702909
rect 362314 702857 362326 702909
rect 362378 702857 362390 702909
rect 362442 702857 362454 702909
rect 362506 702857 362518 702909
rect 362570 702857 362582 702909
rect 362634 702857 362646 702909
rect 362698 702857 362710 702909
rect 362762 702857 362774 702909
rect 362826 702857 362854 702909
rect 362234 702845 362854 702857
rect 362234 702793 362262 702845
rect 362314 702793 362326 702845
rect 362378 702793 362390 702845
rect 362442 702793 362454 702845
rect 362506 702793 362518 702845
rect 362570 702793 362582 702845
rect 362634 702793 362646 702845
rect 362698 702793 362710 702845
rect 362762 702793 362774 702845
rect 362826 702793 362854 702845
rect 362234 702781 362854 702793
rect 362234 702729 362262 702781
rect 362314 702729 362326 702781
rect 362378 702729 362390 702781
rect 362442 702729 362454 702781
rect 362506 702729 362518 702781
rect 362570 702729 362582 702781
rect 362634 702729 362646 702781
rect 362698 702729 362710 702781
rect 362762 702729 362774 702781
rect 362826 702729 362854 702781
rect 362234 702717 362854 702729
rect 252727 702611 252733 702663
rect 252785 702611 252791 702663
rect 324726 702651 324732 702703
rect 324784 702651 324790 702703
rect 362234 702691 362262 702717
rect 360828 702665 362262 702691
rect 362314 702665 362326 702717
rect 362378 702665 362390 702717
rect 362442 702665 362454 702717
rect 362506 702665 362518 702717
rect 362570 702665 362582 702717
rect 362634 702665 362646 702717
rect 362698 702665 362710 702717
rect 362762 702665 362774 702717
rect 362826 702691 362854 702717
rect 434234 702772 434854 702778
rect 434234 702720 434262 702772
rect 434314 702720 434326 702772
rect 434378 702720 434390 702772
rect 434442 702720 434454 702772
rect 434506 702720 434518 702772
rect 434570 702720 434582 702772
rect 434634 702720 434646 702772
rect 434698 702720 434710 702772
rect 434762 702720 434774 702772
rect 434826 702720 434854 702772
rect 434234 702708 434854 702720
rect 362826 702665 362870 702691
rect 360828 702653 362870 702665
rect 324799 702610 325663 702616
rect 252797 702570 253663 702576
rect 252479 702518 252563 702552
rect 252797 702518 253022 702570
rect 253074 702518 253086 702570
rect 253138 702518 253150 702570
rect 253202 702518 253214 702570
rect 253266 702518 253278 702570
rect 253330 702518 253342 702570
rect 253394 702518 253406 702570
rect 253458 702518 253470 702570
rect 253522 702518 253534 702570
rect 253586 702518 253663 702570
rect 324481 702558 324565 702592
rect 324799 702558 325022 702610
rect 325074 702558 325086 702610
rect 325138 702558 325150 702610
rect 325202 702558 325214 702610
rect 325266 702558 325278 702610
rect 325330 702558 325342 702610
rect 325394 702558 325406 702610
rect 325458 702558 325470 702610
rect 325522 702558 325534 702610
rect 325586 702558 325663 702610
rect 360828 702601 362262 702653
rect 362314 702601 362326 702653
rect 362378 702601 362390 702653
rect 362442 702601 362454 702653
rect 362506 702601 362518 702653
rect 362570 702601 362582 702653
rect 362634 702601 362646 702653
rect 362698 702601 362710 702653
rect 362762 702601 362774 702653
rect 362826 702601 362870 702653
rect 360828 702595 362870 702601
rect 434234 702656 434262 702708
rect 434314 702656 434326 702708
rect 434378 702656 434390 702708
rect 434442 702656 434454 702708
rect 434506 702656 434518 702708
rect 434570 702656 434582 702708
rect 434634 702656 434646 702708
rect 434698 702656 434710 702708
rect 434762 702656 434774 702708
rect 434826 702656 434854 702708
rect 434234 702644 434854 702656
rect 324799 702546 325663 702558
rect 434234 702592 434262 702644
rect 434314 702592 434326 702644
rect 434378 702592 434390 702644
rect 434442 702592 434454 702644
rect 434506 702592 434518 702644
rect 434570 702592 434582 702644
rect 434634 702592 434646 702644
rect 434698 702592 434710 702644
rect 434762 702592 434774 702644
rect 434826 702592 434854 702644
rect 434234 702580 434854 702592
rect 434234 702554 434262 702580
rect 324799 702520 325022 702546
rect 252797 702506 253663 702518
rect 252797 702480 253022 702506
rect 252994 702454 253022 702480
rect 253074 702454 253086 702506
rect 253138 702454 253150 702506
rect 253202 702454 253214 702506
rect 253266 702454 253278 702506
rect 253330 702454 253342 702506
rect 253394 702454 253406 702506
rect 253458 702454 253470 702506
rect 253522 702454 253534 702506
rect 253586 702480 253663 702506
rect 324994 702494 325022 702520
rect 325074 702494 325086 702546
rect 325138 702494 325150 702546
rect 325202 702494 325214 702546
rect 325266 702494 325278 702546
rect 325330 702494 325342 702546
rect 325394 702494 325406 702546
rect 325458 702494 325470 702546
rect 325522 702494 325534 702546
rect 325586 702520 325663 702546
rect 432788 702528 434262 702554
rect 434314 702528 434326 702580
rect 434378 702528 434390 702580
rect 434442 702528 434454 702580
rect 434506 702528 434518 702580
rect 434570 702528 434582 702580
rect 434634 702528 434646 702580
rect 434698 702528 434710 702580
rect 434762 702528 434774 702580
rect 434826 702554 434854 702580
rect 434826 702528 434870 702554
rect 325586 702494 325614 702520
rect 324994 702482 325614 702494
rect 253586 702454 253614 702480
rect 252994 702442 253614 702454
rect 252994 702390 253022 702442
rect 253074 702390 253086 702442
rect 253138 702390 253150 702442
rect 253202 702390 253214 702442
rect 253266 702390 253278 702442
rect 253330 702390 253342 702442
rect 253394 702390 253406 702442
rect 253458 702390 253470 702442
rect 253522 702390 253534 702442
rect 253586 702390 253614 702442
rect 252994 702378 253614 702390
rect 252994 702326 253022 702378
rect 253074 702326 253086 702378
rect 253138 702326 253150 702378
rect 253202 702326 253214 702378
rect 253266 702326 253278 702378
rect 253330 702326 253342 702378
rect 253394 702326 253406 702378
rect 253458 702326 253470 702378
rect 253522 702326 253534 702378
rect 253586 702326 253614 702378
rect 252994 702314 253614 702326
rect 252994 702262 253022 702314
rect 253074 702262 253086 702314
rect 253138 702262 253150 702314
rect 253202 702262 253214 702314
rect 253266 702262 253278 702314
rect 253330 702262 253342 702314
rect 253394 702262 253406 702314
rect 253458 702262 253470 702314
rect 253522 702262 253534 702314
rect 253586 702262 253614 702314
rect 324994 702430 325022 702482
rect 325074 702430 325086 702482
rect 325138 702430 325150 702482
rect 325202 702430 325214 702482
rect 325266 702430 325278 702482
rect 325330 702430 325342 702482
rect 325394 702430 325406 702482
rect 325458 702430 325470 702482
rect 325522 702430 325534 702482
rect 325586 702430 325614 702482
rect 432788 702516 434870 702528
rect 432788 702464 434262 702516
rect 434314 702464 434326 702516
rect 434378 702464 434390 702516
rect 434442 702464 434454 702516
rect 434506 702464 434518 702516
rect 434570 702464 434582 702516
rect 434634 702464 434646 702516
rect 434698 702464 434710 702516
rect 434762 702464 434774 702516
rect 434826 702464 434870 702516
rect 432788 702458 434870 702464
rect 506234 702526 506854 702532
rect 506234 702474 506262 702526
rect 506314 702474 506326 702526
rect 506378 702474 506390 702526
rect 506442 702474 506454 702526
rect 506506 702474 506518 702526
rect 506570 702474 506582 702526
rect 506634 702474 506646 702526
rect 506698 702474 506710 702526
rect 506762 702474 506774 702526
rect 506826 702474 506854 702526
rect 506234 702462 506854 702474
rect 324994 702418 325614 702430
rect 324994 702366 325022 702418
rect 325074 702366 325086 702418
rect 325138 702366 325150 702418
rect 325202 702366 325214 702418
rect 325266 702366 325278 702418
rect 325330 702366 325342 702418
rect 325394 702366 325406 702418
rect 325458 702366 325470 702418
rect 325522 702366 325534 702418
rect 325586 702366 325614 702418
rect 324994 702354 325614 702366
rect 324994 702302 325022 702354
rect 325074 702302 325086 702354
rect 325138 702302 325150 702354
rect 325202 702302 325214 702354
rect 325266 702302 325278 702354
rect 325330 702302 325342 702354
rect 325394 702302 325406 702354
rect 325458 702302 325470 702354
rect 325522 702302 325534 702354
rect 325586 702302 325614 702354
rect 506234 702410 506262 702462
rect 506314 702410 506326 702462
rect 506378 702410 506390 702462
rect 506442 702410 506454 702462
rect 506506 702410 506518 702462
rect 506570 702410 506582 702462
rect 506634 702410 506646 702462
rect 506698 702410 506710 702462
rect 506762 702410 506774 702462
rect 506826 702410 506854 702462
rect 506234 702398 506854 702410
rect 506234 702346 506262 702398
rect 506314 702346 506326 702398
rect 506378 702346 506390 702398
rect 506442 702346 506454 702398
rect 506506 702346 506518 702398
rect 506570 702346 506582 702398
rect 506634 702346 506646 702398
rect 506698 702346 506710 702398
rect 506762 702346 506774 702398
rect 506826 702346 506854 702398
rect 506234 702334 506854 702346
rect 506234 702308 506262 702334
rect 324994 702296 325614 702302
rect 252994 702256 253614 702262
rect 504783 702282 506262 702308
rect 506314 702282 506326 702334
rect 506378 702282 506390 702334
rect 506442 702282 506454 702334
rect 506506 702282 506518 702334
rect 506570 702282 506582 702334
rect 506634 702282 506646 702334
rect 506698 702282 506710 702334
rect 506762 702282 506774 702334
rect 506826 702308 506854 702334
rect 506826 702282 506870 702308
rect 504783 702270 506870 702282
rect 360753 702182 360759 702234
rect 360811 702182 360817 702234
rect 504783 702218 506262 702270
rect 506314 702218 506326 702270
rect 506378 702218 506390 702270
rect 506442 702218 506454 702270
rect 506506 702218 506518 702270
rect 506570 702218 506582 702270
rect 506634 702218 506646 702270
rect 506698 702218 506710 702270
rect 506762 702218 506774 702270
rect 506826 702218 506870 702270
rect 504783 702212 506870 702218
rect 360831 702141 361663 702147
rect 360513 702089 360597 702123
rect 360831 702089 361022 702141
rect 361074 702089 361086 702141
rect 361138 702089 361150 702141
rect 361202 702089 361214 702141
rect 361266 702089 361278 702141
rect 361330 702089 361342 702141
rect 361394 702089 361406 702141
rect 361458 702089 361470 702141
rect 361522 702089 361534 702141
rect 361586 702089 361663 702141
rect 360831 702077 361663 702089
rect 360831 702051 361022 702077
rect 360994 702025 361022 702051
rect 361074 702025 361086 702077
rect 361138 702025 361150 702077
rect 361202 702025 361214 702077
rect 361266 702025 361278 702077
rect 361330 702025 361342 702077
rect 361394 702025 361406 702077
rect 361458 702025 361470 702077
rect 361522 702025 361534 702077
rect 361586 702051 361663 702077
rect 361586 702025 361614 702051
rect 432723 702045 432729 702097
rect 432781 702045 432787 702097
rect 360994 702013 361614 702025
rect 360994 701961 361022 702013
rect 361074 701961 361086 702013
rect 361138 701961 361150 702013
rect 361202 701961 361214 702013
rect 361266 701961 361278 702013
rect 361330 701961 361342 702013
rect 361394 701961 361406 702013
rect 361458 701961 361470 702013
rect 361522 701961 361534 702013
rect 361586 701961 361614 702013
rect 432791 702004 433663 702010
rect 360994 701949 361614 701961
rect 432473 701952 432557 701986
rect 432791 701952 433022 702004
rect 433074 701952 433086 702004
rect 433138 701952 433150 702004
rect 433202 701952 433214 702004
rect 433266 701952 433278 702004
rect 433330 701952 433342 702004
rect 433394 701952 433406 702004
rect 433458 701952 433470 702004
rect 433522 701952 433534 702004
rect 433586 701952 433663 702004
rect 360994 701897 361022 701949
rect 361074 701897 361086 701949
rect 361138 701897 361150 701949
rect 361202 701897 361214 701949
rect 361266 701897 361278 701949
rect 361330 701897 361342 701949
rect 361394 701897 361406 701949
rect 361458 701897 361470 701949
rect 361522 701897 361534 701949
rect 361586 701897 361614 701949
rect 432791 701940 433663 701952
rect 432791 701914 433022 701940
rect 360994 701885 361614 701897
rect 360994 701833 361022 701885
rect 361074 701833 361086 701885
rect 361138 701833 361150 701885
rect 361202 701833 361214 701885
rect 361266 701833 361278 701885
rect 361330 701833 361342 701885
rect 361394 701833 361406 701885
rect 361458 701833 361470 701885
rect 361522 701833 361534 701885
rect 361586 701833 361614 701885
rect 360994 701827 361614 701833
rect 432994 701888 433022 701914
rect 433074 701888 433086 701940
rect 433138 701888 433150 701940
rect 433202 701888 433214 701940
rect 433266 701888 433278 701940
rect 433330 701888 433342 701940
rect 433394 701888 433406 701940
rect 433458 701888 433470 701940
rect 433522 701888 433534 701940
rect 433586 701914 433663 701940
rect 433586 701888 433614 701914
rect 432994 701876 433614 701888
rect 432994 701824 433022 701876
rect 433074 701824 433086 701876
rect 433138 701824 433150 701876
rect 433202 701824 433214 701876
rect 433266 701824 433278 701876
rect 433330 701824 433342 701876
rect 433394 701824 433406 701876
rect 433458 701824 433470 701876
rect 433522 701824 433534 701876
rect 433586 701824 433614 701876
rect 432994 701812 433614 701824
rect 432994 701760 433022 701812
rect 433074 701760 433086 701812
rect 433138 701760 433150 701812
rect 433202 701760 433214 701812
rect 433266 701760 433278 701812
rect 433330 701760 433342 701812
rect 433394 701760 433406 701812
rect 433458 701760 433470 701812
rect 433522 701760 433534 701812
rect 433586 701760 433614 701812
rect 504719 701799 504725 701851
rect 504777 701799 504783 701851
rect 432994 701748 433614 701760
rect 432994 701696 433022 701748
rect 433074 701696 433086 701748
rect 433138 701696 433150 701748
rect 433202 701696 433214 701748
rect 433266 701696 433278 701748
rect 433330 701696 433342 701748
rect 433394 701696 433406 701748
rect 433458 701696 433470 701748
rect 433522 701696 433534 701748
rect 433586 701696 433614 701748
rect 504786 701758 505663 701764
rect 504468 701706 504552 701740
rect 504786 701706 505022 701758
rect 505074 701706 505086 701758
rect 505138 701706 505150 701758
rect 505202 701706 505214 701758
rect 505266 701706 505278 701758
rect 505330 701706 505342 701758
rect 505394 701706 505406 701758
rect 505458 701706 505470 701758
rect 505522 701706 505534 701758
rect 505586 701706 505663 701758
rect 432994 701690 433614 701696
rect 504786 701694 505663 701706
rect 504786 701668 505022 701694
rect 504994 701642 505022 701668
rect 505074 701642 505086 701694
rect 505138 701642 505150 701694
rect 505202 701642 505214 701694
rect 505266 701642 505278 701694
rect 505330 701642 505342 701694
rect 505394 701642 505406 701694
rect 505458 701642 505470 701694
rect 505522 701642 505534 701694
rect 505586 701668 505663 701694
rect 505586 701642 505614 701668
rect 504994 701630 505614 701642
rect 504994 701578 505022 701630
rect 505074 701578 505086 701630
rect 505138 701578 505150 701630
rect 505202 701578 505214 701630
rect 505266 701578 505278 701630
rect 505330 701578 505342 701630
rect 505394 701578 505406 701630
rect 505458 701578 505470 701630
rect 505522 701578 505534 701630
rect 505586 701578 505614 701630
rect 504994 701566 505614 701578
rect 504994 701514 505022 701566
rect 505074 701514 505086 701566
rect 505138 701514 505150 701566
rect 505202 701514 505214 701566
rect 505266 701514 505278 701566
rect 505330 701514 505342 701566
rect 505394 701514 505406 701566
rect 505458 701514 505470 701566
rect 505522 701514 505534 701566
rect 505586 701514 505614 701566
rect 504994 701502 505614 701514
rect 504994 701450 505022 701502
rect 505074 701450 505086 701502
rect 505138 701450 505150 701502
rect 505202 701450 505214 701502
rect 505266 701450 505278 701502
rect 505330 701450 505342 701502
rect 505394 701450 505406 701502
rect 505458 701450 505470 701502
rect 505522 701450 505534 701502
rect 505586 701450 505614 701502
rect 504994 701444 505614 701450
rect 267642 700954 267648 701006
rect 267700 700954 267706 701006
rect 332502 700954 332508 701006
rect 332560 700954 332566 701006
rect 397454 700954 397460 701006
rect 397512 700954 397518 701006
rect 462314 700954 462320 701006
rect 462372 700954 462378 701006
rect 527174 700954 527180 701006
rect 527232 700954 527238 701006
rect 576994 697912 577614 697934
rect 576994 697860 577022 697912
rect 577074 697860 577086 697912
rect 577138 697860 577150 697912
rect 577202 697860 577214 697912
rect 577266 697860 577278 697912
rect 577330 697860 577342 697912
rect 577394 697860 577406 697912
rect 577458 697860 577470 697912
rect 577522 697860 577534 697912
rect 577586 697860 577614 697912
rect 576994 697848 577614 697860
rect 576994 697796 577022 697848
rect 577074 697796 577086 697848
rect 577138 697796 577150 697848
rect 577202 697796 577214 697848
rect 577266 697796 577278 697848
rect 577330 697796 577342 697848
rect 577394 697796 577406 697848
rect 577458 697796 577470 697848
rect 577522 697796 577534 697848
rect 577586 697796 577614 697848
rect 576994 697784 577614 697796
rect 576994 697732 577022 697784
rect 577074 697732 577086 697784
rect 577138 697732 577150 697784
rect 577202 697732 577214 697784
rect 577266 697732 577278 697784
rect 577330 697732 577342 697784
rect 577394 697732 577406 697784
rect 577458 697732 577470 697784
rect 577522 697732 577534 697784
rect 577586 697732 577614 697784
rect 576994 697720 577614 697732
rect 576994 697694 577022 697720
rect 576400 697668 577022 697694
rect 577074 697668 577086 697720
rect 577138 697668 577150 697720
rect 577202 697668 577214 697720
rect 577266 697668 577278 697720
rect 577330 697668 577342 697720
rect 577394 697668 577406 697720
rect 577458 697668 577470 697720
rect 577522 697668 577534 697720
rect 577586 697694 577614 697720
rect 577586 697668 577647 697694
rect 576400 697663 577647 697668
rect 576316 697656 577647 697663
rect 576316 697629 577022 697656
rect 576400 697604 577022 697629
rect 577074 697604 577086 697656
rect 577138 697604 577150 697656
rect 577202 697604 577214 697656
rect 577266 697604 577278 697656
rect 577330 697604 577342 697656
rect 577394 697604 577406 697656
rect 577458 697604 577470 697656
rect 577522 697604 577534 697656
rect 577586 697604 577647 697656
rect 576400 697598 577647 697604
rect 576597 697178 576603 697230
rect 576655 697178 576661 697230
rect 576400 697117 578876 697150
rect 576400 697065 578262 697117
rect 578314 697065 578326 697117
rect 578378 697065 578390 697117
rect 578442 697065 578454 697117
rect 578506 697065 578518 697117
rect 578570 697065 578582 697117
rect 578634 697065 578646 697117
rect 578698 697065 578710 697117
rect 578762 697065 578774 697117
rect 578826 697065 578876 697117
rect 576400 697054 578876 697065
rect 578234 697053 578854 697054
rect 578234 697001 578262 697053
rect 578314 697001 578326 697053
rect 578378 697001 578390 697053
rect 578442 697001 578454 697053
rect 578506 697001 578518 697053
rect 578570 697001 578582 697053
rect 578634 697001 578646 697053
rect 578698 697001 578710 697053
rect 578762 697001 578774 697053
rect 578826 697001 578854 697053
rect 578234 696989 578854 697001
rect 578234 696937 578262 696989
rect 578314 696937 578326 696989
rect 578378 696937 578390 696989
rect 578442 696937 578454 696989
rect 578506 696937 578518 696989
rect 578570 696937 578582 696989
rect 578634 696937 578646 696989
rect 578698 696937 578710 696989
rect 578762 696937 578774 696989
rect 578826 696937 578854 696989
rect 578234 696925 578854 696937
rect 578234 696873 578262 696925
rect 578314 696873 578326 696925
rect 578378 696873 578390 696925
rect 578442 696873 578454 696925
rect 578506 696873 578518 696925
rect 578570 696873 578582 696925
rect 578634 696873 578646 696925
rect 578698 696873 578710 696925
rect 578762 696873 578774 696925
rect 578826 696873 578854 696925
rect 578234 696861 578854 696873
rect 578234 696809 578262 696861
rect 578314 696809 578326 696861
rect 578378 696809 578390 696861
rect 578442 696809 578454 696861
rect 578506 696809 578518 696861
rect 578570 696809 578582 696861
rect 578634 696809 578646 696861
rect 578698 696809 578710 696861
rect 578762 696809 578774 696861
rect 578826 696809 578854 696861
rect 578234 696803 578854 696809
rect 576994 644736 577614 644758
rect 576994 644684 577022 644736
rect 577074 644684 577086 644736
rect 577138 644684 577150 644736
rect 577202 644684 577214 644736
rect 577266 644684 577278 644736
rect 577330 644684 577342 644736
rect 577394 644684 577406 644736
rect 577458 644684 577470 644736
rect 577522 644684 577534 644736
rect 577586 644684 577614 644736
rect 576994 644672 577614 644684
rect 576994 644620 577022 644672
rect 577074 644620 577086 644672
rect 577138 644620 577150 644672
rect 577202 644620 577214 644672
rect 577266 644620 577278 644672
rect 577330 644620 577342 644672
rect 577394 644620 577406 644672
rect 577458 644620 577470 644672
rect 577522 644620 577534 644672
rect 577586 644620 577614 644672
rect 576994 644608 577614 644620
rect 576994 644556 577022 644608
rect 577074 644556 577086 644608
rect 577138 644556 577150 644608
rect 577202 644556 577214 644608
rect 577266 644556 577278 644608
rect 577330 644556 577342 644608
rect 577394 644556 577406 644608
rect 577458 644556 577470 644608
rect 577522 644556 577534 644608
rect 577586 644556 577614 644608
rect 576994 644544 577614 644556
rect 576994 644518 577022 644544
rect 576400 644492 577022 644518
rect 577074 644492 577086 644544
rect 577138 644492 577150 644544
rect 577202 644492 577214 644544
rect 577266 644492 577278 644544
rect 577330 644492 577342 644544
rect 577394 644492 577406 644544
rect 577458 644492 577470 644544
rect 577522 644492 577534 644544
rect 577586 644518 577614 644544
rect 577586 644492 577647 644518
rect 576400 644487 577647 644492
rect 576316 644480 577647 644487
rect 576316 644453 577022 644480
rect 576400 644428 577022 644453
rect 577074 644428 577086 644480
rect 577138 644428 577150 644480
rect 577202 644428 577214 644480
rect 577266 644428 577278 644480
rect 577330 644428 577342 644480
rect 577394 644428 577406 644480
rect 577458 644428 577470 644480
rect 577522 644428 577534 644480
rect 577586 644428 577647 644480
rect 576400 644422 577647 644428
rect 576597 644002 576603 644054
rect 576655 644002 576661 644054
rect 576400 643941 578876 643974
rect 576400 643889 578262 643941
rect 578314 643889 578326 643941
rect 578378 643889 578390 643941
rect 578442 643889 578454 643941
rect 578506 643889 578518 643941
rect 578570 643889 578582 643941
rect 578634 643889 578646 643941
rect 578698 643889 578710 643941
rect 578762 643889 578774 643941
rect 578826 643889 578876 643941
rect 576400 643878 578876 643889
rect 578234 643877 578854 643878
rect 578234 643825 578262 643877
rect 578314 643825 578326 643877
rect 578378 643825 578390 643877
rect 578442 643825 578454 643877
rect 578506 643825 578518 643877
rect 578570 643825 578582 643877
rect 578634 643825 578646 643877
rect 578698 643825 578710 643877
rect 578762 643825 578774 643877
rect 578826 643825 578854 643877
rect 578234 643813 578854 643825
rect 578234 643761 578262 643813
rect 578314 643761 578326 643813
rect 578378 643761 578390 643813
rect 578442 643761 578454 643813
rect 578506 643761 578518 643813
rect 578570 643761 578582 643813
rect 578634 643761 578646 643813
rect 578698 643761 578710 643813
rect 578762 643761 578774 643813
rect 578826 643761 578854 643813
rect 578234 643749 578854 643761
rect 578234 643697 578262 643749
rect 578314 643697 578326 643749
rect 578378 643697 578390 643749
rect 578442 643697 578454 643749
rect 578506 643697 578518 643749
rect 578570 643697 578582 643749
rect 578634 643697 578646 643749
rect 578698 643697 578710 643749
rect 578762 643697 578774 643749
rect 578826 643697 578854 643749
rect 578234 643685 578854 643697
rect 578234 643633 578262 643685
rect 578314 643633 578326 643685
rect 578378 643633 578390 643685
rect 578442 643633 578454 643685
rect 578506 643633 578518 643685
rect 578570 643633 578582 643685
rect 578634 643633 578646 643685
rect 578698 643633 578710 643685
rect 578762 643633 578774 643685
rect 578826 643633 578854 643685
rect 578234 643627 578854 643633
rect 576994 591696 577614 591718
rect 576994 591644 577022 591696
rect 577074 591644 577086 591696
rect 577138 591644 577150 591696
rect 577202 591644 577214 591696
rect 577266 591644 577278 591696
rect 577330 591644 577342 591696
rect 577394 591644 577406 591696
rect 577458 591644 577470 591696
rect 577522 591644 577534 591696
rect 577586 591644 577614 591696
rect 576994 591632 577614 591644
rect 576994 591580 577022 591632
rect 577074 591580 577086 591632
rect 577138 591580 577150 591632
rect 577202 591580 577214 591632
rect 577266 591580 577278 591632
rect 577330 591580 577342 591632
rect 577394 591580 577406 591632
rect 577458 591580 577470 591632
rect 577522 591580 577534 591632
rect 577586 591580 577614 591632
rect 576994 591568 577614 591580
rect 576994 591516 577022 591568
rect 577074 591516 577086 591568
rect 577138 591516 577150 591568
rect 577202 591516 577214 591568
rect 577266 591516 577278 591568
rect 577330 591516 577342 591568
rect 577394 591516 577406 591568
rect 577458 591516 577470 591568
rect 577522 591516 577534 591568
rect 577586 591516 577614 591568
rect 576994 591504 577614 591516
rect 576994 591478 577022 591504
rect 576400 591452 577022 591478
rect 577074 591452 577086 591504
rect 577138 591452 577150 591504
rect 577202 591452 577214 591504
rect 577266 591452 577278 591504
rect 577330 591452 577342 591504
rect 577394 591452 577406 591504
rect 577458 591452 577470 591504
rect 577522 591452 577534 591504
rect 577586 591478 577614 591504
rect 577586 591452 577647 591478
rect 576400 591447 577647 591452
rect 576316 591440 577647 591447
rect 576316 591413 577022 591440
rect 576400 591388 577022 591413
rect 577074 591388 577086 591440
rect 577138 591388 577150 591440
rect 577202 591388 577214 591440
rect 577266 591388 577278 591440
rect 577330 591388 577342 591440
rect 577394 591388 577406 591440
rect 577458 591388 577470 591440
rect 577522 591388 577534 591440
rect 577586 591388 577647 591440
rect 576400 591382 577647 591388
rect 576597 590962 576603 591014
rect 576655 590962 576661 591014
rect 576400 590901 578876 590934
rect 576400 590849 578262 590901
rect 578314 590849 578326 590901
rect 578378 590849 578390 590901
rect 578442 590849 578454 590901
rect 578506 590849 578518 590901
rect 578570 590849 578582 590901
rect 578634 590849 578646 590901
rect 578698 590849 578710 590901
rect 578762 590849 578774 590901
rect 578826 590849 578876 590901
rect 576400 590838 578876 590849
rect 578234 590837 578854 590838
rect 578234 590785 578262 590837
rect 578314 590785 578326 590837
rect 578378 590785 578390 590837
rect 578442 590785 578454 590837
rect 578506 590785 578518 590837
rect 578570 590785 578582 590837
rect 578634 590785 578646 590837
rect 578698 590785 578710 590837
rect 578762 590785 578774 590837
rect 578826 590785 578854 590837
rect 578234 590773 578854 590785
rect 578234 590721 578262 590773
rect 578314 590721 578326 590773
rect 578378 590721 578390 590773
rect 578442 590721 578454 590773
rect 578506 590721 578518 590773
rect 578570 590721 578582 590773
rect 578634 590721 578646 590773
rect 578698 590721 578710 590773
rect 578762 590721 578774 590773
rect 578826 590721 578854 590773
rect 578234 590709 578854 590721
rect 578234 590657 578262 590709
rect 578314 590657 578326 590709
rect 578378 590657 578390 590709
rect 578442 590657 578454 590709
rect 578506 590657 578518 590709
rect 578570 590657 578582 590709
rect 578634 590657 578646 590709
rect 578698 590657 578710 590709
rect 578762 590657 578774 590709
rect 578826 590657 578854 590709
rect 578234 590645 578854 590657
rect 578234 590593 578262 590645
rect 578314 590593 578326 590645
rect 578378 590593 578390 590645
rect 578442 590593 578454 590645
rect 578506 590593 578518 590645
rect 578570 590593 578582 590645
rect 578634 590593 578646 590645
rect 578698 590593 578710 590645
rect 578762 590593 578774 590645
rect 578826 590593 578854 590645
rect 578234 590587 578854 590593
rect 504994 554604 505614 554626
rect 504994 554552 505022 554604
rect 505074 554552 505086 554604
rect 505138 554552 505150 554604
rect 505202 554552 505214 554604
rect 505266 554552 505278 554604
rect 505330 554552 505342 554604
rect 505394 554552 505406 554604
rect 505458 554552 505470 554604
rect 505522 554552 505534 554604
rect 505586 554552 505614 554604
rect 504994 554540 505614 554552
rect 504994 554488 505022 554540
rect 505074 554488 505086 554540
rect 505138 554488 505150 554540
rect 505202 554488 505214 554540
rect 505266 554488 505278 554540
rect 505330 554488 505342 554540
rect 505394 554488 505406 554540
rect 505458 554488 505470 554540
rect 505522 554488 505534 554540
rect 505586 554488 505614 554540
rect 504994 554476 505614 554488
rect 504994 554424 505022 554476
rect 505074 554424 505086 554476
rect 505138 554424 505150 554476
rect 505202 554424 505214 554476
rect 505266 554424 505278 554476
rect 505330 554424 505342 554476
rect 505394 554424 505406 554476
rect 505458 554424 505470 554476
rect 505522 554424 505534 554476
rect 505586 554424 505614 554476
rect 504994 554412 505614 554424
rect 504994 554386 505022 554412
rect 504306 554360 505022 554386
rect 505074 554360 505086 554412
rect 505138 554360 505150 554412
rect 505202 554360 505214 554412
rect 505266 554360 505278 554412
rect 505330 554360 505342 554412
rect 505394 554360 505406 554412
rect 505458 554360 505470 554412
rect 505522 554360 505534 554412
rect 505586 554386 505614 554412
rect 505586 554360 505647 554386
rect 504306 554355 505647 554360
rect 504222 554348 505647 554355
rect 504222 554321 505022 554348
rect 504306 554296 505022 554321
rect 505074 554296 505086 554348
rect 505138 554296 505150 554348
rect 505202 554296 505214 554348
rect 505266 554296 505278 554348
rect 505330 554296 505342 554348
rect 505394 554296 505406 554348
rect 505458 554296 505470 554348
rect 505522 554296 505534 554348
rect 505586 554296 505647 554348
rect 504306 554290 505647 554296
rect 504507 554049 504565 554055
rect 504507 554015 504519 554049
rect 504553 554046 504565 554049
rect 536098 554046 536104 554058
rect 504553 554018 536104 554046
rect 504553 554015 504565 554018
rect 504507 554009 504565 554015
rect 536098 554006 536104 554018
rect 536156 554006 536162 554058
rect 504306 553809 506876 553842
rect 504306 553757 506262 553809
rect 506314 553757 506326 553809
rect 506378 553757 506390 553809
rect 506442 553757 506454 553809
rect 506506 553757 506518 553809
rect 506570 553757 506582 553809
rect 506634 553757 506646 553809
rect 506698 553757 506710 553809
rect 506762 553757 506774 553809
rect 506826 553757 506876 553809
rect 504306 553746 506876 553757
rect 506234 553745 506854 553746
rect 506234 553693 506262 553745
rect 506314 553693 506326 553745
rect 506378 553693 506390 553745
rect 506442 553693 506454 553745
rect 506506 553693 506518 553745
rect 506570 553693 506582 553745
rect 506634 553693 506646 553745
rect 506698 553693 506710 553745
rect 506762 553693 506774 553745
rect 506826 553693 506854 553745
rect 506234 553681 506854 553693
rect 506234 553629 506262 553681
rect 506314 553629 506326 553681
rect 506378 553629 506390 553681
rect 506442 553629 506454 553681
rect 506506 553629 506518 553681
rect 506570 553629 506582 553681
rect 506634 553629 506646 553681
rect 506698 553629 506710 553681
rect 506762 553629 506774 553681
rect 506826 553629 506854 553681
rect 506234 553617 506854 553629
rect 506234 553565 506262 553617
rect 506314 553565 506326 553617
rect 506378 553565 506390 553617
rect 506442 553565 506454 553617
rect 506506 553565 506518 553617
rect 506570 553565 506582 553617
rect 506634 553565 506646 553617
rect 506698 553565 506710 553617
rect 506762 553565 506774 553617
rect 506826 553565 506854 553617
rect 506234 553553 506854 553565
rect 506234 553501 506262 553553
rect 506314 553501 506326 553553
rect 506378 553501 506390 553553
rect 506442 553501 506454 553553
rect 506506 553501 506518 553553
rect 506570 553501 506582 553553
rect 506634 553501 506646 553553
rect 506698 553501 506710 553553
rect 506762 553501 506774 553553
rect 506826 553501 506854 553553
rect 506234 553495 506854 553501
rect 576994 538520 577614 538542
rect 576994 538468 577022 538520
rect 577074 538468 577086 538520
rect 577138 538468 577150 538520
rect 577202 538468 577214 538520
rect 577266 538468 577278 538520
rect 577330 538468 577342 538520
rect 577394 538468 577406 538520
rect 577458 538468 577470 538520
rect 577522 538468 577534 538520
rect 577586 538468 577614 538520
rect 576994 538456 577614 538468
rect 576994 538404 577022 538456
rect 577074 538404 577086 538456
rect 577138 538404 577150 538456
rect 577202 538404 577214 538456
rect 577266 538404 577278 538456
rect 577330 538404 577342 538456
rect 577394 538404 577406 538456
rect 577458 538404 577470 538456
rect 577522 538404 577534 538456
rect 577586 538404 577614 538456
rect 576994 538392 577614 538404
rect 576994 538340 577022 538392
rect 577074 538340 577086 538392
rect 577138 538340 577150 538392
rect 577202 538340 577214 538392
rect 577266 538340 577278 538392
rect 577330 538340 577342 538392
rect 577394 538340 577406 538392
rect 577458 538340 577470 538392
rect 577522 538340 577534 538392
rect 577586 538340 577614 538392
rect 576994 538328 577614 538340
rect 576994 538302 577022 538328
rect 576400 538276 577022 538302
rect 577074 538276 577086 538328
rect 577138 538276 577150 538328
rect 577202 538276 577214 538328
rect 577266 538276 577278 538328
rect 577330 538276 577342 538328
rect 577394 538276 577406 538328
rect 577458 538276 577470 538328
rect 577522 538276 577534 538328
rect 577586 538302 577614 538328
rect 577586 538276 577647 538302
rect 576400 538271 577647 538276
rect 576316 538264 577647 538271
rect 576316 538237 577022 538264
rect 576400 538212 577022 538237
rect 577074 538212 577086 538264
rect 577138 538212 577150 538264
rect 577202 538212 577214 538264
rect 577266 538212 577278 538264
rect 577330 538212 577342 538264
rect 577394 538212 577406 538264
rect 577458 538212 577470 538264
rect 577522 538212 577534 538264
rect 577586 538212 577647 538264
rect 576400 538206 577647 538212
rect 576597 537786 576603 537838
rect 576655 537786 576661 537838
rect 576400 537725 578876 537758
rect 576400 537673 578262 537725
rect 578314 537673 578326 537725
rect 578378 537673 578390 537725
rect 578442 537673 578454 537725
rect 578506 537673 578518 537725
rect 578570 537673 578582 537725
rect 578634 537673 578646 537725
rect 578698 537673 578710 537725
rect 578762 537673 578774 537725
rect 578826 537673 578876 537725
rect 576400 537662 578876 537673
rect 578234 537661 578854 537662
rect 578234 537609 578262 537661
rect 578314 537609 578326 537661
rect 578378 537609 578390 537661
rect 578442 537609 578454 537661
rect 578506 537609 578518 537661
rect 578570 537609 578582 537661
rect 578634 537609 578646 537661
rect 578698 537609 578710 537661
rect 578762 537609 578774 537661
rect 578826 537609 578854 537661
rect 578234 537597 578854 537609
rect 578234 537545 578262 537597
rect 578314 537545 578326 537597
rect 578378 537545 578390 537597
rect 578442 537545 578454 537597
rect 578506 537545 578518 537597
rect 578570 537545 578582 537597
rect 578634 537545 578646 537597
rect 578698 537545 578710 537597
rect 578762 537545 578774 537597
rect 578826 537545 578854 537597
rect 578234 537533 578854 537545
rect 578234 537481 578262 537533
rect 578314 537481 578326 537533
rect 578378 537481 578390 537533
rect 578442 537481 578454 537533
rect 578506 537481 578518 537533
rect 578570 537481 578582 537533
rect 578634 537481 578646 537533
rect 578698 537481 578710 537533
rect 578762 537481 578774 537533
rect 578826 537481 578854 537533
rect 578234 537469 578854 537481
rect 578234 537417 578262 537469
rect 578314 537417 578326 537469
rect 578378 537417 578390 537469
rect 578442 537417 578454 537469
rect 578506 537417 578518 537469
rect 578570 537417 578582 537469
rect 578634 537417 578646 537469
rect 578698 537417 578710 537469
rect 578762 537417 578774 537469
rect 578826 537417 578854 537469
rect 578234 537411 578854 537417
rect 576994 485344 577614 485366
rect 576994 485292 577022 485344
rect 577074 485292 577086 485344
rect 577138 485292 577150 485344
rect 577202 485292 577214 485344
rect 577266 485292 577278 485344
rect 577330 485292 577342 485344
rect 577394 485292 577406 485344
rect 577458 485292 577470 485344
rect 577522 485292 577534 485344
rect 577586 485292 577614 485344
rect 576994 485280 577614 485292
rect 576994 485228 577022 485280
rect 577074 485228 577086 485280
rect 577138 485228 577150 485280
rect 577202 485228 577214 485280
rect 577266 485228 577278 485280
rect 577330 485228 577342 485280
rect 577394 485228 577406 485280
rect 577458 485228 577470 485280
rect 577522 485228 577534 485280
rect 577586 485228 577614 485280
rect 576994 485216 577614 485228
rect 576994 485164 577022 485216
rect 577074 485164 577086 485216
rect 577138 485164 577150 485216
rect 577202 485164 577214 485216
rect 577266 485164 577278 485216
rect 577330 485164 577342 485216
rect 577394 485164 577406 485216
rect 577458 485164 577470 485216
rect 577522 485164 577534 485216
rect 577586 485164 577614 485216
rect 576994 485152 577614 485164
rect 576994 485126 577022 485152
rect 576400 485100 577022 485126
rect 577074 485100 577086 485152
rect 577138 485100 577150 485152
rect 577202 485100 577214 485152
rect 577266 485100 577278 485152
rect 577330 485100 577342 485152
rect 577394 485100 577406 485152
rect 577458 485100 577470 485152
rect 577522 485100 577534 485152
rect 577586 485126 577614 485152
rect 577586 485100 577647 485126
rect 576400 485095 577647 485100
rect 576316 485088 577647 485095
rect 576316 485061 577022 485088
rect 576400 485036 577022 485061
rect 577074 485036 577086 485088
rect 577138 485036 577150 485088
rect 577202 485036 577214 485088
rect 577266 485036 577278 485088
rect 577330 485036 577342 485088
rect 577394 485036 577406 485088
rect 577458 485036 577470 485088
rect 577522 485036 577534 485088
rect 577586 485036 577647 485088
rect 576400 485030 577647 485036
rect 576597 484610 576603 484662
rect 576655 484610 576661 484662
rect 576400 484549 578876 484582
rect 576400 484497 578262 484549
rect 578314 484497 578326 484549
rect 578378 484497 578390 484549
rect 578442 484497 578454 484549
rect 578506 484497 578518 484549
rect 578570 484497 578582 484549
rect 578634 484497 578646 484549
rect 578698 484497 578710 484549
rect 578762 484497 578774 484549
rect 578826 484497 578876 484549
rect 576400 484486 578876 484497
rect 578234 484485 578854 484486
rect 578234 484433 578262 484485
rect 578314 484433 578326 484485
rect 578378 484433 578390 484485
rect 578442 484433 578454 484485
rect 578506 484433 578518 484485
rect 578570 484433 578582 484485
rect 578634 484433 578646 484485
rect 578698 484433 578710 484485
rect 578762 484433 578774 484485
rect 578826 484433 578854 484485
rect 578234 484421 578854 484433
rect 578234 484369 578262 484421
rect 578314 484369 578326 484421
rect 578378 484369 578390 484421
rect 578442 484369 578454 484421
rect 578506 484369 578518 484421
rect 578570 484369 578582 484421
rect 578634 484369 578646 484421
rect 578698 484369 578710 484421
rect 578762 484369 578774 484421
rect 578826 484369 578854 484421
rect 578234 484357 578854 484369
rect 578234 484305 578262 484357
rect 578314 484305 578326 484357
rect 578378 484305 578390 484357
rect 578442 484305 578454 484357
rect 578506 484305 578518 484357
rect 578570 484305 578582 484357
rect 578634 484305 578646 484357
rect 578698 484305 578710 484357
rect 578762 484305 578774 484357
rect 578826 484305 578854 484357
rect 578234 484293 578854 484305
rect 578234 484241 578262 484293
rect 578314 484241 578326 484293
rect 578378 484241 578390 484293
rect 578442 484241 578454 484293
rect 578506 484241 578518 484293
rect 578570 484241 578582 484293
rect 578634 484241 578646 484293
rect 578698 484241 578710 484293
rect 578762 484241 578774 484293
rect 578826 484241 578854 484293
rect 578234 484235 578854 484241
rect 471698 453298 471704 453350
rect 471756 453338 471762 453350
rect 580166 453338 580172 453350
rect 471756 453310 580172 453338
rect 471756 453298 471762 453310
rect 580166 453298 580172 453310
rect 580224 453298 580230 453350
rect 470234 451487 470854 451493
rect 470234 451435 470262 451487
rect 470314 451435 470326 451487
rect 470378 451435 470390 451487
rect 470442 451435 470454 451487
rect 470506 451435 470518 451487
rect 470570 451435 470582 451487
rect 470634 451435 470646 451487
rect 470698 451435 470710 451487
rect 470762 451435 470774 451487
rect 470826 451435 470854 451487
rect 470234 451423 470854 451435
rect 470234 451371 470262 451423
rect 470314 451371 470326 451423
rect 470378 451371 470390 451423
rect 470442 451371 470454 451423
rect 470506 451371 470518 451423
rect 470570 451371 470582 451423
rect 470634 451371 470646 451423
rect 470698 451371 470710 451423
rect 470762 451371 470774 451423
rect 470826 451371 470854 451423
rect 470234 451359 470854 451371
rect 470234 451307 470262 451359
rect 470314 451307 470326 451359
rect 470378 451307 470390 451359
rect 470442 451307 470454 451359
rect 470506 451307 470518 451359
rect 470570 451307 470582 451359
rect 470634 451307 470646 451359
rect 470698 451307 470710 451359
rect 470762 451307 470774 451359
rect 470826 451307 470854 451359
rect 470234 451295 470854 451307
rect 470234 451243 470262 451295
rect 470314 451243 470326 451295
rect 470378 451243 470390 451295
rect 470442 451243 470454 451295
rect 470506 451243 470518 451295
rect 470570 451243 470582 451295
rect 470634 451243 470646 451295
rect 470698 451243 470710 451295
rect 470762 451243 470774 451295
rect 470826 451243 470854 451295
rect 470234 451231 470854 451243
rect 470234 451179 470262 451231
rect 470314 451179 470326 451231
rect 470378 451179 470390 451231
rect 470442 451179 470454 451231
rect 470506 451179 470518 451231
rect 470570 451179 470582 451231
rect 470634 451179 470646 451231
rect 470698 451179 470710 451231
rect 470762 451179 470774 451231
rect 470826 451179 470854 451231
rect 470234 451173 470854 451179
rect 471624 450482 471652 450664
rect 471698 450482 471704 450494
rect 471624 450454 471704 450482
rect 471698 450442 471704 450454
rect 471756 450442 471762 450494
rect 468994 450401 469614 450407
rect 468994 450349 469022 450401
rect 469074 450349 469086 450401
rect 469138 450349 469150 450401
rect 469202 450349 469214 450401
rect 469266 450349 469278 450401
rect 469330 450349 469342 450401
rect 469394 450349 469406 450401
rect 469458 450349 469470 450401
rect 469522 450349 469534 450401
rect 469586 450349 469614 450401
rect 468994 450337 469614 450349
rect 468994 450285 469022 450337
rect 469074 450285 469086 450337
rect 469138 450285 469150 450337
rect 469202 450285 469214 450337
rect 469266 450285 469278 450337
rect 469330 450285 469342 450337
rect 469394 450285 469406 450337
rect 469458 450285 469470 450337
rect 469522 450285 469534 450337
rect 469586 450285 469614 450337
rect 468994 450273 469614 450285
rect 468994 450221 469022 450273
rect 469074 450221 469086 450273
rect 469138 450221 469150 450273
rect 469202 450221 469214 450273
rect 469266 450221 469278 450273
rect 469330 450221 469342 450273
rect 469394 450221 469406 450273
rect 469458 450221 469470 450273
rect 469522 450221 469534 450273
rect 469586 450221 469614 450273
rect 468994 450209 469614 450221
rect 468994 450157 469022 450209
rect 469074 450157 469086 450209
rect 469138 450157 469150 450209
rect 469202 450157 469214 450209
rect 469266 450157 469278 450209
rect 469330 450157 469342 450209
rect 469394 450157 469406 450209
rect 469458 450157 469470 450209
rect 469522 450157 469534 450209
rect 469586 450157 469614 450209
rect 468994 450145 469614 450157
rect 468994 450093 469022 450145
rect 469074 450093 469086 450145
rect 469138 450093 469150 450145
rect 469202 450093 469214 450145
rect 469266 450093 469278 450145
rect 469330 450093 469342 450145
rect 469394 450093 469406 450145
rect 469458 450093 469470 450145
rect 469522 450093 469534 450145
rect 469586 450093 469614 450145
rect 468994 450087 469614 450093
rect 475378 449438 475384 449490
rect 475436 449438 475442 449490
rect 478690 449438 478696 449490
rect 478748 449438 478754 449490
rect 482002 449438 482008 449490
rect 482060 449438 482066 449490
rect 485314 449438 485320 449490
rect 485372 449438 485378 449490
rect 488644 449394 488672 449464
rect 491938 449394 491944 449406
rect 488644 449366 491944 449394
rect 491938 449354 491944 449366
rect 491996 449354 492002 449406
rect 470234 449316 470854 449322
rect 470234 449264 470262 449316
rect 470314 449264 470326 449316
rect 470378 449264 470390 449316
rect 470442 449264 470454 449316
rect 470506 449264 470518 449316
rect 470570 449264 470582 449316
rect 470634 449264 470646 449316
rect 470698 449264 470710 449316
rect 470762 449264 470774 449316
rect 470826 449264 470854 449316
rect 470234 449252 470854 449264
rect 470234 449200 470262 449252
rect 470314 449200 470326 449252
rect 470378 449200 470390 449252
rect 470442 449200 470454 449252
rect 470506 449200 470518 449252
rect 470570 449200 470582 449252
rect 470634 449200 470646 449252
rect 470698 449200 470710 449252
rect 470762 449200 470774 449252
rect 470826 449200 470854 449252
rect 470234 449188 470854 449200
rect 470234 449136 470262 449188
rect 470314 449136 470326 449188
rect 470378 449136 470390 449188
rect 470442 449136 470454 449188
rect 470506 449136 470518 449188
rect 470570 449136 470582 449188
rect 470634 449136 470646 449188
rect 470698 449136 470710 449188
rect 470762 449136 470774 449188
rect 470826 449136 470854 449188
rect 470234 449124 470854 449136
rect 470234 449072 470262 449124
rect 470314 449072 470326 449124
rect 470378 449072 470390 449124
rect 470442 449072 470454 449124
rect 470506 449072 470518 449124
rect 470570 449072 470582 449124
rect 470634 449072 470646 449124
rect 470698 449072 470710 449124
rect 470762 449072 470774 449124
rect 470826 449072 470854 449124
rect 470234 449060 470854 449072
rect 470234 449008 470262 449060
rect 470314 449008 470326 449060
rect 470378 449008 470390 449060
rect 470442 449008 470454 449060
rect 470506 449008 470518 449060
rect 470570 449008 470582 449060
rect 470634 449008 470646 449060
rect 470698 449008 470710 449060
rect 470762 449008 470774 449060
rect 470826 449008 470854 449060
rect 470234 449002 470854 449008
rect 478690 446226 478696 446278
rect 478748 446266 478754 446278
rect 478748 446238 480254 446266
rect 478748 446226 478754 446238
rect 480226 445926 480254 446238
rect 515398 445926 515404 445938
rect 480226 445898 515404 445926
rect 515398 445886 515404 445898
rect 515456 445886 515462 445938
rect 482002 445818 482008 445870
rect 482060 445818 482066 445870
rect 485314 445818 485320 445870
rect 485372 445858 485378 445870
rect 523678 445858 523684 445870
rect 485372 445830 523684 445858
rect 485372 445818 485378 445830
rect 523678 445818 523684 445830
rect 523736 445818 523742 445870
rect 482020 445790 482048 445818
rect 520918 445790 520924 445802
rect 482020 445762 520924 445790
rect 520918 445750 520924 445762
rect 520976 445750 520982 445802
rect 475378 445682 475384 445734
rect 475436 445722 475442 445734
rect 535454 445722 535460 445734
rect 475436 445694 535460 445722
rect 475436 445682 475442 445694
rect 535454 445682 535460 445694
rect 535512 445682 535518 445734
rect 546954 445138 546960 445190
rect 547012 445178 547018 445190
rect 547506 445178 547512 445190
rect 547012 445150 547512 445178
rect 547012 445138 547018 445150
rect 547506 445138 547512 445150
rect 547564 445138 547570 445190
rect 490558 442962 490564 443014
rect 490616 443002 490622 443014
rect 535454 443002 535460 443014
rect 490616 442974 535460 443002
rect 490616 442962 490622 442974
rect 535454 442962 535460 442974
rect 535512 442962 535518 443014
rect 493318 441602 493324 441654
rect 493376 441642 493382 441654
rect 535454 441642 535460 441654
rect 493376 441614 535460 441642
rect 493376 441602 493382 441614
rect 535454 441602 535460 441614
rect 535512 441602 535518 441654
rect 494698 440242 494704 440294
rect 494756 440282 494762 440294
rect 535454 440282 535460 440294
rect 494756 440254 535460 440282
rect 494756 440242 494762 440254
rect 535454 440242 535460 440254
rect 535512 440242 535518 440294
rect 496078 438882 496084 438934
rect 496136 438922 496142 438934
rect 535454 438922 535460 438934
rect 496136 438894 535460 438922
rect 496136 438882 496142 438894
rect 535454 438882 535460 438894
rect 535512 438882 535518 438934
rect 497458 437454 497464 437506
rect 497516 437494 497522 437506
rect 535454 437494 535460 437506
rect 497516 437466 535460 437494
rect 497516 437454 497522 437466
rect 535454 437454 535460 437466
rect 535512 437454 535518 437506
rect 498838 436094 498844 436146
rect 498896 436134 498902 436146
rect 535454 436134 535460 436146
rect 498896 436106 535460 436134
rect 498896 436094 498902 436106
rect 535454 436094 535460 436106
rect 535512 436094 535518 436146
rect 500218 434734 500224 434786
rect 500276 434774 500282 434786
rect 535454 434774 535460 434786
rect 500276 434746 535460 434774
rect 500276 434734 500282 434746
rect 535454 434734 535460 434746
rect 535512 434734 535518 434786
rect 501598 433306 501604 433358
rect 501656 433346 501662 433358
rect 535454 433346 535460 433358
rect 501656 433318 535460 433346
rect 501656 433306 501662 433318
rect 535454 433306 535460 433318
rect 535512 433306 535518 433358
rect 470234 433088 470854 433094
rect 470234 433036 470262 433088
rect 470314 433036 470326 433088
rect 470378 433036 470390 433088
rect 470442 433036 470454 433088
rect 470506 433036 470518 433088
rect 470570 433036 470582 433088
rect 470634 433036 470646 433088
rect 470698 433036 470710 433088
rect 470762 433036 470774 433088
rect 470826 433036 470854 433088
rect 470234 433024 470854 433036
rect 470234 432972 470262 433024
rect 470314 432972 470326 433024
rect 470378 432972 470390 433024
rect 470442 432972 470454 433024
rect 470506 432972 470518 433024
rect 470570 432972 470582 433024
rect 470634 432972 470646 433024
rect 470698 432972 470710 433024
rect 470762 432972 470774 433024
rect 470826 432972 470854 433024
rect 470234 432960 470854 432972
rect 470234 432908 470262 432960
rect 470314 432908 470326 432960
rect 470378 432908 470390 432960
rect 470442 432908 470454 432960
rect 470506 432908 470518 432960
rect 470570 432908 470582 432960
rect 470634 432908 470646 432960
rect 470698 432908 470710 432960
rect 470762 432908 470774 432960
rect 470826 432908 470854 432960
rect 470234 432896 470854 432908
rect 470234 432844 470262 432896
rect 470314 432844 470326 432896
rect 470378 432844 470390 432896
rect 470442 432844 470454 432896
rect 470506 432844 470518 432896
rect 470570 432844 470582 432896
rect 470634 432844 470646 432896
rect 470698 432844 470710 432896
rect 470762 432844 470774 432896
rect 470826 432844 470854 432896
rect 470234 432832 470854 432844
rect 470234 432780 470262 432832
rect 470314 432780 470326 432832
rect 470378 432780 470390 432832
rect 470442 432780 470454 432832
rect 470506 432780 470518 432832
rect 470570 432780 470582 432832
rect 470634 432780 470646 432832
rect 470698 432780 470710 432832
rect 470762 432780 470774 432832
rect 470826 432780 470854 432832
rect 470234 432774 470854 432780
rect 576994 432304 577614 432310
rect 471612 432292 471664 432298
rect 471612 432234 471664 432240
rect 576994 432252 577022 432304
rect 577074 432252 577086 432304
rect 577138 432252 577150 432304
rect 577202 432252 577214 432304
rect 577266 432252 577278 432304
rect 577330 432252 577342 432304
rect 577394 432252 577406 432304
rect 577458 432252 577470 432304
rect 577522 432252 577534 432304
rect 577586 432252 577614 432304
rect 576994 432240 577614 432252
rect 576994 432188 577022 432240
rect 577074 432188 577086 432240
rect 577138 432188 577150 432240
rect 577202 432188 577214 432240
rect 577266 432188 577278 432240
rect 577330 432188 577342 432240
rect 577394 432188 577406 432240
rect 577458 432188 577470 432240
rect 577522 432188 577534 432240
rect 577586 432188 577614 432240
rect 576994 432176 577614 432188
rect 576994 432124 577022 432176
rect 577074 432124 577086 432176
rect 577138 432124 577150 432176
rect 577202 432124 577214 432176
rect 577266 432124 577278 432176
rect 577330 432124 577342 432176
rect 577394 432124 577406 432176
rect 577458 432124 577470 432176
rect 577522 432124 577534 432176
rect 577586 432124 577614 432176
rect 576994 432112 577614 432124
rect 576994 432086 577022 432112
rect 576400 432060 577022 432086
rect 577074 432060 577086 432112
rect 577138 432060 577150 432112
rect 577202 432060 577214 432112
rect 577266 432060 577278 432112
rect 577330 432060 577342 432112
rect 577394 432060 577406 432112
rect 577458 432060 577470 432112
rect 577522 432060 577534 432112
rect 577586 432086 577614 432112
rect 577586 432060 577647 432086
rect 576400 432055 577647 432060
rect 576316 432048 577647 432055
rect 576316 432021 577022 432048
rect 468994 432001 469614 432007
rect 468994 431949 469022 432001
rect 469074 431949 469086 432001
rect 469138 431949 469150 432001
rect 469202 431949 469214 432001
rect 469266 431949 469278 432001
rect 469330 431949 469342 432001
rect 469394 431949 469406 432001
rect 469458 431949 469470 432001
rect 469522 431949 469534 432001
rect 469586 431949 469614 432001
rect 468994 431937 469614 431949
rect 502978 431946 502984 431998
rect 503036 431986 503042 431998
rect 535454 431986 535460 431998
rect 503036 431958 535460 431986
rect 503036 431946 503042 431958
rect 535454 431946 535460 431958
rect 535512 431946 535518 431998
rect 576400 431996 577022 432021
rect 577074 431996 577086 432048
rect 577138 431996 577150 432048
rect 577202 431996 577214 432048
rect 577266 431996 577278 432048
rect 577330 431996 577342 432048
rect 577394 431996 577406 432048
rect 577458 431996 577470 432048
rect 577522 431996 577534 432048
rect 577586 431996 577647 432048
rect 576400 431990 577647 431996
rect 468994 431885 469022 431937
rect 469074 431885 469086 431937
rect 469138 431885 469150 431937
rect 469202 431885 469214 431937
rect 469266 431885 469278 431937
rect 469330 431885 469342 431937
rect 469394 431885 469406 431937
rect 469458 431885 469470 431937
rect 469522 431885 469534 431937
rect 469586 431885 469614 431937
rect 468994 431873 469614 431885
rect 468994 431821 469022 431873
rect 469074 431821 469086 431873
rect 469138 431821 469150 431873
rect 469202 431821 469214 431873
rect 469266 431821 469278 431873
rect 469330 431821 469342 431873
rect 469394 431821 469406 431873
rect 469458 431821 469470 431873
rect 469522 431821 469534 431873
rect 469586 431821 469614 431873
rect 468994 431809 469614 431821
rect 468994 431757 469022 431809
rect 469074 431757 469086 431809
rect 469138 431757 469150 431809
rect 469202 431757 469214 431809
rect 469266 431757 469278 431809
rect 469330 431757 469342 431809
rect 469394 431757 469406 431809
rect 469458 431757 469470 431809
rect 469522 431757 469534 431809
rect 469586 431757 469614 431809
rect 468994 431745 469614 431757
rect 468994 431693 469022 431745
rect 469074 431693 469086 431745
rect 469138 431693 469150 431745
rect 469202 431693 469214 431745
rect 469266 431693 469278 431745
rect 469330 431693 469342 431745
rect 469394 431693 469406 431745
rect 469458 431693 469470 431745
rect 469522 431693 469534 431745
rect 469586 431693 469614 431745
rect 468994 431687 469614 431693
rect 576597 431570 576603 431622
rect 576655 431570 576661 431622
rect 576400 431509 578876 431542
rect 576400 431457 578262 431509
rect 578314 431457 578326 431509
rect 578378 431457 578390 431509
rect 578442 431457 578454 431509
rect 578506 431457 578518 431509
rect 578570 431457 578582 431509
rect 578634 431457 578646 431509
rect 578698 431457 578710 431509
rect 578762 431457 578774 431509
rect 578826 431457 578876 431509
rect 478966 431451 478972 431454
rect 478931 431445 478972 431451
rect 478931 431411 478943 431445
rect 478931 431405 478972 431411
rect 478966 431402 478972 431405
rect 479024 431402 479030 431454
rect 485774 431402 485780 431454
rect 485832 431451 485838 431454
rect 485832 431445 485877 431451
rect 576400 431446 578876 431457
rect 485865 431411 485877 431445
rect 485832 431405 485877 431411
rect 578234 431445 578854 431446
rect 485832 431402 485838 431405
rect 578234 431393 578262 431445
rect 578314 431393 578326 431445
rect 578378 431393 578390 431445
rect 578442 431393 578454 431445
rect 578506 431393 578518 431445
rect 578570 431393 578582 431445
rect 578634 431393 578646 431445
rect 578698 431393 578710 431445
rect 578762 431393 578774 431445
rect 578826 431393 578854 431445
rect 578234 431381 578854 431393
rect 578234 431329 578262 431381
rect 578314 431329 578326 431381
rect 578378 431329 578390 431381
rect 578442 431329 578454 431381
rect 578506 431329 578518 431381
rect 578570 431329 578582 431381
rect 578634 431329 578646 431381
rect 578698 431329 578710 431381
rect 578762 431329 578774 431381
rect 578826 431329 578854 431381
rect 578234 431317 578854 431329
rect 578234 431265 578262 431317
rect 578314 431265 578326 431317
rect 578378 431265 578390 431317
rect 578442 431265 578454 431317
rect 578506 431265 578518 431317
rect 578570 431265 578582 431317
rect 578634 431265 578646 431317
rect 578698 431265 578710 431317
rect 578762 431265 578774 431317
rect 578826 431265 578854 431317
rect 578234 431253 578854 431265
rect 578234 431201 578262 431253
rect 578314 431201 578326 431253
rect 578378 431201 578390 431253
rect 578442 431201 578454 431253
rect 578506 431201 578518 431253
rect 578570 431201 578582 431253
rect 578634 431201 578646 431253
rect 578698 431201 578710 431253
rect 578762 431201 578774 431253
rect 578826 431201 578854 431253
rect 578234 431195 578854 431201
rect 475470 431037 475476 431089
rect 475528 431037 475534 431089
rect 482370 431037 482376 431089
rect 482428 431037 482434 431089
rect 489302 431049 489592 431077
rect 489564 431034 489592 431049
rect 492030 431034 492036 431046
rect 489564 431006 492036 431034
rect 492030 430994 492036 431006
rect 492088 430994 492094 431046
rect 470234 430916 470854 430922
rect 470234 430864 470262 430916
rect 470314 430864 470326 430916
rect 470378 430864 470390 430916
rect 470442 430864 470454 430916
rect 470506 430864 470518 430916
rect 470570 430864 470582 430916
rect 470634 430864 470646 430916
rect 470698 430864 470710 430916
rect 470762 430864 470774 430916
rect 470826 430864 470854 430916
rect 470234 430852 470854 430864
rect 470234 430800 470262 430852
rect 470314 430800 470326 430852
rect 470378 430800 470390 430852
rect 470442 430800 470454 430852
rect 470506 430800 470518 430852
rect 470570 430800 470582 430852
rect 470634 430800 470646 430852
rect 470698 430800 470710 430852
rect 470762 430800 470774 430852
rect 470826 430800 470854 430852
rect 470234 430788 470854 430800
rect 470234 430736 470262 430788
rect 470314 430736 470326 430788
rect 470378 430736 470390 430788
rect 470442 430736 470454 430788
rect 470506 430736 470518 430788
rect 470570 430736 470582 430788
rect 470634 430736 470646 430788
rect 470698 430736 470710 430788
rect 470762 430736 470774 430788
rect 470826 430736 470854 430788
rect 470234 430724 470854 430736
rect 470234 430672 470262 430724
rect 470314 430672 470326 430724
rect 470378 430672 470390 430724
rect 470442 430672 470454 430724
rect 470506 430672 470518 430724
rect 470570 430672 470582 430724
rect 470634 430672 470646 430724
rect 470698 430672 470710 430724
rect 470762 430672 470774 430724
rect 470826 430672 470854 430724
rect 470234 430660 470854 430672
rect 470234 430608 470262 430660
rect 470314 430608 470326 430660
rect 470378 430608 470390 430660
rect 470442 430608 470454 430660
rect 470506 430608 470518 430660
rect 470570 430608 470582 430660
rect 470634 430608 470646 430660
rect 470698 430608 470710 430660
rect 470762 430608 470774 430660
rect 470826 430608 470854 430660
rect 470234 430602 470854 430608
rect 475470 429090 475476 429142
rect 475528 429130 475534 429142
rect 490558 429130 490564 429142
rect 475528 429102 490564 429130
rect 475528 429090 475534 429102
rect 490558 429090 490564 429102
rect 490616 429090 490622 429142
rect 482370 427798 482376 427850
rect 482428 427838 482434 427850
rect 522298 427838 522304 427850
rect 482428 427810 522304 427838
rect 482428 427798 482434 427810
rect 522298 427798 522304 427810
rect 522356 427798 522362 427850
rect 470234 412088 470854 412094
rect 470234 412036 470262 412088
rect 470314 412036 470326 412088
rect 470378 412036 470390 412088
rect 470442 412036 470454 412088
rect 470506 412036 470518 412088
rect 470570 412036 470582 412088
rect 470634 412036 470646 412088
rect 470698 412036 470710 412088
rect 470762 412036 470774 412088
rect 470826 412036 470854 412088
rect 470234 412024 470854 412036
rect 470234 411972 470262 412024
rect 470314 411972 470326 412024
rect 470378 411972 470390 412024
rect 470442 411972 470454 412024
rect 470506 411972 470518 412024
rect 470570 411972 470582 412024
rect 470634 411972 470646 412024
rect 470698 411972 470710 412024
rect 470762 411972 470774 412024
rect 470826 411972 470854 412024
rect 470234 411960 470854 411972
rect 470234 411908 470262 411960
rect 470314 411908 470326 411960
rect 470378 411908 470390 411960
rect 470442 411908 470454 411960
rect 470506 411908 470518 411960
rect 470570 411908 470582 411960
rect 470634 411908 470646 411960
rect 470698 411908 470710 411960
rect 470762 411908 470774 411960
rect 470826 411908 470854 411960
rect 470234 411896 470854 411908
rect 470234 411844 470262 411896
rect 470314 411844 470326 411896
rect 470378 411844 470390 411896
rect 470442 411844 470454 411896
rect 470506 411844 470518 411896
rect 470570 411844 470582 411896
rect 470634 411844 470646 411896
rect 470698 411844 470710 411896
rect 470762 411844 470774 411896
rect 470826 411844 470854 411896
rect 470234 411832 470854 411844
rect 470234 411780 470262 411832
rect 470314 411780 470326 411832
rect 470378 411780 470390 411832
rect 470442 411780 470454 411832
rect 470506 411780 470518 411832
rect 470570 411780 470582 411832
rect 470634 411780 470646 411832
rect 470698 411780 470710 411832
rect 470762 411780 470774 411832
rect 470826 411780 470854 411832
rect 470234 411774 470854 411780
rect 471238 411206 471244 411258
rect 471296 411246 471302 411258
rect 471624 411246 471652 411265
rect 471296 411218 471652 411246
rect 473722 411234 473728 411286
rect 473780 411234 473786 411286
rect 471296 411206 471302 411218
rect 468994 411002 469614 411008
rect 468994 410950 469022 411002
rect 469074 410950 469086 411002
rect 469138 410950 469150 411002
rect 469202 410950 469214 411002
rect 469266 410950 469278 411002
rect 469330 410950 469342 411002
rect 469394 410950 469406 411002
rect 469458 410950 469470 411002
rect 469522 410950 469534 411002
rect 469586 410950 469614 411002
rect 468994 410938 469614 410950
rect 468994 410886 469022 410938
rect 469074 410886 469086 410938
rect 469138 410886 469150 410938
rect 469202 410886 469214 410938
rect 469266 410886 469278 410938
rect 469330 410886 469342 410938
rect 469394 410886 469406 410938
rect 469458 410886 469470 410938
rect 469522 410886 469534 410938
rect 469586 410886 469614 410938
rect 468994 410874 469614 410886
rect 468994 410822 469022 410874
rect 469074 410822 469086 410874
rect 469138 410822 469150 410874
rect 469202 410822 469214 410874
rect 469266 410822 469278 410874
rect 469330 410822 469342 410874
rect 469394 410822 469406 410874
rect 469458 410822 469470 410874
rect 469522 410822 469534 410874
rect 469586 410822 469614 410874
rect 468994 410810 469614 410822
rect 468994 410758 469022 410810
rect 469074 410758 469086 410810
rect 469138 410758 469150 410810
rect 469202 410758 469214 410810
rect 469266 410758 469278 410810
rect 469330 410758 469342 410810
rect 469394 410758 469406 410810
rect 469458 410758 469470 410810
rect 469522 410758 469534 410810
rect 469586 410758 469614 410810
rect 468994 410746 469614 410758
rect 468994 410694 469022 410746
rect 469074 410694 469086 410746
rect 469138 410694 469150 410746
rect 469202 410694 469214 410746
rect 469266 410694 469278 410746
rect 469330 410694 469342 410746
rect 469394 410694 469406 410746
rect 469458 410694 469470 410746
rect 469522 410694 469534 410746
rect 469586 410694 469614 410746
rect 468994 410688 469614 410694
rect 477788 410442 478472 410447
rect 477788 410419 478420 410442
rect 478414 410390 478420 410419
rect 478472 410390 478478 410442
rect 478598 410439 478604 410442
rect 478569 410433 478604 410439
rect 478569 410399 478581 410433
rect 478569 410393 478604 410399
rect 478598 410390 478604 410393
rect 478656 410390 478662 410442
rect 485130 410439 485136 410442
rect 485099 410433 485136 410439
rect 485099 410399 485111 410433
rect 485099 410393 485136 410399
rect 485130 410390 485136 410393
rect 485188 410390 485194 410442
rect 475286 410038 475292 410090
rect 475344 410038 475350 410090
rect 481818 410038 481824 410090
rect 481876 410038 481882 410090
rect 488382 410050 488672 410078
rect 488644 410022 488672 410050
rect 490742 410022 490748 410034
rect 488644 409994 490748 410022
rect 490742 409982 490748 409994
rect 490800 409982 490806 410034
rect 470234 409916 470854 409922
rect 470234 409864 470262 409916
rect 470314 409864 470326 409916
rect 470378 409864 470390 409916
rect 470442 409864 470454 409916
rect 470506 409864 470518 409916
rect 470570 409864 470582 409916
rect 470634 409864 470646 409916
rect 470698 409864 470710 409916
rect 470762 409864 470774 409916
rect 470826 409864 470854 409916
rect 470234 409852 470854 409864
rect 470234 409800 470262 409852
rect 470314 409800 470326 409852
rect 470378 409800 470390 409852
rect 470442 409800 470454 409852
rect 470506 409800 470518 409852
rect 470570 409800 470582 409852
rect 470634 409800 470646 409852
rect 470698 409800 470710 409852
rect 470762 409800 470774 409852
rect 470826 409800 470854 409852
rect 470234 409788 470854 409800
rect 470234 409736 470262 409788
rect 470314 409736 470326 409788
rect 470378 409736 470390 409788
rect 470442 409736 470454 409788
rect 470506 409736 470518 409788
rect 470570 409736 470582 409788
rect 470634 409736 470646 409788
rect 470698 409736 470710 409788
rect 470762 409736 470774 409788
rect 470826 409736 470854 409788
rect 515398 409778 515404 409830
rect 515456 409818 515462 409830
rect 535454 409818 535460 409830
rect 515456 409790 535460 409818
rect 515456 409778 515462 409790
rect 535454 409778 535460 409790
rect 535512 409778 535518 409830
rect 470234 409724 470854 409736
rect 470234 409672 470262 409724
rect 470314 409672 470326 409724
rect 470378 409672 470390 409724
rect 470442 409672 470454 409724
rect 470506 409672 470518 409724
rect 470570 409672 470582 409724
rect 470634 409672 470646 409724
rect 470698 409672 470710 409724
rect 470762 409672 470774 409724
rect 470826 409672 470854 409724
rect 470234 409660 470854 409672
rect 470234 409608 470262 409660
rect 470314 409608 470326 409660
rect 470378 409608 470390 409660
rect 470442 409608 470454 409660
rect 470506 409608 470518 409660
rect 470570 409608 470582 409660
rect 470634 409608 470646 409660
rect 470698 409608 470710 409660
rect 470762 409608 470774 409660
rect 470826 409608 470854 409660
rect 470234 409602 470854 409608
rect 475286 408418 475292 408470
rect 475344 408458 475350 408470
rect 493318 408458 493324 408470
rect 475344 408430 493324 408458
rect 475344 408418 475350 408430
rect 493318 408418 493324 408430
rect 493376 408418 493382 408470
rect 547230 408146 547236 408198
rect 547288 408186 547294 408198
rect 547506 408186 547512 408198
rect 547288 408158 547512 408186
rect 547288 408146 547294 408158
rect 547506 408146 547512 408158
rect 547564 408146 547570 408198
rect 478598 407058 478604 407110
rect 478656 407098 478662 407110
rect 535454 407098 535460 407110
rect 478656 407070 535460 407098
rect 478656 407058 478662 407070
rect 535454 407058 535460 407070
rect 535512 407058 535518 407110
rect 515398 404338 515404 404390
rect 515456 404378 515462 404390
rect 535454 404378 535460 404390
rect 515456 404350 535460 404378
rect 515456 404338 515462 404350
rect 535454 404338 535460 404350
rect 535512 404338 535518 404390
rect 516778 402978 516784 403030
rect 516836 403018 516842 403030
rect 535454 403018 535460 403030
rect 516836 402990 535460 403018
rect 516836 402978 516842 402990
rect 535454 402978 535460 402990
rect 535512 402978 535518 403030
rect 518158 398830 518164 398882
rect 518216 398870 518222 398882
rect 535454 398870 535460 398882
rect 518216 398842 535460 398870
rect 518216 398830 518222 398842
rect 535454 398830 535460 398842
rect 535512 398830 535518 398882
rect 519538 396042 519544 396094
rect 519596 396082 519602 396094
rect 535454 396082 535460 396094
rect 519596 396054 535460 396082
rect 519596 396042 519602 396054
rect 535454 396042 535460 396054
rect 535512 396042 535518 396094
rect 470234 391089 470854 391095
rect 470234 391037 470262 391089
rect 470314 391037 470326 391089
rect 470378 391037 470390 391089
rect 470442 391037 470454 391089
rect 470506 391037 470518 391089
rect 470570 391037 470582 391089
rect 470634 391037 470646 391089
rect 470698 391037 470710 391089
rect 470762 391037 470774 391089
rect 470826 391037 470854 391089
rect 470234 391025 470854 391037
rect 470234 390973 470262 391025
rect 470314 390973 470326 391025
rect 470378 390973 470390 391025
rect 470442 390973 470454 391025
rect 470506 390973 470518 391025
rect 470570 390973 470582 391025
rect 470634 390973 470646 391025
rect 470698 390973 470710 391025
rect 470762 390973 470774 391025
rect 470826 390973 470854 391025
rect 470234 390961 470854 390973
rect 470234 390909 470262 390961
rect 470314 390909 470326 390961
rect 470378 390909 470390 390961
rect 470442 390909 470454 390961
rect 470506 390909 470518 390961
rect 470570 390909 470582 390961
rect 470634 390909 470646 390961
rect 470698 390909 470710 390961
rect 470762 390909 470774 390961
rect 470826 390909 470854 390961
rect 470234 390897 470854 390909
rect 470234 390845 470262 390897
rect 470314 390845 470326 390897
rect 470378 390845 470390 390897
rect 470442 390845 470454 390897
rect 470506 390845 470518 390897
rect 470570 390845 470582 390897
rect 470634 390845 470646 390897
rect 470698 390845 470710 390897
rect 470762 390845 470774 390897
rect 470826 390845 470854 390897
rect 470234 390833 470854 390845
rect 470234 390781 470262 390833
rect 470314 390781 470326 390833
rect 470378 390781 470390 390833
rect 470442 390781 470454 390833
rect 470506 390781 470518 390833
rect 470570 390781 470582 390833
rect 470634 390781 470646 390833
rect 470698 390781 470710 390833
rect 470762 390781 470774 390833
rect 470826 390781 470854 390833
rect 470234 390775 470854 390781
rect 471238 390262 471244 390314
rect 471296 390302 471302 390314
rect 471296 390274 471652 390302
rect 471296 390262 471302 390274
rect 471624 390098 471652 390274
rect 471698 390098 471704 390110
rect 471624 390070 471704 390098
rect 471698 390058 471704 390070
rect 471756 390058 471762 390110
rect 468994 390006 469614 390012
rect 468994 389954 469022 390006
rect 469074 389954 469086 390006
rect 469138 389954 469150 390006
rect 469202 389954 469214 390006
rect 469266 389954 469278 390006
rect 469330 389954 469342 390006
rect 469394 389954 469406 390006
rect 469458 389954 469470 390006
rect 469522 389954 469534 390006
rect 469586 389954 469614 390006
rect 468994 389942 469614 389954
rect 468994 389890 469022 389942
rect 469074 389890 469086 389942
rect 469138 389890 469150 389942
rect 469202 389890 469214 389942
rect 469266 389890 469278 389942
rect 469330 389890 469342 389942
rect 469394 389890 469406 389942
rect 469458 389890 469470 389942
rect 469522 389890 469534 389942
rect 469586 389890 469614 389942
rect 468994 389878 469614 389890
rect 468994 389826 469022 389878
rect 469074 389826 469086 389878
rect 469138 389826 469150 389878
rect 469202 389826 469214 389878
rect 469266 389826 469278 389878
rect 469330 389826 469342 389878
rect 469394 389826 469406 389878
rect 469458 389826 469470 389878
rect 469522 389826 469534 389878
rect 469586 389826 469614 389878
rect 468994 389814 469614 389826
rect 468994 389762 469022 389814
rect 469074 389762 469086 389814
rect 469138 389762 469150 389814
rect 469202 389762 469214 389814
rect 469266 389762 469278 389814
rect 469330 389762 469342 389814
rect 469394 389762 469406 389814
rect 469458 389762 469470 389814
rect 469522 389762 469534 389814
rect 469586 389762 469614 389814
rect 468994 389750 469614 389762
rect 468994 389698 469022 389750
rect 469074 389698 469086 389750
rect 469138 389698 469150 389750
rect 469202 389698 469214 389750
rect 469266 389698 469278 389750
rect 469330 389698 469342 389750
rect 469394 389698 469406 389750
rect 469458 389698 469470 389750
rect 469522 389698 469534 389750
rect 469586 389698 469614 389750
rect 468994 389692 469614 389698
rect 479426 389446 479432 389498
rect 479484 389495 479490 389498
rect 479484 389489 479520 389495
rect 479508 389455 479520 389489
rect 479484 389449 479520 389455
rect 490598 389489 490656 389495
rect 490598 389455 490610 389489
rect 490644 389486 490656 389489
rect 493318 389486 493324 389498
rect 490644 389458 493324 389486
rect 490644 389455 490656 389458
rect 490598 389449 490656 389455
rect 479484 389446 479490 389449
rect 493318 389446 493324 389458
rect 493376 389446 493382 389498
rect 475746 389038 475752 389090
rect 475804 389038 475810 389090
rect 483198 389038 483204 389090
rect 483256 389038 483262 389090
rect 486878 389038 486884 389090
rect 486936 389038 486942 389090
rect 470234 388916 470854 388922
rect 470234 388864 470262 388916
rect 470314 388864 470326 388916
rect 470378 388864 470390 388916
rect 470442 388864 470454 388916
rect 470506 388864 470518 388916
rect 470570 388864 470582 388916
rect 470634 388864 470646 388916
rect 470698 388864 470710 388916
rect 470762 388864 470774 388916
rect 470826 388864 470854 388916
rect 470234 388852 470854 388864
rect 470234 388800 470262 388852
rect 470314 388800 470326 388852
rect 470378 388800 470390 388852
rect 470442 388800 470454 388852
rect 470506 388800 470518 388852
rect 470570 388800 470582 388852
rect 470634 388800 470646 388852
rect 470698 388800 470710 388852
rect 470762 388800 470774 388852
rect 470826 388800 470854 388852
rect 470234 388788 470854 388800
rect 470234 388736 470262 388788
rect 470314 388736 470326 388788
rect 470378 388736 470390 388788
rect 470442 388736 470454 388788
rect 470506 388736 470518 388788
rect 470570 388736 470582 388788
rect 470634 388736 470646 388788
rect 470698 388736 470710 388788
rect 470762 388736 470774 388788
rect 470826 388736 470854 388788
rect 470234 388724 470854 388736
rect 470234 388672 470262 388724
rect 470314 388672 470326 388724
rect 470378 388672 470390 388724
rect 470442 388672 470454 388724
rect 470506 388672 470518 388724
rect 470570 388672 470582 388724
rect 470634 388672 470646 388724
rect 470698 388672 470710 388724
rect 470762 388672 470774 388724
rect 470826 388672 470854 388724
rect 470234 388660 470854 388672
rect 470234 388608 470262 388660
rect 470314 388608 470326 388660
rect 470378 388608 470390 388660
rect 470442 388608 470454 388660
rect 470506 388608 470518 388660
rect 470570 388608 470582 388660
rect 470634 388608 470646 388660
rect 470698 388608 470710 388660
rect 470762 388608 470774 388660
rect 470826 388608 470854 388660
rect 470234 388602 470854 388608
rect 475746 387746 475752 387798
rect 475804 387746 475810 387798
rect 479426 387746 479432 387798
rect 479484 387786 479490 387798
rect 515398 387786 515404 387798
rect 479484 387758 515404 387786
rect 479484 387746 479490 387758
rect 515398 387746 515404 387758
rect 515456 387746 515462 387798
rect 475764 387718 475792 387746
rect 494698 387718 494704 387730
rect 475764 387690 494704 387718
rect 494698 387678 494704 387690
rect 494756 387678 494762 387730
rect 483198 386386 483204 386438
rect 483256 386426 483262 386438
rect 484302 386426 484308 386438
rect 483256 386398 484308 386426
rect 483256 386386 483262 386398
rect 484302 386386 484308 386398
rect 484360 386386 484366 386438
rect 576994 379128 577614 379134
rect 576994 379076 577022 379128
rect 577074 379076 577086 379128
rect 577138 379076 577150 379128
rect 577202 379076 577214 379128
rect 577266 379076 577278 379128
rect 577330 379076 577342 379128
rect 577394 379076 577406 379128
rect 577458 379076 577470 379128
rect 577522 379076 577534 379128
rect 577586 379076 577614 379128
rect 576994 379064 577614 379076
rect 576994 379012 577022 379064
rect 577074 379012 577086 379064
rect 577138 379012 577150 379064
rect 577202 379012 577214 379064
rect 577266 379012 577278 379064
rect 577330 379012 577342 379064
rect 577394 379012 577406 379064
rect 577458 379012 577470 379064
rect 577522 379012 577534 379064
rect 577586 379012 577614 379064
rect 576994 379000 577614 379012
rect 576994 378948 577022 379000
rect 577074 378948 577086 379000
rect 577138 378948 577150 379000
rect 577202 378948 577214 379000
rect 577266 378948 577278 379000
rect 577330 378948 577342 379000
rect 577394 378948 577406 379000
rect 577458 378948 577470 379000
rect 577522 378948 577534 379000
rect 577586 378948 577614 379000
rect 576994 378936 577614 378948
rect 576994 378910 577022 378936
rect 576400 378884 577022 378910
rect 577074 378884 577086 378936
rect 577138 378884 577150 378936
rect 577202 378884 577214 378936
rect 577266 378884 577278 378936
rect 577330 378884 577342 378936
rect 577394 378884 577406 378936
rect 577458 378884 577470 378936
rect 577522 378884 577534 378936
rect 577586 378910 577614 378936
rect 577586 378884 577647 378910
rect 576400 378879 577647 378884
rect 576316 378872 577647 378879
rect 576316 378845 577022 378872
rect 576400 378820 577022 378845
rect 577074 378820 577086 378872
rect 577138 378820 577150 378872
rect 577202 378820 577214 378872
rect 577266 378820 577278 378872
rect 577330 378820 577342 378872
rect 577394 378820 577406 378872
rect 577458 378820 577470 378872
rect 577522 378820 577534 378872
rect 577586 378820 577647 378872
rect 576400 378814 577647 378820
rect 576597 378394 576603 378446
rect 576655 378394 576661 378446
rect 576400 378333 578876 378366
rect 576400 378281 578262 378333
rect 578314 378281 578326 378333
rect 578378 378281 578390 378333
rect 578442 378281 578454 378333
rect 578506 378281 578518 378333
rect 578570 378281 578582 378333
rect 578634 378281 578646 378333
rect 578698 378281 578710 378333
rect 578762 378281 578774 378333
rect 578826 378281 578876 378333
rect 576400 378270 578876 378281
rect 578234 378269 578854 378270
rect 578234 378217 578262 378269
rect 578314 378217 578326 378269
rect 578378 378217 578390 378269
rect 578442 378217 578454 378269
rect 578506 378217 578518 378269
rect 578570 378217 578582 378269
rect 578634 378217 578646 378269
rect 578698 378217 578710 378269
rect 578762 378217 578774 378269
rect 578826 378217 578854 378269
rect 578234 378205 578854 378217
rect 578234 378153 578262 378205
rect 578314 378153 578326 378205
rect 578378 378153 578390 378205
rect 578442 378153 578454 378205
rect 578506 378153 578518 378205
rect 578570 378153 578582 378205
rect 578634 378153 578646 378205
rect 578698 378153 578710 378205
rect 578762 378153 578774 378205
rect 578826 378153 578854 378205
rect 578234 378141 578854 378153
rect 578234 378089 578262 378141
rect 578314 378089 578326 378141
rect 578378 378089 578390 378141
rect 578442 378089 578454 378141
rect 578506 378089 578518 378141
rect 578570 378089 578582 378141
rect 578634 378089 578646 378141
rect 578698 378089 578710 378141
rect 578762 378089 578774 378141
rect 578826 378089 578854 378141
rect 578234 378077 578854 378089
rect 578234 378025 578262 378077
rect 578314 378025 578326 378077
rect 578378 378025 578390 378077
rect 578442 378025 578454 378077
rect 578506 378025 578518 378077
rect 578570 378025 578582 378077
rect 578634 378025 578646 378077
rect 578698 378025 578710 378077
rect 578762 378025 578774 378077
rect 578826 378025 578854 378077
rect 578234 378019 578854 378025
rect 520918 373942 520924 373994
rect 520976 373982 520982 373994
rect 535454 373982 535460 373994
rect 520976 373954 535460 373982
rect 520976 373942 520982 373954
rect 535454 373942 535460 373954
rect 535512 373942 535518 373994
rect 547046 373262 547052 373314
rect 547104 373302 547110 373314
rect 547506 373302 547512 373314
rect 547104 373274 547512 373302
rect 547104 373262 547110 373274
rect 547506 373262 547512 373274
rect 547564 373262 547570 373314
rect 522298 372514 522304 372566
rect 522356 372554 522362 372566
rect 535454 372554 535460 372566
rect 522356 372526 535460 372554
rect 522356 372514 522362 372526
rect 535454 372514 535460 372526
rect 535512 372514 535518 372566
rect 484302 369794 484308 369846
rect 484360 369834 484366 369846
rect 535454 369834 535460 369846
rect 484360 369806 535460 369834
rect 484360 369794 484366 369806
rect 535454 369794 535460 369806
rect 535512 369794 535518 369846
rect 520918 367074 520924 367126
rect 520976 367114 520982 367126
rect 535454 367114 535460 367126
rect 520976 367086 535460 367114
rect 520976 367074 520982 367086
rect 535454 367074 535460 367086
rect 535512 367074 535518 367126
rect 515398 365714 515404 365766
rect 515456 365754 515462 365766
rect 535454 365754 535460 365766
rect 515456 365726 535460 365754
rect 515456 365714 515462 365726
rect 535454 365714 535460 365726
rect 535512 365714 535518 365766
rect 522298 361566 522304 361618
rect 522356 361606 522362 361618
rect 535454 361606 535460 361618
rect 522356 361578 535460 361606
rect 522356 361566 522362 361578
rect 535454 361566 535460 361578
rect 535512 361566 535518 361618
rect 470234 358489 470854 358495
rect 470234 358437 470262 358489
rect 470314 358437 470326 358489
rect 470378 358437 470390 358489
rect 470442 358437 470454 358489
rect 470506 358437 470518 358489
rect 470570 358437 470582 358489
rect 470634 358437 470646 358489
rect 470698 358437 470710 358489
rect 470762 358437 470774 358489
rect 470826 358437 470854 358489
rect 470234 358425 470854 358437
rect 470234 358373 470262 358425
rect 470314 358373 470326 358425
rect 470378 358373 470390 358425
rect 470442 358373 470454 358425
rect 470506 358373 470518 358425
rect 470570 358373 470582 358425
rect 470634 358373 470646 358425
rect 470698 358373 470710 358425
rect 470762 358373 470774 358425
rect 470826 358373 470854 358425
rect 470234 358361 470854 358373
rect 470234 358309 470262 358361
rect 470314 358309 470326 358361
rect 470378 358309 470390 358361
rect 470442 358309 470454 358361
rect 470506 358309 470518 358361
rect 470570 358309 470582 358361
rect 470634 358309 470646 358361
rect 470698 358309 470710 358361
rect 470762 358309 470774 358361
rect 470826 358309 470854 358361
rect 470234 358297 470854 358309
rect 470234 358245 470262 358297
rect 470314 358245 470326 358297
rect 470378 358245 470390 358297
rect 470442 358245 470454 358297
rect 470506 358245 470518 358297
rect 470570 358245 470582 358297
rect 470634 358245 470646 358297
rect 470698 358245 470710 358297
rect 470762 358245 470774 358297
rect 470826 358245 470854 358297
rect 470234 358233 470854 358245
rect 470234 358181 470262 358233
rect 470314 358181 470326 358233
rect 470378 358181 470390 358233
rect 470442 358181 470454 358233
rect 470506 358181 470518 358233
rect 470570 358181 470582 358233
rect 470634 358181 470646 358233
rect 470698 358181 470710 358233
rect 470762 358181 470774 358233
rect 470826 358181 470854 358233
rect 470234 358175 470854 358181
rect 471698 357554 471704 357606
rect 471756 357594 471762 357606
rect 473648 357594 473676 357666
rect 475102 357622 475108 357674
rect 475160 357622 475166 357674
rect 478874 357633 478880 357685
rect 478932 357633 478938 357685
rect 481818 357633 481824 357685
rect 481876 357633 481882 357685
rect 484946 357633 484952 357685
rect 485004 357633 485010 357685
rect 471756 357566 473676 357594
rect 471756 357554 471762 357566
rect 468994 357403 469614 357409
rect 468994 357351 469022 357403
rect 469074 357351 469086 357403
rect 469138 357351 469150 357403
rect 469202 357351 469214 357403
rect 469266 357351 469278 357403
rect 469330 357351 469342 357403
rect 469394 357351 469406 357403
rect 469458 357351 469470 357403
rect 469522 357351 469534 357403
rect 469586 357351 469614 357403
rect 468994 357339 469614 357351
rect 468994 357287 469022 357339
rect 469074 357287 469086 357339
rect 469138 357287 469150 357339
rect 469202 357287 469214 357339
rect 469266 357287 469278 357339
rect 469330 357287 469342 357339
rect 469394 357287 469406 357339
rect 469458 357287 469470 357339
rect 469522 357287 469534 357339
rect 469586 357287 469614 357339
rect 468994 357275 469614 357287
rect 468994 357223 469022 357275
rect 469074 357223 469086 357275
rect 469138 357223 469150 357275
rect 469202 357223 469214 357275
rect 469266 357223 469278 357275
rect 469330 357223 469342 357275
rect 469394 357223 469406 357275
rect 469458 357223 469470 357275
rect 469522 357223 469534 357275
rect 469586 357223 469614 357275
rect 468994 357211 469614 357223
rect 468994 357159 469022 357211
rect 469074 357159 469086 357211
rect 469138 357159 469150 357211
rect 469202 357159 469214 357211
rect 469266 357159 469278 357211
rect 469330 357159 469342 357211
rect 469394 357159 469406 357211
rect 469458 357159 469470 357211
rect 469522 357159 469534 357211
rect 469586 357159 469614 357211
rect 468994 357147 469614 357159
rect 468994 357095 469022 357147
rect 469074 357095 469086 357147
rect 469138 357095 469150 357147
rect 469202 357095 469214 357147
rect 469266 357095 469278 357147
rect 469330 357095 469342 357147
rect 469394 357095 469406 357147
rect 469458 357095 469470 357147
rect 469522 357095 469534 357147
rect 469586 357095 469614 357147
rect 468994 357089 469614 357095
rect 477034 356806 477040 356858
rect 477092 356855 477098 356858
rect 480162 356855 480168 356858
rect 477092 356849 477137 356855
rect 477125 356815 477137 356849
rect 477092 356809 477137 356815
rect 480131 356849 480168 356855
rect 480131 356815 480143 356849
rect 480131 356809 480168 356815
rect 477092 356806 477098 356809
rect 480162 356806 480168 356809
rect 480220 356806 480226 356858
rect 483198 356437 483204 356489
rect 483256 356437 483262 356489
rect 486234 356437 486240 356489
rect 486292 356437 486298 356489
rect 489288 356438 489316 356463
rect 492122 356438 492128 356450
rect 489288 356410 492128 356438
rect 492122 356398 492128 356410
rect 492180 356398 492186 356450
rect 470234 356316 470854 356322
rect 470234 356264 470262 356316
rect 470314 356264 470326 356316
rect 470378 356264 470390 356316
rect 470442 356264 470454 356316
rect 470506 356264 470518 356316
rect 470570 356264 470582 356316
rect 470634 356264 470646 356316
rect 470698 356264 470710 356316
rect 470762 356264 470774 356316
rect 470826 356264 470854 356316
rect 470234 356252 470854 356264
rect 470234 356200 470262 356252
rect 470314 356200 470326 356252
rect 470378 356200 470390 356252
rect 470442 356200 470454 356252
rect 470506 356200 470518 356252
rect 470570 356200 470582 356252
rect 470634 356200 470646 356252
rect 470698 356200 470710 356252
rect 470762 356200 470774 356252
rect 470826 356200 470854 356252
rect 470234 356188 470854 356200
rect 470234 356136 470262 356188
rect 470314 356136 470326 356188
rect 470378 356136 470390 356188
rect 470442 356136 470454 356188
rect 470506 356136 470518 356188
rect 470570 356136 470582 356188
rect 470634 356136 470646 356188
rect 470698 356136 470710 356188
rect 470762 356136 470774 356188
rect 470826 356136 470854 356188
rect 470234 356124 470854 356136
rect 470234 356072 470262 356124
rect 470314 356072 470326 356124
rect 470378 356072 470390 356124
rect 470442 356072 470454 356124
rect 470506 356072 470518 356124
rect 470570 356072 470582 356124
rect 470634 356072 470646 356124
rect 470698 356072 470710 356124
rect 470762 356072 470774 356124
rect 470826 356072 470854 356124
rect 470234 356060 470854 356072
rect 470234 356008 470262 356060
rect 470314 356008 470326 356060
rect 470378 356008 470390 356060
rect 470442 356008 470454 356060
rect 470506 356008 470518 356060
rect 470570 356008 470582 356060
rect 470634 356008 470646 356060
rect 470698 356008 470710 356060
rect 470762 356008 470774 356060
rect 470826 356008 470854 356060
rect 470234 356002 470854 356008
rect 483198 354630 483204 354682
rect 483256 354670 483262 354682
rect 520918 354670 520924 354682
rect 483256 354642 520924 354670
rect 483256 354630 483262 354642
rect 520918 354630 520924 354642
rect 520976 354630 520982 354682
rect 480162 354562 480168 354614
rect 480220 354602 480226 354614
rect 516778 354602 516784 354614
rect 480220 354574 516784 354602
rect 480220 354562 480226 354574
rect 516778 354562 516784 354574
rect 516836 354562 516842 354614
rect 477126 354494 477132 354546
rect 477184 354534 477190 354546
rect 496078 354534 496084 354546
rect 477184 354506 496084 354534
rect 477184 354494 477190 354506
rect 496078 354494 496084 354506
rect 496136 354494 496142 354546
rect 486234 353610 486240 353662
rect 486292 353650 486298 353662
rect 486292 353622 489914 353650
rect 486292 353610 486298 353622
rect 489886 353310 489914 353622
rect 525058 353310 525064 353322
rect 489886 353282 525064 353310
rect 525058 353270 525064 353282
rect 525116 353270 525122 353322
rect 547138 344974 547144 345026
rect 547196 345014 547202 345026
rect 547506 345014 547512 345026
rect 547196 344986 547512 345014
rect 547196 344974 547202 344986
rect 547506 344974 547512 344986
rect 547564 344974 547570 345026
rect 470234 342488 470854 342494
rect 470234 342436 470262 342488
rect 470314 342436 470326 342488
rect 470378 342436 470390 342488
rect 470442 342436 470454 342488
rect 470506 342436 470518 342488
rect 470570 342436 470582 342488
rect 470634 342436 470646 342488
rect 470698 342436 470710 342488
rect 470762 342436 470774 342488
rect 470826 342436 470854 342488
rect 470234 342424 470854 342436
rect 470234 342372 470262 342424
rect 470314 342372 470326 342424
rect 470378 342372 470390 342424
rect 470442 342372 470454 342424
rect 470506 342372 470518 342424
rect 470570 342372 470582 342424
rect 470634 342372 470646 342424
rect 470698 342372 470710 342424
rect 470762 342372 470774 342424
rect 470826 342372 470854 342424
rect 470234 342360 470854 342372
rect 470234 342308 470262 342360
rect 470314 342308 470326 342360
rect 470378 342308 470390 342360
rect 470442 342308 470454 342360
rect 470506 342308 470518 342360
rect 470570 342308 470582 342360
rect 470634 342308 470646 342360
rect 470698 342308 470710 342360
rect 470762 342308 470774 342360
rect 470826 342308 470854 342360
rect 470234 342296 470854 342308
rect 470234 342244 470262 342296
rect 470314 342244 470326 342296
rect 470378 342244 470390 342296
rect 470442 342244 470454 342296
rect 470506 342244 470518 342296
rect 470570 342244 470582 342296
rect 470634 342244 470646 342296
rect 470698 342244 470710 342296
rect 470762 342244 470774 342296
rect 470826 342244 470854 342296
rect 470234 342232 470854 342244
rect 470234 342180 470262 342232
rect 470314 342180 470326 342232
rect 470378 342180 470390 342232
rect 470442 342180 470454 342232
rect 470506 342180 470518 342232
rect 470570 342180 470582 342232
rect 470634 342180 470646 342232
rect 470698 342180 470710 342232
rect 470762 342180 470774 342232
rect 470826 342180 470854 342232
rect 470234 342174 470854 342180
rect 471698 341778 471704 341830
rect 471756 341778 471762 341830
rect 471238 341710 471244 341762
rect 471296 341750 471302 341762
rect 471716 341750 471744 341778
rect 471296 341722 471744 341750
rect 471296 341710 471302 341722
rect 471716 341665 471744 341722
rect 468994 341401 469614 341407
rect 468994 341349 469022 341401
rect 469074 341349 469086 341401
rect 469138 341349 469150 341401
rect 469202 341349 469214 341401
rect 469266 341349 469278 341401
rect 469330 341349 469342 341401
rect 469394 341349 469406 341401
rect 469458 341349 469470 341401
rect 469522 341349 469534 341401
rect 469586 341349 469614 341401
rect 468994 341337 469614 341349
rect 468994 341285 469022 341337
rect 469074 341285 469086 341337
rect 469138 341285 469150 341337
rect 469202 341285 469214 341337
rect 469266 341285 469278 341337
rect 469330 341285 469342 341337
rect 469394 341285 469406 341337
rect 469458 341285 469470 341337
rect 469522 341285 469534 341337
rect 469586 341285 469614 341337
rect 468994 341273 469614 341285
rect 468994 341221 469022 341273
rect 469074 341221 469086 341273
rect 469138 341221 469150 341273
rect 469202 341221 469214 341273
rect 469266 341221 469278 341273
rect 469330 341221 469342 341273
rect 469394 341221 469406 341273
rect 469458 341221 469470 341273
rect 469522 341221 469534 341273
rect 469586 341221 469614 341273
rect 468994 341209 469614 341221
rect 468994 341157 469022 341209
rect 469074 341157 469086 341209
rect 469138 341157 469150 341209
rect 469202 341157 469214 341209
rect 469266 341157 469278 341209
rect 469330 341157 469342 341209
rect 469394 341157 469406 341209
rect 469458 341157 469470 341209
rect 469522 341157 469534 341209
rect 469586 341157 469614 341209
rect 468994 341145 469614 341157
rect 468994 341093 469022 341145
rect 469074 341093 469086 341145
rect 469138 341093 469150 341145
rect 469202 341093 469214 341145
rect 469266 341093 469278 341145
rect 469330 341093 469342 341145
rect 469394 341093 469406 341145
rect 469458 341093 469470 341145
rect 469522 341093 469534 341145
rect 469586 341093 469614 341145
rect 468994 341087 469614 341093
rect 484394 340894 484400 340946
rect 484452 340934 484458 340946
rect 484452 340906 484624 340934
rect 484452 340894 484458 340906
rect 482094 340875 482100 340878
rect 482063 340869 482100 340875
rect 474642 340805 474648 340857
rect 474700 340805 474706 340857
rect 482063 340835 482075 340869
rect 482063 340829 482100 340835
rect 482094 340826 482100 340829
rect 482152 340826 482158 340878
rect 484596 340866 484624 340906
rect 484563 340838 484624 340866
rect 484563 340833 484610 340838
rect 484563 340819 484624 340833
rect 484394 340486 484400 340538
rect 484452 340526 484458 340538
rect 484596 340526 484624 340819
rect 484452 340498 484624 340526
rect 484452 340486 484458 340498
rect 485590 340480 485596 340492
rect 485438 340452 485596 340480
rect 485590 340440 485596 340452
rect 485648 340440 485654 340492
rect 475470 340399 475476 340402
rect 475430 340393 475476 340399
rect 475430 340359 475442 340393
rect 475430 340353 475476 340359
rect 475470 340350 475476 340353
rect 475528 340350 475534 340402
rect 478782 340399 478788 340402
rect 478747 340393 478788 340399
rect 478747 340359 478759 340393
rect 478747 340353 478788 340359
rect 478782 340350 478788 340353
rect 478840 340350 478846 340402
rect 488736 340390 488764 340466
rect 492214 340390 492220 340402
rect 488736 340362 492220 340390
rect 492214 340350 492220 340362
rect 492272 340350 492278 340402
rect 470234 340316 470854 340322
rect 470234 340264 470262 340316
rect 470314 340264 470326 340316
rect 470378 340264 470390 340316
rect 470442 340264 470454 340316
rect 470506 340264 470518 340316
rect 470570 340264 470582 340316
rect 470634 340264 470646 340316
rect 470698 340264 470710 340316
rect 470762 340264 470774 340316
rect 470826 340264 470854 340316
rect 470234 340252 470854 340264
rect 470234 340200 470262 340252
rect 470314 340200 470326 340252
rect 470378 340200 470390 340252
rect 470442 340200 470454 340252
rect 470506 340200 470518 340252
rect 470570 340200 470582 340252
rect 470634 340200 470646 340252
rect 470698 340200 470710 340252
rect 470762 340200 470774 340252
rect 470826 340200 470854 340252
rect 470234 340188 470854 340200
rect 470234 340136 470262 340188
rect 470314 340136 470326 340188
rect 470378 340136 470390 340188
rect 470442 340136 470454 340188
rect 470506 340136 470518 340188
rect 470570 340136 470582 340188
rect 470634 340136 470646 340188
rect 470698 340136 470710 340188
rect 470762 340136 470774 340188
rect 470826 340136 470854 340188
rect 470234 340124 470854 340136
rect 470234 340072 470262 340124
rect 470314 340072 470326 340124
rect 470378 340072 470390 340124
rect 470442 340072 470454 340124
rect 470506 340072 470518 340124
rect 470570 340072 470582 340124
rect 470634 340072 470646 340124
rect 470698 340072 470710 340124
rect 470762 340072 470774 340124
rect 470826 340072 470854 340124
rect 470234 340060 470854 340072
rect 470234 340008 470262 340060
rect 470314 340008 470326 340060
rect 470378 340008 470390 340060
rect 470442 340008 470454 340060
rect 470506 340008 470518 340060
rect 470570 340008 470582 340060
rect 470634 340008 470646 340060
rect 470698 340008 470710 340060
rect 470762 340008 470774 340060
rect 470826 340008 470854 340060
rect 470234 340002 470854 340008
rect 475470 339398 475476 339450
rect 475528 339398 475534 339450
rect 478782 339398 478788 339450
rect 478840 339438 478846 339450
rect 536374 339438 536380 339450
rect 478840 339410 536380 339438
rect 478840 339398 478846 339410
rect 536374 339398 536380 339410
rect 536432 339398 536438 339450
rect 475488 339302 475516 339398
rect 482094 339330 482100 339382
rect 482152 339370 482158 339382
rect 515398 339370 515404 339382
rect 482152 339342 515404 339370
rect 482152 339330 482158 339342
rect 515398 339330 515404 339342
rect 515456 339330 515462 339382
rect 497458 339302 497464 339314
rect 475488 339274 497464 339302
rect 497458 339262 497464 339274
rect 497516 339262 497522 339314
rect 523678 338038 523684 338090
rect 523736 338078 523742 338090
rect 535454 338078 535460 338090
rect 523736 338050 535460 338078
rect 523736 338038 523742 338050
rect 535454 338038 535460 338050
rect 535512 338038 535518 338090
rect 546954 337698 546960 337750
rect 547012 337738 547018 337750
rect 547506 337738 547512 337750
rect 547012 337710 547512 337738
rect 547012 337698 547018 337710
rect 547506 337698 547512 337710
rect 547564 337698 547570 337750
rect 525058 332530 525064 332582
rect 525116 332570 525122 332582
rect 535454 332570 535460 332582
rect 525116 332542 535460 332570
rect 525116 332530 525122 332542
rect 535454 332530 535460 332542
rect 535512 332530 535518 332582
rect 485682 331170 485688 331222
rect 485740 331210 485746 331222
rect 535454 331210 535460 331222
rect 485740 331182 535460 331210
rect 485740 331170 485746 331182
rect 535454 331170 535460 331182
rect 535512 331170 535518 331222
rect 576994 325952 577614 325958
rect 576994 325900 577022 325952
rect 577074 325900 577086 325952
rect 577138 325900 577150 325952
rect 577202 325900 577214 325952
rect 577266 325900 577278 325952
rect 577330 325900 577342 325952
rect 577394 325900 577406 325952
rect 577458 325900 577470 325952
rect 577522 325900 577534 325952
rect 577586 325900 577614 325952
rect 576994 325888 577614 325900
rect 576994 325836 577022 325888
rect 577074 325836 577086 325888
rect 577138 325836 577150 325888
rect 577202 325836 577214 325888
rect 577266 325836 577278 325888
rect 577330 325836 577342 325888
rect 577394 325836 577406 325888
rect 577458 325836 577470 325888
rect 577522 325836 577534 325888
rect 577586 325836 577614 325888
rect 576994 325824 577614 325836
rect 576994 325772 577022 325824
rect 577074 325772 577086 325824
rect 577138 325772 577150 325824
rect 577202 325772 577214 325824
rect 577266 325772 577278 325824
rect 577330 325772 577342 325824
rect 577394 325772 577406 325824
rect 577458 325772 577470 325824
rect 577522 325772 577534 325824
rect 577586 325772 577614 325824
rect 576994 325760 577614 325772
rect 576994 325734 577022 325760
rect 523678 325662 523684 325714
rect 523736 325702 523742 325714
rect 535454 325702 535460 325714
rect 523736 325674 535460 325702
rect 523736 325662 523742 325674
rect 535454 325662 535460 325674
rect 535512 325662 535518 325714
rect 576400 325708 577022 325734
rect 577074 325708 577086 325760
rect 577138 325708 577150 325760
rect 577202 325708 577214 325760
rect 577266 325708 577278 325760
rect 577330 325708 577342 325760
rect 577394 325708 577406 325760
rect 577458 325708 577470 325760
rect 577522 325708 577534 325760
rect 577586 325734 577614 325760
rect 577586 325708 577647 325734
rect 576400 325703 577647 325708
rect 576316 325696 577647 325703
rect 576316 325669 577022 325696
rect 576400 325644 577022 325669
rect 577074 325644 577086 325696
rect 577138 325644 577150 325696
rect 577202 325644 577214 325696
rect 577266 325644 577278 325696
rect 577330 325644 577342 325696
rect 577394 325644 577406 325696
rect 577458 325644 577470 325696
rect 577522 325644 577534 325696
rect 577586 325644 577647 325696
rect 576400 325638 577647 325644
rect 576597 325218 576603 325270
rect 576655 325218 576661 325270
rect 576400 325157 578876 325190
rect 576400 325105 578262 325157
rect 578314 325105 578326 325157
rect 578378 325105 578390 325157
rect 578442 325105 578454 325157
rect 578506 325105 578518 325157
rect 578570 325105 578582 325157
rect 578634 325105 578646 325157
rect 578698 325105 578710 325157
rect 578762 325105 578774 325157
rect 578826 325105 578876 325157
rect 576400 325094 578876 325105
rect 578234 325093 578854 325094
rect 578234 325041 578262 325093
rect 578314 325041 578326 325093
rect 578378 325041 578390 325093
rect 578442 325041 578454 325093
rect 578506 325041 578518 325093
rect 578570 325041 578582 325093
rect 578634 325041 578646 325093
rect 578698 325041 578710 325093
rect 578762 325041 578774 325093
rect 578826 325041 578854 325093
rect 578234 325029 578854 325041
rect 578234 324977 578262 325029
rect 578314 324977 578326 325029
rect 578378 324977 578390 325029
rect 578442 324977 578454 325029
rect 578506 324977 578518 325029
rect 578570 324977 578582 325029
rect 578634 324977 578646 325029
rect 578698 324977 578710 325029
rect 578762 324977 578774 325029
rect 578826 324977 578854 325029
rect 578234 324965 578854 324977
rect 578234 324913 578262 324965
rect 578314 324913 578326 324965
rect 578378 324913 578390 324965
rect 578442 324913 578454 324965
rect 578506 324913 578518 324965
rect 578570 324913 578582 324965
rect 578634 324913 578646 324965
rect 578698 324913 578710 324965
rect 578762 324913 578774 324965
rect 578826 324913 578854 324965
rect 578234 324901 578854 324913
rect 578234 324849 578262 324901
rect 578314 324849 578326 324901
rect 578378 324849 578390 324901
rect 578442 324849 578454 324901
rect 578506 324849 578518 324901
rect 578570 324849 578582 324901
rect 578634 324849 578646 324901
rect 578698 324849 578710 324901
rect 578762 324849 578774 324901
rect 578826 324849 578854 324901
rect 578234 324843 578854 324849
rect 470234 322488 470854 322494
rect 470234 322436 470262 322488
rect 470314 322436 470326 322488
rect 470378 322436 470390 322488
rect 470442 322436 470454 322488
rect 470506 322436 470518 322488
rect 470570 322436 470582 322488
rect 470634 322436 470646 322488
rect 470698 322436 470710 322488
rect 470762 322436 470774 322488
rect 470826 322436 470854 322488
rect 470234 322424 470854 322436
rect 470234 322372 470262 322424
rect 470314 322372 470326 322424
rect 470378 322372 470390 322424
rect 470442 322372 470454 322424
rect 470506 322372 470518 322424
rect 470570 322372 470582 322424
rect 470634 322372 470646 322424
rect 470698 322372 470710 322424
rect 470762 322372 470774 322424
rect 470826 322372 470854 322424
rect 470234 322360 470854 322372
rect 470234 322308 470262 322360
rect 470314 322308 470326 322360
rect 470378 322308 470390 322360
rect 470442 322308 470454 322360
rect 470506 322308 470518 322360
rect 470570 322308 470582 322360
rect 470634 322308 470646 322360
rect 470698 322308 470710 322360
rect 470762 322308 470774 322360
rect 470826 322308 470854 322360
rect 470234 322296 470854 322308
rect 470234 322244 470262 322296
rect 470314 322244 470326 322296
rect 470378 322244 470390 322296
rect 470442 322244 470454 322296
rect 470506 322244 470518 322296
rect 470570 322244 470582 322296
rect 470634 322244 470646 322296
rect 470698 322244 470710 322296
rect 470762 322244 470774 322296
rect 470826 322244 470854 322296
rect 470234 322232 470854 322244
rect 470234 322180 470262 322232
rect 470314 322180 470326 322232
rect 470378 322180 470390 322232
rect 470442 322180 470454 322232
rect 470506 322180 470518 322232
rect 470570 322180 470582 322232
rect 470634 322180 470646 322232
rect 470698 322180 470710 322232
rect 470762 322180 470774 322232
rect 470826 322180 470854 322232
rect 470234 322174 470854 322180
rect 471238 321582 471244 321634
rect 471296 321622 471302 321634
rect 471624 321622 471652 321665
rect 471296 321594 471652 321622
rect 471296 321582 471302 321594
rect 468994 321401 469614 321407
rect 468994 321349 469022 321401
rect 469074 321349 469086 321401
rect 469138 321349 469150 321401
rect 469202 321349 469214 321401
rect 469266 321349 469278 321401
rect 469330 321349 469342 321401
rect 469394 321349 469406 321401
rect 469458 321349 469470 321401
rect 469522 321349 469534 321401
rect 469586 321349 469614 321401
rect 468994 321337 469614 321349
rect 468994 321285 469022 321337
rect 469074 321285 469086 321337
rect 469138 321285 469150 321337
rect 469202 321285 469214 321337
rect 469266 321285 469278 321337
rect 469330 321285 469342 321337
rect 469394 321285 469406 321337
rect 469458 321285 469470 321337
rect 469522 321285 469534 321337
rect 469586 321285 469614 321337
rect 468994 321273 469614 321285
rect 468994 321221 469022 321273
rect 469074 321221 469086 321273
rect 469138 321221 469150 321273
rect 469202 321221 469214 321273
rect 469266 321221 469278 321273
rect 469330 321221 469342 321273
rect 469394 321221 469406 321273
rect 469458 321221 469470 321273
rect 469522 321221 469534 321273
rect 469586 321221 469614 321273
rect 468994 321209 469614 321221
rect 468994 321157 469022 321209
rect 469074 321157 469086 321209
rect 469138 321157 469150 321209
rect 469202 321157 469214 321209
rect 469266 321157 469278 321209
rect 469330 321157 469342 321209
rect 469394 321157 469406 321209
rect 469458 321157 469470 321209
rect 469522 321157 469534 321209
rect 469586 321157 469614 321209
rect 468994 321145 469614 321157
rect 468994 321093 469022 321145
rect 469074 321093 469086 321145
rect 469138 321093 469150 321145
rect 469202 321093 469214 321145
rect 469266 321093 469278 321145
rect 469330 321093 469342 321145
rect 469394 321093 469406 321145
rect 469458 321093 469470 321145
rect 469522 321093 469534 321145
rect 469586 321093 469614 321145
rect 468994 321087 469614 321093
rect 475470 320437 475476 320489
rect 475528 320437 475534 320489
rect 482370 320426 482376 320478
rect 482428 320426 482434 320478
rect 478927 320401 478985 320407
rect 478927 320367 478939 320401
rect 478973 320398 478985 320401
rect 479058 320398 479064 320410
rect 478973 320370 479064 320398
rect 478973 320367 478985 320370
rect 478927 320361 478985 320367
rect 479058 320358 479064 320370
rect 479116 320358 479122 320410
rect 485815 320401 485873 320407
rect 485815 320367 485827 320401
rect 485861 320398 485873 320401
rect 485958 320398 485964 320410
rect 485861 320370 485964 320398
rect 485861 320367 485873 320370
rect 485815 320361 485873 320367
rect 485958 320358 485964 320370
rect 486016 320358 486022 320410
rect 489288 320398 489316 320463
rect 492306 320398 492312 320410
rect 489288 320370 492312 320398
rect 492306 320358 492312 320370
rect 492364 320358 492370 320410
rect 470234 320316 470854 320322
rect 470234 320264 470262 320316
rect 470314 320264 470326 320316
rect 470378 320264 470390 320316
rect 470442 320264 470454 320316
rect 470506 320264 470518 320316
rect 470570 320264 470582 320316
rect 470634 320264 470646 320316
rect 470698 320264 470710 320316
rect 470762 320264 470774 320316
rect 470826 320264 470854 320316
rect 470234 320252 470854 320264
rect 470234 320200 470262 320252
rect 470314 320200 470326 320252
rect 470378 320200 470390 320252
rect 470442 320200 470454 320252
rect 470506 320200 470518 320252
rect 470570 320200 470582 320252
rect 470634 320200 470646 320252
rect 470698 320200 470710 320252
rect 470762 320200 470774 320252
rect 470826 320200 470854 320252
rect 470234 320188 470854 320200
rect 470234 320136 470262 320188
rect 470314 320136 470326 320188
rect 470378 320136 470390 320188
rect 470442 320136 470454 320188
rect 470506 320136 470518 320188
rect 470570 320136 470582 320188
rect 470634 320136 470646 320188
rect 470698 320136 470710 320188
rect 470762 320136 470774 320188
rect 470826 320136 470854 320188
rect 470234 320124 470854 320136
rect 470234 320072 470262 320124
rect 470314 320072 470326 320124
rect 470378 320072 470390 320124
rect 470442 320072 470454 320124
rect 470506 320072 470518 320124
rect 470570 320072 470582 320124
rect 470634 320072 470646 320124
rect 470698 320072 470710 320124
rect 470762 320072 470774 320124
rect 470826 320072 470854 320124
rect 470234 320060 470854 320072
rect 470234 320008 470262 320060
rect 470314 320008 470326 320060
rect 470378 320008 470390 320060
rect 470442 320008 470454 320060
rect 470506 320008 470518 320060
rect 470570 320008 470582 320060
rect 470634 320008 470646 320060
rect 470698 320008 470710 320060
rect 470762 320008 470774 320060
rect 470826 320008 470854 320060
rect 470234 320002 470854 320008
rect 475470 318726 475476 318778
rect 475528 318726 475534 318778
rect 479058 318726 479064 318778
rect 479116 318766 479122 318778
rect 536282 318766 536288 318778
rect 479116 318738 536288 318766
rect 479116 318726 479122 318738
rect 536282 318726 536288 318738
rect 536340 318726 536346 318778
rect 475488 318562 475516 318726
rect 482370 318658 482376 318710
rect 482428 318698 482434 318710
rect 536558 318698 536564 318710
rect 482428 318670 536564 318698
rect 482428 318658 482434 318670
rect 536558 318658 536564 318670
rect 536616 318658 536622 318710
rect 485958 318590 485964 318642
rect 486016 318630 486022 318642
rect 536006 318630 536012 318642
rect 486016 318602 536012 318630
rect 486016 318590 486022 318602
rect 536006 318590 536012 318602
rect 536064 318590 536070 318642
rect 498838 318562 498844 318574
rect 475488 318534 498844 318562
rect 498838 318522 498844 318534
rect 498896 318522 498902 318574
rect 470234 307088 470854 307094
rect 470234 307036 470262 307088
rect 470314 307036 470326 307088
rect 470378 307036 470390 307088
rect 470442 307036 470454 307088
rect 470506 307036 470518 307088
rect 470570 307036 470582 307088
rect 470634 307036 470646 307088
rect 470698 307036 470710 307088
rect 470762 307036 470774 307088
rect 470826 307036 470854 307088
rect 470234 307024 470854 307036
rect 470234 306972 470262 307024
rect 470314 306972 470326 307024
rect 470378 306972 470390 307024
rect 470442 306972 470454 307024
rect 470506 306972 470518 307024
rect 470570 306972 470582 307024
rect 470634 306972 470646 307024
rect 470698 306972 470710 307024
rect 470762 306972 470774 307024
rect 470826 306972 470854 307024
rect 470234 306960 470854 306972
rect 470234 306908 470262 306960
rect 470314 306908 470326 306960
rect 470378 306908 470390 306960
rect 470442 306908 470454 306960
rect 470506 306908 470518 306960
rect 470570 306908 470582 306960
rect 470634 306908 470646 306960
rect 470698 306908 470710 306960
rect 470762 306908 470774 306960
rect 470826 306908 470854 306960
rect 470234 306896 470854 306908
rect 470234 306844 470262 306896
rect 470314 306844 470326 306896
rect 470378 306844 470390 306896
rect 470442 306844 470454 306896
rect 470506 306844 470518 306896
rect 470570 306844 470582 306896
rect 470634 306844 470646 306896
rect 470698 306844 470710 306896
rect 470762 306844 470774 306896
rect 470826 306844 470854 306896
rect 470234 306832 470854 306844
rect 470234 306780 470262 306832
rect 470314 306780 470326 306832
rect 470378 306780 470390 306832
rect 470442 306780 470454 306832
rect 470506 306780 470518 306832
rect 470570 306780 470582 306832
rect 470634 306780 470646 306832
rect 470698 306780 470710 306832
rect 470762 306780 470774 306832
rect 470826 306780 470854 306832
rect 470234 306774 470854 306780
rect 471238 306282 471244 306334
rect 471296 306322 471302 306334
rect 471296 306294 471652 306322
rect 471296 306282 471302 306294
rect 471624 306266 471652 306294
rect 473722 306234 473728 306286
rect 473780 306234 473786 306286
rect 468994 306003 469614 306009
rect 468994 305951 469022 306003
rect 469074 305951 469086 306003
rect 469138 305951 469150 306003
rect 469202 305951 469214 306003
rect 469266 305951 469278 306003
rect 469330 305951 469342 306003
rect 469394 305951 469406 306003
rect 469458 305951 469470 306003
rect 469522 305951 469534 306003
rect 469586 305951 469614 306003
rect 468994 305939 469614 305951
rect 468994 305887 469022 305939
rect 469074 305887 469086 305939
rect 469138 305887 469150 305939
rect 469202 305887 469214 305939
rect 469266 305887 469278 305939
rect 469330 305887 469342 305939
rect 469394 305887 469406 305939
rect 469458 305887 469470 305939
rect 469522 305887 469534 305939
rect 469586 305887 469614 305939
rect 468994 305875 469614 305887
rect 468994 305823 469022 305875
rect 469074 305823 469086 305875
rect 469138 305823 469150 305875
rect 469202 305823 469214 305875
rect 469266 305823 469278 305875
rect 469330 305823 469342 305875
rect 469394 305823 469406 305875
rect 469458 305823 469470 305875
rect 469522 305823 469534 305875
rect 469586 305823 469614 305875
rect 468994 305811 469614 305823
rect 468994 305759 469022 305811
rect 469074 305759 469086 305811
rect 469138 305759 469150 305811
rect 469202 305759 469214 305811
rect 469266 305759 469278 305811
rect 469330 305759 469342 305811
rect 469394 305759 469406 305811
rect 469458 305759 469470 305811
rect 469522 305759 469534 305811
rect 469586 305759 469614 305811
rect 468994 305747 469614 305759
rect 468994 305695 469022 305747
rect 469074 305695 469086 305747
rect 469138 305695 469150 305747
rect 469202 305695 469214 305747
rect 469266 305695 469278 305747
rect 469330 305695 469342 305747
rect 469394 305695 469406 305747
rect 469458 305695 469470 305747
rect 469522 305695 469534 305747
rect 469586 305695 469614 305747
rect 468994 305689 469614 305695
rect 478598 305447 478604 305450
rect 478568 305441 478604 305447
rect 478568 305407 478580 305441
rect 478568 305401 478604 305407
rect 478598 305398 478604 305401
rect 478656 305398 478662 305450
rect 485130 305447 485136 305450
rect 485098 305441 485136 305447
rect 485098 305407 485110 305441
rect 485098 305401 485136 305407
rect 485130 305398 485136 305401
rect 485188 305398 485194 305450
rect 475286 305038 475292 305090
rect 475344 305038 475350 305090
rect 481818 305038 481824 305090
rect 481876 305038 481882 305090
rect 488382 305050 488672 305078
rect 488644 305030 488672 305050
rect 490558 305030 490564 305042
rect 488644 305002 490564 305030
rect 490558 304990 490564 305002
rect 490616 304990 490622 305042
rect 470234 304916 470854 304922
rect 470234 304864 470262 304916
rect 470314 304864 470326 304916
rect 470378 304864 470390 304916
rect 470442 304864 470454 304916
rect 470506 304864 470518 304916
rect 470570 304864 470582 304916
rect 470634 304864 470646 304916
rect 470698 304864 470710 304916
rect 470762 304864 470774 304916
rect 470826 304864 470854 304916
rect 470234 304852 470854 304864
rect 470234 304800 470262 304852
rect 470314 304800 470326 304852
rect 470378 304800 470390 304852
rect 470442 304800 470454 304852
rect 470506 304800 470518 304852
rect 470570 304800 470582 304852
rect 470634 304800 470646 304852
rect 470698 304800 470710 304852
rect 470762 304800 470774 304852
rect 470826 304800 470854 304852
rect 470234 304788 470854 304800
rect 470234 304736 470262 304788
rect 470314 304736 470326 304788
rect 470378 304736 470390 304788
rect 470442 304736 470454 304788
rect 470506 304736 470518 304788
rect 470570 304736 470582 304788
rect 470634 304736 470646 304788
rect 470698 304736 470710 304788
rect 470762 304736 470774 304788
rect 470826 304736 470854 304788
rect 470234 304724 470854 304736
rect 470234 304672 470262 304724
rect 470314 304672 470326 304724
rect 470378 304672 470390 304724
rect 470442 304672 470454 304724
rect 470506 304672 470518 304724
rect 470570 304672 470582 304724
rect 470634 304672 470646 304724
rect 470698 304672 470710 304724
rect 470762 304672 470774 304724
rect 470826 304672 470854 304724
rect 470234 304660 470854 304672
rect 470234 304608 470262 304660
rect 470314 304608 470326 304660
rect 470378 304608 470390 304660
rect 470442 304608 470454 304660
rect 470506 304608 470518 304660
rect 470570 304608 470582 304660
rect 470634 304608 470646 304660
rect 470698 304608 470710 304660
rect 470762 304608 470774 304660
rect 470826 304608 470854 304660
rect 470234 304602 470854 304608
rect 547046 303698 547052 303750
rect 547104 303738 547110 303750
rect 547506 303738 547512 303750
rect 547104 303710 547512 303738
rect 547104 303698 547110 303710
rect 547506 303698 547512 303710
rect 547564 303698 547570 303750
rect 485056 303642 485268 303670
rect 475286 303562 475292 303614
rect 475344 303562 475350 303614
rect 478598 303562 478604 303614
rect 478656 303602 478662 303614
rect 478656 303574 480254 303602
rect 478656 303562 478662 303574
rect 475304 303398 475332 303562
rect 480226 303466 480254 303574
rect 481818 303562 481824 303614
rect 481876 303602 481882 303614
rect 485056 303602 485084 303642
rect 481876 303574 485084 303602
rect 481876 303562 481882 303574
rect 485130 303562 485136 303614
rect 485188 303562 485194 303614
rect 485240 303602 485268 303642
rect 536466 303602 536472 303614
rect 485240 303574 536472 303602
rect 536466 303562 536472 303574
rect 536524 303562 536530 303614
rect 485148 303534 485176 303562
rect 536650 303534 536656 303546
rect 485148 303506 536656 303534
rect 536650 303494 536656 303506
rect 536708 303494 536714 303546
rect 518158 303466 518164 303478
rect 480226 303438 518164 303466
rect 518158 303426 518164 303438
rect 518216 303426 518222 303478
rect 500218 303398 500224 303410
rect 475304 303370 500224 303398
rect 500218 303358 500224 303370
rect 500276 303358 500282 303410
rect 491938 300774 491944 300826
rect 491996 300814 492002 300826
rect 535454 300814 535460 300826
rect 491996 300786 535460 300814
rect 491996 300774 492002 300786
rect 535454 300774 535460 300786
rect 535512 300774 535518 300826
rect 492030 299414 492036 299466
rect 492088 299454 492094 299466
rect 535454 299454 535460 299466
rect 492088 299426 535460 299454
rect 492088 299414 492094 299426
rect 535454 299414 535460 299426
rect 535512 299414 535518 299466
rect 490742 298054 490748 298106
rect 490800 298094 490806 298106
rect 535454 298094 535460 298106
rect 490800 298066 535460 298094
rect 490800 298054 490806 298066
rect 535454 298054 535460 298066
rect 535512 298054 535518 298106
rect 492122 296626 492128 296678
rect 492180 296666 492186 296678
rect 535546 296666 535552 296678
rect 492180 296638 535552 296666
rect 492180 296626 492186 296638
rect 535546 296626 535552 296638
rect 535604 296626 535610 296678
rect 493318 296558 493324 296610
rect 493376 296598 493382 296610
rect 535454 296598 535460 296610
rect 493376 296570 535460 296598
rect 493376 296558 493382 296570
rect 535454 296558 535460 296570
rect 535512 296558 535518 296610
rect 492214 295266 492220 295318
rect 492272 295306 492278 295318
rect 535454 295306 535460 295318
rect 492272 295278 535460 295306
rect 492272 295266 492278 295278
rect 535454 295266 535460 295278
rect 535512 295266 535518 295318
rect 492306 293906 492312 293958
rect 492364 293946 492370 293958
rect 535546 293946 535552 293958
rect 492364 293918 535552 293946
rect 492364 293906 492370 293918
rect 535546 293906 535552 293918
rect 535604 293906 535610 293958
rect 490558 292478 490564 292530
rect 490616 292518 490622 292530
rect 535454 292518 535460 292530
rect 490616 292490 535460 292518
rect 490616 292478 490622 292490
rect 535454 292478 535460 292490
rect 535512 292478 535518 292530
rect 492950 289826 492956 289878
rect 493008 289866 493014 289878
rect 535454 289866 535460 289878
rect 493008 289838 535460 289866
rect 493008 289826 493014 289838
rect 535454 289826 535460 289838
rect 535512 289826 535518 289878
rect 491938 288398 491944 288450
rect 491996 288438 492002 288450
rect 535454 288438 535460 288450
rect 491996 288410 535460 288438
rect 491996 288398 492002 288410
rect 535454 288398 535460 288410
rect 535512 288398 535518 288450
rect 470234 287489 470854 287495
rect 470234 287437 470262 287489
rect 470314 287437 470326 287489
rect 470378 287437 470390 287489
rect 470442 287437 470454 287489
rect 470506 287437 470518 287489
rect 470570 287437 470582 287489
rect 470634 287437 470646 287489
rect 470698 287437 470710 287489
rect 470762 287437 470774 287489
rect 470826 287437 470854 287489
rect 470234 287425 470854 287437
rect 470234 287373 470262 287425
rect 470314 287373 470326 287425
rect 470378 287373 470390 287425
rect 470442 287373 470454 287425
rect 470506 287373 470518 287425
rect 470570 287373 470582 287425
rect 470634 287373 470646 287425
rect 470698 287373 470710 287425
rect 470762 287373 470774 287425
rect 470826 287373 470854 287425
rect 470234 287361 470854 287373
rect 470234 287309 470262 287361
rect 470314 287309 470326 287361
rect 470378 287309 470390 287361
rect 470442 287309 470454 287361
rect 470506 287309 470518 287361
rect 470570 287309 470582 287361
rect 470634 287309 470646 287361
rect 470698 287309 470710 287361
rect 470762 287309 470774 287361
rect 470826 287309 470854 287361
rect 470234 287297 470854 287309
rect 470234 287245 470262 287297
rect 470314 287245 470326 287297
rect 470378 287245 470390 287297
rect 470442 287245 470454 287297
rect 470506 287245 470518 287297
rect 470570 287245 470582 287297
rect 470634 287245 470646 287297
rect 470698 287245 470710 287297
rect 470762 287245 470774 287297
rect 470826 287245 470854 287297
rect 470234 287233 470854 287245
rect 470234 287181 470262 287233
rect 470314 287181 470326 287233
rect 470378 287181 470390 287233
rect 470442 287181 470454 287233
rect 470506 287181 470518 287233
rect 470570 287181 470582 287233
rect 470634 287181 470646 287233
rect 470698 287181 470710 287233
rect 470762 287181 470774 287233
rect 470826 287181 470854 287233
rect 470234 287175 470854 287181
rect 488632 286682 488684 286688
rect 471238 286630 471244 286682
rect 471296 286670 471302 286682
rect 471296 286642 471652 286670
rect 471296 286630 471302 286642
rect 471624 286534 471652 286642
rect 484946 286630 484952 286682
rect 485004 286630 485010 286682
rect 488632 286624 488684 286630
rect 471698 286534 471704 286546
rect 471624 286506 471704 286534
rect 471698 286494 471704 286506
rect 471756 286494 471762 286546
rect 468994 286404 469614 286410
rect 468994 286352 469022 286404
rect 469074 286352 469086 286404
rect 469138 286352 469150 286404
rect 469202 286352 469214 286404
rect 469266 286352 469278 286404
rect 469330 286352 469342 286404
rect 469394 286352 469406 286404
rect 469458 286352 469470 286404
rect 469522 286352 469534 286404
rect 469586 286352 469614 286404
rect 468994 286340 469614 286352
rect 468994 286288 469022 286340
rect 469074 286288 469086 286340
rect 469138 286288 469150 286340
rect 469202 286288 469214 286340
rect 469266 286288 469278 286340
rect 469330 286288 469342 286340
rect 469394 286288 469406 286340
rect 469458 286288 469470 286340
rect 469522 286288 469534 286340
rect 469586 286288 469614 286340
rect 468994 286276 469614 286288
rect 468994 286224 469022 286276
rect 469074 286224 469086 286276
rect 469138 286224 469150 286276
rect 469202 286224 469214 286276
rect 469266 286224 469278 286276
rect 469330 286224 469342 286276
rect 469394 286224 469406 286276
rect 469458 286224 469470 286276
rect 469522 286224 469534 286276
rect 469586 286224 469614 286276
rect 468994 286212 469614 286224
rect 468994 286160 469022 286212
rect 469074 286160 469086 286212
rect 469138 286160 469150 286212
rect 469202 286160 469214 286212
rect 469266 286160 469278 286212
rect 469330 286160 469342 286212
rect 469394 286160 469406 286212
rect 469458 286160 469470 286212
rect 469522 286160 469534 286212
rect 469586 286160 469614 286212
rect 468994 286148 469614 286160
rect 468994 286096 469022 286148
rect 469074 286096 469086 286148
rect 469138 286096 469150 286148
rect 469202 286096 469214 286148
rect 469266 286096 469278 286148
rect 469330 286096 469342 286148
rect 469394 286096 469406 286148
rect 469458 286096 469470 286148
rect 469522 286096 469534 286148
rect 469586 286096 469614 286148
rect 468994 286090 469614 286096
rect 490598 285993 490656 285999
rect 490598 285959 490610 285993
rect 490644 285990 490656 285993
rect 490644 285962 490880 285990
rect 490644 285959 490656 285962
rect 490598 285953 490656 285959
rect 479426 285814 479432 285866
rect 479484 285863 479490 285866
rect 479484 285857 479520 285863
rect 479508 285823 479520 285857
rect 479484 285817 479520 285823
rect 479484 285814 479490 285817
rect 490852 285650 490880 285962
rect 492950 285650 492956 285662
rect 490852 285622 492956 285650
rect 492950 285610 492956 285622
rect 493008 285610 493014 285662
rect 475746 285438 475752 285490
rect 475804 285438 475810 285490
rect 483198 285438 483204 285490
rect 483256 285438 483262 285490
rect 486878 285438 486884 285490
rect 486936 285438 486942 285490
rect 470234 285316 470854 285322
rect 470234 285264 470262 285316
rect 470314 285264 470326 285316
rect 470378 285264 470390 285316
rect 470442 285264 470454 285316
rect 470506 285264 470518 285316
rect 470570 285264 470582 285316
rect 470634 285264 470646 285316
rect 470698 285264 470710 285316
rect 470762 285264 470774 285316
rect 470826 285264 470854 285316
rect 470234 285252 470854 285264
rect 470234 285200 470262 285252
rect 470314 285200 470326 285252
rect 470378 285200 470390 285252
rect 470442 285200 470454 285252
rect 470506 285200 470518 285252
rect 470570 285200 470582 285252
rect 470634 285200 470646 285252
rect 470698 285200 470710 285252
rect 470762 285200 470774 285252
rect 470826 285200 470854 285252
rect 470234 285188 470854 285200
rect 470234 285136 470262 285188
rect 470314 285136 470326 285188
rect 470378 285136 470390 285188
rect 470442 285136 470454 285188
rect 470506 285136 470518 285188
rect 470570 285136 470582 285188
rect 470634 285136 470646 285188
rect 470698 285136 470710 285188
rect 470762 285136 470774 285188
rect 470826 285136 470854 285188
rect 470234 285124 470854 285136
rect 470234 285072 470262 285124
rect 470314 285072 470326 285124
rect 470378 285072 470390 285124
rect 470442 285072 470454 285124
rect 470506 285072 470518 285124
rect 470570 285072 470582 285124
rect 470634 285072 470646 285124
rect 470698 285072 470710 285124
rect 470762 285072 470774 285124
rect 470826 285072 470854 285124
rect 470234 285060 470854 285072
rect 470234 285008 470262 285060
rect 470314 285008 470326 285060
rect 470378 285008 470390 285060
rect 470442 285008 470454 285060
rect 470506 285008 470518 285060
rect 470570 285008 470582 285060
rect 470634 285008 470646 285060
rect 470698 285008 470710 285060
rect 470762 285008 470774 285060
rect 470826 285008 470854 285060
rect 470234 285002 470854 285008
rect 475746 284250 475752 284302
rect 475804 284250 475810 284302
rect 479426 284250 479432 284302
rect 479484 284290 479490 284302
rect 536098 284290 536104 284302
rect 479484 284262 536104 284290
rect 479484 284250 479490 284262
rect 536098 284250 536104 284262
rect 536156 284250 536162 284302
rect 475764 284086 475792 284250
rect 483198 284182 483204 284234
rect 483256 284182 483262 284234
rect 522298 284222 522304 284234
rect 485746 284194 522304 284222
rect 483216 284154 483244 284182
rect 485746 284154 485774 284194
rect 522298 284182 522304 284194
rect 522356 284182 522362 284234
rect 483216 284126 485774 284154
rect 486878 284114 486884 284166
rect 486936 284154 486942 284166
rect 523678 284154 523684 284166
rect 486936 284126 523684 284154
rect 486936 284114 486942 284126
rect 523678 284114 523684 284126
rect 523736 284114 523742 284166
rect 501598 284086 501604 284098
rect 475764 284058 501604 284086
rect 501598 284046 501604 284058
rect 501656 284046 501662 284098
rect 576994 272912 577614 272918
rect 576994 272860 577022 272912
rect 577074 272860 577086 272912
rect 577138 272860 577150 272912
rect 577202 272860 577214 272912
rect 577266 272860 577278 272912
rect 577330 272860 577342 272912
rect 577394 272860 577406 272912
rect 577458 272860 577470 272912
rect 577522 272860 577534 272912
rect 577586 272860 577614 272912
rect 576994 272848 577614 272860
rect 576994 272796 577022 272848
rect 577074 272796 577086 272848
rect 577138 272796 577150 272848
rect 577202 272796 577214 272848
rect 577266 272796 577278 272848
rect 577330 272796 577342 272848
rect 577394 272796 577406 272848
rect 577458 272796 577470 272848
rect 577522 272796 577534 272848
rect 577586 272796 577614 272848
rect 576994 272784 577614 272796
rect 576994 272732 577022 272784
rect 577074 272732 577086 272784
rect 577138 272732 577150 272784
rect 577202 272732 577214 272784
rect 577266 272732 577278 272784
rect 577330 272732 577342 272784
rect 577394 272732 577406 272784
rect 577458 272732 577470 272784
rect 577522 272732 577534 272784
rect 577586 272732 577614 272784
rect 576994 272720 577614 272732
rect 576994 272694 577022 272720
rect 576400 272668 577022 272694
rect 577074 272668 577086 272720
rect 577138 272668 577150 272720
rect 577202 272668 577214 272720
rect 577266 272668 577278 272720
rect 577330 272668 577342 272720
rect 577394 272668 577406 272720
rect 577458 272668 577470 272720
rect 577522 272668 577534 272720
rect 577586 272694 577614 272720
rect 577586 272668 577647 272694
rect 576400 272663 577647 272668
rect 576316 272656 577647 272663
rect 576316 272629 577022 272656
rect 576400 272604 577022 272629
rect 577074 272604 577086 272656
rect 577138 272604 577150 272656
rect 577202 272604 577214 272656
rect 577266 272604 577278 272656
rect 577330 272604 577342 272656
rect 577394 272604 577406 272656
rect 577458 272604 577470 272656
rect 577522 272604 577534 272656
rect 577586 272604 577647 272656
rect 576400 272598 577647 272604
rect 576597 272178 576603 272230
rect 576655 272178 576661 272230
rect 576400 272117 578876 272150
rect 576400 272065 578262 272117
rect 578314 272065 578326 272117
rect 578378 272065 578390 272117
rect 578442 272065 578454 272117
rect 578506 272065 578518 272117
rect 578570 272065 578582 272117
rect 578634 272065 578646 272117
rect 578698 272065 578710 272117
rect 578762 272065 578774 272117
rect 578826 272065 578876 272117
rect 576400 272054 578876 272065
rect 578234 272053 578854 272054
rect 578234 272001 578262 272053
rect 578314 272001 578326 272053
rect 578378 272001 578390 272053
rect 578442 272001 578454 272053
rect 578506 272001 578518 272053
rect 578570 272001 578582 272053
rect 578634 272001 578646 272053
rect 578698 272001 578710 272053
rect 578762 272001 578774 272053
rect 578826 272001 578854 272053
rect 578234 271989 578854 272001
rect 578234 271937 578262 271989
rect 578314 271937 578326 271989
rect 578378 271937 578390 271989
rect 578442 271937 578454 271989
rect 578506 271937 578518 271989
rect 578570 271937 578582 271989
rect 578634 271937 578646 271989
rect 578698 271937 578710 271989
rect 578762 271937 578774 271989
rect 578826 271937 578854 271989
rect 578234 271925 578854 271937
rect 578234 271873 578262 271925
rect 578314 271873 578326 271925
rect 578378 271873 578390 271925
rect 578442 271873 578454 271925
rect 578506 271873 578518 271925
rect 578570 271873 578582 271925
rect 578634 271873 578646 271925
rect 578698 271873 578710 271925
rect 578762 271873 578774 271925
rect 578826 271873 578854 271925
rect 578234 271861 578854 271873
rect 578234 271809 578262 271861
rect 578314 271809 578326 271861
rect 578378 271809 578390 271861
rect 578442 271809 578454 271861
rect 578506 271809 578518 271861
rect 578570 271809 578582 271861
rect 578634 271809 578646 271861
rect 578698 271809 578710 271861
rect 578762 271809 578774 271861
rect 578826 271809 578854 271861
rect 578234 271803 578854 271809
rect 471698 269086 471704 269138
rect 471756 269126 471762 269138
rect 473630 269126 473636 269138
rect 471756 269098 473636 269126
rect 471756 269086 471762 269098
rect 473630 269086 473636 269098
rect 473688 269086 473694 269138
rect 470234 267489 470854 267495
rect 470234 267437 470262 267489
rect 470314 267437 470326 267489
rect 470378 267437 470390 267489
rect 470442 267437 470454 267489
rect 470506 267437 470518 267489
rect 470570 267437 470582 267489
rect 470634 267437 470646 267489
rect 470698 267437 470710 267489
rect 470762 267437 470774 267489
rect 470826 267437 470854 267489
rect 470234 267425 470854 267437
rect 470234 267373 470262 267425
rect 470314 267373 470326 267425
rect 470378 267373 470390 267425
rect 470442 267373 470454 267425
rect 470506 267373 470518 267425
rect 470570 267373 470582 267425
rect 470634 267373 470646 267425
rect 470698 267373 470710 267425
rect 470762 267373 470774 267425
rect 470826 267373 470854 267425
rect 470234 267361 470854 267373
rect 470234 267309 470262 267361
rect 470314 267309 470326 267361
rect 470378 267309 470390 267361
rect 470442 267309 470454 267361
rect 470506 267309 470518 267361
rect 470570 267309 470582 267361
rect 470634 267309 470646 267361
rect 470698 267309 470710 267361
rect 470762 267309 470774 267361
rect 470826 267309 470854 267361
rect 470234 267297 470854 267309
rect 470234 267245 470262 267297
rect 470314 267245 470326 267297
rect 470378 267245 470390 267297
rect 470442 267245 470454 267297
rect 470506 267245 470518 267297
rect 470570 267245 470582 267297
rect 470634 267245 470646 267297
rect 470698 267245 470710 267297
rect 470762 267245 470774 267297
rect 470826 267245 470854 267297
rect 470234 267233 470854 267245
rect 470234 267181 470262 267233
rect 470314 267181 470326 267233
rect 470378 267181 470390 267233
rect 470442 267181 470454 267233
rect 470506 267181 470518 267233
rect 470570 267181 470582 267233
rect 470634 267181 470646 267233
rect 470698 267181 470710 267233
rect 470762 267181 470774 267233
rect 470826 267181 470854 267233
rect 470234 267175 470854 267181
rect 473630 266641 473636 266693
rect 473688 266641 473694 266693
rect 468994 266403 469614 266409
rect 468994 266351 469022 266403
rect 469074 266351 469086 266403
rect 469138 266351 469150 266403
rect 469202 266351 469214 266403
rect 469266 266351 469278 266403
rect 469330 266351 469342 266403
rect 469394 266351 469406 266403
rect 469458 266351 469470 266403
rect 469522 266351 469534 266403
rect 469586 266351 469614 266403
rect 468994 266339 469614 266351
rect 468994 266287 469022 266339
rect 469074 266287 469086 266339
rect 469138 266287 469150 266339
rect 469202 266287 469214 266339
rect 469266 266287 469278 266339
rect 469330 266287 469342 266339
rect 469394 266287 469406 266339
rect 469458 266287 469470 266339
rect 469522 266287 469534 266339
rect 469586 266287 469614 266339
rect 468994 266275 469614 266287
rect 468994 266223 469022 266275
rect 469074 266223 469086 266275
rect 469138 266223 469150 266275
rect 469202 266223 469214 266275
rect 469266 266223 469278 266275
rect 469330 266223 469342 266275
rect 469394 266223 469406 266275
rect 469458 266223 469470 266275
rect 469522 266223 469534 266275
rect 469586 266223 469614 266275
rect 468994 266211 469614 266223
rect 468994 266159 469022 266211
rect 469074 266159 469086 266211
rect 469138 266159 469150 266211
rect 469202 266159 469214 266211
rect 469266 266159 469278 266211
rect 469330 266159 469342 266211
rect 469394 266159 469406 266211
rect 469458 266159 469470 266211
rect 469522 266159 469534 266211
rect 469586 266159 469614 266211
rect 468994 266147 469614 266159
rect 468994 266095 469022 266147
rect 469074 266095 469086 266147
rect 469138 266095 469150 266147
rect 469202 266095 469214 266147
rect 469266 266095 469278 266147
rect 469330 266095 469342 266147
rect 469394 266095 469406 266147
rect 469458 266095 469470 266147
rect 469522 266095 469534 266147
rect 469586 266095 469614 266147
rect 468994 266089 469614 266095
rect 491938 265998 491944 266010
rect 489288 265970 491944 265998
rect 477126 265871 477132 265874
rect 477089 265865 477132 265871
rect 477089 265831 477101 265865
rect 477089 265825 477132 265831
rect 477126 265822 477132 265825
rect 477184 265822 477190 265874
rect 489288 265733 489316 265970
rect 491938 265958 491944 265970
rect 491996 265958 492002 266010
rect 480162 265437 480168 265489
rect 480220 265437 480226 265489
rect 483198 265437 483204 265489
rect 483256 265437 483262 265489
rect 486234 265437 486240 265489
rect 486292 265437 486298 265489
rect 470234 265316 470854 265322
rect 470234 265264 470262 265316
rect 470314 265264 470326 265316
rect 470378 265264 470390 265316
rect 470442 265264 470454 265316
rect 470506 265264 470518 265316
rect 470570 265264 470582 265316
rect 470634 265264 470646 265316
rect 470698 265264 470710 265316
rect 470762 265264 470774 265316
rect 470826 265264 470854 265316
rect 470234 265252 470854 265264
rect 470234 265200 470262 265252
rect 470314 265200 470326 265252
rect 470378 265200 470390 265252
rect 470442 265200 470454 265252
rect 470506 265200 470518 265252
rect 470570 265200 470582 265252
rect 470634 265200 470646 265252
rect 470698 265200 470710 265252
rect 470762 265200 470774 265252
rect 470826 265200 470854 265252
rect 470234 265188 470854 265200
rect 470234 265136 470262 265188
rect 470314 265136 470326 265188
rect 470378 265136 470390 265188
rect 470442 265136 470454 265188
rect 470506 265136 470518 265188
rect 470570 265136 470582 265188
rect 470634 265136 470646 265188
rect 470698 265136 470710 265188
rect 470762 265136 470774 265188
rect 470826 265136 470854 265188
rect 470234 265124 470854 265136
rect 470234 265072 470262 265124
rect 470314 265072 470326 265124
rect 470378 265072 470390 265124
rect 470442 265072 470454 265124
rect 470506 265072 470518 265124
rect 470570 265072 470582 265124
rect 470634 265072 470646 265124
rect 470698 265072 470710 265124
rect 470762 265072 470774 265124
rect 470826 265072 470854 265124
rect 470234 265060 470854 265072
rect 470234 265008 470262 265060
rect 470314 265008 470326 265060
rect 470378 265008 470390 265060
rect 470442 265008 470454 265060
rect 470506 265008 470518 265060
rect 470570 265008 470582 265060
rect 470634 265008 470646 265060
rect 470698 265008 470710 265060
rect 470762 265008 470774 265060
rect 470826 265008 470854 265060
rect 470234 265002 470854 265008
rect 494716 263590 494928 263618
rect 477126 263510 477132 263562
rect 477184 263510 477190 263562
rect 480162 263510 480168 263562
rect 480220 263550 480226 263562
rect 480220 263510 480254 263550
rect 483198 263510 483204 263562
rect 483256 263510 483262 263562
rect 486234 263510 486240 263562
rect 486292 263550 486298 263562
rect 494716 263550 494744 263590
rect 486292 263522 494744 263550
rect 494900 263550 494928 263590
rect 494900 263522 495020 263550
rect 486292 263510 486298 263522
rect 477144 263346 477172 263510
rect 480226 263414 480254 263510
rect 483216 263482 483244 263510
rect 494790 263482 494796 263494
rect 483216 263454 494796 263482
rect 494790 263442 494796 263454
rect 494848 263442 494854 263494
rect 494992 263482 495020 263522
rect 495066 263510 495072 263562
rect 495124 263550 495130 263562
rect 536190 263550 536196 263562
rect 495124 263522 536196 263550
rect 495124 263510 495130 263522
rect 536190 263510 536196 263522
rect 536248 263510 536254 263562
rect 536374 263482 536380 263494
rect 494992 263454 536380 263482
rect 536374 263442 536380 263454
rect 536432 263442 536438 263494
rect 519538 263414 519544 263426
rect 480226 263386 519544 263414
rect 519538 263374 519544 263386
rect 519596 263374 519602 263426
rect 502978 263346 502984 263358
rect 477144 263318 502984 263346
rect 502978 263306 502984 263318
rect 503036 263306 503042 263358
rect 576994 233065 577614 233071
rect 576994 233013 577022 233065
rect 577074 233013 577086 233065
rect 577138 233013 577150 233065
rect 577202 233013 577214 233065
rect 577266 233013 577278 233065
rect 577330 233013 577342 233065
rect 577394 233013 577406 233065
rect 577458 233013 577470 233065
rect 577522 233013 577534 233065
rect 577586 233013 577614 233065
rect 576994 233001 577614 233013
rect 576994 232949 577022 233001
rect 577074 232949 577086 233001
rect 577138 232949 577150 233001
rect 577202 232949 577214 233001
rect 577266 232949 577278 233001
rect 577330 232949 577342 233001
rect 577394 232949 577406 233001
rect 577458 232949 577470 233001
rect 577522 232949 577534 233001
rect 577586 232949 577614 233001
rect 576994 232937 577614 232949
rect 576994 232885 577022 232937
rect 577074 232885 577086 232937
rect 577138 232885 577150 232937
rect 577202 232885 577214 232937
rect 577266 232885 577278 232937
rect 577330 232885 577342 232937
rect 577394 232885 577406 232937
rect 577458 232885 577470 232937
rect 577522 232885 577534 232937
rect 577586 232885 577614 232937
rect 576994 232873 577614 232885
rect 576994 232847 577022 232873
rect 576400 232821 577022 232847
rect 577074 232821 577086 232873
rect 577138 232821 577150 232873
rect 577202 232821 577214 232873
rect 577266 232821 577278 232873
rect 577330 232821 577342 232873
rect 577394 232821 577406 232873
rect 577458 232821 577470 232873
rect 577522 232821 577534 232873
rect 577586 232847 577614 232873
rect 577586 232821 577647 232847
rect 576400 232816 577647 232821
rect 576316 232809 577647 232816
rect 576316 232782 577022 232809
rect 576400 232757 577022 232782
rect 577074 232757 577086 232809
rect 577138 232757 577150 232809
rect 577202 232757 577214 232809
rect 577266 232757 577278 232809
rect 577330 232757 577342 232809
rect 577394 232757 577406 232809
rect 577458 232757 577470 232809
rect 577522 232757 577534 232809
rect 577586 232757 577647 232809
rect 576400 232751 577647 232757
rect 576597 232331 576603 232383
rect 576655 232331 576661 232383
rect 576400 232270 578876 232303
rect 576400 232218 578262 232270
rect 578314 232218 578326 232270
rect 578378 232218 578390 232270
rect 578442 232218 578454 232270
rect 578506 232218 578518 232270
rect 578570 232218 578582 232270
rect 578634 232218 578646 232270
rect 578698 232218 578710 232270
rect 578762 232218 578774 232270
rect 578826 232218 578876 232270
rect 576400 232207 578876 232218
rect 578234 232206 578854 232207
rect 578234 232154 578262 232206
rect 578314 232154 578326 232206
rect 578378 232154 578390 232206
rect 578442 232154 578454 232206
rect 578506 232154 578518 232206
rect 578570 232154 578582 232206
rect 578634 232154 578646 232206
rect 578698 232154 578710 232206
rect 578762 232154 578774 232206
rect 578826 232154 578854 232206
rect 578234 232142 578854 232154
rect 578234 232090 578262 232142
rect 578314 232090 578326 232142
rect 578378 232090 578390 232142
rect 578442 232090 578454 232142
rect 578506 232090 578518 232142
rect 578570 232090 578582 232142
rect 578634 232090 578646 232142
rect 578698 232090 578710 232142
rect 578762 232090 578774 232142
rect 578826 232090 578854 232142
rect 578234 232078 578854 232090
rect 578234 232026 578262 232078
rect 578314 232026 578326 232078
rect 578378 232026 578390 232078
rect 578442 232026 578454 232078
rect 578506 232026 578518 232078
rect 578570 232026 578582 232078
rect 578634 232026 578646 232078
rect 578698 232026 578710 232078
rect 578762 232026 578774 232078
rect 578826 232026 578854 232078
rect 578234 232014 578854 232026
rect 578234 231962 578262 232014
rect 578314 231962 578326 232014
rect 578378 231962 578390 232014
rect 578442 231962 578454 232014
rect 578506 231962 578518 232014
rect 578570 231962 578582 232014
rect 578634 231962 578646 232014
rect 578698 231962 578710 232014
rect 578762 231962 578774 232014
rect 578826 231962 578854 232014
rect 578234 231956 578854 231962
<< via1 >>
rect 254262 703286 254314 703338
rect 254326 703286 254378 703338
rect 254390 703286 254442 703338
rect 254454 703286 254506 703338
rect 254518 703286 254570 703338
rect 254582 703286 254634 703338
rect 254646 703286 254698 703338
rect 254710 703286 254762 703338
rect 254774 703286 254826 703338
rect 254262 703222 254314 703274
rect 254326 703222 254378 703274
rect 254390 703222 254442 703274
rect 254454 703222 254506 703274
rect 254518 703222 254570 703274
rect 254582 703222 254634 703274
rect 254646 703222 254698 703274
rect 254710 703222 254762 703274
rect 254774 703222 254826 703274
rect 254262 703158 254314 703210
rect 254326 703158 254378 703210
rect 254390 703158 254442 703210
rect 254454 703158 254506 703210
rect 254518 703158 254570 703210
rect 254582 703158 254634 703210
rect 254646 703158 254698 703210
rect 254710 703158 254762 703210
rect 254774 703158 254826 703210
rect 326262 703326 326314 703378
rect 326326 703326 326378 703378
rect 326390 703326 326442 703378
rect 326454 703326 326506 703378
rect 326518 703326 326570 703378
rect 326582 703326 326634 703378
rect 326646 703326 326698 703378
rect 326710 703326 326762 703378
rect 326774 703326 326826 703378
rect 326262 703262 326314 703314
rect 326326 703262 326378 703314
rect 326390 703262 326442 703314
rect 326454 703262 326506 703314
rect 326518 703262 326570 703314
rect 326582 703262 326634 703314
rect 326646 703262 326698 703314
rect 326710 703262 326762 703314
rect 326774 703262 326826 703314
rect 326262 703198 326314 703250
rect 326326 703198 326378 703250
rect 326390 703198 326442 703250
rect 326454 703198 326506 703250
rect 326518 703198 326570 703250
rect 326582 703198 326634 703250
rect 326646 703198 326698 703250
rect 326710 703198 326762 703250
rect 326774 703198 326826 703250
rect 254262 703094 254314 703146
rect 254326 703094 254378 703146
rect 254390 703094 254442 703146
rect 254454 703094 254506 703146
rect 254518 703094 254570 703146
rect 254582 703094 254634 703146
rect 254646 703094 254698 703146
rect 254710 703094 254762 703146
rect 254774 703094 254826 703146
rect 326262 703134 326314 703186
rect 326326 703134 326378 703186
rect 326390 703134 326442 703186
rect 326454 703134 326506 703186
rect 326518 703134 326570 703186
rect 326582 703134 326634 703186
rect 326646 703134 326698 703186
rect 326710 703134 326762 703186
rect 326774 703134 326826 703186
rect 254262 703030 254314 703082
rect 254326 703030 254378 703082
rect 254390 703030 254442 703082
rect 254454 703030 254506 703082
rect 254518 703030 254570 703082
rect 254582 703030 254634 703082
rect 254646 703030 254698 703082
rect 254710 703030 254762 703082
rect 254774 703030 254826 703082
rect 326262 703070 326314 703122
rect 326326 703070 326378 703122
rect 326390 703070 326442 703122
rect 326454 703070 326506 703122
rect 326518 703070 326570 703122
rect 326582 703070 326634 703122
rect 326646 703070 326698 703122
rect 326710 703070 326762 703122
rect 326774 703070 326826 703122
rect 362262 702857 362314 702909
rect 362326 702857 362378 702909
rect 362390 702857 362442 702909
rect 362454 702857 362506 702909
rect 362518 702857 362570 702909
rect 362582 702857 362634 702909
rect 362646 702857 362698 702909
rect 362710 702857 362762 702909
rect 362774 702857 362826 702909
rect 362262 702793 362314 702845
rect 362326 702793 362378 702845
rect 362390 702793 362442 702845
rect 362454 702793 362506 702845
rect 362518 702793 362570 702845
rect 362582 702793 362634 702845
rect 362646 702793 362698 702845
rect 362710 702793 362762 702845
rect 362774 702793 362826 702845
rect 362262 702729 362314 702781
rect 362326 702729 362378 702781
rect 362390 702729 362442 702781
rect 362454 702729 362506 702781
rect 362518 702729 362570 702781
rect 362582 702729 362634 702781
rect 362646 702729 362698 702781
rect 362710 702729 362762 702781
rect 362774 702729 362826 702781
rect 252733 702652 252785 702663
rect 252733 702618 252742 702652
rect 252742 702618 252776 702652
rect 252776 702618 252785 702652
rect 252733 702611 252785 702618
rect 324732 702692 324784 702703
rect 324732 702658 324741 702692
rect 324741 702658 324775 702692
rect 324775 702658 324784 702692
rect 324732 702651 324784 702658
rect 362262 702665 362314 702717
rect 362326 702665 362378 702717
rect 362390 702665 362442 702717
rect 362454 702665 362506 702717
rect 362518 702665 362570 702717
rect 362582 702665 362634 702717
rect 362646 702665 362698 702717
rect 362710 702665 362762 702717
rect 362774 702665 362826 702717
rect 434262 702720 434314 702772
rect 434326 702720 434378 702772
rect 434390 702720 434442 702772
rect 434454 702720 434506 702772
rect 434518 702720 434570 702772
rect 434582 702720 434634 702772
rect 434646 702720 434698 702772
rect 434710 702720 434762 702772
rect 434774 702720 434826 702772
rect 253022 702518 253074 702570
rect 253086 702518 253138 702570
rect 253150 702518 253202 702570
rect 253214 702518 253266 702570
rect 253278 702518 253330 702570
rect 253342 702518 253394 702570
rect 253406 702518 253458 702570
rect 253470 702518 253522 702570
rect 253534 702518 253586 702570
rect 325022 702558 325074 702610
rect 325086 702558 325138 702610
rect 325150 702558 325202 702610
rect 325214 702558 325266 702610
rect 325278 702558 325330 702610
rect 325342 702558 325394 702610
rect 325406 702558 325458 702610
rect 325470 702558 325522 702610
rect 325534 702558 325586 702610
rect 362262 702601 362314 702653
rect 362326 702601 362378 702653
rect 362390 702601 362442 702653
rect 362454 702601 362506 702653
rect 362518 702601 362570 702653
rect 362582 702601 362634 702653
rect 362646 702601 362698 702653
rect 362710 702601 362762 702653
rect 362774 702601 362826 702653
rect 434262 702656 434314 702708
rect 434326 702656 434378 702708
rect 434390 702656 434442 702708
rect 434454 702656 434506 702708
rect 434518 702656 434570 702708
rect 434582 702656 434634 702708
rect 434646 702656 434698 702708
rect 434710 702656 434762 702708
rect 434774 702656 434826 702708
rect 434262 702592 434314 702644
rect 434326 702592 434378 702644
rect 434390 702592 434442 702644
rect 434454 702592 434506 702644
rect 434518 702592 434570 702644
rect 434582 702592 434634 702644
rect 434646 702592 434698 702644
rect 434710 702592 434762 702644
rect 434774 702592 434826 702644
rect 253022 702454 253074 702506
rect 253086 702454 253138 702506
rect 253150 702454 253202 702506
rect 253214 702454 253266 702506
rect 253278 702454 253330 702506
rect 253342 702454 253394 702506
rect 253406 702454 253458 702506
rect 253470 702454 253522 702506
rect 253534 702454 253586 702506
rect 325022 702494 325074 702546
rect 325086 702494 325138 702546
rect 325150 702494 325202 702546
rect 325214 702494 325266 702546
rect 325278 702494 325330 702546
rect 325342 702494 325394 702546
rect 325406 702494 325458 702546
rect 325470 702494 325522 702546
rect 325534 702494 325586 702546
rect 434262 702528 434314 702580
rect 434326 702528 434378 702580
rect 434390 702528 434442 702580
rect 434454 702528 434506 702580
rect 434518 702528 434570 702580
rect 434582 702528 434634 702580
rect 434646 702528 434698 702580
rect 434710 702528 434762 702580
rect 434774 702528 434826 702580
rect 253022 702390 253074 702442
rect 253086 702390 253138 702442
rect 253150 702390 253202 702442
rect 253214 702390 253266 702442
rect 253278 702390 253330 702442
rect 253342 702390 253394 702442
rect 253406 702390 253458 702442
rect 253470 702390 253522 702442
rect 253534 702390 253586 702442
rect 253022 702326 253074 702378
rect 253086 702326 253138 702378
rect 253150 702326 253202 702378
rect 253214 702326 253266 702378
rect 253278 702326 253330 702378
rect 253342 702326 253394 702378
rect 253406 702326 253458 702378
rect 253470 702326 253522 702378
rect 253534 702326 253586 702378
rect 253022 702262 253074 702314
rect 253086 702262 253138 702314
rect 253150 702262 253202 702314
rect 253214 702262 253266 702314
rect 253278 702262 253330 702314
rect 253342 702262 253394 702314
rect 253406 702262 253458 702314
rect 253470 702262 253522 702314
rect 253534 702262 253586 702314
rect 325022 702430 325074 702482
rect 325086 702430 325138 702482
rect 325150 702430 325202 702482
rect 325214 702430 325266 702482
rect 325278 702430 325330 702482
rect 325342 702430 325394 702482
rect 325406 702430 325458 702482
rect 325470 702430 325522 702482
rect 325534 702430 325586 702482
rect 434262 702464 434314 702516
rect 434326 702464 434378 702516
rect 434390 702464 434442 702516
rect 434454 702464 434506 702516
rect 434518 702464 434570 702516
rect 434582 702464 434634 702516
rect 434646 702464 434698 702516
rect 434710 702464 434762 702516
rect 434774 702464 434826 702516
rect 506262 702474 506314 702526
rect 506326 702474 506378 702526
rect 506390 702474 506442 702526
rect 506454 702474 506506 702526
rect 506518 702474 506570 702526
rect 506582 702474 506634 702526
rect 506646 702474 506698 702526
rect 506710 702474 506762 702526
rect 506774 702474 506826 702526
rect 325022 702366 325074 702418
rect 325086 702366 325138 702418
rect 325150 702366 325202 702418
rect 325214 702366 325266 702418
rect 325278 702366 325330 702418
rect 325342 702366 325394 702418
rect 325406 702366 325458 702418
rect 325470 702366 325522 702418
rect 325534 702366 325586 702418
rect 325022 702302 325074 702354
rect 325086 702302 325138 702354
rect 325150 702302 325202 702354
rect 325214 702302 325266 702354
rect 325278 702302 325330 702354
rect 325342 702302 325394 702354
rect 325406 702302 325458 702354
rect 325470 702302 325522 702354
rect 325534 702302 325586 702354
rect 506262 702410 506314 702462
rect 506326 702410 506378 702462
rect 506390 702410 506442 702462
rect 506454 702410 506506 702462
rect 506518 702410 506570 702462
rect 506582 702410 506634 702462
rect 506646 702410 506698 702462
rect 506710 702410 506762 702462
rect 506774 702410 506826 702462
rect 506262 702346 506314 702398
rect 506326 702346 506378 702398
rect 506390 702346 506442 702398
rect 506454 702346 506506 702398
rect 506518 702346 506570 702398
rect 506582 702346 506634 702398
rect 506646 702346 506698 702398
rect 506710 702346 506762 702398
rect 506774 702346 506826 702398
rect 506262 702282 506314 702334
rect 506326 702282 506378 702334
rect 506390 702282 506442 702334
rect 506454 702282 506506 702334
rect 506518 702282 506570 702334
rect 506582 702282 506634 702334
rect 506646 702282 506698 702334
rect 506710 702282 506762 702334
rect 506774 702282 506826 702334
rect 360759 702223 360811 702234
rect 360759 702189 360768 702223
rect 360768 702189 360802 702223
rect 360802 702189 360811 702223
rect 360759 702182 360811 702189
rect 506262 702218 506314 702270
rect 506326 702218 506378 702270
rect 506390 702218 506442 702270
rect 506454 702218 506506 702270
rect 506518 702218 506570 702270
rect 506582 702218 506634 702270
rect 506646 702218 506698 702270
rect 506710 702218 506762 702270
rect 506774 702218 506826 702270
rect 361022 702089 361074 702141
rect 361086 702089 361138 702141
rect 361150 702089 361202 702141
rect 361214 702089 361266 702141
rect 361278 702089 361330 702141
rect 361342 702089 361394 702141
rect 361406 702089 361458 702141
rect 361470 702089 361522 702141
rect 361534 702089 361586 702141
rect 361022 702025 361074 702077
rect 361086 702025 361138 702077
rect 361150 702025 361202 702077
rect 361214 702025 361266 702077
rect 361278 702025 361330 702077
rect 361342 702025 361394 702077
rect 361406 702025 361458 702077
rect 361470 702025 361522 702077
rect 361534 702025 361586 702077
rect 432729 702086 432781 702097
rect 432729 702052 432738 702086
rect 432738 702052 432772 702086
rect 432772 702052 432781 702086
rect 432729 702045 432781 702052
rect 361022 701961 361074 702013
rect 361086 701961 361138 702013
rect 361150 701961 361202 702013
rect 361214 701961 361266 702013
rect 361278 701961 361330 702013
rect 361342 701961 361394 702013
rect 361406 701961 361458 702013
rect 361470 701961 361522 702013
rect 361534 701961 361586 702013
rect 433022 701952 433074 702004
rect 433086 701952 433138 702004
rect 433150 701952 433202 702004
rect 433214 701952 433266 702004
rect 433278 701952 433330 702004
rect 433342 701952 433394 702004
rect 433406 701952 433458 702004
rect 433470 701952 433522 702004
rect 433534 701952 433586 702004
rect 361022 701897 361074 701949
rect 361086 701897 361138 701949
rect 361150 701897 361202 701949
rect 361214 701897 361266 701949
rect 361278 701897 361330 701949
rect 361342 701897 361394 701949
rect 361406 701897 361458 701949
rect 361470 701897 361522 701949
rect 361534 701897 361586 701949
rect 361022 701833 361074 701885
rect 361086 701833 361138 701885
rect 361150 701833 361202 701885
rect 361214 701833 361266 701885
rect 361278 701833 361330 701885
rect 361342 701833 361394 701885
rect 361406 701833 361458 701885
rect 361470 701833 361522 701885
rect 361534 701833 361586 701885
rect 433022 701888 433074 701940
rect 433086 701888 433138 701940
rect 433150 701888 433202 701940
rect 433214 701888 433266 701940
rect 433278 701888 433330 701940
rect 433342 701888 433394 701940
rect 433406 701888 433458 701940
rect 433470 701888 433522 701940
rect 433534 701888 433586 701940
rect 433022 701824 433074 701876
rect 433086 701824 433138 701876
rect 433150 701824 433202 701876
rect 433214 701824 433266 701876
rect 433278 701824 433330 701876
rect 433342 701824 433394 701876
rect 433406 701824 433458 701876
rect 433470 701824 433522 701876
rect 433534 701824 433586 701876
rect 433022 701760 433074 701812
rect 433086 701760 433138 701812
rect 433150 701760 433202 701812
rect 433214 701760 433266 701812
rect 433278 701760 433330 701812
rect 433342 701760 433394 701812
rect 433406 701760 433458 701812
rect 433470 701760 433522 701812
rect 433534 701760 433586 701812
rect 504725 701840 504777 701851
rect 504725 701806 504734 701840
rect 504734 701806 504768 701840
rect 504768 701806 504777 701840
rect 504725 701799 504777 701806
rect 433022 701696 433074 701748
rect 433086 701696 433138 701748
rect 433150 701696 433202 701748
rect 433214 701696 433266 701748
rect 433278 701696 433330 701748
rect 433342 701696 433394 701748
rect 433406 701696 433458 701748
rect 433470 701696 433522 701748
rect 433534 701696 433586 701748
rect 505022 701706 505074 701758
rect 505086 701706 505138 701758
rect 505150 701706 505202 701758
rect 505214 701706 505266 701758
rect 505278 701706 505330 701758
rect 505342 701706 505394 701758
rect 505406 701706 505458 701758
rect 505470 701706 505522 701758
rect 505534 701706 505586 701758
rect 505022 701642 505074 701694
rect 505086 701642 505138 701694
rect 505150 701642 505202 701694
rect 505214 701642 505266 701694
rect 505278 701642 505330 701694
rect 505342 701642 505394 701694
rect 505406 701642 505458 701694
rect 505470 701642 505522 701694
rect 505534 701642 505586 701694
rect 505022 701578 505074 701630
rect 505086 701578 505138 701630
rect 505150 701578 505202 701630
rect 505214 701578 505266 701630
rect 505278 701578 505330 701630
rect 505342 701578 505394 701630
rect 505406 701578 505458 701630
rect 505470 701578 505522 701630
rect 505534 701578 505586 701630
rect 505022 701514 505074 701566
rect 505086 701514 505138 701566
rect 505150 701514 505202 701566
rect 505214 701514 505266 701566
rect 505278 701514 505330 701566
rect 505342 701514 505394 701566
rect 505406 701514 505458 701566
rect 505470 701514 505522 701566
rect 505534 701514 505586 701566
rect 505022 701450 505074 701502
rect 505086 701450 505138 701502
rect 505150 701450 505202 701502
rect 505214 701450 505266 701502
rect 505278 701450 505330 701502
rect 505342 701450 505394 701502
rect 505406 701450 505458 701502
rect 505470 701450 505522 701502
rect 505534 701450 505586 701502
rect 267648 700954 267700 701006
rect 332508 700954 332560 701006
rect 397460 700954 397512 701006
rect 462320 700954 462372 701006
rect 527180 700954 527232 701006
rect 577022 697860 577074 697912
rect 577086 697860 577138 697912
rect 577150 697860 577202 697912
rect 577214 697860 577266 697912
rect 577278 697860 577330 697912
rect 577342 697860 577394 697912
rect 577406 697860 577458 697912
rect 577470 697860 577522 697912
rect 577534 697860 577586 697912
rect 577022 697796 577074 697848
rect 577086 697796 577138 697848
rect 577150 697796 577202 697848
rect 577214 697796 577266 697848
rect 577278 697796 577330 697848
rect 577342 697796 577394 697848
rect 577406 697796 577458 697848
rect 577470 697796 577522 697848
rect 577534 697796 577586 697848
rect 577022 697732 577074 697784
rect 577086 697732 577138 697784
rect 577150 697732 577202 697784
rect 577214 697732 577266 697784
rect 577278 697732 577330 697784
rect 577342 697732 577394 697784
rect 577406 697732 577458 697784
rect 577470 697732 577522 697784
rect 577534 697732 577586 697784
rect 577022 697668 577074 697720
rect 577086 697668 577138 697720
rect 577150 697668 577202 697720
rect 577214 697668 577266 697720
rect 577278 697668 577330 697720
rect 577342 697668 577394 697720
rect 577406 697668 577458 697720
rect 577470 697668 577522 697720
rect 577534 697668 577586 697720
rect 577022 697604 577074 697656
rect 577086 697604 577138 697656
rect 577150 697604 577202 697656
rect 577214 697604 577266 697656
rect 577278 697604 577330 697656
rect 577342 697604 577394 697656
rect 577406 697604 577458 697656
rect 577470 697604 577522 697656
rect 577534 697604 577586 697656
rect 576603 697221 576655 697230
rect 576603 697187 576613 697221
rect 576613 697187 576647 697221
rect 576647 697187 576655 697221
rect 576603 697178 576655 697187
rect 578262 697065 578314 697117
rect 578326 697065 578378 697117
rect 578390 697065 578442 697117
rect 578454 697065 578506 697117
rect 578518 697065 578570 697117
rect 578582 697065 578634 697117
rect 578646 697065 578698 697117
rect 578710 697065 578762 697117
rect 578774 697065 578826 697117
rect 578262 697001 578314 697053
rect 578326 697001 578378 697053
rect 578390 697001 578442 697053
rect 578454 697001 578506 697053
rect 578518 697001 578570 697053
rect 578582 697001 578634 697053
rect 578646 697001 578698 697053
rect 578710 697001 578762 697053
rect 578774 697001 578826 697053
rect 578262 696937 578314 696989
rect 578326 696937 578378 696989
rect 578390 696937 578442 696989
rect 578454 696937 578506 696989
rect 578518 696937 578570 696989
rect 578582 696937 578634 696989
rect 578646 696937 578698 696989
rect 578710 696937 578762 696989
rect 578774 696937 578826 696989
rect 578262 696873 578314 696925
rect 578326 696873 578378 696925
rect 578390 696873 578442 696925
rect 578454 696873 578506 696925
rect 578518 696873 578570 696925
rect 578582 696873 578634 696925
rect 578646 696873 578698 696925
rect 578710 696873 578762 696925
rect 578774 696873 578826 696925
rect 578262 696809 578314 696861
rect 578326 696809 578378 696861
rect 578390 696809 578442 696861
rect 578454 696809 578506 696861
rect 578518 696809 578570 696861
rect 578582 696809 578634 696861
rect 578646 696809 578698 696861
rect 578710 696809 578762 696861
rect 578774 696809 578826 696861
rect 577022 644684 577074 644736
rect 577086 644684 577138 644736
rect 577150 644684 577202 644736
rect 577214 644684 577266 644736
rect 577278 644684 577330 644736
rect 577342 644684 577394 644736
rect 577406 644684 577458 644736
rect 577470 644684 577522 644736
rect 577534 644684 577586 644736
rect 577022 644620 577074 644672
rect 577086 644620 577138 644672
rect 577150 644620 577202 644672
rect 577214 644620 577266 644672
rect 577278 644620 577330 644672
rect 577342 644620 577394 644672
rect 577406 644620 577458 644672
rect 577470 644620 577522 644672
rect 577534 644620 577586 644672
rect 577022 644556 577074 644608
rect 577086 644556 577138 644608
rect 577150 644556 577202 644608
rect 577214 644556 577266 644608
rect 577278 644556 577330 644608
rect 577342 644556 577394 644608
rect 577406 644556 577458 644608
rect 577470 644556 577522 644608
rect 577534 644556 577586 644608
rect 577022 644492 577074 644544
rect 577086 644492 577138 644544
rect 577150 644492 577202 644544
rect 577214 644492 577266 644544
rect 577278 644492 577330 644544
rect 577342 644492 577394 644544
rect 577406 644492 577458 644544
rect 577470 644492 577522 644544
rect 577534 644492 577586 644544
rect 577022 644428 577074 644480
rect 577086 644428 577138 644480
rect 577150 644428 577202 644480
rect 577214 644428 577266 644480
rect 577278 644428 577330 644480
rect 577342 644428 577394 644480
rect 577406 644428 577458 644480
rect 577470 644428 577522 644480
rect 577534 644428 577586 644480
rect 576603 644045 576655 644054
rect 576603 644011 576613 644045
rect 576613 644011 576647 644045
rect 576647 644011 576655 644045
rect 576603 644002 576655 644011
rect 578262 643889 578314 643941
rect 578326 643889 578378 643941
rect 578390 643889 578442 643941
rect 578454 643889 578506 643941
rect 578518 643889 578570 643941
rect 578582 643889 578634 643941
rect 578646 643889 578698 643941
rect 578710 643889 578762 643941
rect 578774 643889 578826 643941
rect 578262 643825 578314 643877
rect 578326 643825 578378 643877
rect 578390 643825 578442 643877
rect 578454 643825 578506 643877
rect 578518 643825 578570 643877
rect 578582 643825 578634 643877
rect 578646 643825 578698 643877
rect 578710 643825 578762 643877
rect 578774 643825 578826 643877
rect 578262 643761 578314 643813
rect 578326 643761 578378 643813
rect 578390 643761 578442 643813
rect 578454 643761 578506 643813
rect 578518 643761 578570 643813
rect 578582 643761 578634 643813
rect 578646 643761 578698 643813
rect 578710 643761 578762 643813
rect 578774 643761 578826 643813
rect 578262 643697 578314 643749
rect 578326 643697 578378 643749
rect 578390 643697 578442 643749
rect 578454 643697 578506 643749
rect 578518 643697 578570 643749
rect 578582 643697 578634 643749
rect 578646 643697 578698 643749
rect 578710 643697 578762 643749
rect 578774 643697 578826 643749
rect 578262 643633 578314 643685
rect 578326 643633 578378 643685
rect 578390 643633 578442 643685
rect 578454 643633 578506 643685
rect 578518 643633 578570 643685
rect 578582 643633 578634 643685
rect 578646 643633 578698 643685
rect 578710 643633 578762 643685
rect 578774 643633 578826 643685
rect 577022 591644 577074 591696
rect 577086 591644 577138 591696
rect 577150 591644 577202 591696
rect 577214 591644 577266 591696
rect 577278 591644 577330 591696
rect 577342 591644 577394 591696
rect 577406 591644 577458 591696
rect 577470 591644 577522 591696
rect 577534 591644 577586 591696
rect 577022 591580 577074 591632
rect 577086 591580 577138 591632
rect 577150 591580 577202 591632
rect 577214 591580 577266 591632
rect 577278 591580 577330 591632
rect 577342 591580 577394 591632
rect 577406 591580 577458 591632
rect 577470 591580 577522 591632
rect 577534 591580 577586 591632
rect 577022 591516 577074 591568
rect 577086 591516 577138 591568
rect 577150 591516 577202 591568
rect 577214 591516 577266 591568
rect 577278 591516 577330 591568
rect 577342 591516 577394 591568
rect 577406 591516 577458 591568
rect 577470 591516 577522 591568
rect 577534 591516 577586 591568
rect 577022 591452 577074 591504
rect 577086 591452 577138 591504
rect 577150 591452 577202 591504
rect 577214 591452 577266 591504
rect 577278 591452 577330 591504
rect 577342 591452 577394 591504
rect 577406 591452 577458 591504
rect 577470 591452 577522 591504
rect 577534 591452 577586 591504
rect 577022 591388 577074 591440
rect 577086 591388 577138 591440
rect 577150 591388 577202 591440
rect 577214 591388 577266 591440
rect 577278 591388 577330 591440
rect 577342 591388 577394 591440
rect 577406 591388 577458 591440
rect 577470 591388 577522 591440
rect 577534 591388 577586 591440
rect 576603 591005 576655 591014
rect 576603 590971 576613 591005
rect 576613 590971 576647 591005
rect 576647 590971 576655 591005
rect 576603 590962 576655 590971
rect 578262 590849 578314 590901
rect 578326 590849 578378 590901
rect 578390 590849 578442 590901
rect 578454 590849 578506 590901
rect 578518 590849 578570 590901
rect 578582 590849 578634 590901
rect 578646 590849 578698 590901
rect 578710 590849 578762 590901
rect 578774 590849 578826 590901
rect 578262 590785 578314 590837
rect 578326 590785 578378 590837
rect 578390 590785 578442 590837
rect 578454 590785 578506 590837
rect 578518 590785 578570 590837
rect 578582 590785 578634 590837
rect 578646 590785 578698 590837
rect 578710 590785 578762 590837
rect 578774 590785 578826 590837
rect 578262 590721 578314 590773
rect 578326 590721 578378 590773
rect 578390 590721 578442 590773
rect 578454 590721 578506 590773
rect 578518 590721 578570 590773
rect 578582 590721 578634 590773
rect 578646 590721 578698 590773
rect 578710 590721 578762 590773
rect 578774 590721 578826 590773
rect 578262 590657 578314 590709
rect 578326 590657 578378 590709
rect 578390 590657 578442 590709
rect 578454 590657 578506 590709
rect 578518 590657 578570 590709
rect 578582 590657 578634 590709
rect 578646 590657 578698 590709
rect 578710 590657 578762 590709
rect 578774 590657 578826 590709
rect 578262 590593 578314 590645
rect 578326 590593 578378 590645
rect 578390 590593 578442 590645
rect 578454 590593 578506 590645
rect 578518 590593 578570 590645
rect 578582 590593 578634 590645
rect 578646 590593 578698 590645
rect 578710 590593 578762 590645
rect 578774 590593 578826 590645
rect 505022 554552 505074 554604
rect 505086 554552 505138 554604
rect 505150 554552 505202 554604
rect 505214 554552 505266 554604
rect 505278 554552 505330 554604
rect 505342 554552 505394 554604
rect 505406 554552 505458 554604
rect 505470 554552 505522 554604
rect 505534 554552 505586 554604
rect 505022 554488 505074 554540
rect 505086 554488 505138 554540
rect 505150 554488 505202 554540
rect 505214 554488 505266 554540
rect 505278 554488 505330 554540
rect 505342 554488 505394 554540
rect 505406 554488 505458 554540
rect 505470 554488 505522 554540
rect 505534 554488 505586 554540
rect 505022 554424 505074 554476
rect 505086 554424 505138 554476
rect 505150 554424 505202 554476
rect 505214 554424 505266 554476
rect 505278 554424 505330 554476
rect 505342 554424 505394 554476
rect 505406 554424 505458 554476
rect 505470 554424 505522 554476
rect 505534 554424 505586 554476
rect 505022 554360 505074 554412
rect 505086 554360 505138 554412
rect 505150 554360 505202 554412
rect 505214 554360 505266 554412
rect 505278 554360 505330 554412
rect 505342 554360 505394 554412
rect 505406 554360 505458 554412
rect 505470 554360 505522 554412
rect 505534 554360 505586 554412
rect 505022 554296 505074 554348
rect 505086 554296 505138 554348
rect 505150 554296 505202 554348
rect 505214 554296 505266 554348
rect 505278 554296 505330 554348
rect 505342 554296 505394 554348
rect 505406 554296 505458 554348
rect 505470 554296 505522 554348
rect 505534 554296 505586 554348
rect 536104 554006 536156 554058
rect 506262 553757 506314 553809
rect 506326 553757 506378 553809
rect 506390 553757 506442 553809
rect 506454 553757 506506 553809
rect 506518 553757 506570 553809
rect 506582 553757 506634 553809
rect 506646 553757 506698 553809
rect 506710 553757 506762 553809
rect 506774 553757 506826 553809
rect 506262 553693 506314 553745
rect 506326 553693 506378 553745
rect 506390 553693 506442 553745
rect 506454 553693 506506 553745
rect 506518 553693 506570 553745
rect 506582 553693 506634 553745
rect 506646 553693 506698 553745
rect 506710 553693 506762 553745
rect 506774 553693 506826 553745
rect 506262 553629 506314 553681
rect 506326 553629 506378 553681
rect 506390 553629 506442 553681
rect 506454 553629 506506 553681
rect 506518 553629 506570 553681
rect 506582 553629 506634 553681
rect 506646 553629 506698 553681
rect 506710 553629 506762 553681
rect 506774 553629 506826 553681
rect 506262 553565 506314 553617
rect 506326 553565 506378 553617
rect 506390 553565 506442 553617
rect 506454 553565 506506 553617
rect 506518 553565 506570 553617
rect 506582 553565 506634 553617
rect 506646 553565 506698 553617
rect 506710 553565 506762 553617
rect 506774 553565 506826 553617
rect 506262 553501 506314 553553
rect 506326 553501 506378 553553
rect 506390 553501 506442 553553
rect 506454 553501 506506 553553
rect 506518 553501 506570 553553
rect 506582 553501 506634 553553
rect 506646 553501 506698 553553
rect 506710 553501 506762 553553
rect 506774 553501 506826 553553
rect 577022 538468 577074 538520
rect 577086 538468 577138 538520
rect 577150 538468 577202 538520
rect 577214 538468 577266 538520
rect 577278 538468 577330 538520
rect 577342 538468 577394 538520
rect 577406 538468 577458 538520
rect 577470 538468 577522 538520
rect 577534 538468 577586 538520
rect 577022 538404 577074 538456
rect 577086 538404 577138 538456
rect 577150 538404 577202 538456
rect 577214 538404 577266 538456
rect 577278 538404 577330 538456
rect 577342 538404 577394 538456
rect 577406 538404 577458 538456
rect 577470 538404 577522 538456
rect 577534 538404 577586 538456
rect 577022 538340 577074 538392
rect 577086 538340 577138 538392
rect 577150 538340 577202 538392
rect 577214 538340 577266 538392
rect 577278 538340 577330 538392
rect 577342 538340 577394 538392
rect 577406 538340 577458 538392
rect 577470 538340 577522 538392
rect 577534 538340 577586 538392
rect 577022 538276 577074 538328
rect 577086 538276 577138 538328
rect 577150 538276 577202 538328
rect 577214 538276 577266 538328
rect 577278 538276 577330 538328
rect 577342 538276 577394 538328
rect 577406 538276 577458 538328
rect 577470 538276 577522 538328
rect 577534 538276 577586 538328
rect 577022 538212 577074 538264
rect 577086 538212 577138 538264
rect 577150 538212 577202 538264
rect 577214 538212 577266 538264
rect 577278 538212 577330 538264
rect 577342 538212 577394 538264
rect 577406 538212 577458 538264
rect 577470 538212 577522 538264
rect 577534 538212 577586 538264
rect 576603 537829 576655 537838
rect 576603 537795 576613 537829
rect 576613 537795 576647 537829
rect 576647 537795 576655 537829
rect 576603 537786 576655 537795
rect 578262 537673 578314 537725
rect 578326 537673 578378 537725
rect 578390 537673 578442 537725
rect 578454 537673 578506 537725
rect 578518 537673 578570 537725
rect 578582 537673 578634 537725
rect 578646 537673 578698 537725
rect 578710 537673 578762 537725
rect 578774 537673 578826 537725
rect 578262 537609 578314 537661
rect 578326 537609 578378 537661
rect 578390 537609 578442 537661
rect 578454 537609 578506 537661
rect 578518 537609 578570 537661
rect 578582 537609 578634 537661
rect 578646 537609 578698 537661
rect 578710 537609 578762 537661
rect 578774 537609 578826 537661
rect 578262 537545 578314 537597
rect 578326 537545 578378 537597
rect 578390 537545 578442 537597
rect 578454 537545 578506 537597
rect 578518 537545 578570 537597
rect 578582 537545 578634 537597
rect 578646 537545 578698 537597
rect 578710 537545 578762 537597
rect 578774 537545 578826 537597
rect 578262 537481 578314 537533
rect 578326 537481 578378 537533
rect 578390 537481 578442 537533
rect 578454 537481 578506 537533
rect 578518 537481 578570 537533
rect 578582 537481 578634 537533
rect 578646 537481 578698 537533
rect 578710 537481 578762 537533
rect 578774 537481 578826 537533
rect 578262 537417 578314 537469
rect 578326 537417 578378 537469
rect 578390 537417 578442 537469
rect 578454 537417 578506 537469
rect 578518 537417 578570 537469
rect 578582 537417 578634 537469
rect 578646 537417 578698 537469
rect 578710 537417 578762 537469
rect 578774 537417 578826 537469
rect 577022 485292 577074 485344
rect 577086 485292 577138 485344
rect 577150 485292 577202 485344
rect 577214 485292 577266 485344
rect 577278 485292 577330 485344
rect 577342 485292 577394 485344
rect 577406 485292 577458 485344
rect 577470 485292 577522 485344
rect 577534 485292 577586 485344
rect 577022 485228 577074 485280
rect 577086 485228 577138 485280
rect 577150 485228 577202 485280
rect 577214 485228 577266 485280
rect 577278 485228 577330 485280
rect 577342 485228 577394 485280
rect 577406 485228 577458 485280
rect 577470 485228 577522 485280
rect 577534 485228 577586 485280
rect 577022 485164 577074 485216
rect 577086 485164 577138 485216
rect 577150 485164 577202 485216
rect 577214 485164 577266 485216
rect 577278 485164 577330 485216
rect 577342 485164 577394 485216
rect 577406 485164 577458 485216
rect 577470 485164 577522 485216
rect 577534 485164 577586 485216
rect 577022 485100 577074 485152
rect 577086 485100 577138 485152
rect 577150 485100 577202 485152
rect 577214 485100 577266 485152
rect 577278 485100 577330 485152
rect 577342 485100 577394 485152
rect 577406 485100 577458 485152
rect 577470 485100 577522 485152
rect 577534 485100 577586 485152
rect 577022 485036 577074 485088
rect 577086 485036 577138 485088
rect 577150 485036 577202 485088
rect 577214 485036 577266 485088
rect 577278 485036 577330 485088
rect 577342 485036 577394 485088
rect 577406 485036 577458 485088
rect 577470 485036 577522 485088
rect 577534 485036 577586 485088
rect 576603 484653 576655 484662
rect 576603 484619 576613 484653
rect 576613 484619 576647 484653
rect 576647 484619 576655 484653
rect 576603 484610 576655 484619
rect 578262 484497 578314 484549
rect 578326 484497 578378 484549
rect 578390 484497 578442 484549
rect 578454 484497 578506 484549
rect 578518 484497 578570 484549
rect 578582 484497 578634 484549
rect 578646 484497 578698 484549
rect 578710 484497 578762 484549
rect 578774 484497 578826 484549
rect 578262 484433 578314 484485
rect 578326 484433 578378 484485
rect 578390 484433 578442 484485
rect 578454 484433 578506 484485
rect 578518 484433 578570 484485
rect 578582 484433 578634 484485
rect 578646 484433 578698 484485
rect 578710 484433 578762 484485
rect 578774 484433 578826 484485
rect 578262 484369 578314 484421
rect 578326 484369 578378 484421
rect 578390 484369 578442 484421
rect 578454 484369 578506 484421
rect 578518 484369 578570 484421
rect 578582 484369 578634 484421
rect 578646 484369 578698 484421
rect 578710 484369 578762 484421
rect 578774 484369 578826 484421
rect 578262 484305 578314 484357
rect 578326 484305 578378 484357
rect 578390 484305 578442 484357
rect 578454 484305 578506 484357
rect 578518 484305 578570 484357
rect 578582 484305 578634 484357
rect 578646 484305 578698 484357
rect 578710 484305 578762 484357
rect 578774 484305 578826 484357
rect 578262 484241 578314 484293
rect 578326 484241 578378 484293
rect 578390 484241 578442 484293
rect 578454 484241 578506 484293
rect 578518 484241 578570 484293
rect 578582 484241 578634 484293
rect 578646 484241 578698 484293
rect 578710 484241 578762 484293
rect 578774 484241 578826 484293
rect 471704 453298 471756 453350
rect 580172 453298 580224 453350
rect 470262 451435 470314 451487
rect 470326 451435 470378 451487
rect 470390 451435 470442 451487
rect 470454 451435 470506 451487
rect 470518 451435 470570 451487
rect 470582 451435 470634 451487
rect 470646 451435 470698 451487
rect 470710 451435 470762 451487
rect 470774 451435 470826 451487
rect 470262 451371 470314 451423
rect 470326 451371 470378 451423
rect 470390 451371 470442 451423
rect 470454 451371 470506 451423
rect 470518 451371 470570 451423
rect 470582 451371 470634 451423
rect 470646 451371 470698 451423
rect 470710 451371 470762 451423
rect 470774 451371 470826 451423
rect 470262 451307 470314 451359
rect 470326 451307 470378 451359
rect 470390 451307 470442 451359
rect 470454 451307 470506 451359
rect 470518 451307 470570 451359
rect 470582 451307 470634 451359
rect 470646 451307 470698 451359
rect 470710 451307 470762 451359
rect 470774 451307 470826 451359
rect 470262 451243 470314 451295
rect 470326 451243 470378 451295
rect 470390 451243 470442 451295
rect 470454 451243 470506 451295
rect 470518 451243 470570 451295
rect 470582 451243 470634 451295
rect 470646 451243 470698 451295
rect 470710 451243 470762 451295
rect 470774 451243 470826 451295
rect 470262 451179 470314 451231
rect 470326 451179 470378 451231
rect 470390 451179 470442 451231
rect 470454 451179 470506 451231
rect 470518 451179 470570 451231
rect 470582 451179 470634 451231
rect 470646 451179 470698 451231
rect 470710 451179 470762 451231
rect 470774 451179 470826 451231
rect 471704 450442 471756 450494
rect 469022 450349 469074 450401
rect 469086 450349 469138 450401
rect 469150 450349 469202 450401
rect 469214 450349 469266 450401
rect 469278 450349 469330 450401
rect 469342 450349 469394 450401
rect 469406 450349 469458 450401
rect 469470 450349 469522 450401
rect 469534 450349 469586 450401
rect 469022 450285 469074 450337
rect 469086 450285 469138 450337
rect 469150 450285 469202 450337
rect 469214 450285 469266 450337
rect 469278 450285 469330 450337
rect 469342 450285 469394 450337
rect 469406 450285 469458 450337
rect 469470 450285 469522 450337
rect 469534 450285 469586 450337
rect 469022 450221 469074 450273
rect 469086 450221 469138 450273
rect 469150 450221 469202 450273
rect 469214 450221 469266 450273
rect 469278 450221 469330 450273
rect 469342 450221 469394 450273
rect 469406 450221 469458 450273
rect 469470 450221 469522 450273
rect 469534 450221 469586 450273
rect 469022 450157 469074 450209
rect 469086 450157 469138 450209
rect 469150 450157 469202 450209
rect 469214 450157 469266 450209
rect 469278 450157 469330 450209
rect 469342 450157 469394 450209
rect 469406 450157 469458 450209
rect 469470 450157 469522 450209
rect 469534 450157 469586 450209
rect 469022 450093 469074 450145
rect 469086 450093 469138 450145
rect 469150 450093 469202 450145
rect 469214 450093 469266 450145
rect 469278 450093 469330 450145
rect 469342 450093 469394 450145
rect 469406 450093 469458 450145
rect 469470 450093 469522 450145
rect 469534 450093 469586 450145
rect 475384 449438 475436 449490
rect 478696 449438 478748 449490
rect 482008 449438 482060 449490
rect 485320 449438 485372 449490
rect 491944 449354 491996 449406
rect 470262 449264 470314 449316
rect 470326 449264 470378 449316
rect 470390 449264 470442 449316
rect 470454 449264 470506 449316
rect 470518 449264 470570 449316
rect 470582 449264 470634 449316
rect 470646 449264 470698 449316
rect 470710 449264 470762 449316
rect 470774 449264 470826 449316
rect 470262 449200 470314 449252
rect 470326 449200 470378 449252
rect 470390 449200 470442 449252
rect 470454 449200 470506 449252
rect 470518 449200 470570 449252
rect 470582 449200 470634 449252
rect 470646 449200 470698 449252
rect 470710 449200 470762 449252
rect 470774 449200 470826 449252
rect 470262 449136 470314 449188
rect 470326 449136 470378 449188
rect 470390 449136 470442 449188
rect 470454 449136 470506 449188
rect 470518 449136 470570 449188
rect 470582 449136 470634 449188
rect 470646 449136 470698 449188
rect 470710 449136 470762 449188
rect 470774 449136 470826 449188
rect 470262 449072 470314 449124
rect 470326 449072 470378 449124
rect 470390 449072 470442 449124
rect 470454 449072 470506 449124
rect 470518 449072 470570 449124
rect 470582 449072 470634 449124
rect 470646 449072 470698 449124
rect 470710 449072 470762 449124
rect 470774 449072 470826 449124
rect 470262 449008 470314 449060
rect 470326 449008 470378 449060
rect 470390 449008 470442 449060
rect 470454 449008 470506 449060
rect 470518 449008 470570 449060
rect 470582 449008 470634 449060
rect 470646 449008 470698 449060
rect 470710 449008 470762 449060
rect 470774 449008 470826 449060
rect 478696 446226 478748 446278
rect 515404 445886 515456 445938
rect 482008 445818 482060 445870
rect 485320 445818 485372 445870
rect 523684 445818 523736 445870
rect 520924 445750 520976 445802
rect 475384 445682 475436 445734
rect 535460 445682 535512 445734
rect 546960 445138 547012 445190
rect 547512 445138 547564 445190
rect 490564 442962 490616 443014
rect 535460 442962 535512 443014
rect 493324 441602 493376 441654
rect 535460 441602 535512 441654
rect 494704 440242 494756 440294
rect 535460 440242 535512 440294
rect 496084 438882 496136 438934
rect 535460 438882 535512 438934
rect 497464 437454 497516 437506
rect 535460 437454 535512 437506
rect 498844 436094 498896 436146
rect 535460 436094 535512 436146
rect 500224 434734 500276 434786
rect 535460 434734 535512 434786
rect 501604 433306 501656 433358
rect 535460 433306 535512 433358
rect 470262 433036 470314 433088
rect 470326 433036 470378 433088
rect 470390 433036 470442 433088
rect 470454 433036 470506 433088
rect 470518 433036 470570 433088
rect 470582 433036 470634 433088
rect 470646 433036 470698 433088
rect 470710 433036 470762 433088
rect 470774 433036 470826 433088
rect 470262 432972 470314 433024
rect 470326 432972 470378 433024
rect 470390 432972 470442 433024
rect 470454 432972 470506 433024
rect 470518 432972 470570 433024
rect 470582 432972 470634 433024
rect 470646 432972 470698 433024
rect 470710 432972 470762 433024
rect 470774 432972 470826 433024
rect 470262 432908 470314 432960
rect 470326 432908 470378 432960
rect 470390 432908 470442 432960
rect 470454 432908 470506 432960
rect 470518 432908 470570 432960
rect 470582 432908 470634 432960
rect 470646 432908 470698 432960
rect 470710 432908 470762 432960
rect 470774 432908 470826 432960
rect 470262 432844 470314 432896
rect 470326 432844 470378 432896
rect 470390 432844 470442 432896
rect 470454 432844 470506 432896
rect 470518 432844 470570 432896
rect 470582 432844 470634 432896
rect 470646 432844 470698 432896
rect 470710 432844 470762 432896
rect 470774 432844 470826 432896
rect 470262 432780 470314 432832
rect 470326 432780 470378 432832
rect 470390 432780 470442 432832
rect 470454 432780 470506 432832
rect 470518 432780 470570 432832
rect 470582 432780 470634 432832
rect 470646 432780 470698 432832
rect 470710 432780 470762 432832
rect 470774 432780 470826 432832
rect 471612 432240 471664 432292
rect 577022 432252 577074 432304
rect 577086 432252 577138 432304
rect 577150 432252 577202 432304
rect 577214 432252 577266 432304
rect 577278 432252 577330 432304
rect 577342 432252 577394 432304
rect 577406 432252 577458 432304
rect 577470 432252 577522 432304
rect 577534 432252 577586 432304
rect 577022 432188 577074 432240
rect 577086 432188 577138 432240
rect 577150 432188 577202 432240
rect 577214 432188 577266 432240
rect 577278 432188 577330 432240
rect 577342 432188 577394 432240
rect 577406 432188 577458 432240
rect 577470 432188 577522 432240
rect 577534 432188 577586 432240
rect 577022 432124 577074 432176
rect 577086 432124 577138 432176
rect 577150 432124 577202 432176
rect 577214 432124 577266 432176
rect 577278 432124 577330 432176
rect 577342 432124 577394 432176
rect 577406 432124 577458 432176
rect 577470 432124 577522 432176
rect 577534 432124 577586 432176
rect 577022 432060 577074 432112
rect 577086 432060 577138 432112
rect 577150 432060 577202 432112
rect 577214 432060 577266 432112
rect 577278 432060 577330 432112
rect 577342 432060 577394 432112
rect 577406 432060 577458 432112
rect 577470 432060 577522 432112
rect 577534 432060 577586 432112
rect 469022 431949 469074 432001
rect 469086 431949 469138 432001
rect 469150 431949 469202 432001
rect 469214 431949 469266 432001
rect 469278 431949 469330 432001
rect 469342 431949 469394 432001
rect 469406 431949 469458 432001
rect 469470 431949 469522 432001
rect 469534 431949 469586 432001
rect 502984 431946 503036 431998
rect 535460 431946 535512 431998
rect 577022 431996 577074 432048
rect 577086 431996 577138 432048
rect 577150 431996 577202 432048
rect 577214 431996 577266 432048
rect 577278 431996 577330 432048
rect 577342 431996 577394 432048
rect 577406 431996 577458 432048
rect 577470 431996 577522 432048
rect 577534 431996 577586 432048
rect 469022 431885 469074 431937
rect 469086 431885 469138 431937
rect 469150 431885 469202 431937
rect 469214 431885 469266 431937
rect 469278 431885 469330 431937
rect 469342 431885 469394 431937
rect 469406 431885 469458 431937
rect 469470 431885 469522 431937
rect 469534 431885 469586 431937
rect 469022 431821 469074 431873
rect 469086 431821 469138 431873
rect 469150 431821 469202 431873
rect 469214 431821 469266 431873
rect 469278 431821 469330 431873
rect 469342 431821 469394 431873
rect 469406 431821 469458 431873
rect 469470 431821 469522 431873
rect 469534 431821 469586 431873
rect 469022 431757 469074 431809
rect 469086 431757 469138 431809
rect 469150 431757 469202 431809
rect 469214 431757 469266 431809
rect 469278 431757 469330 431809
rect 469342 431757 469394 431809
rect 469406 431757 469458 431809
rect 469470 431757 469522 431809
rect 469534 431757 469586 431809
rect 469022 431693 469074 431745
rect 469086 431693 469138 431745
rect 469150 431693 469202 431745
rect 469214 431693 469266 431745
rect 469278 431693 469330 431745
rect 469342 431693 469394 431745
rect 469406 431693 469458 431745
rect 469470 431693 469522 431745
rect 469534 431693 469586 431745
rect 576603 431613 576655 431622
rect 576603 431579 576613 431613
rect 576613 431579 576647 431613
rect 576647 431579 576655 431613
rect 576603 431570 576655 431579
rect 578262 431457 578314 431509
rect 578326 431457 578378 431509
rect 578390 431457 578442 431509
rect 578454 431457 578506 431509
rect 578518 431457 578570 431509
rect 578582 431457 578634 431509
rect 578646 431457 578698 431509
rect 578710 431457 578762 431509
rect 578774 431457 578826 431509
rect 478972 431445 479024 431454
rect 478972 431411 478977 431445
rect 478977 431411 479024 431445
rect 478972 431402 479024 431411
rect 485780 431445 485832 431454
rect 485780 431411 485831 431445
rect 485831 431411 485832 431445
rect 485780 431402 485832 431411
rect 578262 431393 578314 431445
rect 578326 431393 578378 431445
rect 578390 431393 578442 431445
rect 578454 431393 578506 431445
rect 578518 431393 578570 431445
rect 578582 431393 578634 431445
rect 578646 431393 578698 431445
rect 578710 431393 578762 431445
rect 578774 431393 578826 431445
rect 578262 431329 578314 431381
rect 578326 431329 578378 431381
rect 578390 431329 578442 431381
rect 578454 431329 578506 431381
rect 578518 431329 578570 431381
rect 578582 431329 578634 431381
rect 578646 431329 578698 431381
rect 578710 431329 578762 431381
rect 578774 431329 578826 431381
rect 578262 431265 578314 431317
rect 578326 431265 578378 431317
rect 578390 431265 578442 431317
rect 578454 431265 578506 431317
rect 578518 431265 578570 431317
rect 578582 431265 578634 431317
rect 578646 431265 578698 431317
rect 578710 431265 578762 431317
rect 578774 431265 578826 431317
rect 578262 431201 578314 431253
rect 578326 431201 578378 431253
rect 578390 431201 578442 431253
rect 578454 431201 578506 431253
rect 578518 431201 578570 431253
rect 578582 431201 578634 431253
rect 578646 431201 578698 431253
rect 578710 431201 578762 431253
rect 578774 431201 578826 431253
rect 475476 431037 475528 431089
rect 482376 431037 482428 431089
rect 492036 430994 492088 431046
rect 470262 430864 470314 430916
rect 470326 430864 470378 430916
rect 470390 430864 470442 430916
rect 470454 430864 470506 430916
rect 470518 430864 470570 430916
rect 470582 430864 470634 430916
rect 470646 430864 470698 430916
rect 470710 430864 470762 430916
rect 470774 430864 470826 430916
rect 470262 430800 470314 430852
rect 470326 430800 470378 430852
rect 470390 430800 470442 430852
rect 470454 430800 470506 430852
rect 470518 430800 470570 430852
rect 470582 430800 470634 430852
rect 470646 430800 470698 430852
rect 470710 430800 470762 430852
rect 470774 430800 470826 430852
rect 470262 430736 470314 430788
rect 470326 430736 470378 430788
rect 470390 430736 470442 430788
rect 470454 430736 470506 430788
rect 470518 430736 470570 430788
rect 470582 430736 470634 430788
rect 470646 430736 470698 430788
rect 470710 430736 470762 430788
rect 470774 430736 470826 430788
rect 470262 430672 470314 430724
rect 470326 430672 470378 430724
rect 470390 430672 470442 430724
rect 470454 430672 470506 430724
rect 470518 430672 470570 430724
rect 470582 430672 470634 430724
rect 470646 430672 470698 430724
rect 470710 430672 470762 430724
rect 470774 430672 470826 430724
rect 470262 430608 470314 430660
rect 470326 430608 470378 430660
rect 470390 430608 470442 430660
rect 470454 430608 470506 430660
rect 470518 430608 470570 430660
rect 470582 430608 470634 430660
rect 470646 430608 470698 430660
rect 470710 430608 470762 430660
rect 470774 430608 470826 430660
rect 475476 429090 475528 429142
rect 490564 429090 490616 429142
rect 482376 427798 482428 427850
rect 522304 427798 522356 427850
rect 470262 412036 470314 412088
rect 470326 412036 470378 412088
rect 470390 412036 470442 412088
rect 470454 412036 470506 412088
rect 470518 412036 470570 412088
rect 470582 412036 470634 412088
rect 470646 412036 470698 412088
rect 470710 412036 470762 412088
rect 470774 412036 470826 412088
rect 470262 411972 470314 412024
rect 470326 411972 470378 412024
rect 470390 411972 470442 412024
rect 470454 411972 470506 412024
rect 470518 411972 470570 412024
rect 470582 411972 470634 412024
rect 470646 411972 470698 412024
rect 470710 411972 470762 412024
rect 470774 411972 470826 412024
rect 470262 411908 470314 411960
rect 470326 411908 470378 411960
rect 470390 411908 470442 411960
rect 470454 411908 470506 411960
rect 470518 411908 470570 411960
rect 470582 411908 470634 411960
rect 470646 411908 470698 411960
rect 470710 411908 470762 411960
rect 470774 411908 470826 411960
rect 470262 411844 470314 411896
rect 470326 411844 470378 411896
rect 470390 411844 470442 411896
rect 470454 411844 470506 411896
rect 470518 411844 470570 411896
rect 470582 411844 470634 411896
rect 470646 411844 470698 411896
rect 470710 411844 470762 411896
rect 470774 411844 470826 411896
rect 470262 411780 470314 411832
rect 470326 411780 470378 411832
rect 470390 411780 470442 411832
rect 470454 411780 470506 411832
rect 470518 411780 470570 411832
rect 470582 411780 470634 411832
rect 470646 411780 470698 411832
rect 470710 411780 470762 411832
rect 470774 411780 470826 411832
rect 471244 411206 471296 411258
rect 473728 411234 473780 411286
rect 469022 410950 469074 411002
rect 469086 410950 469138 411002
rect 469150 410950 469202 411002
rect 469214 410950 469266 411002
rect 469278 410950 469330 411002
rect 469342 410950 469394 411002
rect 469406 410950 469458 411002
rect 469470 410950 469522 411002
rect 469534 410950 469586 411002
rect 469022 410886 469074 410938
rect 469086 410886 469138 410938
rect 469150 410886 469202 410938
rect 469214 410886 469266 410938
rect 469278 410886 469330 410938
rect 469342 410886 469394 410938
rect 469406 410886 469458 410938
rect 469470 410886 469522 410938
rect 469534 410886 469586 410938
rect 469022 410822 469074 410874
rect 469086 410822 469138 410874
rect 469150 410822 469202 410874
rect 469214 410822 469266 410874
rect 469278 410822 469330 410874
rect 469342 410822 469394 410874
rect 469406 410822 469458 410874
rect 469470 410822 469522 410874
rect 469534 410822 469586 410874
rect 469022 410758 469074 410810
rect 469086 410758 469138 410810
rect 469150 410758 469202 410810
rect 469214 410758 469266 410810
rect 469278 410758 469330 410810
rect 469342 410758 469394 410810
rect 469406 410758 469458 410810
rect 469470 410758 469522 410810
rect 469534 410758 469586 410810
rect 469022 410694 469074 410746
rect 469086 410694 469138 410746
rect 469150 410694 469202 410746
rect 469214 410694 469266 410746
rect 469278 410694 469330 410746
rect 469342 410694 469394 410746
rect 469406 410694 469458 410746
rect 469470 410694 469522 410746
rect 469534 410694 469586 410746
rect 478420 410390 478472 410442
rect 478604 410433 478656 410442
rect 478604 410399 478615 410433
rect 478615 410399 478656 410433
rect 478604 410390 478656 410399
rect 485136 410433 485188 410442
rect 485136 410399 485145 410433
rect 485145 410399 485188 410433
rect 485136 410390 485188 410399
rect 475292 410038 475344 410090
rect 481824 410038 481876 410090
rect 490748 409982 490800 410034
rect 470262 409864 470314 409916
rect 470326 409864 470378 409916
rect 470390 409864 470442 409916
rect 470454 409864 470506 409916
rect 470518 409864 470570 409916
rect 470582 409864 470634 409916
rect 470646 409864 470698 409916
rect 470710 409864 470762 409916
rect 470774 409864 470826 409916
rect 470262 409800 470314 409852
rect 470326 409800 470378 409852
rect 470390 409800 470442 409852
rect 470454 409800 470506 409852
rect 470518 409800 470570 409852
rect 470582 409800 470634 409852
rect 470646 409800 470698 409852
rect 470710 409800 470762 409852
rect 470774 409800 470826 409852
rect 470262 409736 470314 409788
rect 470326 409736 470378 409788
rect 470390 409736 470442 409788
rect 470454 409736 470506 409788
rect 470518 409736 470570 409788
rect 470582 409736 470634 409788
rect 470646 409736 470698 409788
rect 470710 409736 470762 409788
rect 470774 409736 470826 409788
rect 515404 409778 515456 409830
rect 535460 409778 535512 409830
rect 470262 409672 470314 409724
rect 470326 409672 470378 409724
rect 470390 409672 470442 409724
rect 470454 409672 470506 409724
rect 470518 409672 470570 409724
rect 470582 409672 470634 409724
rect 470646 409672 470698 409724
rect 470710 409672 470762 409724
rect 470774 409672 470826 409724
rect 470262 409608 470314 409660
rect 470326 409608 470378 409660
rect 470390 409608 470442 409660
rect 470454 409608 470506 409660
rect 470518 409608 470570 409660
rect 470582 409608 470634 409660
rect 470646 409608 470698 409660
rect 470710 409608 470762 409660
rect 470774 409608 470826 409660
rect 475292 408418 475344 408470
rect 493324 408418 493376 408470
rect 547236 408146 547288 408198
rect 547512 408146 547564 408198
rect 478604 407058 478656 407110
rect 535460 407058 535512 407110
rect 515404 404338 515456 404390
rect 535460 404338 535512 404390
rect 516784 402978 516836 403030
rect 535460 402978 535512 403030
rect 518164 398830 518216 398882
rect 535460 398830 535512 398882
rect 519544 396042 519596 396094
rect 535460 396042 535512 396094
rect 470262 391037 470314 391089
rect 470326 391037 470378 391089
rect 470390 391037 470442 391089
rect 470454 391037 470506 391089
rect 470518 391037 470570 391089
rect 470582 391037 470634 391089
rect 470646 391037 470698 391089
rect 470710 391037 470762 391089
rect 470774 391037 470826 391089
rect 470262 390973 470314 391025
rect 470326 390973 470378 391025
rect 470390 390973 470442 391025
rect 470454 390973 470506 391025
rect 470518 390973 470570 391025
rect 470582 390973 470634 391025
rect 470646 390973 470698 391025
rect 470710 390973 470762 391025
rect 470774 390973 470826 391025
rect 470262 390909 470314 390961
rect 470326 390909 470378 390961
rect 470390 390909 470442 390961
rect 470454 390909 470506 390961
rect 470518 390909 470570 390961
rect 470582 390909 470634 390961
rect 470646 390909 470698 390961
rect 470710 390909 470762 390961
rect 470774 390909 470826 390961
rect 470262 390845 470314 390897
rect 470326 390845 470378 390897
rect 470390 390845 470442 390897
rect 470454 390845 470506 390897
rect 470518 390845 470570 390897
rect 470582 390845 470634 390897
rect 470646 390845 470698 390897
rect 470710 390845 470762 390897
rect 470774 390845 470826 390897
rect 470262 390781 470314 390833
rect 470326 390781 470378 390833
rect 470390 390781 470442 390833
rect 470454 390781 470506 390833
rect 470518 390781 470570 390833
rect 470582 390781 470634 390833
rect 470646 390781 470698 390833
rect 470710 390781 470762 390833
rect 470774 390781 470826 390833
rect 471244 390262 471296 390314
rect 471704 390058 471756 390110
rect 469022 389954 469074 390006
rect 469086 389954 469138 390006
rect 469150 389954 469202 390006
rect 469214 389954 469266 390006
rect 469278 389954 469330 390006
rect 469342 389954 469394 390006
rect 469406 389954 469458 390006
rect 469470 389954 469522 390006
rect 469534 389954 469586 390006
rect 469022 389890 469074 389942
rect 469086 389890 469138 389942
rect 469150 389890 469202 389942
rect 469214 389890 469266 389942
rect 469278 389890 469330 389942
rect 469342 389890 469394 389942
rect 469406 389890 469458 389942
rect 469470 389890 469522 389942
rect 469534 389890 469586 389942
rect 469022 389826 469074 389878
rect 469086 389826 469138 389878
rect 469150 389826 469202 389878
rect 469214 389826 469266 389878
rect 469278 389826 469330 389878
rect 469342 389826 469394 389878
rect 469406 389826 469458 389878
rect 469470 389826 469522 389878
rect 469534 389826 469586 389878
rect 469022 389762 469074 389814
rect 469086 389762 469138 389814
rect 469150 389762 469202 389814
rect 469214 389762 469266 389814
rect 469278 389762 469330 389814
rect 469342 389762 469394 389814
rect 469406 389762 469458 389814
rect 469470 389762 469522 389814
rect 469534 389762 469586 389814
rect 469022 389698 469074 389750
rect 469086 389698 469138 389750
rect 469150 389698 469202 389750
rect 469214 389698 469266 389750
rect 469278 389698 469330 389750
rect 469342 389698 469394 389750
rect 469406 389698 469458 389750
rect 469470 389698 469522 389750
rect 469534 389698 469586 389750
rect 479432 389489 479484 389498
rect 479432 389455 479474 389489
rect 479474 389455 479484 389489
rect 479432 389446 479484 389455
rect 493324 389446 493376 389498
rect 475752 389038 475804 389090
rect 483204 389038 483256 389090
rect 486884 389038 486936 389090
rect 470262 388864 470314 388916
rect 470326 388864 470378 388916
rect 470390 388864 470442 388916
rect 470454 388864 470506 388916
rect 470518 388864 470570 388916
rect 470582 388864 470634 388916
rect 470646 388864 470698 388916
rect 470710 388864 470762 388916
rect 470774 388864 470826 388916
rect 470262 388800 470314 388852
rect 470326 388800 470378 388852
rect 470390 388800 470442 388852
rect 470454 388800 470506 388852
rect 470518 388800 470570 388852
rect 470582 388800 470634 388852
rect 470646 388800 470698 388852
rect 470710 388800 470762 388852
rect 470774 388800 470826 388852
rect 470262 388736 470314 388788
rect 470326 388736 470378 388788
rect 470390 388736 470442 388788
rect 470454 388736 470506 388788
rect 470518 388736 470570 388788
rect 470582 388736 470634 388788
rect 470646 388736 470698 388788
rect 470710 388736 470762 388788
rect 470774 388736 470826 388788
rect 470262 388672 470314 388724
rect 470326 388672 470378 388724
rect 470390 388672 470442 388724
rect 470454 388672 470506 388724
rect 470518 388672 470570 388724
rect 470582 388672 470634 388724
rect 470646 388672 470698 388724
rect 470710 388672 470762 388724
rect 470774 388672 470826 388724
rect 470262 388608 470314 388660
rect 470326 388608 470378 388660
rect 470390 388608 470442 388660
rect 470454 388608 470506 388660
rect 470518 388608 470570 388660
rect 470582 388608 470634 388660
rect 470646 388608 470698 388660
rect 470710 388608 470762 388660
rect 470774 388608 470826 388660
rect 475752 387746 475804 387798
rect 479432 387746 479484 387798
rect 515404 387746 515456 387798
rect 494704 387678 494756 387730
rect 483204 386386 483256 386438
rect 484308 386386 484360 386438
rect 577022 379076 577074 379128
rect 577086 379076 577138 379128
rect 577150 379076 577202 379128
rect 577214 379076 577266 379128
rect 577278 379076 577330 379128
rect 577342 379076 577394 379128
rect 577406 379076 577458 379128
rect 577470 379076 577522 379128
rect 577534 379076 577586 379128
rect 577022 379012 577074 379064
rect 577086 379012 577138 379064
rect 577150 379012 577202 379064
rect 577214 379012 577266 379064
rect 577278 379012 577330 379064
rect 577342 379012 577394 379064
rect 577406 379012 577458 379064
rect 577470 379012 577522 379064
rect 577534 379012 577586 379064
rect 577022 378948 577074 379000
rect 577086 378948 577138 379000
rect 577150 378948 577202 379000
rect 577214 378948 577266 379000
rect 577278 378948 577330 379000
rect 577342 378948 577394 379000
rect 577406 378948 577458 379000
rect 577470 378948 577522 379000
rect 577534 378948 577586 379000
rect 577022 378884 577074 378936
rect 577086 378884 577138 378936
rect 577150 378884 577202 378936
rect 577214 378884 577266 378936
rect 577278 378884 577330 378936
rect 577342 378884 577394 378936
rect 577406 378884 577458 378936
rect 577470 378884 577522 378936
rect 577534 378884 577586 378936
rect 577022 378820 577074 378872
rect 577086 378820 577138 378872
rect 577150 378820 577202 378872
rect 577214 378820 577266 378872
rect 577278 378820 577330 378872
rect 577342 378820 577394 378872
rect 577406 378820 577458 378872
rect 577470 378820 577522 378872
rect 577534 378820 577586 378872
rect 576603 378437 576655 378446
rect 576603 378403 576613 378437
rect 576613 378403 576647 378437
rect 576647 378403 576655 378437
rect 576603 378394 576655 378403
rect 578262 378281 578314 378333
rect 578326 378281 578378 378333
rect 578390 378281 578442 378333
rect 578454 378281 578506 378333
rect 578518 378281 578570 378333
rect 578582 378281 578634 378333
rect 578646 378281 578698 378333
rect 578710 378281 578762 378333
rect 578774 378281 578826 378333
rect 578262 378217 578314 378269
rect 578326 378217 578378 378269
rect 578390 378217 578442 378269
rect 578454 378217 578506 378269
rect 578518 378217 578570 378269
rect 578582 378217 578634 378269
rect 578646 378217 578698 378269
rect 578710 378217 578762 378269
rect 578774 378217 578826 378269
rect 578262 378153 578314 378205
rect 578326 378153 578378 378205
rect 578390 378153 578442 378205
rect 578454 378153 578506 378205
rect 578518 378153 578570 378205
rect 578582 378153 578634 378205
rect 578646 378153 578698 378205
rect 578710 378153 578762 378205
rect 578774 378153 578826 378205
rect 578262 378089 578314 378141
rect 578326 378089 578378 378141
rect 578390 378089 578442 378141
rect 578454 378089 578506 378141
rect 578518 378089 578570 378141
rect 578582 378089 578634 378141
rect 578646 378089 578698 378141
rect 578710 378089 578762 378141
rect 578774 378089 578826 378141
rect 578262 378025 578314 378077
rect 578326 378025 578378 378077
rect 578390 378025 578442 378077
rect 578454 378025 578506 378077
rect 578518 378025 578570 378077
rect 578582 378025 578634 378077
rect 578646 378025 578698 378077
rect 578710 378025 578762 378077
rect 578774 378025 578826 378077
rect 520924 373942 520976 373994
rect 535460 373942 535512 373994
rect 547052 373262 547104 373314
rect 547512 373262 547564 373314
rect 522304 372514 522356 372566
rect 535460 372514 535512 372566
rect 484308 369794 484360 369846
rect 535460 369794 535512 369846
rect 520924 367074 520976 367126
rect 535460 367074 535512 367126
rect 515404 365714 515456 365766
rect 535460 365714 535512 365766
rect 522304 361566 522356 361618
rect 535460 361566 535512 361618
rect 470262 358437 470314 358489
rect 470326 358437 470378 358489
rect 470390 358437 470442 358489
rect 470454 358437 470506 358489
rect 470518 358437 470570 358489
rect 470582 358437 470634 358489
rect 470646 358437 470698 358489
rect 470710 358437 470762 358489
rect 470774 358437 470826 358489
rect 470262 358373 470314 358425
rect 470326 358373 470378 358425
rect 470390 358373 470442 358425
rect 470454 358373 470506 358425
rect 470518 358373 470570 358425
rect 470582 358373 470634 358425
rect 470646 358373 470698 358425
rect 470710 358373 470762 358425
rect 470774 358373 470826 358425
rect 470262 358309 470314 358361
rect 470326 358309 470378 358361
rect 470390 358309 470442 358361
rect 470454 358309 470506 358361
rect 470518 358309 470570 358361
rect 470582 358309 470634 358361
rect 470646 358309 470698 358361
rect 470710 358309 470762 358361
rect 470774 358309 470826 358361
rect 470262 358245 470314 358297
rect 470326 358245 470378 358297
rect 470390 358245 470442 358297
rect 470454 358245 470506 358297
rect 470518 358245 470570 358297
rect 470582 358245 470634 358297
rect 470646 358245 470698 358297
rect 470710 358245 470762 358297
rect 470774 358245 470826 358297
rect 470262 358181 470314 358233
rect 470326 358181 470378 358233
rect 470390 358181 470442 358233
rect 470454 358181 470506 358233
rect 470518 358181 470570 358233
rect 470582 358181 470634 358233
rect 470646 358181 470698 358233
rect 470710 358181 470762 358233
rect 470774 358181 470826 358233
rect 471704 357554 471756 357606
rect 475108 357622 475160 357674
rect 478880 357633 478932 357685
rect 481824 357633 481876 357685
rect 484952 357633 485004 357685
rect 469022 357351 469074 357403
rect 469086 357351 469138 357403
rect 469150 357351 469202 357403
rect 469214 357351 469266 357403
rect 469278 357351 469330 357403
rect 469342 357351 469394 357403
rect 469406 357351 469458 357403
rect 469470 357351 469522 357403
rect 469534 357351 469586 357403
rect 469022 357287 469074 357339
rect 469086 357287 469138 357339
rect 469150 357287 469202 357339
rect 469214 357287 469266 357339
rect 469278 357287 469330 357339
rect 469342 357287 469394 357339
rect 469406 357287 469458 357339
rect 469470 357287 469522 357339
rect 469534 357287 469586 357339
rect 469022 357223 469074 357275
rect 469086 357223 469138 357275
rect 469150 357223 469202 357275
rect 469214 357223 469266 357275
rect 469278 357223 469330 357275
rect 469342 357223 469394 357275
rect 469406 357223 469458 357275
rect 469470 357223 469522 357275
rect 469534 357223 469586 357275
rect 469022 357159 469074 357211
rect 469086 357159 469138 357211
rect 469150 357159 469202 357211
rect 469214 357159 469266 357211
rect 469278 357159 469330 357211
rect 469342 357159 469394 357211
rect 469406 357159 469458 357211
rect 469470 357159 469522 357211
rect 469534 357159 469586 357211
rect 469022 357095 469074 357147
rect 469086 357095 469138 357147
rect 469150 357095 469202 357147
rect 469214 357095 469266 357147
rect 469278 357095 469330 357147
rect 469342 357095 469394 357147
rect 469406 357095 469458 357147
rect 469470 357095 469522 357147
rect 469534 357095 469586 357147
rect 477040 356849 477092 356858
rect 477040 356815 477091 356849
rect 477091 356815 477092 356849
rect 477040 356806 477092 356815
rect 480168 356849 480220 356858
rect 480168 356815 480177 356849
rect 480177 356815 480220 356849
rect 480168 356806 480220 356815
rect 483204 356437 483256 356489
rect 486240 356437 486292 356489
rect 492128 356398 492180 356450
rect 470262 356264 470314 356316
rect 470326 356264 470378 356316
rect 470390 356264 470442 356316
rect 470454 356264 470506 356316
rect 470518 356264 470570 356316
rect 470582 356264 470634 356316
rect 470646 356264 470698 356316
rect 470710 356264 470762 356316
rect 470774 356264 470826 356316
rect 470262 356200 470314 356252
rect 470326 356200 470378 356252
rect 470390 356200 470442 356252
rect 470454 356200 470506 356252
rect 470518 356200 470570 356252
rect 470582 356200 470634 356252
rect 470646 356200 470698 356252
rect 470710 356200 470762 356252
rect 470774 356200 470826 356252
rect 470262 356136 470314 356188
rect 470326 356136 470378 356188
rect 470390 356136 470442 356188
rect 470454 356136 470506 356188
rect 470518 356136 470570 356188
rect 470582 356136 470634 356188
rect 470646 356136 470698 356188
rect 470710 356136 470762 356188
rect 470774 356136 470826 356188
rect 470262 356072 470314 356124
rect 470326 356072 470378 356124
rect 470390 356072 470442 356124
rect 470454 356072 470506 356124
rect 470518 356072 470570 356124
rect 470582 356072 470634 356124
rect 470646 356072 470698 356124
rect 470710 356072 470762 356124
rect 470774 356072 470826 356124
rect 470262 356008 470314 356060
rect 470326 356008 470378 356060
rect 470390 356008 470442 356060
rect 470454 356008 470506 356060
rect 470518 356008 470570 356060
rect 470582 356008 470634 356060
rect 470646 356008 470698 356060
rect 470710 356008 470762 356060
rect 470774 356008 470826 356060
rect 483204 354630 483256 354682
rect 520924 354630 520976 354682
rect 480168 354562 480220 354614
rect 516784 354562 516836 354614
rect 477132 354494 477184 354546
rect 496084 354494 496136 354546
rect 486240 353610 486292 353662
rect 525064 353270 525116 353322
rect 547144 344974 547196 345026
rect 547512 344974 547564 345026
rect 470262 342436 470314 342488
rect 470326 342436 470378 342488
rect 470390 342436 470442 342488
rect 470454 342436 470506 342488
rect 470518 342436 470570 342488
rect 470582 342436 470634 342488
rect 470646 342436 470698 342488
rect 470710 342436 470762 342488
rect 470774 342436 470826 342488
rect 470262 342372 470314 342424
rect 470326 342372 470378 342424
rect 470390 342372 470442 342424
rect 470454 342372 470506 342424
rect 470518 342372 470570 342424
rect 470582 342372 470634 342424
rect 470646 342372 470698 342424
rect 470710 342372 470762 342424
rect 470774 342372 470826 342424
rect 470262 342308 470314 342360
rect 470326 342308 470378 342360
rect 470390 342308 470442 342360
rect 470454 342308 470506 342360
rect 470518 342308 470570 342360
rect 470582 342308 470634 342360
rect 470646 342308 470698 342360
rect 470710 342308 470762 342360
rect 470774 342308 470826 342360
rect 470262 342244 470314 342296
rect 470326 342244 470378 342296
rect 470390 342244 470442 342296
rect 470454 342244 470506 342296
rect 470518 342244 470570 342296
rect 470582 342244 470634 342296
rect 470646 342244 470698 342296
rect 470710 342244 470762 342296
rect 470774 342244 470826 342296
rect 470262 342180 470314 342232
rect 470326 342180 470378 342232
rect 470390 342180 470442 342232
rect 470454 342180 470506 342232
rect 470518 342180 470570 342232
rect 470582 342180 470634 342232
rect 470646 342180 470698 342232
rect 470710 342180 470762 342232
rect 470774 342180 470826 342232
rect 471704 341778 471756 341830
rect 471244 341710 471296 341762
rect 469022 341349 469074 341401
rect 469086 341349 469138 341401
rect 469150 341349 469202 341401
rect 469214 341349 469266 341401
rect 469278 341349 469330 341401
rect 469342 341349 469394 341401
rect 469406 341349 469458 341401
rect 469470 341349 469522 341401
rect 469534 341349 469586 341401
rect 469022 341285 469074 341337
rect 469086 341285 469138 341337
rect 469150 341285 469202 341337
rect 469214 341285 469266 341337
rect 469278 341285 469330 341337
rect 469342 341285 469394 341337
rect 469406 341285 469458 341337
rect 469470 341285 469522 341337
rect 469534 341285 469586 341337
rect 469022 341221 469074 341273
rect 469086 341221 469138 341273
rect 469150 341221 469202 341273
rect 469214 341221 469266 341273
rect 469278 341221 469330 341273
rect 469342 341221 469394 341273
rect 469406 341221 469458 341273
rect 469470 341221 469522 341273
rect 469534 341221 469586 341273
rect 469022 341157 469074 341209
rect 469086 341157 469138 341209
rect 469150 341157 469202 341209
rect 469214 341157 469266 341209
rect 469278 341157 469330 341209
rect 469342 341157 469394 341209
rect 469406 341157 469458 341209
rect 469470 341157 469522 341209
rect 469534 341157 469586 341209
rect 469022 341093 469074 341145
rect 469086 341093 469138 341145
rect 469150 341093 469202 341145
rect 469214 341093 469266 341145
rect 469278 341093 469330 341145
rect 469342 341093 469394 341145
rect 469406 341093 469458 341145
rect 469470 341093 469522 341145
rect 469534 341093 469586 341145
rect 484400 340894 484452 340946
rect 482100 340869 482152 340878
rect 474648 340805 474700 340857
rect 482100 340835 482109 340869
rect 482109 340835 482152 340869
rect 482100 340826 482152 340835
rect 484400 340486 484452 340538
rect 485596 340440 485648 340492
rect 475476 340350 475528 340402
rect 478788 340393 478840 340402
rect 478788 340359 478793 340393
rect 478793 340359 478840 340393
rect 478788 340350 478840 340359
rect 492220 340350 492272 340402
rect 470262 340264 470314 340316
rect 470326 340264 470378 340316
rect 470390 340264 470442 340316
rect 470454 340264 470506 340316
rect 470518 340264 470570 340316
rect 470582 340264 470634 340316
rect 470646 340264 470698 340316
rect 470710 340264 470762 340316
rect 470774 340264 470826 340316
rect 470262 340200 470314 340252
rect 470326 340200 470378 340252
rect 470390 340200 470442 340252
rect 470454 340200 470506 340252
rect 470518 340200 470570 340252
rect 470582 340200 470634 340252
rect 470646 340200 470698 340252
rect 470710 340200 470762 340252
rect 470774 340200 470826 340252
rect 470262 340136 470314 340188
rect 470326 340136 470378 340188
rect 470390 340136 470442 340188
rect 470454 340136 470506 340188
rect 470518 340136 470570 340188
rect 470582 340136 470634 340188
rect 470646 340136 470698 340188
rect 470710 340136 470762 340188
rect 470774 340136 470826 340188
rect 470262 340072 470314 340124
rect 470326 340072 470378 340124
rect 470390 340072 470442 340124
rect 470454 340072 470506 340124
rect 470518 340072 470570 340124
rect 470582 340072 470634 340124
rect 470646 340072 470698 340124
rect 470710 340072 470762 340124
rect 470774 340072 470826 340124
rect 470262 340008 470314 340060
rect 470326 340008 470378 340060
rect 470390 340008 470442 340060
rect 470454 340008 470506 340060
rect 470518 340008 470570 340060
rect 470582 340008 470634 340060
rect 470646 340008 470698 340060
rect 470710 340008 470762 340060
rect 470774 340008 470826 340060
rect 475476 339398 475528 339450
rect 478788 339398 478840 339450
rect 536380 339398 536432 339450
rect 482100 339330 482152 339382
rect 515404 339330 515456 339382
rect 497464 339262 497516 339314
rect 523684 338038 523736 338090
rect 535460 338038 535512 338090
rect 546960 337698 547012 337750
rect 547512 337698 547564 337750
rect 525064 332530 525116 332582
rect 535460 332530 535512 332582
rect 485688 331170 485740 331222
rect 535460 331170 535512 331222
rect 577022 325900 577074 325952
rect 577086 325900 577138 325952
rect 577150 325900 577202 325952
rect 577214 325900 577266 325952
rect 577278 325900 577330 325952
rect 577342 325900 577394 325952
rect 577406 325900 577458 325952
rect 577470 325900 577522 325952
rect 577534 325900 577586 325952
rect 577022 325836 577074 325888
rect 577086 325836 577138 325888
rect 577150 325836 577202 325888
rect 577214 325836 577266 325888
rect 577278 325836 577330 325888
rect 577342 325836 577394 325888
rect 577406 325836 577458 325888
rect 577470 325836 577522 325888
rect 577534 325836 577586 325888
rect 577022 325772 577074 325824
rect 577086 325772 577138 325824
rect 577150 325772 577202 325824
rect 577214 325772 577266 325824
rect 577278 325772 577330 325824
rect 577342 325772 577394 325824
rect 577406 325772 577458 325824
rect 577470 325772 577522 325824
rect 577534 325772 577586 325824
rect 523684 325662 523736 325714
rect 535460 325662 535512 325714
rect 577022 325708 577074 325760
rect 577086 325708 577138 325760
rect 577150 325708 577202 325760
rect 577214 325708 577266 325760
rect 577278 325708 577330 325760
rect 577342 325708 577394 325760
rect 577406 325708 577458 325760
rect 577470 325708 577522 325760
rect 577534 325708 577586 325760
rect 577022 325644 577074 325696
rect 577086 325644 577138 325696
rect 577150 325644 577202 325696
rect 577214 325644 577266 325696
rect 577278 325644 577330 325696
rect 577342 325644 577394 325696
rect 577406 325644 577458 325696
rect 577470 325644 577522 325696
rect 577534 325644 577586 325696
rect 576603 325261 576655 325270
rect 576603 325227 576613 325261
rect 576613 325227 576647 325261
rect 576647 325227 576655 325261
rect 576603 325218 576655 325227
rect 578262 325105 578314 325157
rect 578326 325105 578378 325157
rect 578390 325105 578442 325157
rect 578454 325105 578506 325157
rect 578518 325105 578570 325157
rect 578582 325105 578634 325157
rect 578646 325105 578698 325157
rect 578710 325105 578762 325157
rect 578774 325105 578826 325157
rect 578262 325041 578314 325093
rect 578326 325041 578378 325093
rect 578390 325041 578442 325093
rect 578454 325041 578506 325093
rect 578518 325041 578570 325093
rect 578582 325041 578634 325093
rect 578646 325041 578698 325093
rect 578710 325041 578762 325093
rect 578774 325041 578826 325093
rect 578262 324977 578314 325029
rect 578326 324977 578378 325029
rect 578390 324977 578442 325029
rect 578454 324977 578506 325029
rect 578518 324977 578570 325029
rect 578582 324977 578634 325029
rect 578646 324977 578698 325029
rect 578710 324977 578762 325029
rect 578774 324977 578826 325029
rect 578262 324913 578314 324965
rect 578326 324913 578378 324965
rect 578390 324913 578442 324965
rect 578454 324913 578506 324965
rect 578518 324913 578570 324965
rect 578582 324913 578634 324965
rect 578646 324913 578698 324965
rect 578710 324913 578762 324965
rect 578774 324913 578826 324965
rect 578262 324849 578314 324901
rect 578326 324849 578378 324901
rect 578390 324849 578442 324901
rect 578454 324849 578506 324901
rect 578518 324849 578570 324901
rect 578582 324849 578634 324901
rect 578646 324849 578698 324901
rect 578710 324849 578762 324901
rect 578774 324849 578826 324901
rect 470262 322436 470314 322488
rect 470326 322436 470378 322488
rect 470390 322436 470442 322488
rect 470454 322436 470506 322488
rect 470518 322436 470570 322488
rect 470582 322436 470634 322488
rect 470646 322436 470698 322488
rect 470710 322436 470762 322488
rect 470774 322436 470826 322488
rect 470262 322372 470314 322424
rect 470326 322372 470378 322424
rect 470390 322372 470442 322424
rect 470454 322372 470506 322424
rect 470518 322372 470570 322424
rect 470582 322372 470634 322424
rect 470646 322372 470698 322424
rect 470710 322372 470762 322424
rect 470774 322372 470826 322424
rect 470262 322308 470314 322360
rect 470326 322308 470378 322360
rect 470390 322308 470442 322360
rect 470454 322308 470506 322360
rect 470518 322308 470570 322360
rect 470582 322308 470634 322360
rect 470646 322308 470698 322360
rect 470710 322308 470762 322360
rect 470774 322308 470826 322360
rect 470262 322244 470314 322296
rect 470326 322244 470378 322296
rect 470390 322244 470442 322296
rect 470454 322244 470506 322296
rect 470518 322244 470570 322296
rect 470582 322244 470634 322296
rect 470646 322244 470698 322296
rect 470710 322244 470762 322296
rect 470774 322244 470826 322296
rect 470262 322180 470314 322232
rect 470326 322180 470378 322232
rect 470390 322180 470442 322232
rect 470454 322180 470506 322232
rect 470518 322180 470570 322232
rect 470582 322180 470634 322232
rect 470646 322180 470698 322232
rect 470710 322180 470762 322232
rect 470774 322180 470826 322232
rect 471244 321582 471296 321634
rect 469022 321349 469074 321401
rect 469086 321349 469138 321401
rect 469150 321349 469202 321401
rect 469214 321349 469266 321401
rect 469278 321349 469330 321401
rect 469342 321349 469394 321401
rect 469406 321349 469458 321401
rect 469470 321349 469522 321401
rect 469534 321349 469586 321401
rect 469022 321285 469074 321337
rect 469086 321285 469138 321337
rect 469150 321285 469202 321337
rect 469214 321285 469266 321337
rect 469278 321285 469330 321337
rect 469342 321285 469394 321337
rect 469406 321285 469458 321337
rect 469470 321285 469522 321337
rect 469534 321285 469586 321337
rect 469022 321221 469074 321273
rect 469086 321221 469138 321273
rect 469150 321221 469202 321273
rect 469214 321221 469266 321273
rect 469278 321221 469330 321273
rect 469342 321221 469394 321273
rect 469406 321221 469458 321273
rect 469470 321221 469522 321273
rect 469534 321221 469586 321273
rect 469022 321157 469074 321209
rect 469086 321157 469138 321209
rect 469150 321157 469202 321209
rect 469214 321157 469266 321209
rect 469278 321157 469330 321209
rect 469342 321157 469394 321209
rect 469406 321157 469458 321209
rect 469470 321157 469522 321209
rect 469534 321157 469586 321209
rect 469022 321093 469074 321145
rect 469086 321093 469138 321145
rect 469150 321093 469202 321145
rect 469214 321093 469266 321145
rect 469278 321093 469330 321145
rect 469342 321093 469394 321145
rect 469406 321093 469458 321145
rect 469470 321093 469522 321145
rect 469534 321093 469586 321145
rect 475476 320437 475528 320489
rect 482376 320426 482428 320478
rect 479064 320358 479116 320410
rect 485964 320358 486016 320410
rect 492312 320358 492364 320410
rect 470262 320264 470314 320316
rect 470326 320264 470378 320316
rect 470390 320264 470442 320316
rect 470454 320264 470506 320316
rect 470518 320264 470570 320316
rect 470582 320264 470634 320316
rect 470646 320264 470698 320316
rect 470710 320264 470762 320316
rect 470774 320264 470826 320316
rect 470262 320200 470314 320252
rect 470326 320200 470378 320252
rect 470390 320200 470442 320252
rect 470454 320200 470506 320252
rect 470518 320200 470570 320252
rect 470582 320200 470634 320252
rect 470646 320200 470698 320252
rect 470710 320200 470762 320252
rect 470774 320200 470826 320252
rect 470262 320136 470314 320188
rect 470326 320136 470378 320188
rect 470390 320136 470442 320188
rect 470454 320136 470506 320188
rect 470518 320136 470570 320188
rect 470582 320136 470634 320188
rect 470646 320136 470698 320188
rect 470710 320136 470762 320188
rect 470774 320136 470826 320188
rect 470262 320072 470314 320124
rect 470326 320072 470378 320124
rect 470390 320072 470442 320124
rect 470454 320072 470506 320124
rect 470518 320072 470570 320124
rect 470582 320072 470634 320124
rect 470646 320072 470698 320124
rect 470710 320072 470762 320124
rect 470774 320072 470826 320124
rect 470262 320008 470314 320060
rect 470326 320008 470378 320060
rect 470390 320008 470442 320060
rect 470454 320008 470506 320060
rect 470518 320008 470570 320060
rect 470582 320008 470634 320060
rect 470646 320008 470698 320060
rect 470710 320008 470762 320060
rect 470774 320008 470826 320060
rect 475476 318726 475528 318778
rect 479064 318726 479116 318778
rect 536288 318726 536340 318778
rect 482376 318658 482428 318710
rect 536564 318658 536616 318710
rect 485964 318590 486016 318642
rect 536012 318590 536064 318642
rect 498844 318522 498896 318574
rect 470262 307036 470314 307088
rect 470326 307036 470378 307088
rect 470390 307036 470442 307088
rect 470454 307036 470506 307088
rect 470518 307036 470570 307088
rect 470582 307036 470634 307088
rect 470646 307036 470698 307088
rect 470710 307036 470762 307088
rect 470774 307036 470826 307088
rect 470262 306972 470314 307024
rect 470326 306972 470378 307024
rect 470390 306972 470442 307024
rect 470454 306972 470506 307024
rect 470518 306972 470570 307024
rect 470582 306972 470634 307024
rect 470646 306972 470698 307024
rect 470710 306972 470762 307024
rect 470774 306972 470826 307024
rect 470262 306908 470314 306960
rect 470326 306908 470378 306960
rect 470390 306908 470442 306960
rect 470454 306908 470506 306960
rect 470518 306908 470570 306960
rect 470582 306908 470634 306960
rect 470646 306908 470698 306960
rect 470710 306908 470762 306960
rect 470774 306908 470826 306960
rect 470262 306844 470314 306896
rect 470326 306844 470378 306896
rect 470390 306844 470442 306896
rect 470454 306844 470506 306896
rect 470518 306844 470570 306896
rect 470582 306844 470634 306896
rect 470646 306844 470698 306896
rect 470710 306844 470762 306896
rect 470774 306844 470826 306896
rect 470262 306780 470314 306832
rect 470326 306780 470378 306832
rect 470390 306780 470442 306832
rect 470454 306780 470506 306832
rect 470518 306780 470570 306832
rect 470582 306780 470634 306832
rect 470646 306780 470698 306832
rect 470710 306780 470762 306832
rect 470774 306780 470826 306832
rect 471244 306282 471296 306334
rect 473728 306234 473780 306286
rect 469022 305951 469074 306003
rect 469086 305951 469138 306003
rect 469150 305951 469202 306003
rect 469214 305951 469266 306003
rect 469278 305951 469330 306003
rect 469342 305951 469394 306003
rect 469406 305951 469458 306003
rect 469470 305951 469522 306003
rect 469534 305951 469586 306003
rect 469022 305887 469074 305939
rect 469086 305887 469138 305939
rect 469150 305887 469202 305939
rect 469214 305887 469266 305939
rect 469278 305887 469330 305939
rect 469342 305887 469394 305939
rect 469406 305887 469458 305939
rect 469470 305887 469522 305939
rect 469534 305887 469586 305939
rect 469022 305823 469074 305875
rect 469086 305823 469138 305875
rect 469150 305823 469202 305875
rect 469214 305823 469266 305875
rect 469278 305823 469330 305875
rect 469342 305823 469394 305875
rect 469406 305823 469458 305875
rect 469470 305823 469522 305875
rect 469534 305823 469586 305875
rect 469022 305759 469074 305811
rect 469086 305759 469138 305811
rect 469150 305759 469202 305811
rect 469214 305759 469266 305811
rect 469278 305759 469330 305811
rect 469342 305759 469394 305811
rect 469406 305759 469458 305811
rect 469470 305759 469522 305811
rect 469534 305759 469586 305811
rect 469022 305695 469074 305747
rect 469086 305695 469138 305747
rect 469150 305695 469202 305747
rect 469214 305695 469266 305747
rect 469278 305695 469330 305747
rect 469342 305695 469394 305747
rect 469406 305695 469458 305747
rect 469470 305695 469522 305747
rect 469534 305695 469586 305747
rect 478604 305441 478656 305450
rect 478604 305407 478614 305441
rect 478614 305407 478656 305441
rect 478604 305398 478656 305407
rect 485136 305441 485188 305450
rect 485136 305407 485144 305441
rect 485144 305407 485188 305441
rect 485136 305398 485188 305407
rect 475292 305038 475344 305090
rect 481824 305038 481876 305090
rect 490564 304990 490616 305042
rect 470262 304864 470314 304916
rect 470326 304864 470378 304916
rect 470390 304864 470442 304916
rect 470454 304864 470506 304916
rect 470518 304864 470570 304916
rect 470582 304864 470634 304916
rect 470646 304864 470698 304916
rect 470710 304864 470762 304916
rect 470774 304864 470826 304916
rect 470262 304800 470314 304852
rect 470326 304800 470378 304852
rect 470390 304800 470442 304852
rect 470454 304800 470506 304852
rect 470518 304800 470570 304852
rect 470582 304800 470634 304852
rect 470646 304800 470698 304852
rect 470710 304800 470762 304852
rect 470774 304800 470826 304852
rect 470262 304736 470314 304788
rect 470326 304736 470378 304788
rect 470390 304736 470442 304788
rect 470454 304736 470506 304788
rect 470518 304736 470570 304788
rect 470582 304736 470634 304788
rect 470646 304736 470698 304788
rect 470710 304736 470762 304788
rect 470774 304736 470826 304788
rect 470262 304672 470314 304724
rect 470326 304672 470378 304724
rect 470390 304672 470442 304724
rect 470454 304672 470506 304724
rect 470518 304672 470570 304724
rect 470582 304672 470634 304724
rect 470646 304672 470698 304724
rect 470710 304672 470762 304724
rect 470774 304672 470826 304724
rect 470262 304608 470314 304660
rect 470326 304608 470378 304660
rect 470390 304608 470442 304660
rect 470454 304608 470506 304660
rect 470518 304608 470570 304660
rect 470582 304608 470634 304660
rect 470646 304608 470698 304660
rect 470710 304608 470762 304660
rect 470774 304608 470826 304660
rect 547052 303698 547104 303750
rect 547512 303698 547564 303750
rect 475292 303562 475344 303614
rect 478604 303562 478656 303614
rect 481824 303562 481876 303614
rect 485136 303562 485188 303614
rect 536472 303562 536524 303614
rect 536656 303494 536708 303546
rect 518164 303426 518216 303478
rect 500224 303358 500276 303410
rect 491944 300774 491996 300826
rect 535460 300774 535512 300826
rect 492036 299414 492088 299466
rect 535460 299414 535512 299466
rect 490748 298054 490800 298106
rect 535460 298054 535512 298106
rect 492128 296626 492180 296678
rect 535552 296626 535604 296678
rect 493324 296558 493376 296610
rect 535460 296558 535512 296610
rect 492220 295266 492272 295318
rect 535460 295266 535512 295318
rect 492312 293906 492364 293958
rect 535552 293906 535604 293958
rect 490564 292478 490616 292530
rect 535460 292478 535512 292530
rect 492956 289826 493008 289878
rect 535460 289826 535512 289878
rect 491944 288398 491996 288450
rect 535460 288398 535512 288450
rect 470262 287437 470314 287489
rect 470326 287437 470378 287489
rect 470390 287437 470442 287489
rect 470454 287437 470506 287489
rect 470518 287437 470570 287489
rect 470582 287437 470634 287489
rect 470646 287437 470698 287489
rect 470710 287437 470762 287489
rect 470774 287437 470826 287489
rect 470262 287373 470314 287425
rect 470326 287373 470378 287425
rect 470390 287373 470442 287425
rect 470454 287373 470506 287425
rect 470518 287373 470570 287425
rect 470582 287373 470634 287425
rect 470646 287373 470698 287425
rect 470710 287373 470762 287425
rect 470774 287373 470826 287425
rect 470262 287309 470314 287361
rect 470326 287309 470378 287361
rect 470390 287309 470442 287361
rect 470454 287309 470506 287361
rect 470518 287309 470570 287361
rect 470582 287309 470634 287361
rect 470646 287309 470698 287361
rect 470710 287309 470762 287361
rect 470774 287309 470826 287361
rect 470262 287245 470314 287297
rect 470326 287245 470378 287297
rect 470390 287245 470442 287297
rect 470454 287245 470506 287297
rect 470518 287245 470570 287297
rect 470582 287245 470634 287297
rect 470646 287245 470698 287297
rect 470710 287245 470762 287297
rect 470774 287245 470826 287297
rect 470262 287181 470314 287233
rect 470326 287181 470378 287233
rect 470390 287181 470442 287233
rect 470454 287181 470506 287233
rect 470518 287181 470570 287233
rect 470582 287181 470634 287233
rect 470646 287181 470698 287233
rect 470710 287181 470762 287233
rect 470774 287181 470826 287233
rect 471244 286630 471296 286682
rect 484952 286630 485004 286682
rect 488632 286630 488684 286682
rect 471704 286494 471756 286546
rect 469022 286352 469074 286404
rect 469086 286352 469138 286404
rect 469150 286352 469202 286404
rect 469214 286352 469266 286404
rect 469278 286352 469330 286404
rect 469342 286352 469394 286404
rect 469406 286352 469458 286404
rect 469470 286352 469522 286404
rect 469534 286352 469586 286404
rect 469022 286288 469074 286340
rect 469086 286288 469138 286340
rect 469150 286288 469202 286340
rect 469214 286288 469266 286340
rect 469278 286288 469330 286340
rect 469342 286288 469394 286340
rect 469406 286288 469458 286340
rect 469470 286288 469522 286340
rect 469534 286288 469586 286340
rect 469022 286224 469074 286276
rect 469086 286224 469138 286276
rect 469150 286224 469202 286276
rect 469214 286224 469266 286276
rect 469278 286224 469330 286276
rect 469342 286224 469394 286276
rect 469406 286224 469458 286276
rect 469470 286224 469522 286276
rect 469534 286224 469586 286276
rect 469022 286160 469074 286212
rect 469086 286160 469138 286212
rect 469150 286160 469202 286212
rect 469214 286160 469266 286212
rect 469278 286160 469330 286212
rect 469342 286160 469394 286212
rect 469406 286160 469458 286212
rect 469470 286160 469522 286212
rect 469534 286160 469586 286212
rect 469022 286096 469074 286148
rect 469086 286096 469138 286148
rect 469150 286096 469202 286148
rect 469214 286096 469266 286148
rect 469278 286096 469330 286148
rect 469342 286096 469394 286148
rect 469406 286096 469458 286148
rect 469470 286096 469522 286148
rect 469534 286096 469586 286148
rect 479432 285857 479484 285866
rect 479432 285823 479474 285857
rect 479474 285823 479484 285857
rect 479432 285814 479484 285823
rect 492956 285610 493008 285662
rect 475752 285438 475804 285490
rect 483204 285438 483256 285490
rect 486884 285438 486936 285490
rect 470262 285264 470314 285316
rect 470326 285264 470378 285316
rect 470390 285264 470442 285316
rect 470454 285264 470506 285316
rect 470518 285264 470570 285316
rect 470582 285264 470634 285316
rect 470646 285264 470698 285316
rect 470710 285264 470762 285316
rect 470774 285264 470826 285316
rect 470262 285200 470314 285252
rect 470326 285200 470378 285252
rect 470390 285200 470442 285252
rect 470454 285200 470506 285252
rect 470518 285200 470570 285252
rect 470582 285200 470634 285252
rect 470646 285200 470698 285252
rect 470710 285200 470762 285252
rect 470774 285200 470826 285252
rect 470262 285136 470314 285188
rect 470326 285136 470378 285188
rect 470390 285136 470442 285188
rect 470454 285136 470506 285188
rect 470518 285136 470570 285188
rect 470582 285136 470634 285188
rect 470646 285136 470698 285188
rect 470710 285136 470762 285188
rect 470774 285136 470826 285188
rect 470262 285072 470314 285124
rect 470326 285072 470378 285124
rect 470390 285072 470442 285124
rect 470454 285072 470506 285124
rect 470518 285072 470570 285124
rect 470582 285072 470634 285124
rect 470646 285072 470698 285124
rect 470710 285072 470762 285124
rect 470774 285072 470826 285124
rect 470262 285008 470314 285060
rect 470326 285008 470378 285060
rect 470390 285008 470442 285060
rect 470454 285008 470506 285060
rect 470518 285008 470570 285060
rect 470582 285008 470634 285060
rect 470646 285008 470698 285060
rect 470710 285008 470762 285060
rect 470774 285008 470826 285060
rect 475752 284250 475804 284302
rect 479432 284250 479484 284302
rect 536104 284250 536156 284302
rect 483204 284182 483256 284234
rect 522304 284182 522356 284234
rect 486884 284114 486936 284166
rect 523684 284114 523736 284166
rect 501604 284046 501656 284098
rect 577022 272860 577074 272912
rect 577086 272860 577138 272912
rect 577150 272860 577202 272912
rect 577214 272860 577266 272912
rect 577278 272860 577330 272912
rect 577342 272860 577394 272912
rect 577406 272860 577458 272912
rect 577470 272860 577522 272912
rect 577534 272860 577586 272912
rect 577022 272796 577074 272848
rect 577086 272796 577138 272848
rect 577150 272796 577202 272848
rect 577214 272796 577266 272848
rect 577278 272796 577330 272848
rect 577342 272796 577394 272848
rect 577406 272796 577458 272848
rect 577470 272796 577522 272848
rect 577534 272796 577586 272848
rect 577022 272732 577074 272784
rect 577086 272732 577138 272784
rect 577150 272732 577202 272784
rect 577214 272732 577266 272784
rect 577278 272732 577330 272784
rect 577342 272732 577394 272784
rect 577406 272732 577458 272784
rect 577470 272732 577522 272784
rect 577534 272732 577586 272784
rect 577022 272668 577074 272720
rect 577086 272668 577138 272720
rect 577150 272668 577202 272720
rect 577214 272668 577266 272720
rect 577278 272668 577330 272720
rect 577342 272668 577394 272720
rect 577406 272668 577458 272720
rect 577470 272668 577522 272720
rect 577534 272668 577586 272720
rect 577022 272604 577074 272656
rect 577086 272604 577138 272656
rect 577150 272604 577202 272656
rect 577214 272604 577266 272656
rect 577278 272604 577330 272656
rect 577342 272604 577394 272656
rect 577406 272604 577458 272656
rect 577470 272604 577522 272656
rect 577534 272604 577586 272656
rect 576603 272221 576655 272230
rect 576603 272187 576613 272221
rect 576613 272187 576647 272221
rect 576647 272187 576655 272221
rect 576603 272178 576655 272187
rect 578262 272065 578314 272117
rect 578326 272065 578378 272117
rect 578390 272065 578442 272117
rect 578454 272065 578506 272117
rect 578518 272065 578570 272117
rect 578582 272065 578634 272117
rect 578646 272065 578698 272117
rect 578710 272065 578762 272117
rect 578774 272065 578826 272117
rect 578262 272001 578314 272053
rect 578326 272001 578378 272053
rect 578390 272001 578442 272053
rect 578454 272001 578506 272053
rect 578518 272001 578570 272053
rect 578582 272001 578634 272053
rect 578646 272001 578698 272053
rect 578710 272001 578762 272053
rect 578774 272001 578826 272053
rect 578262 271937 578314 271989
rect 578326 271937 578378 271989
rect 578390 271937 578442 271989
rect 578454 271937 578506 271989
rect 578518 271937 578570 271989
rect 578582 271937 578634 271989
rect 578646 271937 578698 271989
rect 578710 271937 578762 271989
rect 578774 271937 578826 271989
rect 578262 271873 578314 271925
rect 578326 271873 578378 271925
rect 578390 271873 578442 271925
rect 578454 271873 578506 271925
rect 578518 271873 578570 271925
rect 578582 271873 578634 271925
rect 578646 271873 578698 271925
rect 578710 271873 578762 271925
rect 578774 271873 578826 271925
rect 578262 271809 578314 271861
rect 578326 271809 578378 271861
rect 578390 271809 578442 271861
rect 578454 271809 578506 271861
rect 578518 271809 578570 271861
rect 578582 271809 578634 271861
rect 578646 271809 578698 271861
rect 578710 271809 578762 271861
rect 578774 271809 578826 271861
rect 471704 269086 471756 269138
rect 473636 269086 473688 269138
rect 470262 267437 470314 267489
rect 470326 267437 470378 267489
rect 470390 267437 470442 267489
rect 470454 267437 470506 267489
rect 470518 267437 470570 267489
rect 470582 267437 470634 267489
rect 470646 267437 470698 267489
rect 470710 267437 470762 267489
rect 470774 267437 470826 267489
rect 470262 267373 470314 267425
rect 470326 267373 470378 267425
rect 470390 267373 470442 267425
rect 470454 267373 470506 267425
rect 470518 267373 470570 267425
rect 470582 267373 470634 267425
rect 470646 267373 470698 267425
rect 470710 267373 470762 267425
rect 470774 267373 470826 267425
rect 470262 267309 470314 267361
rect 470326 267309 470378 267361
rect 470390 267309 470442 267361
rect 470454 267309 470506 267361
rect 470518 267309 470570 267361
rect 470582 267309 470634 267361
rect 470646 267309 470698 267361
rect 470710 267309 470762 267361
rect 470774 267309 470826 267361
rect 470262 267245 470314 267297
rect 470326 267245 470378 267297
rect 470390 267245 470442 267297
rect 470454 267245 470506 267297
rect 470518 267245 470570 267297
rect 470582 267245 470634 267297
rect 470646 267245 470698 267297
rect 470710 267245 470762 267297
rect 470774 267245 470826 267297
rect 470262 267181 470314 267233
rect 470326 267181 470378 267233
rect 470390 267181 470442 267233
rect 470454 267181 470506 267233
rect 470518 267181 470570 267233
rect 470582 267181 470634 267233
rect 470646 267181 470698 267233
rect 470710 267181 470762 267233
rect 470774 267181 470826 267233
rect 473636 266641 473688 266693
rect 469022 266351 469074 266403
rect 469086 266351 469138 266403
rect 469150 266351 469202 266403
rect 469214 266351 469266 266403
rect 469278 266351 469330 266403
rect 469342 266351 469394 266403
rect 469406 266351 469458 266403
rect 469470 266351 469522 266403
rect 469534 266351 469586 266403
rect 469022 266287 469074 266339
rect 469086 266287 469138 266339
rect 469150 266287 469202 266339
rect 469214 266287 469266 266339
rect 469278 266287 469330 266339
rect 469342 266287 469394 266339
rect 469406 266287 469458 266339
rect 469470 266287 469522 266339
rect 469534 266287 469586 266339
rect 469022 266223 469074 266275
rect 469086 266223 469138 266275
rect 469150 266223 469202 266275
rect 469214 266223 469266 266275
rect 469278 266223 469330 266275
rect 469342 266223 469394 266275
rect 469406 266223 469458 266275
rect 469470 266223 469522 266275
rect 469534 266223 469586 266275
rect 469022 266159 469074 266211
rect 469086 266159 469138 266211
rect 469150 266159 469202 266211
rect 469214 266159 469266 266211
rect 469278 266159 469330 266211
rect 469342 266159 469394 266211
rect 469406 266159 469458 266211
rect 469470 266159 469522 266211
rect 469534 266159 469586 266211
rect 469022 266095 469074 266147
rect 469086 266095 469138 266147
rect 469150 266095 469202 266147
rect 469214 266095 469266 266147
rect 469278 266095 469330 266147
rect 469342 266095 469394 266147
rect 469406 266095 469458 266147
rect 469470 266095 469522 266147
rect 469534 266095 469586 266147
rect 477132 265865 477184 265874
rect 477132 265831 477135 265865
rect 477135 265831 477184 265865
rect 477132 265822 477184 265831
rect 491944 265958 491996 266010
rect 480168 265437 480220 265489
rect 483204 265437 483256 265489
rect 486240 265437 486292 265489
rect 470262 265264 470314 265316
rect 470326 265264 470378 265316
rect 470390 265264 470442 265316
rect 470454 265264 470506 265316
rect 470518 265264 470570 265316
rect 470582 265264 470634 265316
rect 470646 265264 470698 265316
rect 470710 265264 470762 265316
rect 470774 265264 470826 265316
rect 470262 265200 470314 265252
rect 470326 265200 470378 265252
rect 470390 265200 470442 265252
rect 470454 265200 470506 265252
rect 470518 265200 470570 265252
rect 470582 265200 470634 265252
rect 470646 265200 470698 265252
rect 470710 265200 470762 265252
rect 470774 265200 470826 265252
rect 470262 265136 470314 265188
rect 470326 265136 470378 265188
rect 470390 265136 470442 265188
rect 470454 265136 470506 265188
rect 470518 265136 470570 265188
rect 470582 265136 470634 265188
rect 470646 265136 470698 265188
rect 470710 265136 470762 265188
rect 470774 265136 470826 265188
rect 470262 265072 470314 265124
rect 470326 265072 470378 265124
rect 470390 265072 470442 265124
rect 470454 265072 470506 265124
rect 470518 265072 470570 265124
rect 470582 265072 470634 265124
rect 470646 265072 470698 265124
rect 470710 265072 470762 265124
rect 470774 265072 470826 265124
rect 470262 265008 470314 265060
rect 470326 265008 470378 265060
rect 470390 265008 470442 265060
rect 470454 265008 470506 265060
rect 470518 265008 470570 265060
rect 470582 265008 470634 265060
rect 470646 265008 470698 265060
rect 470710 265008 470762 265060
rect 470774 265008 470826 265060
rect 477132 263510 477184 263562
rect 480168 263510 480220 263562
rect 483204 263510 483256 263562
rect 486240 263510 486292 263562
rect 494796 263442 494848 263494
rect 495072 263510 495124 263562
rect 536196 263510 536248 263562
rect 536380 263442 536432 263494
rect 519544 263374 519596 263426
rect 502984 263306 503036 263358
rect 577022 233013 577074 233065
rect 577086 233013 577138 233065
rect 577150 233013 577202 233065
rect 577214 233013 577266 233065
rect 577278 233013 577330 233065
rect 577342 233013 577394 233065
rect 577406 233013 577458 233065
rect 577470 233013 577522 233065
rect 577534 233013 577586 233065
rect 577022 232949 577074 233001
rect 577086 232949 577138 233001
rect 577150 232949 577202 233001
rect 577214 232949 577266 233001
rect 577278 232949 577330 233001
rect 577342 232949 577394 233001
rect 577406 232949 577458 233001
rect 577470 232949 577522 233001
rect 577534 232949 577586 233001
rect 577022 232885 577074 232937
rect 577086 232885 577138 232937
rect 577150 232885 577202 232937
rect 577214 232885 577266 232937
rect 577278 232885 577330 232937
rect 577342 232885 577394 232937
rect 577406 232885 577458 232937
rect 577470 232885 577522 232937
rect 577534 232885 577586 232937
rect 577022 232821 577074 232873
rect 577086 232821 577138 232873
rect 577150 232821 577202 232873
rect 577214 232821 577266 232873
rect 577278 232821 577330 232873
rect 577342 232821 577394 232873
rect 577406 232821 577458 232873
rect 577470 232821 577522 232873
rect 577534 232821 577586 232873
rect 577022 232757 577074 232809
rect 577086 232757 577138 232809
rect 577150 232757 577202 232809
rect 577214 232757 577266 232809
rect 577278 232757 577330 232809
rect 577342 232757 577394 232809
rect 577406 232757 577458 232809
rect 577470 232757 577522 232809
rect 577534 232757 577586 232809
rect 576603 232374 576655 232383
rect 576603 232340 576613 232374
rect 576613 232340 576647 232374
rect 576647 232340 576655 232374
rect 576603 232331 576655 232340
rect 578262 232218 578314 232270
rect 578326 232218 578378 232270
rect 578390 232218 578442 232270
rect 578454 232218 578506 232270
rect 578518 232218 578570 232270
rect 578582 232218 578634 232270
rect 578646 232218 578698 232270
rect 578710 232218 578762 232270
rect 578774 232218 578826 232270
rect 578262 232154 578314 232206
rect 578326 232154 578378 232206
rect 578390 232154 578442 232206
rect 578454 232154 578506 232206
rect 578518 232154 578570 232206
rect 578582 232154 578634 232206
rect 578646 232154 578698 232206
rect 578710 232154 578762 232206
rect 578774 232154 578826 232206
rect 578262 232090 578314 232142
rect 578326 232090 578378 232142
rect 578390 232090 578442 232142
rect 578454 232090 578506 232142
rect 578518 232090 578570 232142
rect 578582 232090 578634 232142
rect 578646 232090 578698 232142
rect 578710 232090 578762 232142
rect 578774 232090 578826 232142
rect 578262 232026 578314 232078
rect 578326 232026 578378 232078
rect 578390 232026 578442 232078
rect 578454 232026 578506 232078
rect 578518 232026 578570 232078
rect 578582 232026 578634 232078
rect 578646 232026 578698 232078
rect 578710 232026 578762 232078
rect 578774 232026 578826 232078
rect 578262 231962 578314 232014
rect 578326 231962 578378 232014
rect 578390 231962 578442 232014
rect 578454 231962 578506 232014
rect 578518 231962 578570 232014
rect 578582 231962 578634 232014
rect 578646 231962 578698 232014
rect 578710 231962 578762 232014
rect 578774 231962 578826 232014
<< metal2 >>
rect 8086 703522 8198 704962
rect 24278 703522 24390 704962
rect 40470 703522 40582 704962
rect 56754 703522 56866 704962
rect 72946 703522 73058 704962
rect 89138 703522 89250 704962
rect 105422 703522 105534 704962
rect 121614 703522 121726 704962
rect 137806 703522 137918 704962
rect 154090 703522 154202 704962
rect 170282 703522 170394 704962
rect 186474 703522 186586 704962
rect 202758 703522 202870 704962
rect 218950 703522 219062 704962
rect 235142 703522 235254 704962
rect 251426 703522 251538 704962
rect 267618 703522 267730 704962
rect 283810 703522 283922 704962
rect 300094 703522 300206 704962
rect 316286 703522 316398 704962
rect 332478 703522 332590 704962
rect 348762 703522 348874 704962
rect 364954 703522 365066 704962
rect 381146 703522 381258 704962
rect 397430 703522 397542 704962
rect 413622 703522 413734 704962
rect 429814 703522 429926 704962
rect 446098 703522 446210 704962
rect 462290 703522 462402 704962
rect 478482 703522 478594 704962
rect 494766 703522 494878 704962
rect 510958 703522 511070 704962
rect 527150 703522 527262 704962
rect 543434 703522 543546 704962
rect 559626 703522 559738 704962
rect 575818 703522 575930 704962
rect 254262 703338 254826 703344
rect 254314 703332 254326 703338
rect 254378 703332 254390 703338
rect 254442 703332 254454 703338
rect 254506 703332 254518 703338
rect 254570 703332 254582 703338
rect 254634 703332 254646 703338
rect 254698 703332 254710 703338
rect 254762 703332 254774 703338
rect 254506 703286 254516 703332
rect 254572 703286 254582 703332
rect 254262 703276 254276 703286
rect 254332 703276 254356 703286
rect 254412 703276 254436 703286
rect 254492 703276 254516 703286
rect 254572 703276 254596 703286
rect 254652 703276 254676 703286
rect 254732 703276 254756 703286
rect 254812 703276 254826 703286
rect 254262 703274 254826 703276
rect 254314 703252 254326 703274
rect 254378 703252 254390 703274
rect 254442 703252 254454 703274
rect 254506 703252 254518 703274
rect 254570 703252 254582 703274
rect 254634 703252 254646 703274
rect 254698 703252 254710 703274
rect 254762 703252 254774 703274
rect 254506 703222 254516 703252
rect 254572 703222 254582 703252
rect 254262 703210 254276 703222
rect 254332 703210 254356 703222
rect 254412 703210 254436 703222
rect 254492 703210 254516 703222
rect 254572 703210 254596 703222
rect 254652 703210 254676 703222
rect 254732 703210 254756 703222
rect 254812 703210 254826 703222
rect 254506 703196 254516 703210
rect 254572 703196 254582 703210
rect 254314 703172 254326 703196
rect 254378 703172 254390 703196
rect 254442 703172 254454 703196
rect 254506 703172 254518 703196
rect 254570 703172 254582 703196
rect 254634 703172 254646 703196
rect 254698 703172 254710 703196
rect 254762 703172 254774 703196
rect 254506 703158 254516 703172
rect 254572 703158 254582 703172
rect 254262 703146 254276 703158
rect 254332 703146 254356 703158
rect 254412 703146 254436 703158
rect 254492 703146 254516 703158
rect 254572 703146 254596 703158
rect 254652 703146 254676 703158
rect 254732 703146 254756 703158
rect 254812 703146 254826 703158
rect 254506 703116 254516 703146
rect 254572 703116 254582 703146
rect 254314 703094 254326 703116
rect 254378 703094 254390 703116
rect 254442 703094 254454 703116
rect 254506 703094 254518 703116
rect 254570 703094 254582 703116
rect 254634 703094 254646 703116
rect 254698 703094 254710 703116
rect 254762 703094 254774 703116
rect 254262 703092 254826 703094
rect 254262 703082 254276 703092
rect 254332 703082 254356 703092
rect 254412 703082 254436 703092
rect 254492 703082 254516 703092
rect 254572 703082 254596 703092
rect 254652 703082 254676 703092
rect 254732 703082 254756 703092
rect 254812 703082 254826 703092
rect 254506 703036 254516 703082
rect 254572 703036 254582 703082
rect 254314 703030 254326 703036
rect 254378 703030 254390 703036
rect 254442 703030 254454 703036
rect 254506 703030 254518 703036
rect 254570 703030 254582 703036
rect 254634 703030 254646 703036
rect 254698 703030 254710 703036
rect 254762 703030 254774 703036
rect 254262 703024 254826 703030
rect 252733 702663 252784 702669
rect 252727 702611 252733 702663
rect 252785 702652 252791 702663
rect 267660 702652 267688 703522
rect 252785 702619 267688 702652
rect 252785 702611 252791 702619
rect 252733 702605 252784 702611
rect 253022 702570 253586 702576
rect 253074 702564 253086 702570
rect 253138 702564 253150 702570
rect 253202 702564 253214 702570
rect 253266 702564 253278 702570
rect 253330 702564 253342 702570
rect 253394 702564 253406 702570
rect 253458 702564 253470 702570
rect 253522 702564 253534 702570
rect 253266 702518 253276 702564
rect 253332 702518 253342 702564
rect 253022 702508 253036 702518
rect 253092 702508 253116 702518
rect 253172 702508 253196 702518
rect 253252 702508 253276 702518
rect 253332 702508 253356 702518
rect 253412 702508 253436 702518
rect 253492 702508 253516 702518
rect 253572 702508 253586 702518
rect 253022 702506 253586 702508
rect 253074 702484 253086 702506
rect 253138 702484 253150 702506
rect 253202 702484 253214 702506
rect 253266 702484 253278 702506
rect 253330 702484 253342 702506
rect 253394 702484 253406 702506
rect 253458 702484 253470 702506
rect 253522 702484 253534 702506
rect 253266 702454 253276 702484
rect 253332 702454 253342 702484
rect 253022 702442 253036 702454
rect 253092 702442 253116 702454
rect 253172 702442 253196 702454
rect 253252 702442 253276 702454
rect 253332 702442 253356 702454
rect 253412 702442 253436 702454
rect 253492 702442 253516 702454
rect 253572 702442 253586 702454
rect 253266 702428 253276 702442
rect 253332 702428 253342 702442
rect 253074 702404 253086 702428
rect 253138 702404 253150 702428
rect 253202 702404 253214 702428
rect 253266 702404 253278 702428
rect 253330 702404 253342 702428
rect 253394 702404 253406 702428
rect 253458 702404 253470 702428
rect 253522 702404 253534 702428
rect 253266 702390 253276 702404
rect 253332 702390 253342 702404
rect 253022 702378 253036 702390
rect 253092 702378 253116 702390
rect 253172 702378 253196 702390
rect 253252 702378 253276 702390
rect 253332 702378 253356 702390
rect 253412 702378 253436 702390
rect 253492 702378 253516 702390
rect 253572 702378 253586 702390
rect 253266 702348 253276 702378
rect 253332 702348 253342 702378
rect 253074 702326 253086 702348
rect 253138 702326 253150 702348
rect 253202 702326 253214 702348
rect 253266 702326 253278 702348
rect 253330 702326 253342 702348
rect 253394 702326 253406 702348
rect 253458 702326 253470 702348
rect 253522 702326 253534 702348
rect 253022 702324 253586 702326
rect 253022 702314 253036 702324
rect 253092 702314 253116 702324
rect 253172 702314 253196 702324
rect 253252 702314 253276 702324
rect 253332 702314 253356 702324
rect 253412 702314 253436 702324
rect 253492 702314 253516 702324
rect 253572 702314 253586 702324
rect 253266 702268 253276 702314
rect 253332 702268 253342 702314
rect 253074 702262 253086 702268
rect 253138 702262 253150 702268
rect 253202 702262 253214 702268
rect 253266 702262 253278 702268
rect 253330 702262 253342 702268
rect 253394 702262 253406 702268
rect 253458 702262 253470 702268
rect 253522 702262 253534 702268
rect 253022 702256 253586 702262
rect 267660 701012 267688 702619
rect 267648 701006 267700 701012
rect 267648 700948 267700 700954
rect 283852 700371 283880 703522
rect 326262 703378 326826 703384
rect 326314 703372 326326 703378
rect 326378 703372 326390 703378
rect 326442 703372 326454 703378
rect 326506 703372 326518 703378
rect 326570 703372 326582 703378
rect 326634 703372 326646 703378
rect 326698 703372 326710 703378
rect 326762 703372 326774 703378
rect 326506 703326 326516 703372
rect 326572 703326 326582 703372
rect 326262 703316 326276 703326
rect 326332 703316 326356 703326
rect 326412 703316 326436 703326
rect 326492 703316 326516 703326
rect 326572 703316 326596 703326
rect 326652 703316 326676 703326
rect 326732 703316 326756 703326
rect 326812 703316 326826 703326
rect 326262 703314 326826 703316
rect 326314 703292 326326 703314
rect 326378 703292 326390 703314
rect 326442 703292 326454 703314
rect 326506 703292 326518 703314
rect 326570 703292 326582 703314
rect 326634 703292 326646 703314
rect 326698 703292 326710 703314
rect 326762 703292 326774 703314
rect 326506 703262 326516 703292
rect 326572 703262 326582 703292
rect 326262 703250 326276 703262
rect 326332 703250 326356 703262
rect 326412 703250 326436 703262
rect 326492 703250 326516 703262
rect 326572 703250 326596 703262
rect 326652 703250 326676 703262
rect 326732 703250 326756 703262
rect 326812 703250 326826 703262
rect 326506 703236 326516 703250
rect 326572 703236 326582 703250
rect 326314 703212 326326 703236
rect 326378 703212 326390 703236
rect 326442 703212 326454 703236
rect 326506 703212 326518 703236
rect 326570 703212 326582 703236
rect 326634 703212 326646 703236
rect 326698 703212 326710 703236
rect 326762 703212 326774 703236
rect 326506 703198 326516 703212
rect 326572 703198 326582 703212
rect 326262 703186 326276 703198
rect 326332 703186 326356 703198
rect 326412 703186 326436 703198
rect 326492 703186 326516 703198
rect 326572 703186 326596 703198
rect 326652 703186 326676 703198
rect 326732 703186 326756 703198
rect 326812 703186 326826 703198
rect 326506 703156 326516 703186
rect 326572 703156 326582 703186
rect 326314 703134 326326 703156
rect 326378 703134 326390 703156
rect 326442 703134 326454 703156
rect 326506 703134 326518 703156
rect 326570 703134 326582 703156
rect 326634 703134 326646 703156
rect 326698 703134 326710 703156
rect 326762 703134 326774 703156
rect 326262 703132 326826 703134
rect 326262 703122 326276 703132
rect 326332 703122 326356 703132
rect 326412 703122 326436 703132
rect 326492 703122 326516 703132
rect 326572 703122 326596 703132
rect 326652 703122 326676 703132
rect 326732 703122 326756 703132
rect 326812 703122 326826 703132
rect 326506 703076 326516 703122
rect 326572 703076 326582 703122
rect 326314 703070 326326 703076
rect 326378 703070 326390 703076
rect 326442 703070 326454 703076
rect 326506 703070 326518 703076
rect 326570 703070 326582 703076
rect 326634 703070 326646 703076
rect 326698 703070 326710 703076
rect 326762 703070 326774 703076
rect 326262 703064 326826 703070
rect 324732 702703 324783 702709
rect 324726 702651 324732 702703
rect 324784 702692 324790 702703
rect 332520 702692 332548 703522
rect 324784 702659 332548 702692
rect 324784 702651 324790 702659
rect 324732 702645 324783 702651
rect 325022 702610 325586 702616
rect 325074 702604 325086 702610
rect 325138 702604 325150 702610
rect 325202 702604 325214 702610
rect 325266 702604 325278 702610
rect 325330 702604 325342 702610
rect 325394 702604 325406 702610
rect 325458 702604 325470 702610
rect 325522 702604 325534 702610
rect 325266 702558 325276 702604
rect 325332 702558 325342 702604
rect 325022 702548 325036 702558
rect 325092 702548 325116 702558
rect 325172 702548 325196 702558
rect 325252 702548 325276 702558
rect 325332 702548 325356 702558
rect 325412 702548 325436 702558
rect 325492 702548 325516 702558
rect 325572 702548 325586 702558
rect 325022 702546 325586 702548
rect 325074 702524 325086 702546
rect 325138 702524 325150 702546
rect 325202 702524 325214 702546
rect 325266 702524 325278 702546
rect 325330 702524 325342 702546
rect 325394 702524 325406 702546
rect 325458 702524 325470 702546
rect 325522 702524 325534 702546
rect 325266 702494 325276 702524
rect 325332 702494 325342 702524
rect 325022 702482 325036 702494
rect 325092 702482 325116 702494
rect 325172 702482 325196 702494
rect 325252 702482 325276 702494
rect 325332 702482 325356 702494
rect 325412 702482 325436 702494
rect 325492 702482 325516 702494
rect 325572 702482 325586 702494
rect 325266 702468 325276 702482
rect 325332 702468 325342 702482
rect 325074 702444 325086 702468
rect 325138 702444 325150 702468
rect 325202 702444 325214 702468
rect 325266 702444 325278 702468
rect 325330 702444 325342 702468
rect 325394 702444 325406 702468
rect 325458 702444 325470 702468
rect 325522 702444 325534 702468
rect 325266 702430 325276 702444
rect 325332 702430 325342 702444
rect 325022 702418 325036 702430
rect 325092 702418 325116 702430
rect 325172 702418 325196 702430
rect 325252 702418 325276 702430
rect 325332 702418 325356 702430
rect 325412 702418 325436 702430
rect 325492 702418 325516 702430
rect 325572 702418 325586 702430
rect 325266 702388 325276 702418
rect 325332 702388 325342 702418
rect 325074 702366 325086 702388
rect 325138 702366 325150 702388
rect 325202 702366 325214 702388
rect 325266 702366 325278 702388
rect 325330 702366 325342 702388
rect 325394 702366 325406 702388
rect 325458 702366 325470 702388
rect 325522 702366 325534 702388
rect 325022 702364 325586 702366
rect 325022 702354 325036 702364
rect 325092 702354 325116 702364
rect 325172 702354 325196 702364
rect 325252 702354 325276 702364
rect 325332 702354 325356 702364
rect 325412 702354 325436 702364
rect 325492 702354 325516 702364
rect 325572 702354 325586 702364
rect 325266 702308 325276 702354
rect 325332 702308 325342 702354
rect 325074 702302 325086 702308
rect 325138 702302 325150 702308
rect 325202 702302 325214 702308
rect 325266 702302 325278 702308
rect 325330 702302 325342 702308
rect 325394 702302 325406 702308
rect 325458 702302 325470 702308
rect 325522 702302 325534 702308
rect 325022 702296 325586 702302
rect 332520 701012 332548 702659
rect 332508 701006 332560 701012
rect 332508 700948 332560 700954
rect 348804 700507 348832 703522
rect 362262 702909 362826 702915
rect 362314 702903 362326 702909
rect 362378 702903 362390 702909
rect 362442 702903 362454 702909
rect 362506 702903 362518 702909
rect 362570 702903 362582 702909
rect 362634 702903 362646 702909
rect 362698 702903 362710 702909
rect 362762 702903 362774 702909
rect 362506 702857 362516 702903
rect 362572 702857 362582 702903
rect 362262 702847 362276 702857
rect 362332 702847 362356 702857
rect 362412 702847 362436 702857
rect 362492 702847 362516 702857
rect 362572 702847 362596 702857
rect 362652 702847 362676 702857
rect 362732 702847 362756 702857
rect 362812 702847 362826 702857
rect 362262 702845 362826 702847
rect 362314 702823 362326 702845
rect 362378 702823 362390 702845
rect 362442 702823 362454 702845
rect 362506 702823 362518 702845
rect 362570 702823 362582 702845
rect 362634 702823 362646 702845
rect 362698 702823 362710 702845
rect 362762 702823 362774 702845
rect 362506 702793 362516 702823
rect 362572 702793 362582 702823
rect 362262 702781 362276 702793
rect 362332 702781 362356 702793
rect 362412 702781 362436 702793
rect 362492 702781 362516 702793
rect 362572 702781 362596 702793
rect 362652 702781 362676 702793
rect 362732 702781 362756 702793
rect 362812 702781 362826 702793
rect 362506 702767 362516 702781
rect 362572 702767 362582 702781
rect 362314 702743 362326 702767
rect 362378 702743 362390 702767
rect 362442 702743 362454 702767
rect 362506 702743 362518 702767
rect 362570 702743 362582 702767
rect 362634 702743 362646 702767
rect 362698 702743 362710 702767
rect 362762 702743 362774 702767
rect 362506 702729 362516 702743
rect 362572 702729 362582 702743
rect 362262 702717 362276 702729
rect 362332 702717 362356 702729
rect 362412 702717 362436 702729
rect 362492 702717 362516 702729
rect 362572 702717 362596 702729
rect 362652 702717 362676 702729
rect 362732 702717 362756 702729
rect 362812 702717 362826 702729
rect 362506 702687 362516 702717
rect 362572 702687 362582 702717
rect 362314 702665 362326 702687
rect 362378 702665 362390 702687
rect 362442 702665 362454 702687
rect 362506 702665 362518 702687
rect 362570 702665 362582 702687
rect 362634 702665 362646 702687
rect 362698 702665 362710 702687
rect 362762 702665 362774 702687
rect 362262 702663 362826 702665
rect 362262 702653 362276 702663
rect 362332 702653 362356 702663
rect 362412 702653 362436 702663
rect 362492 702653 362516 702663
rect 362572 702653 362596 702663
rect 362652 702653 362676 702663
rect 362732 702653 362756 702663
rect 362812 702653 362826 702663
rect 362506 702607 362516 702653
rect 362572 702607 362582 702653
rect 362314 702601 362326 702607
rect 362378 702601 362390 702607
rect 362442 702601 362454 702607
rect 362506 702601 362518 702607
rect 362570 702601 362582 702607
rect 362634 702601 362646 702607
rect 362698 702601 362710 702607
rect 362762 702601 362774 702607
rect 362262 702595 362826 702601
rect 360759 702234 360810 702240
rect 360753 702182 360759 702234
rect 360811 702223 360817 702234
rect 397472 702223 397500 703522
rect 360811 702190 397500 702223
rect 360811 702182 360817 702190
rect 360759 702176 360810 702182
rect 361022 702141 361586 702147
rect 361074 702135 361086 702141
rect 361138 702135 361150 702141
rect 361202 702135 361214 702141
rect 361266 702135 361278 702141
rect 361330 702135 361342 702141
rect 361394 702135 361406 702141
rect 361458 702135 361470 702141
rect 361522 702135 361534 702141
rect 361266 702089 361276 702135
rect 361332 702089 361342 702135
rect 361022 702079 361036 702089
rect 361092 702079 361116 702089
rect 361172 702079 361196 702089
rect 361252 702079 361276 702089
rect 361332 702079 361356 702089
rect 361412 702079 361436 702089
rect 361492 702079 361516 702089
rect 361572 702079 361586 702089
rect 361022 702077 361586 702079
rect 361074 702055 361086 702077
rect 361138 702055 361150 702077
rect 361202 702055 361214 702077
rect 361266 702055 361278 702077
rect 361330 702055 361342 702077
rect 361394 702055 361406 702077
rect 361458 702055 361470 702077
rect 361522 702055 361534 702077
rect 361266 702025 361276 702055
rect 361332 702025 361342 702055
rect 361022 702013 361036 702025
rect 361092 702013 361116 702025
rect 361172 702013 361196 702025
rect 361252 702013 361276 702025
rect 361332 702013 361356 702025
rect 361412 702013 361436 702025
rect 361492 702013 361516 702025
rect 361572 702013 361586 702025
rect 361266 701999 361276 702013
rect 361332 701999 361342 702013
rect 361074 701975 361086 701999
rect 361138 701975 361150 701999
rect 361202 701975 361214 701999
rect 361266 701975 361278 701999
rect 361330 701975 361342 701999
rect 361394 701975 361406 701999
rect 361458 701975 361470 701999
rect 361522 701975 361534 701999
rect 361266 701961 361276 701975
rect 361332 701961 361342 701975
rect 361022 701949 361036 701961
rect 361092 701949 361116 701961
rect 361172 701949 361196 701961
rect 361252 701949 361276 701961
rect 361332 701949 361356 701961
rect 361412 701949 361436 701961
rect 361492 701949 361516 701961
rect 361572 701949 361586 701961
rect 361266 701919 361276 701949
rect 361332 701919 361342 701949
rect 361074 701897 361086 701919
rect 361138 701897 361150 701919
rect 361202 701897 361214 701919
rect 361266 701897 361278 701919
rect 361330 701897 361342 701919
rect 361394 701897 361406 701919
rect 361458 701897 361470 701919
rect 361522 701897 361534 701919
rect 361022 701895 361586 701897
rect 361022 701885 361036 701895
rect 361092 701885 361116 701895
rect 361172 701885 361196 701895
rect 361252 701885 361276 701895
rect 361332 701885 361356 701895
rect 361412 701885 361436 701895
rect 361492 701885 361516 701895
rect 361572 701885 361586 701895
rect 361266 701839 361276 701885
rect 361332 701839 361342 701885
rect 361074 701833 361086 701839
rect 361138 701833 361150 701839
rect 361202 701833 361214 701839
rect 361266 701833 361278 701839
rect 361330 701833 361342 701839
rect 361394 701833 361406 701839
rect 361458 701833 361470 701839
rect 361522 701833 361534 701839
rect 361022 701827 361586 701833
rect 397472 701012 397500 702190
rect 397460 701006 397512 701012
rect 397460 700948 397512 700954
rect 413664 700643 413692 703522
rect 434262 702772 434826 702778
rect 434314 702766 434326 702772
rect 434378 702766 434390 702772
rect 434442 702766 434454 702772
rect 434506 702766 434518 702772
rect 434570 702766 434582 702772
rect 434634 702766 434646 702772
rect 434698 702766 434710 702772
rect 434762 702766 434774 702772
rect 434506 702720 434516 702766
rect 434572 702720 434582 702766
rect 434262 702710 434276 702720
rect 434332 702710 434356 702720
rect 434412 702710 434436 702720
rect 434492 702710 434516 702720
rect 434572 702710 434596 702720
rect 434652 702710 434676 702720
rect 434732 702710 434756 702720
rect 434812 702710 434826 702720
rect 434262 702708 434826 702710
rect 434314 702686 434326 702708
rect 434378 702686 434390 702708
rect 434442 702686 434454 702708
rect 434506 702686 434518 702708
rect 434570 702686 434582 702708
rect 434634 702686 434646 702708
rect 434698 702686 434710 702708
rect 434762 702686 434774 702708
rect 434506 702656 434516 702686
rect 434572 702656 434582 702686
rect 434262 702644 434276 702656
rect 434332 702644 434356 702656
rect 434412 702644 434436 702656
rect 434492 702644 434516 702656
rect 434572 702644 434596 702656
rect 434652 702644 434676 702656
rect 434732 702644 434756 702656
rect 434812 702644 434826 702656
rect 434506 702630 434516 702644
rect 434572 702630 434582 702644
rect 434314 702606 434326 702630
rect 434378 702606 434390 702630
rect 434442 702606 434454 702630
rect 434506 702606 434518 702630
rect 434570 702606 434582 702630
rect 434634 702606 434646 702630
rect 434698 702606 434710 702630
rect 434762 702606 434774 702630
rect 434506 702592 434516 702606
rect 434572 702592 434582 702606
rect 434262 702580 434276 702592
rect 434332 702580 434356 702592
rect 434412 702580 434436 702592
rect 434492 702580 434516 702592
rect 434572 702580 434596 702592
rect 434652 702580 434676 702592
rect 434732 702580 434756 702592
rect 434812 702580 434826 702592
rect 434506 702550 434516 702580
rect 434572 702550 434582 702580
rect 434314 702528 434326 702550
rect 434378 702528 434390 702550
rect 434442 702528 434454 702550
rect 434506 702528 434518 702550
rect 434570 702528 434582 702550
rect 434634 702528 434646 702550
rect 434698 702528 434710 702550
rect 434762 702528 434774 702550
rect 434262 702526 434826 702528
rect 434262 702516 434276 702526
rect 434332 702516 434356 702526
rect 434412 702516 434436 702526
rect 434492 702516 434516 702526
rect 434572 702516 434596 702526
rect 434652 702516 434676 702526
rect 434732 702516 434756 702526
rect 434812 702516 434826 702526
rect 434506 702470 434516 702516
rect 434572 702470 434582 702516
rect 434314 702464 434326 702470
rect 434378 702464 434390 702470
rect 434442 702464 434454 702470
rect 434506 702464 434518 702470
rect 434570 702464 434582 702470
rect 434634 702464 434646 702470
rect 434698 702464 434710 702470
rect 434762 702464 434774 702470
rect 434262 702458 434826 702464
rect 432729 702097 432780 702103
rect 432723 702045 432729 702097
rect 432781 702086 432787 702097
rect 462332 702086 462360 703522
rect 432781 702053 462360 702086
rect 432781 702045 432787 702053
rect 432729 702039 432780 702045
rect 433022 702004 433586 702010
rect 433074 701998 433086 702004
rect 433138 701998 433150 702004
rect 433202 701998 433214 702004
rect 433266 701998 433278 702004
rect 433330 701998 433342 702004
rect 433394 701998 433406 702004
rect 433458 701998 433470 702004
rect 433522 701998 433534 702004
rect 433266 701952 433276 701998
rect 433332 701952 433342 701998
rect 433022 701942 433036 701952
rect 433092 701942 433116 701952
rect 433172 701942 433196 701952
rect 433252 701942 433276 701952
rect 433332 701942 433356 701952
rect 433412 701942 433436 701952
rect 433492 701942 433516 701952
rect 433572 701942 433586 701952
rect 433022 701940 433586 701942
rect 433074 701918 433086 701940
rect 433138 701918 433150 701940
rect 433202 701918 433214 701940
rect 433266 701918 433278 701940
rect 433330 701918 433342 701940
rect 433394 701918 433406 701940
rect 433458 701918 433470 701940
rect 433522 701918 433534 701940
rect 433266 701888 433276 701918
rect 433332 701888 433342 701918
rect 433022 701876 433036 701888
rect 433092 701876 433116 701888
rect 433172 701876 433196 701888
rect 433252 701876 433276 701888
rect 433332 701876 433356 701888
rect 433412 701876 433436 701888
rect 433492 701876 433516 701888
rect 433572 701876 433586 701888
rect 433266 701862 433276 701876
rect 433332 701862 433342 701876
rect 433074 701838 433086 701862
rect 433138 701838 433150 701862
rect 433202 701838 433214 701862
rect 433266 701838 433278 701862
rect 433330 701838 433342 701862
rect 433394 701838 433406 701862
rect 433458 701838 433470 701862
rect 433522 701838 433534 701862
rect 433266 701824 433276 701838
rect 433332 701824 433342 701838
rect 433022 701812 433036 701824
rect 433092 701812 433116 701824
rect 433172 701812 433196 701824
rect 433252 701812 433276 701824
rect 433332 701812 433356 701824
rect 433412 701812 433436 701824
rect 433492 701812 433516 701824
rect 433572 701812 433586 701824
rect 433266 701782 433276 701812
rect 433332 701782 433342 701812
rect 433074 701760 433086 701782
rect 433138 701760 433150 701782
rect 433202 701760 433214 701782
rect 433266 701760 433278 701782
rect 433330 701760 433342 701782
rect 433394 701760 433406 701782
rect 433458 701760 433470 701782
rect 433522 701760 433534 701782
rect 433022 701758 433586 701760
rect 433022 701748 433036 701758
rect 433092 701748 433116 701758
rect 433172 701748 433196 701758
rect 433252 701748 433276 701758
rect 433332 701748 433356 701758
rect 433412 701748 433436 701758
rect 433492 701748 433516 701758
rect 433572 701748 433586 701758
rect 433266 701702 433276 701748
rect 433332 701702 433342 701748
rect 433074 701696 433086 701702
rect 433138 701696 433150 701702
rect 433202 701696 433214 701702
rect 433266 701696 433278 701702
rect 433330 701696 433342 701702
rect 433394 701696 433406 701702
rect 433458 701696 433470 701702
rect 433522 701696 433534 701702
rect 433022 701690 433586 701696
rect 462332 701012 462360 702053
rect 462320 701006 462372 701012
rect 462320 700948 462372 700954
rect 478524 700779 478552 703522
rect 506262 702526 506826 702532
rect 506314 702520 506326 702526
rect 506378 702520 506390 702526
rect 506442 702520 506454 702526
rect 506506 702520 506518 702526
rect 506570 702520 506582 702526
rect 506634 702520 506646 702526
rect 506698 702520 506710 702526
rect 506762 702520 506774 702526
rect 506506 702474 506516 702520
rect 506572 702474 506582 702520
rect 506262 702464 506276 702474
rect 506332 702464 506356 702474
rect 506412 702464 506436 702474
rect 506492 702464 506516 702474
rect 506572 702464 506596 702474
rect 506652 702464 506676 702474
rect 506732 702464 506756 702474
rect 506812 702464 506826 702474
rect 506262 702462 506826 702464
rect 506314 702440 506326 702462
rect 506378 702440 506390 702462
rect 506442 702440 506454 702462
rect 506506 702440 506518 702462
rect 506570 702440 506582 702462
rect 506634 702440 506646 702462
rect 506698 702440 506710 702462
rect 506762 702440 506774 702462
rect 506506 702410 506516 702440
rect 506572 702410 506582 702440
rect 506262 702398 506276 702410
rect 506332 702398 506356 702410
rect 506412 702398 506436 702410
rect 506492 702398 506516 702410
rect 506572 702398 506596 702410
rect 506652 702398 506676 702410
rect 506732 702398 506756 702410
rect 506812 702398 506826 702410
rect 506506 702384 506516 702398
rect 506572 702384 506582 702398
rect 506314 702360 506326 702384
rect 506378 702360 506390 702384
rect 506442 702360 506454 702384
rect 506506 702360 506518 702384
rect 506570 702360 506582 702384
rect 506634 702360 506646 702384
rect 506698 702360 506710 702384
rect 506762 702360 506774 702384
rect 506506 702346 506516 702360
rect 506572 702346 506582 702360
rect 506262 702334 506276 702346
rect 506332 702334 506356 702346
rect 506412 702334 506436 702346
rect 506492 702334 506516 702346
rect 506572 702334 506596 702346
rect 506652 702334 506676 702346
rect 506732 702334 506756 702346
rect 506812 702334 506826 702346
rect 506506 702304 506516 702334
rect 506572 702304 506582 702334
rect 506314 702282 506326 702304
rect 506378 702282 506390 702304
rect 506442 702282 506454 702304
rect 506506 702282 506518 702304
rect 506570 702282 506582 702304
rect 506634 702282 506646 702304
rect 506698 702282 506710 702304
rect 506762 702282 506774 702304
rect 506262 702280 506826 702282
rect 506262 702270 506276 702280
rect 506332 702270 506356 702280
rect 506412 702270 506436 702280
rect 506492 702270 506516 702280
rect 506572 702270 506596 702280
rect 506652 702270 506676 702280
rect 506732 702270 506756 702280
rect 506812 702270 506826 702280
rect 506506 702224 506516 702270
rect 506572 702224 506582 702270
rect 506314 702218 506326 702224
rect 506378 702218 506390 702224
rect 506442 702218 506454 702224
rect 506506 702218 506518 702224
rect 506570 702218 506582 702224
rect 506634 702218 506646 702224
rect 506698 702218 506710 702224
rect 506762 702218 506774 702224
rect 506262 702212 506826 702218
rect 504725 701851 504776 701857
rect 504719 701799 504725 701851
rect 504777 701840 504783 701851
rect 527192 701840 527220 703522
rect 504777 701807 527220 701840
rect 504777 701799 504783 701807
rect 504725 701793 504776 701799
rect 505022 701758 505586 701764
rect 505074 701752 505086 701758
rect 505138 701752 505150 701758
rect 505202 701752 505214 701758
rect 505266 701752 505278 701758
rect 505330 701752 505342 701758
rect 505394 701752 505406 701758
rect 505458 701752 505470 701758
rect 505522 701752 505534 701758
rect 505266 701706 505276 701752
rect 505332 701706 505342 701752
rect 505022 701696 505036 701706
rect 505092 701696 505116 701706
rect 505172 701696 505196 701706
rect 505252 701696 505276 701706
rect 505332 701696 505356 701706
rect 505412 701696 505436 701706
rect 505492 701696 505516 701706
rect 505572 701696 505586 701706
rect 505022 701694 505586 701696
rect 505074 701672 505086 701694
rect 505138 701672 505150 701694
rect 505202 701672 505214 701694
rect 505266 701672 505278 701694
rect 505330 701672 505342 701694
rect 505394 701672 505406 701694
rect 505458 701672 505470 701694
rect 505522 701672 505534 701694
rect 505266 701642 505276 701672
rect 505332 701642 505342 701672
rect 505022 701630 505036 701642
rect 505092 701630 505116 701642
rect 505172 701630 505196 701642
rect 505252 701630 505276 701642
rect 505332 701630 505356 701642
rect 505412 701630 505436 701642
rect 505492 701630 505516 701642
rect 505572 701630 505586 701642
rect 505266 701616 505276 701630
rect 505332 701616 505342 701630
rect 505074 701592 505086 701616
rect 505138 701592 505150 701616
rect 505202 701592 505214 701616
rect 505266 701592 505278 701616
rect 505330 701592 505342 701616
rect 505394 701592 505406 701616
rect 505458 701592 505470 701616
rect 505522 701592 505534 701616
rect 505266 701578 505276 701592
rect 505332 701578 505342 701592
rect 505022 701566 505036 701578
rect 505092 701566 505116 701578
rect 505172 701566 505196 701578
rect 505252 701566 505276 701578
rect 505332 701566 505356 701578
rect 505412 701566 505436 701578
rect 505492 701566 505516 701578
rect 505572 701566 505586 701578
rect 505266 701536 505276 701566
rect 505332 701536 505342 701566
rect 505074 701514 505086 701536
rect 505138 701514 505150 701536
rect 505202 701514 505214 701536
rect 505266 701514 505278 701536
rect 505330 701514 505342 701536
rect 505394 701514 505406 701536
rect 505458 701514 505470 701536
rect 505522 701514 505534 701536
rect 505022 701512 505586 701514
rect 505022 701502 505036 701512
rect 505092 701502 505116 701512
rect 505172 701502 505196 701512
rect 505252 701502 505276 701512
rect 505332 701502 505356 701512
rect 505412 701502 505436 701512
rect 505492 701502 505516 701512
rect 505572 701502 505586 701512
rect 505266 701456 505276 701502
rect 505332 701456 505342 701502
rect 505074 701450 505086 701456
rect 505138 701450 505150 701456
rect 505202 701450 505214 701456
rect 505266 701450 505278 701456
rect 505330 701450 505342 701456
rect 505394 701450 505406 701456
rect 505458 701450 505470 701456
rect 505522 701450 505534 701456
rect 505022 701444 505586 701450
rect 527192 701012 527220 701807
rect 527180 701006 527232 701012
rect 527180 700948 527232 700954
rect 478510 700770 478566 700779
rect 478510 700705 478566 700714
rect 413650 700634 413706 700643
rect 413650 700569 413706 700578
rect 348790 700498 348846 700507
rect 348790 700433 348846 700442
rect 283838 700362 283894 700371
rect 283838 700297 283894 700306
rect 543476 699827 543504 703522
rect 547970 700770 548026 700779
rect 547970 700705 548026 700714
rect 547878 700634 547934 700643
rect 547878 700569 547934 700578
rect 547418 700498 547474 700507
rect 547418 700433 547474 700442
rect 547326 700362 547382 700371
rect 547326 700297 547382 700306
rect 543462 699818 543518 699827
rect 543462 699753 543518 699762
rect 505022 554604 505586 554610
rect 505074 554598 505086 554604
rect 505138 554598 505150 554604
rect 505202 554598 505214 554604
rect 505266 554598 505278 554604
rect 505330 554598 505342 554604
rect 505394 554598 505406 554604
rect 505458 554598 505470 554604
rect 505522 554598 505534 554604
rect 505266 554552 505276 554598
rect 505332 554552 505342 554598
rect 505022 554542 505036 554552
rect 505092 554542 505116 554552
rect 505172 554542 505196 554552
rect 505252 554542 505276 554552
rect 505332 554542 505356 554552
rect 505412 554542 505436 554552
rect 505492 554542 505516 554552
rect 505572 554542 505586 554552
rect 505022 554540 505586 554542
rect 505074 554518 505086 554540
rect 505138 554518 505150 554540
rect 505202 554518 505214 554540
rect 505266 554518 505278 554540
rect 505330 554518 505342 554540
rect 505394 554518 505406 554540
rect 505458 554518 505470 554540
rect 505522 554518 505534 554540
rect 505266 554488 505276 554518
rect 505332 554488 505342 554518
rect 505022 554476 505036 554488
rect 505092 554476 505116 554488
rect 505172 554476 505196 554488
rect 505252 554476 505276 554488
rect 505332 554476 505356 554488
rect 505412 554476 505436 554488
rect 505492 554476 505516 554488
rect 505572 554476 505586 554488
rect 505266 554462 505276 554476
rect 505332 554462 505342 554476
rect 505074 554438 505086 554462
rect 505138 554438 505150 554462
rect 505202 554438 505214 554462
rect 505266 554438 505278 554462
rect 505330 554438 505342 554462
rect 505394 554438 505406 554462
rect 505458 554438 505470 554462
rect 505522 554438 505534 554462
rect 505266 554424 505276 554438
rect 505332 554424 505342 554438
rect 505022 554412 505036 554424
rect 505092 554412 505116 554424
rect 505172 554412 505196 554424
rect 505252 554412 505276 554424
rect 505332 554412 505356 554424
rect 505412 554412 505436 554424
rect 505492 554412 505516 554424
rect 505572 554412 505586 554424
rect 505266 554382 505276 554412
rect 505332 554382 505342 554412
rect 505074 554360 505086 554382
rect 505138 554360 505150 554382
rect 505202 554360 505214 554382
rect 505266 554360 505278 554382
rect 505330 554360 505342 554382
rect 505394 554360 505406 554382
rect 505458 554360 505470 554382
rect 505522 554360 505534 554382
rect 505022 554358 505586 554360
rect 505022 554348 505036 554358
rect 505092 554348 505116 554358
rect 505172 554348 505196 554358
rect 505252 554348 505276 554358
rect 505332 554348 505356 554358
rect 505412 554348 505436 554358
rect 505492 554348 505516 554358
rect 505572 554348 505586 554358
rect 505266 554302 505276 554348
rect 505332 554302 505342 554348
rect 505074 554296 505086 554302
rect 505138 554296 505150 554302
rect 505202 554296 505214 554302
rect 505266 554296 505278 554302
rect 505330 554296 505342 554302
rect 505394 554296 505406 554302
rect 505458 554296 505470 554302
rect 505522 554296 505534 554302
rect 505022 554290 505586 554296
rect 536104 554058 536156 554064
rect 536104 554000 536156 554006
rect 506262 553809 506826 553815
rect 506314 553803 506326 553809
rect 506378 553803 506390 553809
rect 506442 553803 506454 553809
rect 506506 553803 506518 553809
rect 506570 553803 506582 553809
rect 506634 553803 506646 553809
rect 506698 553803 506710 553809
rect 506762 553803 506774 553809
rect 506506 553757 506516 553803
rect 506572 553757 506582 553803
rect 506262 553747 506276 553757
rect 506332 553747 506356 553757
rect 506412 553747 506436 553757
rect 506492 553747 506516 553757
rect 506572 553747 506596 553757
rect 506652 553747 506676 553757
rect 506732 553747 506756 553757
rect 506812 553747 506826 553757
rect 506262 553745 506826 553747
rect 506314 553723 506326 553745
rect 506378 553723 506390 553745
rect 506442 553723 506454 553745
rect 506506 553723 506518 553745
rect 506570 553723 506582 553745
rect 506634 553723 506646 553745
rect 506698 553723 506710 553745
rect 506762 553723 506774 553745
rect 506506 553693 506516 553723
rect 506572 553693 506582 553723
rect 506262 553681 506276 553693
rect 506332 553681 506356 553693
rect 506412 553681 506436 553693
rect 506492 553681 506516 553693
rect 506572 553681 506596 553693
rect 506652 553681 506676 553693
rect 506732 553681 506756 553693
rect 506812 553681 506826 553693
rect 506506 553667 506516 553681
rect 506572 553667 506582 553681
rect 506314 553643 506326 553667
rect 506378 553643 506390 553667
rect 506442 553643 506454 553667
rect 506506 553643 506518 553667
rect 506570 553643 506582 553667
rect 506634 553643 506646 553667
rect 506698 553643 506710 553667
rect 506762 553643 506774 553667
rect 506506 553629 506516 553643
rect 506572 553629 506582 553643
rect 506262 553617 506276 553629
rect 506332 553617 506356 553629
rect 506412 553617 506436 553629
rect 506492 553617 506516 553629
rect 506572 553617 506596 553629
rect 506652 553617 506676 553629
rect 506732 553617 506756 553629
rect 506812 553617 506826 553629
rect 506506 553587 506516 553617
rect 506572 553587 506582 553617
rect 506314 553565 506326 553587
rect 506378 553565 506390 553587
rect 506442 553565 506454 553587
rect 506506 553565 506518 553587
rect 506570 553565 506582 553587
rect 506634 553565 506646 553587
rect 506698 553565 506710 553587
rect 506762 553565 506774 553587
rect 506262 553563 506826 553565
rect 506262 553553 506276 553563
rect 506332 553553 506356 553563
rect 506412 553553 506436 553563
rect 506492 553553 506516 553563
rect 506572 553553 506596 553563
rect 506652 553553 506676 553563
rect 506732 553553 506756 553563
rect 506812 553553 506826 553563
rect 506506 553507 506516 553553
rect 506572 553507 506582 553553
rect 506314 553501 506326 553507
rect 506378 553501 506390 553507
rect 506442 553501 506454 553507
rect 506506 553501 506518 553507
rect 506570 553501 506582 553507
rect 506634 553501 506646 553507
rect 506698 553501 506710 553507
rect 506762 553501 506774 553507
rect 506262 553495 506826 553501
rect 471704 453350 471756 453356
rect 471704 453292 471756 453298
rect 470262 451487 470826 451493
rect 470314 451481 470326 451487
rect 470378 451481 470390 451487
rect 470442 451481 470454 451487
rect 470506 451481 470518 451487
rect 470570 451481 470582 451487
rect 470634 451481 470646 451487
rect 470698 451481 470710 451487
rect 470762 451481 470774 451487
rect 470506 451435 470516 451481
rect 470572 451435 470582 451481
rect 470262 451425 470276 451435
rect 470332 451425 470356 451435
rect 470412 451425 470436 451435
rect 470492 451425 470516 451435
rect 470572 451425 470596 451435
rect 470652 451425 470676 451435
rect 470732 451425 470756 451435
rect 470812 451425 470826 451435
rect 470262 451423 470826 451425
rect 470314 451401 470326 451423
rect 470378 451401 470390 451423
rect 470442 451401 470454 451423
rect 470506 451401 470518 451423
rect 470570 451401 470582 451423
rect 470634 451401 470646 451423
rect 470698 451401 470710 451423
rect 470762 451401 470774 451423
rect 470506 451371 470516 451401
rect 470572 451371 470582 451401
rect 470262 451359 470276 451371
rect 470332 451359 470356 451371
rect 470412 451359 470436 451371
rect 470492 451359 470516 451371
rect 470572 451359 470596 451371
rect 470652 451359 470676 451371
rect 470732 451359 470756 451371
rect 470812 451359 470826 451371
rect 470506 451345 470516 451359
rect 470572 451345 470582 451359
rect 470314 451321 470326 451345
rect 470378 451321 470390 451345
rect 470442 451321 470454 451345
rect 470506 451321 470518 451345
rect 470570 451321 470582 451345
rect 470634 451321 470646 451345
rect 470698 451321 470710 451345
rect 470762 451321 470774 451345
rect 470506 451307 470516 451321
rect 470572 451307 470582 451321
rect 470262 451295 470276 451307
rect 470332 451295 470356 451307
rect 470412 451295 470436 451307
rect 470492 451295 470516 451307
rect 470572 451295 470596 451307
rect 470652 451295 470676 451307
rect 470732 451295 470756 451307
rect 470812 451295 470826 451307
rect 470506 451265 470516 451295
rect 470572 451265 470582 451295
rect 470314 451243 470326 451265
rect 470378 451243 470390 451265
rect 470442 451243 470454 451265
rect 470506 451243 470518 451265
rect 470570 451243 470582 451265
rect 470634 451243 470646 451265
rect 470698 451243 470710 451265
rect 470762 451243 470774 451265
rect 470262 451241 470826 451243
rect 470262 451231 470276 451241
rect 470332 451231 470356 451241
rect 470412 451231 470436 451241
rect 470492 451231 470516 451241
rect 470572 451231 470596 451241
rect 470652 451231 470676 451241
rect 470732 451231 470756 451241
rect 470812 451231 470826 451241
rect 470506 451185 470516 451231
rect 470572 451185 470582 451231
rect 470314 451179 470326 451185
rect 470378 451179 470390 451185
rect 470442 451179 470454 451185
rect 470506 451179 470518 451185
rect 470570 451179 470582 451185
rect 470634 451179 470646 451185
rect 470698 451179 470710 451185
rect 470762 451179 470774 451185
rect 470262 451173 470826 451179
rect 471716 450500 471744 453292
rect 471704 450494 471756 450500
rect 471704 450436 471756 450442
rect 469022 450401 469586 450407
rect 469074 450395 469086 450401
rect 469138 450395 469150 450401
rect 469202 450395 469214 450401
rect 469266 450395 469278 450401
rect 469330 450395 469342 450401
rect 469394 450395 469406 450401
rect 469458 450395 469470 450401
rect 469522 450395 469534 450401
rect 469266 450349 469276 450395
rect 469332 450349 469342 450395
rect 469022 450339 469036 450349
rect 469092 450339 469116 450349
rect 469172 450339 469196 450349
rect 469252 450339 469276 450349
rect 469332 450339 469356 450349
rect 469412 450339 469436 450349
rect 469492 450339 469516 450349
rect 469572 450339 469586 450349
rect 469022 450337 469586 450339
rect 469074 450315 469086 450337
rect 469138 450315 469150 450337
rect 469202 450315 469214 450337
rect 469266 450315 469278 450337
rect 469330 450315 469342 450337
rect 469394 450315 469406 450337
rect 469458 450315 469470 450337
rect 469522 450315 469534 450337
rect 469266 450285 469276 450315
rect 469332 450285 469342 450315
rect 469022 450273 469036 450285
rect 469092 450273 469116 450285
rect 469172 450273 469196 450285
rect 469252 450273 469276 450285
rect 469332 450273 469356 450285
rect 469412 450273 469436 450285
rect 469492 450273 469516 450285
rect 469572 450273 469586 450285
rect 469266 450259 469276 450273
rect 469332 450259 469342 450273
rect 469074 450235 469086 450259
rect 469138 450235 469150 450259
rect 469202 450235 469214 450259
rect 469266 450235 469278 450259
rect 469330 450235 469342 450259
rect 469394 450235 469406 450259
rect 469458 450235 469470 450259
rect 469522 450235 469534 450259
rect 469266 450221 469276 450235
rect 469332 450221 469342 450235
rect 469022 450209 469036 450221
rect 469092 450209 469116 450221
rect 469172 450209 469196 450221
rect 469252 450209 469276 450221
rect 469332 450209 469356 450221
rect 469412 450209 469436 450221
rect 469492 450209 469516 450221
rect 469572 450209 469586 450221
rect 469266 450179 469276 450209
rect 469332 450179 469342 450209
rect 469074 450157 469086 450179
rect 469138 450157 469150 450179
rect 469202 450157 469214 450179
rect 469266 450157 469278 450179
rect 469330 450157 469342 450179
rect 469394 450157 469406 450179
rect 469458 450157 469470 450179
rect 469522 450157 469534 450179
rect 469022 450155 469586 450157
rect 469022 450145 469036 450155
rect 469092 450145 469116 450155
rect 469172 450145 469196 450155
rect 469252 450145 469276 450155
rect 469332 450145 469356 450155
rect 469412 450145 469436 450155
rect 469492 450145 469516 450155
rect 469572 450145 469586 450155
rect 469266 450099 469276 450145
rect 469332 450099 469342 450145
rect 469074 450093 469086 450099
rect 469138 450093 469150 450099
rect 469202 450093 469214 450099
rect 469266 450093 469278 450099
rect 469330 450093 469342 450099
rect 469394 450093 469406 450099
rect 469458 450093 469470 450099
rect 469522 450093 469534 450099
rect 469022 450087 469586 450093
rect 470262 449316 470826 449322
rect 470314 449310 470326 449316
rect 470378 449310 470390 449316
rect 470442 449310 470454 449316
rect 470506 449310 470518 449316
rect 470570 449310 470582 449316
rect 470634 449310 470646 449316
rect 470698 449310 470710 449316
rect 470762 449310 470774 449316
rect 470506 449264 470516 449310
rect 470572 449264 470582 449310
rect 470262 449254 470276 449264
rect 470332 449254 470356 449264
rect 470412 449254 470436 449264
rect 470492 449254 470516 449264
rect 470572 449254 470596 449264
rect 470652 449254 470676 449264
rect 470732 449254 470756 449264
rect 470812 449254 470826 449264
rect 470262 449252 470826 449254
rect 470314 449230 470326 449252
rect 470378 449230 470390 449252
rect 470442 449230 470454 449252
rect 470506 449230 470518 449252
rect 470570 449230 470582 449252
rect 470634 449230 470646 449252
rect 470698 449230 470710 449252
rect 470762 449230 470774 449252
rect 470506 449200 470516 449230
rect 470572 449200 470582 449230
rect 470262 449188 470276 449200
rect 470332 449188 470356 449200
rect 470412 449188 470436 449200
rect 470492 449188 470516 449200
rect 470572 449188 470596 449200
rect 470652 449188 470676 449200
rect 470732 449188 470756 449200
rect 470812 449188 470826 449200
rect 470506 449174 470516 449188
rect 470572 449174 470582 449188
rect 470314 449150 470326 449174
rect 470378 449150 470390 449174
rect 470442 449150 470454 449174
rect 470506 449150 470518 449174
rect 470570 449150 470582 449174
rect 470634 449150 470646 449174
rect 470698 449150 470710 449174
rect 470762 449150 470774 449174
rect 470506 449136 470516 449150
rect 470572 449136 470582 449150
rect 470262 449124 470276 449136
rect 470332 449124 470356 449136
rect 470412 449124 470436 449136
rect 470492 449124 470516 449136
rect 470572 449124 470596 449136
rect 470652 449124 470676 449136
rect 470732 449124 470756 449136
rect 470812 449124 470826 449136
rect 470506 449094 470516 449124
rect 470572 449094 470582 449124
rect 470314 449072 470326 449094
rect 470378 449072 470390 449094
rect 470442 449072 470454 449094
rect 470506 449072 470518 449094
rect 470570 449072 470582 449094
rect 470634 449072 470646 449094
rect 470698 449072 470710 449094
rect 470762 449072 470774 449094
rect 470262 449070 470826 449072
rect 470262 449060 470276 449070
rect 470332 449060 470356 449070
rect 470412 449060 470436 449070
rect 470492 449060 470516 449070
rect 470572 449060 470596 449070
rect 470652 449060 470676 449070
rect 470732 449060 470756 449070
rect 470812 449060 470826 449070
rect 470506 449014 470516 449060
rect 470572 449014 470582 449060
rect 470314 449008 470326 449014
rect 470378 449008 470390 449014
rect 470442 449008 470454 449014
rect 470506 449008 470518 449014
rect 470570 449008 470582 449014
rect 470634 449008 470646 449014
rect 470698 449008 470710 449014
rect 470762 449008 470774 449014
rect 470262 449002 470826 449008
rect 471716 441616 471744 450436
rect 474108 450352 474554 450380
rect 474108 449723 474136 450352
rect 477843 450258 477899 450267
rect 477843 450193 477899 450202
rect 481160 450258 481216 450267
rect 481160 450193 481216 450202
rect 487793 450258 487849 450267
rect 487793 450193 487849 450202
rect 474094 449714 474150 449723
rect 474094 449649 474150 449658
rect 484511 449532 484539 450038
rect 483676 449504 484539 449532
rect 475384 449490 475436 449496
rect 475384 449432 475436 449438
rect 478696 449490 478748 449496
rect 478696 449432 478748 449438
rect 482008 449490 482060 449496
rect 482008 449432 482060 449438
rect 475396 445740 475424 449432
rect 478708 446284 478736 449432
rect 478696 446278 478748 446284
rect 478696 446220 478748 446226
rect 482020 445876 482048 449432
rect 482008 445870 482060 445876
rect 482008 445812 482060 445818
rect 475384 445734 475436 445740
rect 475384 445676 475436 445682
rect 471624 441588 471744 441616
rect 470262 433088 470826 433094
rect 470314 433082 470326 433088
rect 470378 433082 470390 433088
rect 470442 433082 470454 433088
rect 470506 433082 470518 433088
rect 470570 433082 470582 433088
rect 470634 433082 470646 433088
rect 470698 433082 470710 433088
rect 470762 433082 470774 433088
rect 470506 433036 470516 433082
rect 470572 433036 470582 433082
rect 470262 433026 470276 433036
rect 470332 433026 470356 433036
rect 470412 433026 470436 433036
rect 470492 433026 470516 433036
rect 470572 433026 470596 433036
rect 470652 433026 470676 433036
rect 470732 433026 470756 433036
rect 470812 433026 470826 433036
rect 470262 433024 470826 433026
rect 470314 433002 470326 433024
rect 470378 433002 470390 433024
rect 470442 433002 470454 433024
rect 470506 433002 470518 433024
rect 470570 433002 470582 433024
rect 470634 433002 470646 433024
rect 470698 433002 470710 433024
rect 470762 433002 470774 433024
rect 470506 432972 470516 433002
rect 470572 432972 470582 433002
rect 470262 432960 470276 432972
rect 470332 432960 470356 432972
rect 470412 432960 470436 432972
rect 470492 432960 470516 432972
rect 470572 432960 470596 432972
rect 470652 432960 470676 432972
rect 470732 432960 470756 432972
rect 470812 432960 470826 432972
rect 470506 432946 470516 432960
rect 470572 432946 470582 432960
rect 470314 432922 470326 432946
rect 470378 432922 470390 432946
rect 470442 432922 470454 432946
rect 470506 432922 470518 432946
rect 470570 432922 470582 432946
rect 470634 432922 470646 432946
rect 470698 432922 470710 432946
rect 470762 432922 470774 432946
rect 470506 432908 470516 432922
rect 470572 432908 470582 432922
rect 470262 432896 470276 432908
rect 470332 432896 470356 432908
rect 470412 432896 470436 432908
rect 470492 432896 470516 432908
rect 470572 432896 470596 432908
rect 470652 432896 470676 432908
rect 470732 432896 470756 432908
rect 470812 432896 470826 432908
rect 470506 432866 470516 432896
rect 470572 432866 470582 432896
rect 470314 432844 470326 432866
rect 470378 432844 470390 432866
rect 470442 432844 470454 432866
rect 470506 432844 470518 432866
rect 470570 432844 470582 432866
rect 470634 432844 470646 432866
rect 470698 432844 470710 432866
rect 470762 432844 470774 432866
rect 470262 432842 470826 432844
rect 470262 432832 470276 432842
rect 470332 432832 470356 432842
rect 470412 432832 470436 432842
rect 470492 432832 470516 432842
rect 470572 432832 470596 432842
rect 470652 432832 470676 432842
rect 470732 432832 470756 432842
rect 470812 432832 470826 432842
rect 470506 432786 470516 432832
rect 470572 432786 470582 432832
rect 470314 432780 470326 432786
rect 470378 432780 470390 432786
rect 470442 432780 470454 432786
rect 470506 432780 470518 432786
rect 470570 432780 470582 432786
rect 470634 432780 470646 432786
rect 470698 432780 470710 432786
rect 470762 432780 470774 432786
rect 470262 432774 470826 432780
rect 471624 432298 471652 441588
rect 483676 432859 483704 449504
rect 485320 449490 485372 449496
rect 485320 449432 485372 449438
rect 485332 445876 485360 449432
rect 491944 449406 491996 449412
rect 491944 449348 491996 449354
rect 485320 445870 485372 445876
rect 485320 445812 485372 445818
rect 490564 443014 490616 443020
rect 490564 442956 490616 442962
rect 483662 432850 483718 432859
rect 483662 432785 483718 432794
rect 483570 432306 483626 432315
rect 471612 432292 471664 432298
rect 483143 432264 483570 432292
rect 483570 432241 483626 432250
rect 471612 432234 471664 432240
rect 469022 432001 469586 432007
rect 469074 431995 469086 432001
rect 469138 431995 469150 432001
rect 469202 431995 469214 432001
rect 469266 431995 469278 432001
rect 469330 431995 469342 432001
rect 469394 431995 469406 432001
rect 469458 431995 469470 432001
rect 469522 431995 469534 432001
rect 469266 431949 469276 431995
rect 469332 431949 469342 431995
rect 471624 431956 471652 432234
rect 481270 432170 481326 432179
rect 481326 432128 481573 432156
rect 481270 432105 481326 432114
rect 469022 431939 469036 431949
rect 469092 431939 469116 431949
rect 469172 431939 469196 431949
rect 469252 431939 469276 431949
rect 469332 431939 469356 431949
rect 469412 431939 469436 431949
rect 469492 431939 469516 431949
rect 469572 431939 469586 431949
rect 469022 431937 469586 431939
rect 469074 431915 469086 431937
rect 469138 431915 469150 431937
rect 469202 431915 469214 431937
rect 469266 431915 469278 431937
rect 469330 431915 469342 431937
rect 469394 431915 469406 431937
rect 469458 431915 469470 431937
rect 469522 431915 469534 431937
rect 469266 431885 469276 431915
rect 469332 431885 469342 431915
rect 469022 431873 469036 431885
rect 469092 431873 469116 431885
rect 469172 431873 469196 431885
rect 469252 431873 469276 431885
rect 469332 431873 469356 431885
rect 469412 431873 469436 431885
rect 469492 431873 469516 431885
rect 469572 431873 469586 431885
rect 469266 431859 469276 431873
rect 469332 431859 469342 431873
rect 469074 431835 469086 431859
rect 469138 431835 469150 431859
rect 469202 431835 469214 431859
rect 469266 431835 469278 431859
rect 469330 431835 469342 431859
rect 469394 431835 469406 431859
rect 469458 431835 469470 431859
rect 469522 431835 469534 431859
rect 469266 431821 469276 431835
rect 469332 431821 469342 431835
rect 469022 431809 469036 431821
rect 469092 431809 469116 431821
rect 469172 431809 469196 431821
rect 469252 431809 469276 431821
rect 469332 431809 469356 431821
rect 469412 431809 469436 431821
rect 469492 431809 469516 431821
rect 469572 431809 469586 431821
rect 469266 431779 469276 431809
rect 469332 431779 469342 431809
rect 469074 431757 469086 431779
rect 469138 431757 469150 431779
rect 469202 431757 469214 431779
rect 469266 431757 469278 431779
rect 469330 431757 469342 431779
rect 469394 431757 469406 431779
rect 469458 431757 469470 431779
rect 469522 431757 469534 431779
rect 469022 431755 469586 431757
rect 469022 431745 469036 431755
rect 469092 431745 469116 431755
rect 469172 431745 469196 431755
rect 469252 431745 469276 431755
rect 469332 431745 469356 431755
rect 469412 431745 469436 431755
rect 469492 431745 469516 431755
rect 469572 431745 469586 431755
rect 469266 431699 469276 431745
rect 469332 431699 469342 431745
rect 469074 431693 469086 431699
rect 469138 431693 469150 431699
rect 469202 431693 469214 431699
rect 469266 431693 469278 431699
rect 469330 431693 469342 431699
rect 469394 431693 469406 431699
rect 469458 431693 469470 431699
rect 469522 431693 469534 431699
rect 469022 431687 469586 431693
rect 471256 431928 471652 431956
rect 474292 431992 474685 432020
rect 470262 430916 470826 430922
rect 470314 430910 470326 430916
rect 470378 430910 470390 430916
rect 470442 430910 470454 430916
rect 470506 430910 470518 430916
rect 470570 430910 470582 430916
rect 470634 430910 470646 430916
rect 470698 430910 470710 430916
rect 470762 430910 470774 430916
rect 470506 430864 470516 430910
rect 470572 430864 470582 430910
rect 470262 430854 470276 430864
rect 470332 430854 470356 430864
rect 470412 430854 470436 430864
rect 470492 430854 470516 430864
rect 470572 430854 470596 430864
rect 470652 430854 470676 430864
rect 470732 430854 470756 430864
rect 470812 430854 470826 430864
rect 470262 430852 470826 430854
rect 470314 430830 470326 430852
rect 470378 430830 470390 430852
rect 470442 430830 470454 430852
rect 470506 430830 470518 430852
rect 470570 430830 470582 430852
rect 470634 430830 470646 430852
rect 470698 430830 470710 430852
rect 470762 430830 470774 430852
rect 470506 430800 470516 430830
rect 470572 430800 470582 430830
rect 470262 430788 470276 430800
rect 470332 430788 470356 430800
rect 470412 430788 470436 430800
rect 470492 430788 470516 430800
rect 470572 430788 470596 430800
rect 470652 430788 470676 430800
rect 470732 430788 470756 430800
rect 470812 430788 470826 430800
rect 470506 430774 470516 430788
rect 470572 430774 470582 430788
rect 470314 430750 470326 430774
rect 470378 430750 470390 430774
rect 470442 430750 470454 430774
rect 470506 430750 470518 430774
rect 470570 430750 470582 430774
rect 470634 430750 470646 430774
rect 470698 430750 470710 430774
rect 470762 430750 470774 430774
rect 470506 430736 470516 430750
rect 470572 430736 470582 430750
rect 470262 430724 470276 430736
rect 470332 430724 470356 430736
rect 470412 430724 470436 430736
rect 470492 430724 470516 430736
rect 470572 430724 470596 430736
rect 470652 430724 470676 430736
rect 470732 430724 470756 430736
rect 470812 430724 470826 430736
rect 470506 430694 470516 430724
rect 470572 430694 470582 430724
rect 470314 430672 470326 430694
rect 470378 430672 470390 430694
rect 470442 430672 470454 430694
rect 470506 430672 470518 430694
rect 470570 430672 470582 430694
rect 470634 430672 470646 430694
rect 470698 430672 470710 430694
rect 470762 430672 470774 430694
rect 470262 430670 470826 430672
rect 470262 430660 470276 430670
rect 470332 430660 470356 430670
rect 470412 430660 470436 430670
rect 470492 430660 470516 430670
rect 470572 430660 470596 430670
rect 470652 430660 470676 430670
rect 470732 430660 470756 430670
rect 470812 430660 470826 430670
rect 470506 430614 470516 430660
rect 470572 430614 470582 430660
rect 470314 430608 470326 430614
rect 470378 430608 470390 430614
rect 470442 430608 470454 430614
rect 470506 430608 470518 430614
rect 470570 430608 470582 430614
rect 470634 430608 470646 430614
rect 470698 430608 470710 430614
rect 470762 430608 470774 430614
rect 470262 430602 470826 430608
rect 470262 412088 470826 412094
rect 470314 412082 470326 412088
rect 470378 412082 470390 412088
rect 470442 412082 470454 412088
rect 470506 412082 470518 412088
rect 470570 412082 470582 412088
rect 470634 412082 470646 412088
rect 470698 412082 470710 412088
rect 470762 412082 470774 412088
rect 470506 412036 470516 412082
rect 470572 412036 470582 412082
rect 470262 412026 470276 412036
rect 470332 412026 470356 412036
rect 470412 412026 470436 412036
rect 470492 412026 470516 412036
rect 470572 412026 470596 412036
rect 470652 412026 470676 412036
rect 470732 412026 470756 412036
rect 470812 412026 470826 412036
rect 470262 412024 470826 412026
rect 470314 412002 470326 412024
rect 470378 412002 470390 412024
rect 470442 412002 470454 412024
rect 470506 412002 470518 412024
rect 470570 412002 470582 412024
rect 470634 412002 470646 412024
rect 470698 412002 470710 412024
rect 470762 412002 470774 412024
rect 470506 411972 470516 412002
rect 470572 411972 470582 412002
rect 470262 411960 470276 411972
rect 470332 411960 470356 411972
rect 470412 411960 470436 411972
rect 470492 411960 470516 411972
rect 470572 411960 470596 411972
rect 470652 411960 470676 411972
rect 470732 411960 470756 411972
rect 470812 411960 470826 411972
rect 470506 411946 470516 411960
rect 470572 411946 470582 411960
rect 470314 411922 470326 411946
rect 470378 411922 470390 411946
rect 470442 411922 470454 411946
rect 470506 411922 470518 411946
rect 470570 411922 470582 411946
rect 470634 411922 470646 411946
rect 470698 411922 470710 411946
rect 470762 411922 470774 411946
rect 470506 411908 470516 411922
rect 470572 411908 470582 411922
rect 470262 411896 470276 411908
rect 470332 411896 470356 411908
rect 470412 411896 470436 411908
rect 470492 411896 470516 411908
rect 470572 411896 470596 411908
rect 470652 411896 470676 411908
rect 470732 411896 470756 411908
rect 470812 411896 470826 411908
rect 470506 411866 470516 411896
rect 470572 411866 470582 411896
rect 470314 411844 470326 411866
rect 470378 411844 470390 411866
rect 470442 411844 470454 411866
rect 470506 411844 470518 411866
rect 470570 411844 470582 411866
rect 470634 411844 470646 411866
rect 470698 411844 470710 411866
rect 470762 411844 470774 411866
rect 470262 411842 470826 411844
rect 470262 411832 470276 411842
rect 470332 411832 470356 411842
rect 470412 411832 470436 411842
rect 470492 411832 470516 411842
rect 470572 411832 470596 411842
rect 470652 411832 470676 411842
rect 470732 411832 470756 411842
rect 470812 411832 470826 411842
rect 470506 411786 470516 411832
rect 470572 411786 470582 411832
rect 470314 411780 470326 411786
rect 470378 411780 470390 411786
rect 470442 411780 470454 411786
rect 470506 411780 470518 411786
rect 470570 411780 470582 411786
rect 470634 411780 470646 411786
rect 470698 411780 470710 411786
rect 470762 411780 470774 411786
rect 470262 411774 470826 411780
rect 471256 411264 471284 431928
rect 474292 431907 474320 431992
rect 474278 431898 474334 431907
rect 474278 431833 474334 431842
rect 478102 431626 478158 431635
rect 478102 431561 478158 431570
rect 488433 431626 488489 431635
rect 488433 431561 488489 431570
rect 478972 431454 479024 431460
rect 478972 431396 479024 431402
rect 485780 431454 485832 431460
rect 485780 431396 485832 431402
rect 475476 431089 475528 431095
rect 475476 431031 475528 431037
rect 475488 429148 475516 431031
rect 475476 429142 475528 429148
rect 475476 429084 475528 429090
rect 478984 427963 479012 431396
rect 482376 431089 482428 431095
rect 482376 431031 482428 431037
rect 478970 427954 479026 427963
rect 478970 427889 479026 427898
rect 482388 427856 482416 431031
rect 485792 427963 485820 431396
rect 490576 429148 490604 442956
rect 490564 429142 490616 429148
rect 490564 429084 490616 429090
rect 485778 427954 485834 427963
rect 485778 427889 485834 427898
rect 482376 427850 482428 427856
rect 482376 427792 482428 427798
rect 488538 413946 488594 413955
rect 488538 413881 488594 413890
rect 473728 411286 473780 411292
rect 471244 411258 471296 411264
rect 473728 411228 473780 411234
rect 471244 411200 471296 411206
rect 469022 411002 469586 411008
rect 469074 410996 469086 411002
rect 469138 410996 469150 411002
rect 469202 410996 469214 411002
rect 469266 410996 469278 411002
rect 469330 410996 469342 411002
rect 469394 410996 469406 411002
rect 469458 410996 469470 411002
rect 469522 410996 469534 411002
rect 469266 410950 469276 410996
rect 469332 410950 469342 410996
rect 469022 410940 469036 410950
rect 469092 410940 469116 410950
rect 469172 410940 469196 410950
rect 469252 410940 469276 410950
rect 469332 410940 469356 410950
rect 469412 410940 469436 410950
rect 469492 410940 469516 410950
rect 469572 410940 469586 410950
rect 469022 410938 469586 410940
rect 469074 410916 469086 410938
rect 469138 410916 469150 410938
rect 469202 410916 469214 410938
rect 469266 410916 469278 410938
rect 469330 410916 469342 410938
rect 469394 410916 469406 410938
rect 469458 410916 469470 410938
rect 469522 410916 469534 410938
rect 469266 410886 469276 410916
rect 469332 410886 469342 410916
rect 469022 410874 469036 410886
rect 469092 410874 469116 410886
rect 469172 410874 469196 410886
rect 469252 410874 469276 410886
rect 469332 410874 469356 410886
rect 469412 410874 469436 410886
rect 469492 410874 469516 410886
rect 469572 410874 469586 410886
rect 469266 410860 469276 410874
rect 469332 410860 469342 410874
rect 469074 410836 469086 410860
rect 469138 410836 469150 410860
rect 469202 410836 469214 410860
rect 469266 410836 469278 410860
rect 469330 410836 469342 410860
rect 469394 410836 469406 410860
rect 469458 410836 469470 410860
rect 469522 410836 469534 410860
rect 469266 410822 469276 410836
rect 469332 410822 469342 410836
rect 469022 410810 469036 410822
rect 469092 410810 469116 410822
rect 469172 410810 469196 410822
rect 469252 410810 469276 410822
rect 469332 410810 469356 410822
rect 469412 410810 469436 410822
rect 469492 410810 469516 410822
rect 469572 410810 469586 410822
rect 469266 410780 469276 410810
rect 469332 410780 469342 410810
rect 469074 410758 469086 410780
rect 469138 410758 469150 410780
rect 469202 410758 469214 410780
rect 469266 410758 469278 410780
rect 469330 410758 469342 410780
rect 469394 410758 469406 410780
rect 469458 410758 469470 410780
rect 469522 410758 469534 410780
rect 469022 410756 469586 410758
rect 469022 410746 469036 410756
rect 469092 410746 469116 410756
rect 469172 410746 469196 410756
rect 469252 410746 469276 410756
rect 469332 410746 469356 410756
rect 469412 410746 469436 410756
rect 469492 410746 469516 410756
rect 469572 410746 469586 410756
rect 469266 410700 469276 410746
rect 469332 410700 469342 410746
rect 469074 410694 469086 410700
rect 469138 410694 469150 410700
rect 469202 410694 469214 410700
rect 469266 410694 469278 410700
rect 469330 410694 469342 410700
rect 469394 410694 469406 410700
rect 469458 410694 469470 410700
rect 469522 410694 469534 410700
rect 469022 410688 469586 410694
rect 470262 409916 470826 409922
rect 470314 409910 470326 409916
rect 470378 409910 470390 409916
rect 470442 409910 470454 409916
rect 470506 409910 470518 409916
rect 470570 409910 470582 409916
rect 470634 409910 470646 409916
rect 470698 409910 470710 409916
rect 470762 409910 470774 409916
rect 470506 409864 470516 409910
rect 470572 409864 470582 409910
rect 470262 409854 470276 409864
rect 470332 409854 470356 409864
rect 470412 409854 470436 409864
rect 470492 409854 470516 409864
rect 470572 409854 470596 409864
rect 470652 409854 470676 409864
rect 470732 409854 470756 409864
rect 470812 409854 470826 409864
rect 470262 409852 470826 409854
rect 470314 409830 470326 409852
rect 470378 409830 470390 409852
rect 470442 409830 470454 409852
rect 470506 409830 470518 409852
rect 470570 409830 470582 409852
rect 470634 409830 470646 409852
rect 470698 409830 470710 409852
rect 470762 409830 470774 409852
rect 470506 409800 470516 409830
rect 470572 409800 470582 409830
rect 470262 409788 470276 409800
rect 470332 409788 470356 409800
rect 470412 409788 470436 409800
rect 470492 409788 470516 409800
rect 470572 409788 470596 409800
rect 470652 409788 470676 409800
rect 470732 409788 470756 409800
rect 470812 409788 470826 409800
rect 470506 409774 470516 409788
rect 470572 409774 470582 409788
rect 470314 409750 470326 409774
rect 470378 409750 470390 409774
rect 470442 409750 470454 409774
rect 470506 409750 470518 409774
rect 470570 409750 470582 409774
rect 470634 409750 470646 409774
rect 470698 409750 470710 409774
rect 470762 409750 470774 409774
rect 470506 409736 470516 409750
rect 470572 409736 470582 409750
rect 470262 409724 470276 409736
rect 470332 409724 470356 409736
rect 470412 409724 470436 409736
rect 470492 409724 470516 409736
rect 470572 409724 470596 409736
rect 470652 409724 470676 409736
rect 470732 409724 470756 409736
rect 470812 409724 470826 409736
rect 470506 409694 470516 409724
rect 470572 409694 470582 409724
rect 470314 409672 470326 409694
rect 470378 409672 470390 409694
rect 470442 409672 470454 409694
rect 470506 409672 470518 409694
rect 470570 409672 470582 409694
rect 470634 409672 470646 409694
rect 470698 409672 470710 409694
rect 470762 409672 470774 409694
rect 470262 409670 470826 409672
rect 470262 409660 470276 409670
rect 470332 409660 470356 409670
rect 470412 409660 470436 409670
rect 470492 409660 470516 409670
rect 470572 409660 470596 409670
rect 470652 409660 470676 409670
rect 470732 409660 470756 409670
rect 470812 409660 470826 409670
rect 470506 409614 470516 409660
rect 470572 409614 470582 409660
rect 470314 409608 470326 409614
rect 470378 409608 470390 409614
rect 470442 409608 470454 409614
rect 470506 409608 470518 409614
rect 470570 409608 470582 409614
rect 470634 409608 470646 409614
rect 470698 409608 470710 409614
rect 470762 409608 470774 409614
rect 470262 409602 470826 409608
rect 470262 391089 470826 391095
rect 470314 391083 470326 391089
rect 470378 391083 470390 391089
rect 470442 391083 470454 391089
rect 470506 391083 470518 391089
rect 470570 391083 470582 391089
rect 470634 391083 470646 391089
rect 470698 391083 470710 391089
rect 470762 391083 470774 391089
rect 470506 391037 470516 391083
rect 470572 391037 470582 391083
rect 470262 391027 470276 391037
rect 470332 391027 470356 391037
rect 470412 391027 470436 391037
rect 470492 391027 470516 391037
rect 470572 391027 470596 391037
rect 470652 391027 470676 391037
rect 470732 391027 470756 391037
rect 470812 391027 470826 391037
rect 470262 391025 470826 391027
rect 470314 391003 470326 391025
rect 470378 391003 470390 391025
rect 470442 391003 470454 391025
rect 470506 391003 470518 391025
rect 470570 391003 470582 391025
rect 470634 391003 470646 391025
rect 470698 391003 470710 391025
rect 470762 391003 470774 391025
rect 470506 390973 470516 391003
rect 470572 390973 470582 391003
rect 470262 390961 470276 390973
rect 470332 390961 470356 390973
rect 470412 390961 470436 390973
rect 470492 390961 470516 390973
rect 470572 390961 470596 390973
rect 470652 390961 470676 390973
rect 470732 390961 470756 390973
rect 470812 390961 470826 390973
rect 470506 390947 470516 390961
rect 470572 390947 470582 390961
rect 470314 390923 470326 390947
rect 470378 390923 470390 390947
rect 470442 390923 470454 390947
rect 470506 390923 470518 390947
rect 470570 390923 470582 390947
rect 470634 390923 470646 390947
rect 470698 390923 470710 390947
rect 470762 390923 470774 390947
rect 470506 390909 470516 390923
rect 470572 390909 470582 390923
rect 470262 390897 470276 390909
rect 470332 390897 470356 390909
rect 470412 390897 470436 390909
rect 470492 390897 470516 390909
rect 470572 390897 470596 390909
rect 470652 390897 470676 390909
rect 470732 390897 470756 390909
rect 470812 390897 470826 390909
rect 470506 390867 470516 390897
rect 470572 390867 470582 390897
rect 470314 390845 470326 390867
rect 470378 390845 470390 390867
rect 470442 390845 470454 390867
rect 470506 390845 470518 390867
rect 470570 390845 470582 390867
rect 470634 390845 470646 390867
rect 470698 390845 470710 390867
rect 470762 390845 470774 390867
rect 470262 390843 470826 390845
rect 470262 390833 470276 390843
rect 470332 390833 470356 390843
rect 470412 390833 470436 390843
rect 470492 390833 470516 390843
rect 470572 390833 470596 390843
rect 470652 390833 470676 390843
rect 470732 390833 470756 390843
rect 470812 390833 470826 390843
rect 470506 390787 470516 390833
rect 470572 390787 470582 390833
rect 470314 390781 470326 390787
rect 470378 390781 470390 390787
rect 470442 390781 470454 390787
rect 470506 390781 470518 390787
rect 470570 390781 470582 390787
rect 470634 390781 470646 390787
rect 470698 390781 470710 390787
rect 470762 390781 470774 390787
rect 470262 390775 470826 390781
rect 471256 390320 471284 411200
rect 473740 410963 473768 411228
rect 473726 410954 473782 410963
rect 473726 410889 473782 410898
rect 478420 410442 478472 410448
rect 478420 410384 478472 410390
rect 478604 410442 478656 410448
rect 478604 410384 478656 410390
rect 478432 410147 478460 410384
rect 478418 410138 478474 410147
rect 475292 410090 475344 410096
rect 478418 410073 478474 410082
rect 475292 410032 475344 410038
rect 475304 408476 475332 410032
rect 475292 408470 475344 408476
rect 475292 408412 475344 408418
rect 478616 407116 478644 410384
rect 481019 410260 481047 410518
rect 484136 410504 484298 410532
rect 484136 410419 484164 410504
rect 485136 410442 485188 410448
rect 484122 410410 484178 410419
rect 485136 410384 485188 410390
rect 484122 410345 484178 410354
rect 481019 410232 481128 410260
rect 481100 410124 481128 410232
rect 481362 410138 481418 410147
rect 481100 410096 481362 410124
rect 481362 410073 481418 410082
rect 481824 410090 481876 410096
rect 481824 410032 481876 410038
rect 481836 407155 481864 410032
rect 485148 407155 485176 410384
rect 487549 410260 487577 410518
rect 487549 410232 487660 410260
rect 487632 410011 487660 410232
rect 488552 410011 488580 413881
rect 490748 410034 490800 410040
rect 487618 410002 487674 410011
rect 487618 409937 487674 409946
rect 488538 410002 488594 410011
rect 488538 409937 488594 409946
rect 489826 410002 489882 410011
rect 490748 409976 490800 409982
rect 489826 409937 489882 409946
rect 481822 407146 481878 407155
rect 478604 407110 478656 407116
rect 481822 407081 481878 407090
rect 485134 407146 485190 407155
rect 485134 407081 485190 407090
rect 478604 407052 478656 407058
rect 489840 392059 489868 409937
rect 489826 392050 489882 392059
rect 489826 391985 489882 391994
rect 471244 390314 471296 390320
rect 471244 390256 471296 390262
rect 471704 390110 471756 390116
rect 471704 390052 471756 390058
rect 469022 390006 469586 390012
rect 469074 390000 469086 390006
rect 469138 390000 469150 390006
rect 469202 390000 469214 390006
rect 469266 390000 469278 390006
rect 469330 390000 469342 390006
rect 469394 390000 469406 390006
rect 469458 390000 469470 390006
rect 469522 390000 469534 390006
rect 469266 389954 469276 390000
rect 469332 389954 469342 390000
rect 469022 389944 469036 389954
rect 469092 389944 469116 389954
rect 469172 389944 469196 389954
rect 469252 389944 469276 389954
rect 469332 389944 469356 389954
rect 469412 389944 469436 389954
rect 469492 389944 469516 389954
rect 469572 389944 469586 389954
rect 469022 389942 469586 389944
rect 469074 389920 469086 389942
rect 469138 389920 469150 389942
rect 469202 389920 469214 389942
rect 469266 389920 469278 389942
rect 469330 389920 469342 389942
rect 469394 389920 469406 389942
rect 469458 389920 469470 389942
rect 469522 389920 469534 389942
rect 469266 389890 469276 389920
rect 469332 389890 469342 389920
rect 469022 389878 469036 389890
rect 469092 389878 469116 389890
rect 469172 389878 469196 389890
rect 469252 389878 469276 389890
rect 469332 389878 469356 389890
rect 469412 389878 469436 389890
rect 469492 389878 469516 389890
rect 469572 389878 469586 389890
rect 469266 389864 469276 389878
rect 469332 389864 469342 389878
rect 469074 389840 469086 389864
rect 469138 389840 469150 389864
rect 469202 389840 469214 389864
rect 469266 389840 469278 389864
rect 469330 389840 469342 389864
rect 469394 389840 469406 389864
rect 469458 389840 469470 389864
rect 469522 389840 469534 389864
rect 469266 389826 469276 389840
rect 469332 389826 469342 389840
rect 469022 389814 469036 389826
rect 469092 389814 469116 389826
rect 469172 389814 469196 389826
rect 469252 389814 469276 389826
rect 469332 389814 469356 389826
rect 469412 389814 469436 389826
rect 469492 389814 469516 389826
rect 469572 389814 469586 389826
rect 469266 389784 469276 389814
rect 469332 389784 469342 389814
rect 469074 389762 469086 389784
rect 469138 389762 469150 389784
rect 469202 389762 469214 389784
rect 469266 389762 469278 389784
rect 469330 389762 469342 389784
rect 469394 389762 469406 389784
rect 469458 389762 469470 389784
rect 469522 389762 469534 389784
rect 469022 389760 469586 389762
rect 469022 389750 469036 389760
rect 469092 389750 469116 389760
rect 469172 389750 469196 389760
rect 469252 389750 469276 389760
rect 469332 389750 469356 389760
rect 469412 389750 469436 389760
rect 469492 389750 469516 389760
rect 469572 389750 469586 389760
rect 469266 389704 469276 389750
rect 469332 389704 469342 389750
rect 469074 389698 469086 389704
rect 469138 389698 469150 389704
rect 469202 389698 469214 389704
rect 469266 389698 469278 389704
rect 469330 389698 469342 389704
rect 469394 389698 469406 389704
rect 469458 389698 469470 389704
rect 469522 389698 469534 389704
rect 469022 389692 469586 389698
rect 470262 388916 470826 388922
rect 470314 388910 470326 388916
rect 470378 388910 470390 388916
rect 470442 388910 470454 388916
rect 470506 388910 470518 388916
rect 470570 388910 470582 388916
rect 470634 388910 470646 388916
rect 470698 388910 470710 388916
rect 470762 388910 470774 388916
rect 470506 388864 470516 388910
rect 470572 388864 470582 388910
rect 470262 388854 470276 388864
rect 470332 388854 470356 388864
rect 470412 388854 470436 388864
rect 470492 388854 470516 388864
rect 470572 388854 470596 388864
rect 470652 388854 470676 388864
rect 470732 388854 470756 388864
rect 470812 388854 470826 388864
rect 470262 388852 470826 388854
rect 470314 388830 470326 388852
rect 470378 388830 470390 388852
rect 470442 388830 470454 388852
rect 470506 388830 470518 388852
rect 470570 388830 470582 388852
rect 470634 388830 470646 388852
rect 470698 388830 470710 388852
rect 470762 388830 470774 388852
rect 470506 388800 470516 388830
rect 470572 388800 470582 388830
rect 470262 388788 470276 388800
rect 470332 388788 470356 388800
rect 470412 388788 470436 388800
rect 470492 388788 470516 388800
rect 470572 388788 470596 388800
rect 470652 388788 470676 388800
rect 470732 388788 470756 388800
rect 470812 388788 470826 388800
rect 470506 388774 470516 388788
rect 470572 388774 470582 388788
rect 470314 388750 470326 388774
rect 470378 388750 470390 388774
rect 470442 388750 470454 388774
rect 470506 388750 470518 388774
rect 470570 388750 470582 388774
rect 470634 388750 470646 388774
rect 470698 388750 470710 388774
rect 470762 388750 470774 388774
rect 470506 388736 470516 388750
rect 470572 388736 470582 388750
rect 470262 388724 470276 388736
rect 470332 388724 470356 388736
rect 470412 388724 470436 388736
rect 470492 388724 470516 388736
rect 470572 388724 470596 388736
rect 470652 388724 470676 388736
rect 470732 388724 470756 388736
rect 470812 388724 470826 388736
rect 470506 388694 470516 388724
rect 470572 388694 470582 388724
rect 470314 388672 470326 388694
rect 470378 388672 470390 388694
rect 470442 388672 470454 388694
rect 470506 388672 470518 388694
rect 470570 388672 470582 388694
rect 470634 388672 470646 388694
rect 470698 388672 470710 388694
rect 470762 388672 470774 388694
rect 470262 388670 470826 388672
rect 470262 388660 470276 388670
rect 470332 388660 470356 388670
rect 470412 388660 470436 388670
rect 470492 388660 470516 388670
rect 470572 388660 470596 388670
rect 470652 388660 470676 388670
rect 470732 388660 470756 388670
rect 470812 388660 470826 388670
rect 470506 388614 470516 388660
rect 470572 388614 470582 388660
rect 470314 388608 470326 388614
rect 470378 388608 470390 388614
rect 470442 388608 470454 388614
rect 470506 388608 470518 388614
rect 470570 388608 470582 388614
rect 470634 388608 470646 388614
rect 470698 388608 470710 388614
rect 470762 388608 470774 388614
rect 470262 388602 470826 388608
rect 470262 358489 470826 358495
rect 470314 358483 470326 358489
rect 470378 358483 470390 358489
rect 470442 358483 470454 358489
rect 470506 358483 470518 358489
rect 470570 358483 470582 358489
rect 470634 358483 470646 358489
rect 470698 358483 470710 358489
rect 470762 358483 470774 358489
rect 470506 358437 470516 358483
rect 470572 358437 470582 358483
rect 470262 358427 470276 358437
rect 470332 358427 470356 358437
rect 470412 358427 470436 358437
rect 470492 358427 470516 358437
rect 470572 358427 470596 358437
rect 470652 358427 470676 358437
rect 470732 358427 470756 358437
rect 470812 358427 470826 358437
rect 470262 358425 470826 358427
rect 470314 358403 470326 358425
rect 470378 358403 470390 358425
rect 470442 358403 470454 358425
rect 470506 358403 470518 358425
rect 470570 358403 470582 358425
rect 470634 358403 470646 358425
rect 470698 358403 470710 358425
rect 470762 358403 470774 358425
rect 470506 358373 470516 358403
rect 470572 358373 470582 358403
rect 470262 358361 470276 358373
rect 470332 358361 470356 358373
rect 470412 358361 470436 358373
rect 470492 358361 470516 358373
rect 470572 358361 470596 358373
rect 470652 358361 470676 358373
rect 470732 358361 470756 358373
rect 470812 358361 470826 358373
rect 470506 358347 470516 358361
rect 470572 358347 470582 358361
rect 470314 358323 470326 358347
rect 470378 358323 470390 358347
rect 470442 358323 470454 358347
rect 470506 358323 470518 358347
rect 470570 358323 470582 358347
rect 470634 358323 470646 358347
rect 470698 358323 470710 358347
rect 470762 358323 470774 358347
rect 470506 358309 470516 358323
rect 470572 358309 470582 358323
rect 470262 358297 470276 358309
rect 470332 358297 470356 358309
rect 470412 358297 470436 358309
rect 470492 358297 470516 358309
rect 470572 358297 470596 358309
rect 470652 358297 470676 358309
rect 470732 358297 470756 358309
rect 470812 358297 470826 358309
rect 470506 358267 470516 358297
rect 470572 358267 470582 358297
rect 470314 358245 470326 358267
rect 470378 358245 470390 358267
rect 470442 358245 470454 358267
rect 470506 358245 470518 358267
rect 470570 358245 470582 358267
rect 470634 358245 470646 358267
rect 470698 358245 470710 358267
rect 470762 358245 470774 358267
rect 470262 358243 470826 358245
rect 470262 358233 470276 358243
rect 470332 358233 470356 358243
rect 470412 358233 470436 358243
rect 470492 358233 470516 358243
rect 470572 358233 470596 358243
rect 470652 358233 470676 358243
rect 470732 358233 470756 358243
rect 470812 358233 470826 358243
rect 470506 358187 470516 358233
rect 470572 358187 470582 358233
rect 470314 358181 470326 358187
rect 470378 358181 470390 358187
rect 470442 358181 470454 358187
rect 470506 358181 470518 358187
rect 470570 358181 470582 358187
rect 470634 358181 470646 358187
rect 470698 358181 470710 358187
rect 470762 358181 470774 358187
rect 470262 358175 470826 358181
rect 471716 357612 471744 390052
rect 479432 389498 479484 389504
rect 479432 389440 479484 389446
rect 482098 389466 482154 389475
rect 474936 389339 474964 389438
rect 478648 389339 478676 389438
rect 474922 389330 474978 389339
rect 474922 389265 474978 389274
rect 478634 389330 478690 389339
rect 478634 389265 478690 389274
rect 475752 389090 475804 389096
rect 475752 389032 475804 389038
rect 475764 387804 475792 389032
rect 479444 387804 479472 389440
rect 489366 389466 489422 389475
rect 482154 389424 482374 389452
rect 482098 389401 482154 389410
rect 489422 389424 489798 389452
rect 489366 389401 489422 389410
rect 483204 389090 483256 389096
rect 483204 389032 483256 389038
rect 486884 389090 486936 389096
rect 486884 389032 486936 389038
rect 475752 387798 475804 387804
rect 475752 387740 475804 387746
rect 479432 387798 479484 387804
rect 479432 387740 479484 387746
rect 483216 386444 483244 389032
rect 486896 386483 486924 389032
rect 486882 386474 486938 386483
rect 483204 386438 483256 386444
rect 483204 386380 483256 386386
rect 484308 386438 484360 386444
rect 486882 386409 486938 386418
rect 484308 386380 484360 386386
rect 484320 369852 484348 386380
rect 484308 369846 484360 369852
rect 484308 369788 484360 369794
rect 478878 358050 478934 358059
rect 478878 357985 478934 357994
rect 481822 358050 481878 358059
rect 481822 357985 481878 357994
rect 484950 358050 485006 358059
rect 484950 357985 485006 357994
rect 488446 358050 488502 358059
rect 488446 357985 488502 357994
rect 478892 357691 478920 357985
rect 481836 357691 481864 357985
rect 484964 357691 484992 357985
rect 488460 357764 488488 357985
rect 488460 357736 488501 357764
rect 478880 357685 478932 357691
rect 475108 357674 475160 357680
rect 478880 357627 478932 357633
rect 481824 357685 481876 357691
rect 481824 357627 481876 357633
rect 484952 357685 485004 357691
rect 484952 357627 485004 357633
rect 475108 357616 475160 357622
rect 471704 357606 471756 357612
rect 471704 357548 471756 357554
rect 469022 357403 469586 357409
rect 469074 357397 469086 357403
rect 469138 357397 469150 357403
rect 469202 357397 469214 357403
rect 469266 357397 469278 357403
rect 469330 357397 469342 357403
rect 469394 357397 469406 357403
rect 469458 357397 469470 357403
rect 469522 357397 469534 357403
rect 469266 357351 469276 357397
rect 469332 357351 469342 357397
rect 469022 357341 469036 357351
rect 469092 357341 469116 357351
rect 469172 357341 469196 357351
rect 469252 357341 469276 357351
rect 469332 357341 469356 357351
rect 469412 357341 469436 357351
rect 469492 357341 469516 357351
rect 469572 357341 469586 357351
rect 469022 357339 469586 357341
rect 469074 357317 469086 357339
rect 469138 357317 469150 357339
rect 469202 357317 469214 357339
rect 469266 357317 469278 357339
rect 469330 357317 469342 357339
rect 469394 357317 469406 357339
rect 469458 357317 469470 357339
rect 469522 357317 469534 357339
rect 469266 357287 469276 357317
rect 469332 357287 469342 357317
rect 469022 357275 469036 357287
rect 469092 357275 469116 357287
rect 469172 357275 469196 357287
rect 469252 357275 469276 357287
rect 469332 357275 469356 357287
rect 469412 357275 469436 357287
rect 469492 357275 469516 357287
rect 469572 357275 469586 357287
rect 469266 357261 469276 357275
rect 469332 357261 469342 357275
rect 469074 357237 469086 357261
rect 469138 357237 469150 357261
rect 469202 357237 469214 357261
rect 469266 357237 469278 357261
rect 469330 357237 469342 357261
rect 469394 357237 469406 357261
rect 469458 357237 469470 357261
rect 469522 357237 469534 357261
rect 469266 357223 469276 357237
rect 469332 357223 469342 357237
rect 469022 357211 469036 357223
rect 469092 357211 469116 357223
rect 469172 357211 469196 357223
rect 469252 357211 469276 357223
rect 469332 357211 469356 357223
rect 469412 357211 469436 357223
rect 469492 357211 469516 357223
rect 469572 357211 469586 357223
rect 469266 357181 469276 357211
rect 469332 357181 469342 357211
rect 469074 357159 469086 357181
rect 469138 357159 469150 357181
rect 469202 357159 469214 357181
rect 469266 357159 469278 357181
rect 469330 357159 469342 357181
rect 469394 357159 469406 357181
rect 469458 357159 469470 357181
rect 469522 357159 469534 357181
rect 469022 357157 469586 357159
rect 469022 357147 469036 357157
rect 469092 357147 469116 357157
rect 469172 357147 469196 357157
rect 469252 357147 469276 357157
rect 469332 357147 469356 357157
rect 469412 357147 469436 357157
rect 469492 357147 469516 357157
rect 469572 357147 469586 357157
rect 469266 357101 469276 357147
rect 469332 357101 469342 357147
rect 469074 357095 469086 357101
rect 469138 357095 469150 357101
rect 469202 357095 469214 357101
rect 469266 357095 469278 357101
rect 469330 357095 469342 357101
rect 469394 357095 469406 357101
rect 469458 357095 469470 357101
rect 469522 357095 469534 357101
rect 469022 357089 469586 357095
rect 470262 356316 470826 356322
rect 470314 356310 470326 356316
rect 470378 356310 470390 356316
rect 470442 356310 470454 356316
rect 470506 356310 470518 356316
rect 470570 356310 470582 356316
rect 470634 356310 470646 356316
rect 470698 356310 470710 356316
rect 470762 356310 470774 356316
rect 470506 356264 470516 356310
rect 470572 356264 470582 356310
rect 470262 356254 470276 356264
rect 470332 356254 470356 356264
rect 470412 356254 470436 356264
rect 470492 356254 470516 356264
rect 470572 356254 470596 356264
rect 470652 356254 470676 356264
rect 470732 356254 470756 356264
rect 470812 356254 470826 356264
rect 470262 356252 470826 356254
rect 470314 356230 470326 356252
rect 470378 356230 470390 356252
rect 470442 356230 470454 356252
rect 470506 356230 470518 356252
rect 470570 356230 470582 356252
rect 470634 356230 470646 356252
rect 470698 356230 470710 356252
rect 470762 356230 470774 356252
rect 470506 356200 470516 356230
rect 470572 356200 470582 356230
rect 470262 356188 470276 356200
rect 470332 356188 470356 356200
rect 470412 356188 470436 356200
rect 470492 356188 470516 356200
rect 470572 356188 470596 356200
rect 470652 356188 470676 356200
rect 470732 356188 470756 356200
rect 470812 356188 470826 356200
rect 470506 356174 470516 356188
rect 470572 356174 470582 356188
rect 470314 356150 470326 356174
rect 470378 356150 470390 356174
rect 470442 356150 470454 356174
rect 470506 356150 470518 356174
rect 470570 356150 470582 356174
rect 470634 356150 470646 356174
rect 470698 356150 470710 356174
rect 470762 356150 470774 356174
rect 470506 356136 470516 356150
rect 470572 356136 470582 356150
rect 470262 356124 470276 356136
rect 470332 356124 470356 356136
rect 470412 356124 470436 356136
rect 470492 356124 470516 356136
rect 470572 356124 470596 356136
rect 470652 356124 470676 356136
rect 470732 356124 470756 356136
rect 470812 356124 470826 356136
rect 470506 356094 470516 356124
rect 470572 356094 470582 356124
rect 470314 356072 470326 356094
rect 470378 356072 470390 356094
rect 470442 356072 470454 356094
rect 470506 356072 470518 356094
rect 470570 356072 470582 356094
rect 470634 356072 470646 356094
rect 470698 356072 470710 356094
rect 470762 356072 470774 356094
rect 470262 356070 470826 356072
rect 470262 356060 470276 356070
rect 470332 356060 470356 356070
rect 470412 356060 470436 356070
rect 470492 356060 470516 356070
rect 470572 356060 470596 356070
rect 470652 356060 470676 356070
rect 470732 356060 470756 356070
rect 470812 356060 470826 356070
rect 470506 356014 470516 356060
rect 470572 356014 470582 356060
rect 470314 356008 470326 356014
rect 470378 356008 470390 356014
rect 470442 356008 470454 356014
rect 470506 356008 470518 356014
rect 470570 356008 470582 356014
rect 470634 356008 470646 356014
rect 470698 356008 470710 356014
rect 470762 356008 470774 356014
rect 470262 356002 470826 356008
rect 471716 354676 471744 357548
rect 475014 357506 475070 357515
rect 475120 357492 475148 357616
rect 488473 357614 488501 357736
rect 475070 357464 475148 357492
rect 475014 357441 475070 357450
rect 477040 356858 477092 356864
rect 477040 356800 477092 356806
rect 480168 356858 480220 356864
rect 480168 356800 480220 356806
rect 477052 354676 477080 356800
rect 471716 354648 471928 354676
rect 477052 354648 477172 354676
rect 471900 345016 471928 354648
rect 477144 354552 477172 354648
rect 480180 354620 480208 356800
rect 483204 356489 483256 356495
rect 483204 356431 483256 356437
rect 486240 356489 486292 356495
rect 486240 356431 486292 356437
rect 483216 354688 483244 356431
rect 483204 354682 483256 354688
rect 483204 354624 483256 354630
rect 480168 354614 480220 354620
rect 480168 354556 480220 354562
rect 477132 354546 477184 354552
rect 477132 354488 477184 354494
rect 486252 353668 486280 356431
rect 486240 353662 486292 353668
rect 486240 353604 486292 353610
rect 484582 351930 484638 351939
rect 484582 351865 484638 351874
rect 471716 344988 471928 345016
rect 470262 342488 470826 342494
rect 470314 342482 470326 342488
rect 470378 342482 470390 342488
rect 470442 342482 470454 342488
rect 470506 342482 470518 342488
rect 470570 342482 470582 342488
rect 470634 342482 470646 342488
rect 470698 342482 470710 342488
rect 470762 342482 470774 342488
rect 470506 342436 470516 342482
rect 470572 342436 470582 342482
rect 470262 342426 470276 342436
rect 470332 342426 470356 342436
rect 470412 342426 470436 342436
rect 470492 342426 470516 342436
rect 470572 342426 470596 342436
rect 470652 342426 470676 342436
rect 470732 342426 470756 342436
rect 470812 342426 470826 342436
rect 470262 342424 470826 342426
rect 470314 342402 470326 342424
rect 470378 342402 470390 342424
rect 470442 342402 470454 342424
rect 470506 342402 470518 342424
rect 470570 342402 470582 342424
rect 470634 342402 470646 342424
rect 470698 342402 470710 342424
rect 470762 342402 470774 342424
rect 470506 342372 470516 342402
rect 470572 342372 470582 342402
rect 470262 342360 470276 342372
rect 470332 342360 470356 342372
rect 470412 342360 470436 342372
rect 470492 342360 470516 342372
rect 470572 342360 470596 342372
rect 470652 342360 470676 342372
rect 470732 342360 470756 342372
rect 470812 342360 470826 342372
rect 470506 342346 470516 342360
rect 470572 342346 470582 342360
rect 470314 342322 470326 342346
rect 470378 342322 470390 342346
rect 470442 342322 470454 342346
rect 470506 342322 470518 342346
rect 470570 342322 470582 342346
rect 470634 342322 470646 342346
rect 470698 342322 470710 342346
rect 470762 342322 470774 342346
rect 470506 342308 470516 342322
rect 470572 342308 470582 342322
rect 470262 342296 470276 342308
rect 470332 342296 470356 342308
rect 470412 342296 470436 342308
rect 470492 342296 470516 342308
rect 470572 342296 470596 342308
rect 470652 342296 470676 342308
rect 470732 342296 470756 342308
rect 470812 342296 470826 342308
rect 470506 342266 470516 342296
rect 470572 342266 470582 342296
rect 470314 342244 470326 342266
rect 470378 342244 470390 342266
rect 470442 342244 470454 342266
rect 470506 342244 470518 342266
rect 470570 342244 470582 342266
rect 470634 342244 470646 342266
rect 470698 342244 470710 342266
rect 470762 342244 470774 342266
rect 470262 342242 470826 342244
rect 470262 342232 470276 342242
rect 470332 342232 470356 342242
rect 470412 342232 470436 342242
rect 470492 342232 470516 342242
rect 470572 342232 470596 342242
rect 470652 342232 470676 342242
rect 470732 342232 470756 342242
rect 470812 342232 470826 342242
rect 470506 342186 470516 342232
rect 470572 342186 470582 342232
rect 470314 342180 470326 342186
rect 470378 342180 470390 342186
rect 470442 342180 470454 342186
rect 470506 342180 470518 342186
rect 470570 342180 470582 342186
rect 470634 342180 470646 342186
rect 470698 342180 470710 342186
rect 470762 342180 470774 342186
rect 470262 342174 470826 342180
rect 471716 341836 471744 344988
rect 484596 342283 484624 351865
rect 484582 342274 484638 342283
rect 484582 342209 484638 342218
rect 471704 341830 471756 341836
rect 471704 341772 471756 341778
rect 471244 341762 471296 341768
rect 471244 341704 471296 341710
rect 484398 341730 484454 341739
rect 469022 341401 469586 341407
rect 469074 341395 469086 341401
rect 469138 341395 469150 341401
rect 469202 341395 469214 341401
rect 469266 341395 469278 341401
rect 469330 341395 469342 341401
rect 469394 341395 469406 341401
rect 469458 341395 469470 341401
rect 469522 341395 469534 341401
rect 469266 341349 469276 341395
rect 469332 341349 469342 341395
rect 469022 341339 469036 341349
rect 469092 341339 469116 341349
rect 469172 341339 469196 341349
rect 469252 341339 469276 341349
rect 469332 341339 469356 341349
rect 469412 341339 469436 341349
rect 469492 341339 469516 341349
rect 469572 341339 469586 341349
rect 469022 341337 469586 341339
rect 469074 341315 469086 341337
rect 469138 341315 469150 341337
rect 469202 341315 469214 341337
rect 469266 341315 469278 341337
rect 469330 341315 469342 341337
rect 469394 341315 469406 341337
rect 469458 341315 469470 341337
rect 469522 341315 469534 341337
rect 469266 341285 469276 341315
rect 469332 341285 469342 341315
rect 469022 341273 469036 341285
rect 469092 341273 469116 341285
rect 469172 341273 469196 341285
rect 469252 341273 469276 341285
rect 469332 341273 469356 341285
rect 469412 341273 469436 341285
rect 469492 341273 469516 341285
rect 469572 341273 469586 341285
rect 469266 341259 469276 341273
rect 469332 341259 469342 341273
rect 469074 341235 469086 341259
rect 469138 341235 469150 341259
rect 469202 341235 469214 341259
rect 469266 341235 469278 341259
rect 469330 341235 469342 341259
rect 469394 341235 469406 341259
rect 469458 341235 469470 341259
rect 469522 341235 469534 341259
rect 469266 341221 469276 341235
rect 469332 341221 469342 341235
rect 469022 341209 469036 341221
rect 469092 341209 469116 341221
rect 469172 341209 469196 341221
rect 469252 341209 469276 341221
rect 469332 341209 469356 341221
rect 469412 341209 469436 341221
rect 469492 341209 469516 341221
rect 469572 341209 469586 341221
rect 469266 341179 469276 341209
rect 469332 341179 469342 341209
rect 469074 341157 469086 341179
rect 469138 341157 469150 341179
rect 469202 341157 469214 341179
rect 469266 341157 469278 341179
rect 469330 341157 469342 341179
rect 469394 341157 469406 341179
rect 469458 341157 469470 341179
rect 469522 341157 469534 341179
rect 469022 341155 469586 341157
rect 469022 341145 469036 341155
rect 469092 341145 469116 341155
rect 469172 341145 469196 341155
rect 469252 341145 469276 341155
rect 469332 341145 469356 341155
rect 469412 341145 469436 341155
rect 469492 341145 469516 341155
rect 469572 341145 469586 341155
rect 469266 341099 469276 341145
rect 469332 341099 469342 341145
rect 469074 341093 469086 341099
rect 469138 341093 469150 341099
rect 469202 341093 469214 341099
rect 469266 341093 469278 341099
rect 469330 341093 469342 341099
rect 469394 341093 469406 341099
rect 469458 341093 469470 341099
rect 469522 341093 469534 341099
rect 469022 341087 469586 341093
rect 470262 340316 470826 340322
rect 470314 340310 470326 340316
rect 470378 340310 470390 340316
rect 470442 340310 470454 340316
rect 470506 340310 470518 340316
rect 470570 340310 470582 340316
rect 470634 340310 470646 340316
rect 470698 340310 470710 340316
rect 470762 340310 470774 340316
rect 470506 340264 470516 340310
rect 470572 340264 470582 340310
rect 470262 340254 470276 340264
rect 470332 340254 470356 340264
rect 470412 340254 470436 340264
rect 470492 340254 470516 340264
rect 470572 340254 470596 340264
rect 470652 340254 470676 340264
rect 470732 340254 470756 340264
rect 470812 340254 470826 340264
rect 470262 340252 470826 340254
rect 470314 340230 470326 340252
rect 470378 340230 470390 340252
rect 470442 340230 470454 340252
rect 470506 340230 470518 340252
rect 470570 340230 470582 340252
rect 470634 340230 470646 340252
rect 470698 340230 470710 340252
rect 470762 340230 470774 340252
rect 470506 340200 470516 340230
rect 470572 340200 470582 340230
rect 470262 340188 470276 340200
rect 470332 340188 470356 340200
rect 470412 340188 470436 340200
rect 470492 340188 470516 340200
rect 470572 340188 470596 340200
rect 470652 340188 470676 340200
rect 470732 340188 470756 340200
rect 470812 340188 470826 340200
rect 470506 340174 470516 340188
rect 470572 340174 470582 340188
rect 470314 340150 470326 340174
rect 470378 340150 470390 340174
rect 470442 340150 470454 340174
rect 470506 340150 470518 340174
rect 470570 340150 470582 340174
rect 470634 340150 470646 340174
rect 470698 340150 470710 340174
rect 470762 340150 470774 340174
rect 470506 340136 470516 340150
rect 470572 340136 470582 340150
rect 470262 340124 470276 340136
rect 470332 340124 470356 340136
rect 470412 340124 470436 340136
rect 470492 340124 470516 340136
rect 470572 340124 470596 340136
rect 470652 340124 470676 340136
rect 470732 340124 470756 340136
rect 470812 340124 470826 340136
rect 470506 340094 470516 340124
rect 470572 340094 470582 340124
rect 470314 340072 470326 340094
rect 470378 340072 470390 340094
rect 470442 340072 470454 340094
rect 470506 340072 470518 340094
rect 470570 340072 470582 340094
rect 470634 340072 470646 340094
rect 470698 340072 470710 340094
rect 470762 340072 470774 340094
rect 470262 340070 470826 340072
rect 470262 340060 470276 340070
rect 470332 340060 470356 340070
rect 470412 340060 470436 340070
rect 470492 340060 470516 340070
rect 470572 340060 470596 340070
rect 470652 340060 470676 340070
rect 470732 340060 470756 340070
rect 470812 340060 470826 340070
rect 470506 340014 470516 340060
rect 470572 340014 470582 340060
rect 470314 340008 470326 340014
rect 470378 340008 470390 340014
rect 470442 340008 470454 340014
rect 470506 340008 470518 340014
rect 470570 340008 470582 340014
rect 470634 340008 470646 340014
rect 470698 340008 470710 340014
rect 470762 340008 470774 340014
rect 470262 340002 470826 340008
rect 470262 322488 470826 322494
rect 470314 322482 470326 322488
rect 470378 322482 470390 322488
rect 470442 322482 470454 322488
rect 470506 322482 470518 322488
rect 470570 322482 470582 322488
rect 470634 322482 470646 322488
rect 470698 322482 470710 322488
rect 470762 322482 470774 322488
rect 470506 322436 470516 322482
rect 470572 322436 470582 322482
rect 470262 322426 470276 322436
rect 470332 322426 470356 322436
rect 470412 322426 470436 322436
rect 470492 322426 470516 322436
rect 470572 322426 470596 322436
rect 470652 322426 470676 322436
rect 470732 322426 470756 322436
rect 470812 322426 470826 322436
rect 470262 322424 470826 322426
rect 470314 322402 470326 322424
rect 470378 322402 470390 322424
rect 470442 322402 470454 322424
rect 470506 322402 470518 322424
rect 470570 322402 470582 322424
rect 470634 322402 470646 322424
rect 470698 322402 470710 322424
rect 470762 322402 470774 322424
rect 470506 322372 470516 322402
rect 470572 322372 470582 322402
rect 470262 322360 470276 322372
rect 470332 322360 470356 322372
rect 470412 322360 470436 322372
rect 470492 322360 470516 322372
rect 470572 322360 470596 322372
rect 470652 322360 470676 322372
rect 470732 322360 470756 322372
rect 470812 322360 470826 322372
rect 470506 322346 470516 322360
rect 470572 322346 470582 322360
rect 470314 322322 470326 322346
rect 470378 322322 470390 322346
rect 470442 322322 470454 322346
rect 470506 322322 470518 322346
rect 470570 322322 470582 322346
rect 470634 322322 470646 322346
rect 470698 322322 470710 322346
rect 470762 322322 470774 322346
rect 470506 322308 470516 322322
rect 470572 322308 470582 322322
rect 470262 322296 470276 322308
rect 470332 322296 470356 322308
rect 470412 322296 470436 322308
rect 470492 322296 470516 322308
rect 470572 322296 470596 322308
rect 470652 322296 470676 322308
rect 470732 322296 470756 322308
rect 470812 322296 470826 322308
rect 470506 322266 470516 322296
rect 470572 322266 470582 322296
rect 470314 322244 470326 322266
rect 470378 322244 470390 322266
rect 470442 322244 470454 322266
rect 470506 322244 470518 322266
rect 470570 322244 470582 322266
rect 470634 322244 470646 322266
rect 470698 322244 470710 322266
rect 470762 322244 470774 322266
rect 470262 322242 470826 322244
rect 470262 322232 470276 322242
rect 470332 322232 470356 322242
rect 470412 322232 470436 322242
rect 470492 322232 470516 322242
rect 470572 322232 470596 322242
rect 470652 322232 470676 322242
rect 470732 322232 470756 322242
rect 470812 322232 470826 322242
rect 470506 322186 470516 322232
rect 470572 322186 470582 322232
rect 470314 322180 470326 322186
rect 470378 322180 470390 322186
rect 470442 322180 470454 322186
rect 470506 322180 470518 322186
rect 470570 322180 470582 322186
rect 470634 322180 470646 322186
rect 470698 322180 470710 322186
rect 470762 322180 470774 322186
rect 470262 322174 470826 322180
rect 471256 321640 471284 341704
rect 484398 341665 484454 341674
rect 477906 340994 477915 341050
rect 477971 340994 477980 341050
rect 481223 340994 481232 341050
rect 481288 340994 481297 341050
rect 484412 340952 484440 341665
rect 487885 340994 487894 341050
rect 487950 340994 487959 341050
rect 484400 340946 484452 340952
rect 484400 340888 484452 340894
rect 482100 340878 482152 340884
rect 474648 340857 474700 340863
rect 482100 340820 482152 340826
rect 474648 340799 474700 340805
rect 474554 340506 474610 340515
rect 474660 340492 474688 340799
rect 474610 340464 474688 340492
rect 474554 340441 474610 340450
rect 475476 340402 475528 340408
rect 475476 340344 475528 340350
rect 478788 340402 478840 340408
rect 478788 340344 478840 340350
rect 475488 339456 475516 340344
rect 478800 339456 478828 340344
rect 475476 339450 475528 339456
rect 475476 339392 475528 339398
rect 478788 339450 478840 339456
rect 478788 339392 478840 339398
rect 482112 339388 482140 340820
rect 484400 340538 484452 340544
rect 484400 340480 484452 340486
rect 485596 340492 485648 340498
rect 484412 339404 484440 340480
rect 485596 340434 485648 340440
rect 482100 339382 482152 339388
rect 482100 339324 482152 339330
rect 484320 339376 484440 339404
rect 484320 322155 484348 339376
rect 485608 335356 485636 340434
rect 485608 335328 485728 335356
rect 485700 331228 485728 335328
rect 485688 331222 485740 331228
rect 485688 331164 485740 331170
rect 484306 322146 484362 322155
rect 484306 322081 484362 322090
rect 483138 321696 483520 321724
rect 471244 321634 471296 321640
rect 483492 321611 483520 321696
rect 471244 321576 471296 321582
rect 483478 321602 483534 321611
rect 469022 321401 469586 321407
rect 469074 321395 469086 321401
rect 469138 321395 469150 321401
rect 469202 321395 469214 321401
rect 469266 321395 469278 321401
rect 469330 321395 469342 321401
rect 469394 321395 469406 321401
rect 469458 321395 469470 321401
rect 469522 321395 469534 321401
rect 469266 321349 469276 321395
rect 469332 321349 469342 321395
rect 469022 321339 469036 321349
rect 469092 321339 469116 321349
rect 469172 321339 469196 321349
rect 469252 321339 469276 321349
rect 469332 321339 469356 321349
rect 469412 321339 469436 321349
rect 469492 321339 469516 321349
rect 469572 321339 469586 321349
rect 469022 321337 469586 321339
rect 469074 321315 469086 321337
rect 469138 321315 469150 321337
rect 469202 321315 469214 321337
rect 469266 321315 469278 321337
rect 469330 321315 469342 321337
rect 469394 321315 469406 321337
rect 469458 321315 469470 321337
rect 469522 321315 469534 321337
rect 469266 321285 469276 321315
rect 469332 321285 469342 321315
rect 469022 321273 469036 321285
rect 469092 321273 469116 321285
rect 469172 321273 469196 321285
rect 469252 321273 469276 321285
rect 469332 321273 469356 321285
rect 469412 321273 469436 321285
rect 469492 321273 469516 321285
rect 469572 321273 469586 321285
rect 469266 321259 469276 321273
rect 469332 321259 469342 321273
rect 469074 321235 469086 321259
rect 469138 321235 469150 321259
rect 469202 321235 469214 321259
rect 469266 321235 469278 321259
rect 469330 321235 469342 321259
rect 469394 321235 469406 321259
rect 469458 321235 469470 321259
rect 469522 321235 469534 321259
rect 469266 321221 469276 321235
rect 469332 321221 469342 321235
rect 469022 321209 469036 321221
rect 469092 321209 469116 321221
rect 469172 321209 469196 321221
rect 469252 321209 469276 321221
rect 469332 321209 469356 321221
rect 469412 321209 469436 321221
rect 469492 321209 469516 321221
rect 469572 321209 469586 321221
rect 469266 321179 469276 321209
rect 469332 321179 469342 321209
rect 469074 321157 469086 321179
rect 469138 321157 469150 321179
rect 469202 321157 469214 321179
rect 469266 321157 469278 321179
rect 469330 321157 469342 321179
rect 469394 321157 469406 321179
rect 469458 321157 469470 321179
rect 469522 321157 469534 321179
rect 469022 321155 469586 321157
rect 469022 321145 469036 321155
rect 469092 321145 469116 321155
rect 469172 321145 469196 321155
rect 469252 321145 469276 321155
rect 469332 321145 469356 321155
rect 469412 321145 469436 321155
rect 469492 321145 469516 321155
rect 469572 321145 469586 321155
rect 469266 321099 469276 321145
rect 469332 321099 469342 321145
rect 469074 321093 469086 321099
rect 469138 321093 469150 321099
rect 469202 321093 469214 321099
rect 469266 321093 469278 321099
rect 469330 321093 469342 321099
rect 469394 321093 469406 321099
rect 469458 321093 469470 321099
rect 469522 321093 469534 321099
rect 469022 321087 469586 321093
rect 470262 320316 470826 320322
rect 470314 320310 470326 320316
rect 470378 320310 470390 320316
rect 470442 320310 470454 320316
rect 470506 320310 470518 320316
rect 470570 320310 470582 320316
rect 470634 320310 470646 320316
rect 470698 320310 470710 320316
rect 470762 320310 470774 320316
rect 470506 320264 470516 320310
rect 470572 320264 470582 320310
rect 470262 320254 470276 320264
rect 470332 320254 470356 320264
rect 470412 320254 470436 320264
rect 470492 320254 470516 320264
rect 470572 320254 470596 320264
rect 470652 320254 470676 320264
rect 470732 320254 470756 320264
rect 470812 320254 470826 320264
rect 470262 320252 470826 320254
rect 470314 320230 470326 320252
rect 470378 320230 470390 320252
rect 470442 320230 470454 320252
rect 470506 320230 470518 320252
rect 470570 320230 470582 320252
rect 470634 320230 470646 320252
rect 470698 320230 470710 320252
rect 470762 320230 470774 320252
rect 470506 320200 470516 320230
rect 470572 320200 470582 320230
rect 470262 320188 470276 320200
rect 470332 320188 470356 320200
rect 470412 320188 470436 320200
rect 470492 320188 470516 320200
rect 470572 320188 470596 320200
rect 470652 320188 470676 320200
rect 470732 320188 470756 320200
rect 470812 320188 470826 320200
rect 470506 320174 470516 320188
rect 470572 320174 470582 320188
rect 470314 320150 470326 320174
rect 470378 320150 470390 320174
rect 470442 320150 470454 320174
rect 470506 320150 470518 320174
rect 470570 320150 470582 320174
rect 470634 320150 470646 320174
rect 470698 320150 470710 320174
rect 470762 320150 470774 320174
rect 470506 320136 470516 320150
rect 470572 320136 470582 320150
rect 470262 320124 470276 320136
rect 470332 320124 470356 320136
rect 470412 320124 470436 320136
rect 470492 320124 470516 320136
rect 470572 320124 470596 320136
rect 470652 320124 470676 320136
rect 470732 320124 470756 320136
rect 470812 320124 470826 320136
rect 470506 320094 470516 320124
rect 470572 320094 470582 320124
rect 470314 320072 470326 320094
rect 470378 320072 470390 320094
rect 470442 320072 470454 320094
rect 470506 320072 470518 320094
rect 470570 320072 470582 320094
rect 470634 320072 470646 320094
rect 470698 320072 470710 320094
rect 470762 320072 470774 320094
rect 470262 320070 470826 320072
rect 470262 320060 470276 320070
rect 470332 320060 470356 320070
rect 470412 320060 470436 320070
rect 470492 320060 470516 320070
rect 470572 320060 470596 320070
rect 470652 320060 470676 320070
rect 470732 320060 470756 320070
rect 470812 320060 470826 320070
rect 470506 320014 470516 320060
rect 470572 320014 470582 320060
rect 470314 320008 470326 320014
rect 470378 320008 470390 320014
rect 470442 320008 470454 320014
rect 470506 320008 470518 320014
rect 470570 320008 470582 320014
rect 470634 320008 470646 320014
rect 470698 320008 470710 320014
rect 470762 320008 470774 320014
rect 470262 320002 470826 320008
rect 470262 307088 470826 307094
rect 470314 307082 470326 307088
rect 470378 307082 470390 307088
rect 470442 307082 470454 307088
rect 470506 307082 470518 307088
rect 470570 307082 470582 307088
rect 470634 307082 470646 307088
rect 470698 307082 470710 307088
rect 470762 307082 470774 307088
rect 470506 307036 470516 307082
rect 470572 307036 470582 307082
rect 470262 307026 470276 307036
rect 470332 307026 470356 307036
rect 470412 307026 470436 307036
rect 470492 307026 470516 307036
rect 470572 307026 470596 307036
rect 470652 307026 470676 307036
rect 470732 307026 470756 307036
rect 470812 307026 470826 307036
rect 470262 307024 470826 307026
rect 470314 307002 470326 307024
rect 470378 307002 470390 307024
rect 470442 307002 470454 307024
rect 470506 307002 470518 307024
rect 470570 307002 470582 307024
rect 470634 307002 470646 307024
rect 470698 307002 470710 307024
rect 470762 307002 470774 307024
rect 470506 306972 470516 307002
rect 470572 306972 470582 307002
rect 470262 306960 470276 306972
rect 470332 306960 470356 306972
rect 470412 306960 470436 306972
rect 470492 306960 470516 306972
rect 470572 306960 470596 306972
rect 470652 306960 470676 306972
rect 470732 306960 470756 306972
rect 470812 306960 470826 306972
rect 470506 306946 470516 306960
rect 470572 306946 470582 306960
rect 470314 306922 470326 306946
rect 470378 306922 470390 306946
rect 470442 306922 470454 306946
rect 470506 306922 470518 306946
rect 470570 306922 470582 306946
rect 470634 306922 470646 306946
rect 470698 306922 470710 306946
rect 470762 306922 470774 306946
rect 470506 306908 470516 306922
rect 470572 306908 470582 306922
rect 470262 306896 470276 306908
rect 470332 306896 470356 306908
rect 470412 306896 470436 306908
rect 470492 306896 470516 306908
rect 470572 306896 470596 306908
rect 470652 306896 470676 306908
rect 470732 306896 470756 306908
rect 470812 306896 470826 306908
rect 470506 306866 470516 306896
rect 470572 306866 470582 306896
rect 470314 306844 470326 306866
rect 470378 306844 470390 306866
rect 470442 306844 470454 306866
rect 470506 306844 470518 306866
rect 470570 306844 470582 306866
rect 470634 306844 470646 306866
rect 470698 306844 470710 306866
rect 470762 306844 470774 306866
rect 470262 306842 470826 306844
rect 470262 306832 470276 306842
rect 470332 306832 470356 306842
rect 470412 306832 470436 306842
rect 470492 306832 470516 306842
rect 470572 306832 470596 306842
rect 470652 306832 470676 306842
rect 470732 306832 470756 306842
rect 470812 306832 470826 306842
rect 470506 306786 470516 306832
rect 470572 306786 470582 306832
rect 470314 306780 470326 306786
rect 470378 306780 470390 306786
rect 470442 306780 470454 306786
rect 470506 306780 470518 306786
rect 470570 306780 470582 306786
rect 470634 306780 470646 306786
rect 470698 306780 470710 306786
rect 470762 306780 470774 306786
rect 470262 306774 470826 306780
rect 471256 306340 471284 321576
rect 483478 321537 483534 321546
rect 474278 321330 474334 321339
rect 474334 321288 474680 321316
rect 474278 321265 474334 321274
rect 481178 321058 481234 321067
rect 478125 321016 478184 321044
rect 478156 320931 478184 321016
rect 488170 321058 488226 321067
rect 481234 321016 481568 321044
rect 481178 320993 481234 321002
rect 488226 321016 488456 321044
rect 488170 320993 488226 321002
rect 478142 320922 478198 320931
rect 478142 320857 478198 320866
rect 475476 320489 475528 320495
rect 475476 320431 475528 320437
rect 482376 320478 482428 320484
rect 475488 318784 475516 320431
rect 482376 320420 482428 320426
rect 479064 320410 479116 320416
rect 479064 320352 479116 320358
rect 479076 318784 479104 320352
rect 475476 318778 475528 318784
rect 475476 318720 475528 318726
rect 479064 318778 479116 318784
rect 479064 318720 479116 318726
rect 482388 318716 482416 320420
rect 485964 320410 486016 320416
rect 485964 320352 486016 320358
rect 482376 318710 482428 318716
rect 482376 318652 482428 318658
rect 485976 318648 486004 320352
rect 485964 318642 486016 318648
rect 485964 318584 486016 318590
rect 480902 306506 480958 306515
rect 480902 306441 480958 306450
rect 471244 306334 471296 306340
rect 471244 306276 471296 306282
rect 473728 306286 473780 306292
rect 469022 306003 469586 306009
rect 469074 305997 469086 306003
rect 469138 305997 469150 306003
rect 469202 305997 469214 306003
rect 469266 305997 469278 306003
rect 469330 305997 469342 306003
rect 469394 305997 469406 306003
rect 469458 305997 469470 306003
rect 469522 305997 469534 306003
rect 469266 305951 469276 305997
rect 469332 305951 469342 305997
rect 469022 305941 469036 305951
rect 469092 305941 469116 305951
rect 469172 305941 469196 305951
rect 469252 305941 469276 305951
rect 469332 305941 469356 305951
rect 469412 305941 469436 305951
rect 469492 305941 469516 305951
rect 469572 305941 469586 305951
rect 469022 305939 469586 305941
rect 469074 305917 469086 305939
rect 469138 305917 469150 305939
rect 469202 305917 469214 305939
rect 469266 305917 469278 305939
rect 469330 305917 469342 305939
rect 469394 305917 469406 305939
rect 469458 305917 469470 305939
rect 469522 305917 469534 305939
rect 469266 305887 469276 305917
rect 469332 305887 469342 305917
rect 469022 305875 469036 305887
rect 469092 305875 469116 305887
rect 469172 305875 469196 305887
rect 469252 305875 469276 305887
rect 469332 305875 469356 305887
rect 469412 305875 469436 305887
rect 469492 305875 469516 305887
rect 469572 305875 469586 305887
rect 469266 305861 469276 305875
rect 469332 305861 469342 305875
rect 469074 305837 469086 305861
rect 469138 305837 469150 305861
rect 469202 305837 469214 305861
rect 469266 305837 469278 305861
rect 469330 305837 469342 305861
rect 469394 305837 469406 305861
rect 469458 305837 469470 305861
rect 469522 305837 469534 305861
rect 469266 305823 469276 305837
rect 469332 305823 469342 305837
rect 469022 305811 469036 305823
rect 469092 305811 469116 305823
rect 469172 305811 469196 305823
rect 469252 305811 469276 305823
rect 469332 305811 469356 305823
rect 469412 305811 469436 305823
rect 469492 305811 469516 305823
rect 469572 305811 469586 305823
rect 469266 305781 469276 305811
rect 469332 305781 469342 305811
rect 469074 305759 469086 305781
rect 469138 305759 469150 305781
rect 469202 305759 469214 305781
rect 469266 305759 469278 305781
rect 469330 305759 469342 305781
rect 469394 305759 469406 305781
rect 469458 305759 469470 305781
rect 469522 305759 469534 305781
rect 469022 305757 469586 305759
rect 469022 305747 469036 305757
rect 469092 305747 469116 305757
rect 469172 305747 469196 305757
rect 469252 305747 469276 305757
rect 469332 305747 469356 305757
rect 469412 305747 469436 305757
rect 469492 305747 469516 305757
rect 469572 305747 469586 305757
rect 469266 305701 469276 305747
rect 469332 305701 469342 305747
rect 469074 305695 469086 305701
rect 469138 305695 469150 305701
rect 469202 305695 469214 305701
rect 469266 305695 469278 305701
rect 469330 305695 469342 305701
rect 469394 305695 469406 305701
rect 469458 305695 469470 305701
rect 469522 305695 469534 305701
rect 469022 305689 469586 305695
rect 470262 304916 470826 304922
rect 470314 304910 470326 304916
rect 470378 304910 470390 304916
rect 470442 304910 470454 304916
rect 470506 304910 470518 304916
rect 470570 304910 470582 304916
rect 470634 304910 470646 304916
rect 470698 304910 470710 304916
rect 470762 304910 470774 304916
rect 470506 304864 470516 304910
rect 470572 304864 470582 304910
rect 470262 304854 470276 304864
rect 470332 304854 470356 304864
rect 470412 304854 470436 304864
rect 470492 304854 470516 304864
rect 470572 304854 470596 304864
rect 470652 304854 470676 304864
rect 470732 304854 470756 304864
rect 470812 304854 470826 304864
rect 470262 304852 470826 304854
rect 470314 304830 470326 304852
rect 470378 304830 470390 304852
rect 470442 304830 470454 304852
rect 470506 304830 470518 304852
rect 470570 304830 470582 304852
rect 470634 304830 470646 304852
rect 470698 304830 470710 304852
rect 470762 304830 470774 304852
rect 470506 304800 470516 304830
rect 470572 304800 470582 304830
rect 470262 304788 470276 304800
rect 470332 304788 470356 304800
rect 470412 304788 470436 304800
rect 470492 304788 470516 304800
rect 470572 304788 470596 304800
rect 470652 304788 470676 304800
rect 470732 304788 470756 304800
rect 470812 304788 470826 304800
rect 470506 304774 470516 304788
rect 470572 304774 470582 304788
rect 470314 304750 470326 304774
rect 470378 304750 470390 304774
rect 470442 304750 470454 304774
rect 470506 304750 470518 304774
rect 470570 304750 470582 304774
rect 470634 304750 470646 304774
rect 470698 304750 470710 304774
rect 470762 304750 470774 304774
rect 470506 304736 470516 304750
rect 470572 304736 470582 304750
rect 470262 304724 470276 304736
rect 470332 304724 470356 304736
rect 470412 304724 470436 304736
rect 470492 304724 470516 304736
rect 470572 304724 470596 304736
rect 470652 304724 470676 304736
rect 470732 304724 470756 304736
rect 470812 304724 470826 304736
rect 470506 304694 470516 304724
rect 470572 304694 470582 304724
rect 470314 304672 470326 304694
rect 470378 304672 470390 304694
rect 470442 304672 470454 304694
rect 470506 304672 470518 304694
rect 470570 304672 470582 304694
rect 470634 304672 470646 304694
rect 470698 304672 470710 304694
rect 470762 304672 470774 304694
rect 470262 304670 470826 304672
rect 470262 304660 470276 304670
rect 470332 304660 470356 304670
rect 470412 304660 470436 304670
rect 470492 304660 470516 304670
rect 470572 304660 470596 304670
rect 470652 304660 470676 304670
rect 470732 304660 470756 304670
rect 470812 304660 470826 304670
rect 470506 304614 470516 304660
rect 470572 304614 470582 304660
rect 470314 304608 470326 304614
rect 470378 304608 470390 304614
rect 470442 304608 470454 304614
rect 470506 304608 470518 304614
rect 470570 304608 470582 304614
rect 470634 304608 470646 304614
rect 470698 304608 470710 304614
rect 470762 304608 470774 304614
rect 470262 304602 470826 304608
rect 470262 287489 470826 287495
rect 470314 287483 470326 287489
rect 470378 287483 470390 287489
rect 470442 287483 470454 287489
rect 470506 287483 470518 287489
rect 470570 287483 470582 287489
rect 470634 287483 470646 287489
rect 470698 287483 470710 287489
rect 470762 287483 470774 287489
rect 470506 287437 470516 287483
rect 470572 287437 470582 287483
rect 470262 287427 470276 287437
rect 470332 287427 470356 287437
rect 470412 287427 470436 287437
rect 470492 287427 470516 287437
rect 470572 287427 470596 287437
rect 470652 287427 470676 287437
rect 470732 287427 470756 287437
rect 470812 287427 470826 287437
rect 470262 287425 470826 287427
rect 470314 287403 470326 287425
rect 470378 287403 470390 287425
rect 470442 287403 470454 287425
rect 470506 287403 470518 287425
rect 470570 287403 470582 287425
rect 470634 287403 470646 287425
rect 470698 287403 470710 287425
rect 470762 287403 470774 287425
rect 470506 287373 470516 287403
rect 470572 287373 470582 287403
rect 470262 287361 470276 287373
rect 470332 287361 470356 287373
rect 470412 287361 470436 287373
rect 470492 287361 470516 287373
rect 470572 287361 470596 287373
rect 470652 287361 470676 287373
rect 470732 287361 470756 287373
rect 470812 287361 470826 287373
rect 470506 287347 470516 287361
rect 470572 287347 470582 287361
rect 470314 287323 470326 287347
rect 470378 287323 470390 287347
rect 470442 287323 470454 287347
rect 470506 287323 470518 287347
rect 470570 287323 470582 287347
rect 470634 287323 470646 287347
rect 470698 287323 470710 287347
rect 470762 287323 470774 287347
rect 470506 287309 470516 287323
rect 470572 287309 470582 287323
rect 470262 287297 470276 287309
rect 470332 287297 470356 287309
rect 470412 287297 470436 287309
rect 470492 287297 470516 287309
rect 470572 287297 470596 287309
rect 470652 287297 470676 287309
rect 470732 287297 470756 287309
rect 470812 287297 470826 287309
rect 470506 287267 470516 287297
rect 470572 287267 470582 287297
rect 470314 287245 470326 287267
rect 470378 287245 470390 287267
rect 470442 287245 470454 287267
rect 470506 287245 470518 287267
rect 470570 287245 470582 287267
rect 470634 287245 470646 287267
rect 470698 287245 470710 287267
rect 470762 287245 470774 287267
rect 470262 287243 470826 287245
rect 470262 287233 470276 287243
rect 470332 287233 470356 287243
rect 470412 287233 470436 287243
rect 470492 287233 470516 287243
rect 470572 287233 470596 287243
rect 470652 287233 470676 287243
rect 470732 287233 470756 287243
rect 470812 287233 470826 287243
rect 470506 287187 470516 287233
rect 470572 287187 470582 287233
rect 470314 287181 470326 287187
rect 470378 287181 470390 287187
rect 470442 287181 470454 287187
rect 470506 287181 470518 287187
rect 470570 287181 470582 287187
rect 470634 287181 470646 287187
rect 470698 287181 470710 287187
rect 470762 287181 470774 287187
rect 470262 287175 470826 287181
rect 471256 286688 471284 306276
rect 473728 306228 473780 306234
rect 473740 305971 473768 306228
rect 480916 306084 480944 306441
rect 487525 306178 487534 306234
rect 487590 306178 487599 306234
rect 480916 306056 481032 306084
rect 473726 305962 473782 305971
rect 473726 305897 473782 305906
rect 477739 305690 477795 305699
rect 477739 305625 477795 305634
rect 484122 305554 484178 305563
rect 484178 305512 484297 305540
rect 484122 305489 484178 305498
rect 478604 305450 478656 305456
rect 478604 305392 478656 305398
rect 485136 305450 485188 305456
rect 485136 305392 485188 305398
rect 475292 305090 475344 305096
rect 475292 305032 475344 305038
rect 475304 303620 475332 305032
rect 478616 303620 478644 305392
rect 481824 305090 481876 305096
rect 481824 305032 481876 305038
rect 481836 303620 481864 305032
rect 485148 303620 485176 305392
rect 490564 305042 490616 305048
rect 490564 304984 490616 304990
rect 475292 303614 475344 303620
rect 475292 303556 475344 303562
rect 478604 303614 478656 303620
rect 478604 303556 478656 303562
rect 481824 303614 481876 303620
rect 481824 303556 481876 303562
rect 485136 303614 485188 303620
rect 485136 303556 485188 303562
rect 482282 302290 482338 302299
rect 482282 302225 482338 302234
rect 482296 288427 482324 302225
rect 490576 292536 490604 304984
rect 490760 298112 490788 409976
rect 491956 300832 491984 449348
rect 515404 445938 515456 445944
rect 515404 445880 515456 445886
rect 493324 441654 493376 441660
rect 493324 441596 493376 441602
rect 492036 431046 492088 431052
rect 492036 430988 492088 430994
rect 491944 300826 491996 300832
rect 491944 300768 491996 300774
rect 492048 299472 492076 430988
rect 493336 408476 493364 441596
rect 494704 440294 494756 440300
rect 494704 440236 494756 440242
rect 493324 408470 493376 408476
rect 493324 408412 493376 408418
rect 493324 389498 493376 389504
rect 493324 389440 493376 389446
rect 492128 356450 492180 356456
rect 492128 356392 492180 356398
rect 492036 299466 492088 299472
rect 492036 299408 492088 299414
rect 490748 298106 490800 298112
rect 490748 298048 490800 298054
rect 492140 296684 492168 356392
rect 492220 340402 492272 340408
rect 492220 340344 492272 340350
rect 492128 296678 492180 296684
rect 492128 296620 492180 296626
rect 492232 295324 492260 340344
rect 492312 320410 492364 320416
rect 492312 320352 492364 320358
rect 492220 295318 492272 295324
rect 492220 295260 492272 295266
rect 492324 293964 492352 320352
rect 493336 296616 493364 389440
rect 494716 387736 494744 440236
rect 496084 438934 496136 438940
rect 496084 438876 496136 438882
rect 494704 387730 494756 387736
rect 494704 387672 494756 387678
rect 496096 354552 496124 438876
rect 497464 437506 497516 437512
rect 497464 437448 497516 437454
rect 496084 354546 496136 354552
rect 496084 354488 496136 354494
rect 497476 339320 497504 437448
rect 498844 436146 498896 436152
rect 498844 436088 498896 436094
rect 497464 339314 497516 339320
rect 497464 339256 497516 339262
rect 498856 318580 498884 436088
rect 500224 434786 500276 434792
rect 500224 434728 500276 434734
rect 498844 318574 498896 318580
rect 498844 318516 498896 318522
rect 500236 303416 500264 434728
rect 501604 433358 501656 433364
rect 501604 433300 501656 433306
rect 500224 303410 500276 303416
rect 500224 303352 500276 303358
rect 493324 296610 493376 296616
rect 493324 296552 493376 296558
rect 492312 293958 492364 293964
rect 492312 293900 492364 293906
rect 490564 292530 490616 292536
rect 490564 292472 490616 292478
rect 492956 289878 493008 289884
rect 492956 289820 493008 289826
rect 491944 288450 491996 288456
rect 482282 288418 482338 288427
rect 491944 288392 491996 288398
rect 482282 288353 482338 288362
rect 478633 286922 478689 286931
rect 478633 286857 478689 286866
rect 471244 286682 471296 286688
rect 471244 286624 471296 286630
rect 474912 286594 474921 286650
rect 474977 286594 474986 286650
rect 478647 286622 478675 286857
rect 484952 286682 485004 286688
rect 484766 286650 484822 286659
rect 484822 286630 484952 286636
rect 488632 286682 488684 286688
rect 484822 286624 485004 286630
rect 488538 286650 488594 286659
rect 484822 286608 484992 286624
rect 484766 286585 484822 286594
rect 488594 286630 488632 286636
rect 488594 286624 488684 286630
rect 488594 286608 488672 286624
rect 488538 286585 488594 286594
rect 471704 286546 471756 286552
rect 471704 286488 471756 286494
rect 469022 286404 469586 286410
rect 469074 286398 469086 286404
rect 469138 286398 469150 286404
rect 469202 286398 469214 286404
rect 469266 286398 469278 286404
rect 469330 286398 469342 286404
rect 469394 286398 469406 286404
rect 469458 286398 469470 286404
rect 469522 286398 469534 286404
rect 469266 286352 469276 286398
rect 469332 286352 469342 286398
rect 469022 286342 469036 286352
rect 469092 286342 469116 286352
rect 469172 286342 469196 286352
rect 469252 286342 469276 286352
rect 469332 286342 469356 286352
rect 469412 286342 469436 286352
rect 469492 286342 469516 286352
rect 469572 286342 469586 286352
rect 469022 286340 469586 286342
rect 469074 286318 469086 286340
rect 469138 286318 469150 286340
rect 469202 286318 469214 286340
rect 469266 286318 469278 286340
rect 469330 286318 469342 286340
rect 469394 286318 469406 286340
rect 469458 286318 469470 286340
rect 469522 286318 469534 286340
rect 469266 286288 469276 286318
rect 469332 286288 469342 286318
rect 469022 286276 469036 286288
rect 469092 286276 469116 286288
rect 469172 286276 469196 286288
rect 469252 286276 469276 286288
rect 469332 286276 469356 286288
rect 469412 286276 469436 286288
rect 469492 286276 469516 286288
rect 469572 286276 469586 286288
rect 469266 286262 469276 286276
rect 469332 286262 469342 286276
rect 469074 286238 469086 286262
rect 469138 286238 469150 286262
rect 469202 286238 469214 286262
rect 469266 286238 469278 286262
rect 469330 286238 469342 286262
rect 469394 286238 469406 286262
rect 469458 286238 469470 286262
rect 469522 286238 469534 286262
rect 469266 286224 469276 286238
rect 469332 286224 469342 286238
rect 469022 286212 469036 286224
rect 469092 286212 469116 286224
rect 469172 286212 469196 286224
rect 469252 286212 469276 286224
rect 469332 286212 469356 286224
rect 469412 286212 469436 286224
rect 469492 286212 469516 286224
rect 469572 286212 469586 286224
rect 469266 286182 469276 286212
rect 469332 286182 469342 286212
rect 469074 286160 469086 286182
rect 469138 286160 469150 286182
rect 469202 286160 469214 286182
rect 469266 286160 469278 286182
rect 469330 286160 469342 286182
rect 469394 286160 469406 286182
rect 469458 286160 469470 286182
rect 469522 286160 469534 286182
rect 469022 286158 469586 286160
rect 469022 286148 469036 286158
rect 469092 286148 469116 286158
rect 469172 286148 469196 286158
rect 469252 286148 469276 286158
rect 469332 286148 469356 286158
rect 469412 286148 469436 286158
rect 469492 286148 469516 286158
rect 469572 286148 469586 286158
rect 469266 286102 469276 286148
rect 469332 286102 469342 286148
rect 469074 286096 469086 286102
rect 469138 286096 469150 286102
rect 469202 286096 469214 286102
rect 469266 286096 469278 286102
rect 469330 286096 469342 286102
rect 469394 286096 469406 286102
rect 469458 286096 469470 286102
rect 469522 286096 469534 286102
rect 469022 286090 469586 286096
rect 470262 285316 470826 285322
rect 470314 285310 470326 285316
rect 470378 285310 470390 285316
rect 470442 285310 470454 285316
rect 470506 285310 470518 285316
rect 470570 285310 470582 285316
rect 470634 285310 470646 285316
rect 470698 285310 470710 285316
rect 470762 285310 470774 285316
rect 470506 285264 470516 285310
rect 470572 285264 470582 285310
rect 470262 285254 470276 285264
rect 470332 285254 470356 285264
rect 470412 285254 470436 285264
rect 470492 285254 470516 285264
rect 470572 285254 470596 285264
rect 470652 285254 470676 285264
rect 470732 285254 470756 285264
rect 470812 285254 470826 285264
rect 470262 285252 470826 285254
rect 470314 285230 470326 285252
rect 470378 285230 470390 285252
rect 470442 285230 470454 285252
rect 470506 285230 470518 285252
rect 470570 285230 470582 285252
rect 470634 285230 470646 285252
rect 470698 285230 470710 285252
rect 470762 285230 470774 285252
rect 470506 285200 470516 285230
rect 470572 285200 470582 285230
rect 470262 285188 470276 285200
rect 470332 285188 470356 285200
rect 470412 285188 470436 285200
rect 470492 285188 470516 285200
rect 470572 285188 470596 285200
rect 470652 285188 470676 285200
rect 470732 285188 470756 285200
rect 470812 285188 470826 285200
rect 470506 285174 470516 285188
rect 470572 285174 470582 285188
rect 470314 285150 470326 285174
rect 470378 285150 470390 285174
rect 470442 285150 470454 285174
rect 470506 285150 470518 285174
rect 470570 285150 470582 285174
rect 470634 285150 470646 285174
rect 470698 285150 470710 285174
rect 470762 285150 470774 285174
rect 470506 285136 470516 285150
rect 470572 285136 470582 285150
rect 470262 285124 470276 285136
rect 470332 285124 470356 285136
rect 470412 285124 470436 285136
rect 470492 285124 470516 285136
rect 470572 285124 470596 285136
rect 470652 285124 470676 285136
rect 470732 285124 470756 285136
rect 470812 285124 470826 285136
rect 470506 285094 470516 285124
rect 470572 285094 470582 285124
rect 470314 285072 470326 285094
rect 470378 285072 470390 285094
rect 470442 285072 470454 285094
rect 470506 285072 470518 285094
rect 470570 285072 470582 285094
rect 470634 285072 470646 285094
rect 470698 285072 470710 285094
rect 470762 285072 470774 285094
rect 470262 285070 470826 285072
rect 470262 285060 470276 285070
rect 470332 285060 470356 285070
rect 470412 285060 470436 285070
rect 470492 285060 470516 285070
rect 470572 285060 470596 285070
rect 470652 285060 470676 285070
rect 470732 285060 470756 285070
rect 470812 285060 470826 285070
rect 470506 285014 470516 285060
rect 470572 285014 470582 285060
rect 470314 285008 470326 285014
rect 470378 285008 470390 285014
rect 470442 285008 470454 285014
rect 470506 285008 470518 285014
rect 470570 285008 470582 285014
rect 470634 285008 470646 285014
rect 470698 285008 470710 285014
rect 470762 285008 470774 285014
rect 470262 285002 470826 285008
rect 471716 269144 471744 286488
rect 479432 285866 479484 285872
rect 479432 285808 479484 285814
rect 475752 285490 475804 285496
rect 475752 285432 475804 285438
rect 475764 284308 475792 285432
rect 479444 284308 479472 285808
rect 482204 285792 482373 285820
rect 482204 285707 482232 285792
rect 482190 285698 482246 285707
rect 482190 285633 482246 285642
rect 483204 285490 483256 285496
rect 483204 285432 483256 285438
rect 486884 285490 486936 285496
rect 486884 285432 486936 285438
rect 475752 284302 475804 284308
rect 475752 284244 475804 284250
rect 479432 284302 479484 284308
rect 479432 284244 479484 284250
rect 483216 284240 483244 285432
rect 483204 284234 483256 284240
rect 483204 284176 483256 284182
rect 486896 284172 486924 285432
rect 486884 284166 486936 284172
rect 486884 284108 486936 284114
rect 482374 273322 482430 273331
rect 482374 273257 482430 273266
rect 471704 269138 471756 269144
rect 471704 269080 471756 269086
rect 473636 269138 473688 269144
rect 473636 269080 473688 269086
rect 470262 267489 470826 267495
rect 470314 267483 470326 267489
rect 470378 267483 470390 267489
rect 470442 267483 470454 267489
rect 470506 267483 470518 267489
rect 470570 267483 470582 267489
rect 470634 267483 470646 267489
rect 470698 267483 470710 267489
rect 470762 267483 470774 267489
rect 470506 267437 470516 267483
rect 470572 267437 470582 267483
rect 470262 267427 470276 267437
rect 470332 267427 470356 267437
rect 470412 267427 470436 267437
rect 470492 267427 470516 267437
rect 470572 267427 470596 267437
rect 470652 267427 470676 267437
rect 470732 267427 470756 267437
rect 470812 267427 470826 267437
rect 470262 267425 470826 267427
rect 470314 267403 470326 267425
rect 470378 267403 470390 267425
rect 470442 267403 470454 267425
rect 470506 267403 470518 267425
rect 470570 267403 470582 267425
rect 470634 267403 470646 267425
rect 470698 267403 470710 267425
rect 470762 267403 470774 267425
rect 470506 267373 470516 267403
rect 470572 267373 470582 267403
rect 470262 267361 470276 267373
rect 470332 267361 470356 267373
rect 470412 267361 470436 267373
rect 470492 267361 470516 267373
rect 470572 267361 470596 267373
rect 470652 267361 470676 267373
rect 470732 267361 470756 267373
rect 470812 267361 470826 267373
rect 470506 267347 470516 267361
rect 470572 267347 470582 267361
rect 470314 267323 470326 267347
rect 470378 267323 470390 267347
rect 470442 267323 470454 267347
rect 470506 267323 470518 267347
rect 470570 267323 470582 267347
rect 470634 267323 470646 267347
rect 470698 267323 470710 267347
rect 470762 267323 470774 267347
rect 470506 267309 470516 267323
rect 470572 267309 470582 267323
rect 470262 267297 470276 267309
rect 470332 267297 470356 267309
rect 470412 267297 470436 267309
rect 470492 267297 470516 267309
rect 470572 267297 470596 267309
rect 470652 267297 470676 267309
rect 470732 267297 470756 267309
rect 470812 267297 470826 267309
rect 470506 267267 470516 267297
rect 470572 267267 470582 267297
rect 470314 267245 470326 267267
rect 470378 267245 470390 267267
rect 470442 267245 470454 267267
rect 470506 267245 470518 267267
rect 470570 267245 470582 267267
rect 470634 267245 470646 267267
rect 470698 267245 470710 267267
rect 470762 267245 470774 267267
rect 470262 267243 470826 267245
rect 470262 267233 470276 267243
rect 470332 267233 470356 267243
rect 470412 267233 470436 267243
rect 470492 267233 470516 267243
rect 470572 267233 470596 267243
rect 470652 267233 470676 267243
rect 470732 267233 470756 267243
rect 470812 267233 470826 267243
rect 470506 267187 470516 267233
rect 470572 267187 470582 267233
rect 470314 267181 470326 267187
rect 470378 267181 470390 267187
rect 470442 267181 470454 267187
rect 470506 267181 470518 267187
rect 470570 267181 470582 267187
rect 470634 267181 470646 267187
rect 470698 267181 470710 267187
rect 470762 267181 470774 267187
rect 470262 267175 470826 267181
rect 473648 266699 473676 269080
rect 482388 267347 482416 273257
rect 485502 272642 485558 272651
rect 485502 272577 485558 272586
rect 485516 267347 485544 272577
rect 482374 267338 482430 267347
rect 482374 267273 482430 267282
rect 485502 267338 485558 267347
rect 485502 267273 485558 267282
rect 482374 267066 482430 267075
rect 482374 267001 482430 267010
rect 485410 267066 485466 267075
rect 485410 267001 485466 267010
rect 488446 267066 488502 267075
rect 488446 267001 488502 267010
rect 482388 266780 482416 267001
rect 482379 266752 482416 266780
rect 473636 266693 473688 266699
rect 473636 266635 473688 266641
rect 482379 266630 482407 266752
rect 485424 266616 485452 267001
rect 488460 266644 488488 267001
rect 488460 266616 488497 266644
rect 469022 266403 469586 266409
rect 469074 266397 469086 266403
rect 469138 266397 469150 266403
rect 469202 266397 469214 266403
rect 469266 266397 469278 266403
rect 469330 266397 469342 266403
rect 469394 266397 469406 266403
rect 469458 266397 469470 266403
rect 469522 266397 469534 266403
rect 469266 266351 469276 266397
rect 469332 266351 469342 266397
rect 469022 266341 469036 266351
rect 469092 266341 469116 266351
rect 469172 266341 469196 266351
rect 469252 266341 469276 266351
rect 469332 266341 469356 266351
rect 469412 266341 469436 266351
rect 469492 266341 469516 266351
rect 469572 266341 469586 266351
rect 469022 266339 469586 266341
rect 469074 266317 469086 266339
rect 469138 266317 469150 266339
rect 469202 266317 469214 266339
rect 469266 266317 469278 266339
rect 469330 266317 469342 266339
rect 469394 266317 469406 266339
rect 469458 266317 469470 266339
rect 469522 266317 469534 266339
rect 469266 266287 469276 266317
rect 469332 266287 469342 266317
rect 469022 266275 469036 266287
rect 469092 266275 469116 266287
rect 469172 266275 469196 266287
rect 469252 266275 469276 266287
rect 469332 266275 469356 266287
rect 469412 266275 469436 266287
rect 469492 266275 469516 266287
rect 469572 266275 469586 266287
rect 469266 266261 469276 266275
rect 469332 266261 469342 266275
rect 469074 266237 469086 266261
rect 469138 266237 469150 266261
rect 469202 266237 469214 266261
rect 469266 266237 469278 266261
rect 469330 266237 469342 266261
rect 469394 266237 469406 266261
rect 469458 266237 469470 266261
rect 469522 266237 469534 266261
rect 469266 266223 469276 266237
rect 469332 266223 469342 266237
rect 469022 266211 469036 266223
rect 469092 266211 469116 266223
rect 469172 266211 469196 266223
rect 469252 266211 469276 266223
rect 469332 266211 469356 266223
rect 469412 266211 469436 266223
rect 469492 266211 469516 266223
rect 469572 266211 469586 266223
rect 469266 266181 469276 266211
rect 469332 266181 469342 266211
rect 469074 266159 469086 266181
rect 469138 266159 469150 266181
rect 469202 266159 469214 266181
rect 469266 266159 469278 266181
rect 469330 266159 469342 266181
rect 469394 266159 469406 266181
rect 469458 266159 469470 266181
rect 469522 266159 469534 266181
rect 469022 266157 469586 266159
rect 469022 266147 469036 266157
rect 469092 266147 469116 266157
rect 469172 266147 469196 266157
rect 469252 266147 469276 266157
rect 469332 266147 469356 266157
rect 469412 266147 469436 266157
rect 469492 266147 469516 266157
rect 469572 266147 469586 266157
rect 469266 266101 469276 266147
rect 469332 266101 469342 266147
rect 469074 266095 469086 266101
rect 469138 266095 469150 266101
rect 469202 266095 469214 266101
rect 469266 266095 469278 266101
rect 469330 266095 469342 266101
rect 469394 266095 469406 266101
rect 469458 266095 469470 266101
rect 469522 266095 469534 266101
rect 469022 266089 469586 266095
rect 491956 266016 491984 288392
rect 492968 285668 492996 289820
rect 492956 285662 493008 285668
rect 492956 285604 493008 285610
rect 501616 284104 501644 433300
rect 502984 431998 503036 432004
rect 502984 431940 503036 431946
rect 501604 284098 501656 284104
rect 501604 284040 501656 284046
rect 491944 266010 491996 266016
rect 479062 265978 479118 265987
rect 479118 265950 479341 265964
rect 491944 265952 491996 265958
rect 479118 265936 479355 265950
rect 479062 265913 479118 265922
rect 477132 265874 477184 265880
rect 477132 265816 477184 265822
rect 476275 265692 476303 265814
rect 476275 265664 476344 265692
rect 470262 265316 470826 265322
rect 470314 265310 470326 265316
rect 470378 265310 470390 265316
rect 470442 265310 470454 265316
rect 470506 265310 470518 265316
rect 470570 265310 470582 265316
rect 470634 265310 470646 265316
rect 470698 265310 470710 265316
rect 470762 265310 470774 265316
rect 470506 265264 470516 265310
rect 470572 265264 470582 265310
rect 470262 265254 470276 265264
rect 470332 265254 470356 265264
rect 470412 265254 470436 265264
rect 470492 265254 470516 265264
rect 470572 265254 470596 265264
rect 470652 265254 470676 265264
rect 470732 265254 470756 265264
rect 470812 265254 470826 265264
rect 470262 265252 470826 265254
rect 470314 265230 470326 265252
rect 470378 265230 470390 265252
rect 470442 265230 470454 265252
rect 470506 265230 470518 265252
rect 470570 265230 470582 265252
rect 470634 265230 470646 265252
rect 470698 265230 470710 265252
rect 470762 265230 470774 265252
rect 470506 265200 470516 265230
rect 470572 265200 470582 265230
rect 470262 265188 470276 265200
rect 470332 265188 470356 265200
rect 470412 265188 470436 265200
rect 470492 265188 470516 265200
rect 470572 265188 470596 265200
rect 470652 265188 470676 265200
rect 470732 265188 470756 265200
rect 470812 265188 470826 265200
rect 470506 265174 470516 265188
rect 470572 265174 470582 265188
rect 470314 265150 470326 265174
rect 470378 265150 470390 265174
rect 470442 265150 470454 265174
rect 470506 265150 470518 265174
rect 470570 265150 470582 265174
rect 470634 265150 470646 265174
rect 470698 265150 470710 265174
rect 470762 265150 470774 265174
rect 470506 265136 470516 265150
rect 470572 265136 470582 265150
rect 470262 265124 470276 265136
rect 470332 265124 470356 265136
rect 470412 265124 470436 265136
rect 470492 265124 470516 265136
rect 470572 265124 470596 265136
rect 470652 265124 470676 265136
rect 470732 265124 470756 265136
rect 470812 265124 470826 265136
rect 470506 265094 470516 265124
rect 470572 265094 470582 265124
rect 470314 265072 470326 265094
rect 470378 265072 470390 265094
rect 470442 265072 470454 265094
rect 470506 265072 470518 265094
rect 470570 265072 470582 265094
rect 470634 265072 470646 265094
rect 470698 265072 470710 265094
rect 470762 265072 470774 265094
rect 470262 265070 470826 265072
rect 470262 265060 470276 265070
rect 470332 265060 470356 265070
rect 470412 265060 470436 265070
rect 470492 265060 470516 265070
rect 470572 265060 470596 265070
rect 470652 265060 470676 265070
rect 470732 265060 470756 265070
rect 470812 265060 470826 265070
rect 470506 265014 470516 265060
rect 470572 265014 470582 265060
rect 470314 265008 470326 265014
rect 470378 265008 470390 265014
rect 470442 265008 470454 265014
rect 470506 265008 470518 265014
rect 470570 265008 470582 265014
rect 470634 265008 470646 265014
rect 470698 265008 470710 265014
rect 470762 265008 470774 265014
rect 470262 265002 470826 265008
rect 476316 265012 476344 265664
rect 476486 265026 476542 265035
rect 476316 264984 476486 265012
rect 476486 264961 476542 264970
rect 477144 263568 477172 265816
rect 479327 265692 479355 265936
rect 479327 265664 479380 265692
rect 479352 265012 479380 265664
rect 480168 265489 480220 265495
rect 480168 265431 480220 265437
rect 483204 265489 483256 265495
rect 483204 265431 483256 265437
rect 486240 265489 486292 265495
rect 486240 265431 486292 265437
rect 479522 265026 479578 265035
rect 479352 264984 479522 265012
rect 479522 264961 479578 264970
rect 480180 263568 480208 265431
rect 483216 263568 483244 265431
rect 486252 263568 486280 265431
rect 477132 263562 477184 263568
rect 477132 263504 477184 263510
rect 480168 263562 480220 263568
rect 480168 263504 480220 263510
rect 483204 263562 483256 263568
rect 483204 263504 483256 263510
rect 486240 263562 486292 263568
rect 495072 263562 495124 263568
rect 486240 263504 486292 263510
rect 494808 263510 495072 263516
rect 494808 263504 495124 263510
rect 494808 263500 495112 263504
rect 494796 263494 495112 263500
rect 494848 263488 495112 263494
rect 494796 263436 494848 263442
rect 502996 263364 503024 431940
rect 515416 409836 515444 445880
rect 523684 445870 523736 445876
rect 523684 445812 523736 445818
rect 520924 445802 520976 445808
rect 520924 445744 520976 445750
rect 515404 409830 515456 409836
rect 515404 409772 515456 409778
rect 515404 404390 515456 404396
rect 515404 404332 515456 404338
rect 515416 387804 515444 404332
rect 516784 403030 516836 403036
rect 516784 402972 516836 402978
rect 515404 387798 515456 387804
rect 515404 387740 515456 387746
rect 515404 365766 515456 365772
rect 515404 365708 515456 365714
rect 515416 339388 515444 365708
rect 516796 354620 516824 402972
rect 518164 398882 518216 398888
rect 518164 398824 518216 398830
rect 516784 354614 516836 354620
rect 516784 354556 516836 354562
rect 515404 339382 515456 339388
rect 515404 339324 515456 339330
rect 518176 303484 518204 398824
rect 519544 396094 519596 396100
rect 519544 396036 519596 396042
rect 518164 303478 518216 303484
rect 518164 303420 518216 303426
rect 519556 263432 519584 396036
rect 520936 374000 520964 445744
rect 522304 427850 522356 427856
rect 522304 427792 522356 427798
rect 520924 373994 520976 374000
rect 520924 373936 520976 373942
rect 522316 372572 522344 427792
rect 522304 372566 522356 372572
rect 522304 372508 522356 372514
rect 520924 367126 520976 367132
rect 520924 367068 520976 367074
rect 520936 354688 520964 367068
rect 522304 361618 522356 361624
rect 522304 361560 522356 361566
rect 520924 354682 520976 354688
rect 520924 354624 520976 354630
rect 522316 284240 522344 361560
rect 523696 338096 523724 445812
rect 535460 445734 535512 445740
rect 535460 445676 535512 445682
rect 535472 444827 535500 445676
rect 535458 444818 535514 444827
rect 535458 444753 535514 444762
rect 535458 443458 535514 443467
rect 535458 443393 535514 443402
rect 535472 443020 535500 443393
rect 535460 443014 535512 443020
rect 535460 442956 535512 442962
rect 535458 442098 535514 442107
rect 535458 442033 535514 442042
rect 535472 441660 535500 442033
rect 535460 441654 535512 441660
rect 535460 441596 535512 441602
rect 535458 440738 535514 440747
rect 535458 440673 535514 440682
rect 535472 440300 535500 440673
rect 535460 440294 535512 440300
rect 535460 440236 535512 440242
rect 535458 439378 535514 439387
rect 535458 439313 535514 439322
rect 535472 438940 535500 439313
rect 535460 438934 535512 438940
rect 535460 438876 535512 438882
rect 535458 438018 535514 438027
rect 535458 437953 535514 437962
rect 535472 437512 535500 437953
rect 535460 437506 535512 437512
rect 535460 437448 535512 437454
rect 535458 436658 535514 436667
rect 535458 436593 535514 436602
rect 535472 436152 535500 436593
rect 535460 436146 535512 436152
rect 535460 436088 535512 436094
rect 535458 435298 535514 435307
rect 535458 435233 535514 435242
rect 535472 434792 535500 435233
rect 535460 434786 535512 434792
rect 535460 434728 535512 434734
rect 535458 433938 535514 433947
rect 535458 433873 535514 433882
rect 535472 433364 535500 433873
rect 535460 433358 535512 433364
rect 535460 433300 535512 433306
rect 535458 432578 535514 432587
rect 535458 432513 535514 432522
rect 535472 432004 535500 432513
rect 535460 431998 535512 432004
rect 535460 431940 535512 431946
rect 536116 431227 536144 554000
rect 546682 448082 546738 448091
rect 546682 448017 546738 448026
rect 544198 447946 544254 447955
rect 544198 447881 544254 447890
rect 539230 447810 539286 447819
rect 539230 447745 539286 447754
rect 539244 445756 539272 447745
rect 541714 447266 541770 447275
rect 541714 447201 541770 447210
rect 538692 445742 539272 445756
rect 538692 445728 539258 445742
rect 536102 431218 536158 431227
rect 536102 431153 536158 431162
rect 536746 424418 536802 424427
rect 536746 424353 536802 424362
rect 535460 409830 535512 409836
rect 535460 409772 535512 409778
rect 535472 409331 535500 409772
rect 535458 409322 535514 409331
rect 535458 409257 535514 409266
rect 535460 407110 535512 407116
rect 535460 407052 535512 407058
rect 535472 406611 535500 407052
rect 535458 406602 535514 406611
rect 535458 406537 535514 406546
rect 535458 404562 535514 404571
rect 535458 404497 535514 404506
rect 535472 404396 535500 404497
rect 535460 404390 535512 404396
rect 535460 404332 535512 404338
rect 535458 403202 535514 403211
rect 535458 403137 535514 403146
rect 535472 403036 535500 403137
rect 535460 403030 535512 403036
rect 535460 402972 535512 402978
rect 536378 401706 536434 401715
rect 536378 401641 536434 401650
rect 536286 400346 536342 400355
rect 536286 400281 536342 400290
rect 535458 399122 535514 399131
rect 535458 399057 535514 399066
rect 535472 398888 535500 399057
rect 535460 398882 535512 398888
rect 535460 398824 535512 398830
rect 536102 397490 536158 397499
rect 536102 397425 536158 397434
rect 535458 396402 535514 396411
rect 535458 396337 535514 396346
rect 535472 396100 535500 396337
rect 535460 396094 535512 396100
rect 535460 396036 535512 396042
rect 535460 373994 535512 374000
rect 535460 373936 535512 373942
rect 535472 372883 535500 373936
rect 535458 372874 535514 372883
rect 535458 372809 535514 372818
rect 535460 372566 535512 372572
rect 535460 372508 535512 372514
rect 535472 371523 535500 372508
rect 535458 371514 535514 371523
rect 535458 371449 535514 371458
rect 535460 369846 535512 369852
rect 535460 369788 535512 369794
rect 535472 368803 535500 369788
rect 535458 368794 535514 368803
rect 535458 368729 535514 368738
rect 535458 367434 535514 367443
rect 535458 367369 535514 367378
rect 535472 367132 535500 367369
rect 535460 367126 535512 367132
rect 535460 367068 535512 367074
rect 535458 366074 535514 366083
rect 535458 366009 535514 366018
rect 535472 365772 535500 366009
rect 535460 365766 535512 365772
rect 535460 365708 535512 365714
rect 535458 361994 535514 362003
rect 535458 361929 535514 361938
rect 535472 361624 535500 361929
rect 535460 361618 535512 361624
rect 535460 361560 535512 361566
rect 525064 353322 525116 353328
rect 525064 353264 525116 353270
rect 523684 338090 523736 338096
rect 523684 338032 523736 338038
rect 525076 332588 525104 353264
rect 535460 338090 535512 338096
rect 535460 338032 535512 338038
rect 535472 336843 535500 338032
rect 535458 336834 535514 336843
rect 535458 336769 535514 336778
rect 525064 332582 525116 332588
rect 525064 332524 525116 332530
rect 535460 332582 535512 332588
rect 535460 332524 535512 332530
rect 535472 331403 535500 332524
rect 535458 331394 535514 331403
rect 535458 331329 535514 331338
rect 535460 331222 535512 331228
rect 535460 331164 535512 331170
rect 535472 330043 535500 331164
rect 535458 330034 535514 330043
rect 535458 329969 535514 329978
rect 536010 328674 536066 328683
rect 536010 328609 536066 328618
rect 535458 325954 535514 325963
rect 535458 325889 535514 325898
rect 535472 325720 535500 325889
rect 523684 325714 523736 325720
rect 523684 325656 523736 325662
rect 535460 325714 535512 325720
rect 535460 325656 535512 325662
rect 522304 284234 522356 284240
rect 522304 284176 522356 284182
rect 523696 284172 523724 325656
rect 536024 318648 536052 328609
rect 536012 318642 536064 318648
rect 536012 318584 536064 318590
rect 535460 300826 535512 300832
rect 535458 300794 535460 300803
rect 535512 300794 535514 300803
rect 535458 300729 535514 300738
rect 535460 299466 535512 299472
rect 535458 299434 535460 299443
rect 535512 299434 535514 299443
rect 535458 299369 535514 299378
rect 535460 298106 535512 298112
rect 535458 298074 535460 298083
rect 535512 298074 535514 298083
rect 535458 298009 535514 298018
rect 535458 296714 535514 296723
rect 535458 296649 535514 296658
rect 535552 296678 535604 296684
rect 535472 296616 535500 296649
rect 535552 296620 535604 296626
rect 535460 296610 535512 296616
rect 535460 296552 535512 296558
rect 535564 295363 535592 296620
rect 535550 295354 535606 295363
rect 535460 295318 535512 295324
rect 535550 295289 535606 295298
rect 535460 295260 535512 295266
rect 535472 294003 535500 295260
rect 535458 293994 535514 294003
rect 535458 293929 535514 293938
rect 535552 293958 535604 293964
rect 535552 293900 535604 293906
rect 535564 292643 535592 293900
rect 535550 292634 535606 292643
rect 535550 292569 535606 292578
rect 535460 292530 535512 292536
rect 535460 292472 535512 292478
rect 535472 291283 535500 292472
rect 535458 291274 535514 291283
rect 535458 291209 535514 291218
rect 535458 289914 535514 289923
rect 535458 289849 535460 289858
rect 535512 289849 535514 289858
rect 535460 289820 535512 289826
rect 535458 288554 535514 288563
rect 535458 288489 535514 288498
rect 535472 288456 535500 288489
rect 535460 288450 535512 288456
rect 535460 288392 535512 288398
rect 536116 284308 536144 397425
rect 536194 360634 536250 360643
rect 536194 360569 536250 360578
rect 536104 284302 536156 284308
rect 536104 284244 536156 284250
rect 523684 284166 523736 284172
rect 523684 284108 523736 284114
rect 536208 263568 536236 360569
rect 536300 318784 536328 400281
rect 536392 339456 536420 401641
rect 536760 396003 536788 424353
rect 538692 422296 538720 445728
rect 541728 445371 541756 447201
rect 544212 445779 544240 447881
rect 544198 445770 544254 445779
rect 546696 445756 546724 448017
rect 546696 445742 547000 445756
rect 546710 445728 547000 445742
rect 544198 445705 544254 445714
rect 541714 445362 541770 445371
rect 541714 445297 541770 445306
rect 546972 445196 547000 445728
rect 546960 445190 547012 445196
rect 546960 445132 547012 445138
rect 538692 422268 538904 422296
rect 538876 409172 538904 422268
rect 541714 409322 541770 409331
rect 544290 409322 544346 409331
rect 544226 409280 544290 409308
rect 541714 409257 541770 409266
rect 544290 409257 544346 409266
rect 538784 409144 539258 409172
rect 546710 409144 547276 409172
rect 536746 395994 536802 396003
rect 536746 395929 536802 395938
rect 538784 393316 538812 409144
rect 547248 408204 547276 409144
rect 547236 408198 547288 408204
rect 547236 408140 547288 408146
rect 538692 393288 538812 393316
rect 536746 388378 536802 388387
rect 536746 388313 536802 388322
rect 536562 364714 536618 364723
rect 536562 364649 536618 364658
rect 536470 363354 536526 363363
rect 536470 363289 536526 363298
rect 536380 339450 536432 339456
rect 536380 339392 536432 339398
rect 536378 324594 536434 324603
rect 536378 324529 536434 324538
rect 536288 318778 536340 318784
rect 536288 318720 536340 318726
rect 536196 263562 536248 263568
rect 536196 263504 536248 263510
rect 536392 263500 536420 324529
rect 536484 303620 536512 363289
rect 536576 318716 536604 364649
rect 536760 359283 536788 388313
rect 538692 383656 538720 393288
rect 538692 383628 538812 383656
rect 538784 373268 538812 383628
rect 546710 373376 547092 373404
rect 547064 373320 547092 373376
rect 547052 373314 547104 373320
rect 538784 373240 539258 373268
rect 547052 373256 547104 373262
rect 536746 359274 536802 359283
rect 536746 359209 536802 359218
rect 538784 354676 538812 373240
rect 541714 373146 541770 373155
rect 541714 373081 541770 373090
rect 544198 373146 544254 373155
rect 544198 373081 544254 373090
rect 538692 354648 538812 354676
rect 536746 352474 536802 352483
rect 536746 352409 536802 352418
rect 536654 327314 536710 327323
rect 536654 327249 536710 327258
rect 536564 318710 536616 318716
rect 536564 318652 536616 318658
rect 536472 303614 536524 303620
rect 536472 303556 536524 303562
rect 536668 303552 536696 327249
rect 536760 323243 536788 352409
rect 538692 345016 538720 354648
rect 547144 345026 547196 345032
rect 538692 344988 538904 345016
rect 538876 337772 538904 344988
rect 546972 344988 547144 345016
rect 541714 339554 541770 339563
rect 541714 339489 541770 339498
rect 544198 339554 544254 339563
rect 544198 339489 544254 339498
rect 538784 337744 539258 337772
rect 541728 337758 541756 339489
rect 544212 337758 544240 339489
rect 546972 337772 547000 344988
rect 547144 344968 547196 344974
rect 546710 337756 547000 337772
rect 546710 337750 547012 337756
rect 546710 337744 546960 337750
rect 536746 323234 536802 323243
rect 536746 323169 536802 323178
rect 536746 316434 536802 316443
rect 536746 316369 536802 316378
rect 536656 303546 536708 303552
rect 536656 303488 536708 303494
rect 536760 287203 536788 316369
rect 538784 316036 538812 337744
rect 546960 337692 547012 337698
rect 538784 316008 538904 316036
rect 538876 301732 538904 316008
rect 541714 303786 541770 303795
rect 541714 303721 541770 303730
rect 544198 303786 544254 303795
rect 544198 303721 544254 303730
rect 547052 303750 547104 303756
rect 538876 301704 539258 301732
rect 541728 301718 541756 303721
rect 544212 301718 544240 303721
rect 547052 303692 547104 303698
rect 547064 301732 547092 303692
rect 546710 301704 547092 301732
rect 547340 291147 547368 700297
rect 547432 327051 547460 700433
rect 547512 445190 547564 445196
rect 547512 445132 547564 445138
rect 547524 408204 547552 445132
rect 547512 408198 547564 408204
rect 547512 408140 547564 408146
rect 547524 373320 547552 408140
rect 547512 373314 547564 373320
rect 547512 373256 547564 373262
rect 547524 345032 547552 373256
rect 547892 362955 547920 700569
rect 547984 398587 548012 700705
rect 548062 699818 548118 699827
rect 548062 699753 548118 699762
rect 548076 435443 548104 699753
rect 577022 697912 577586 697918
rect 577074 697906 577086 697912
rect 577138 697906 577150 697912
rect 577202 697906 577214 697912
rect 577266 697906 577278 697912
rect 577330 697906 577342 697912
rect 577394 697906 577406 697912
rect 577458 697906 577470 697912
rect 577522 697906 577534 697912
rect 577266 697860 577276 697906
rect 577332 697860 577342 697906
rect 577022 697850 577036 697860
rect 577092 697850 577116 697860
rect 577172 697850 577196 697860
rect 577252 697850 577276 697860
rect 577332 697850 577356 697860
rect 577412 697850 577436 697860
rect 577492 697850 577516 697860
rect 577572 697850 577586 697860
rect 577022 697848 577586 697850
rect 577074 697826 577086 697848
rect 577138 697826 577150 697848
rect 577202 697826 577214 697848
rect 577266 697826 577278 697848
rect 577330 697826 577342 697848
rect 577394 697826 577406 697848
rect 577458 697826 577470 697848
rect 577522 697826 577534 697848
rect 577266 697796 577276 697826
rect 577332 697796 577342 697826
rect 577022 697784 577036 697796
rect 577092 697784 577116 697796
rect 577172 697784 577196 697796
rect 577252 697784 577276 697796
rect 577332 697784 577356 697796
rect 577412 697784 577436 697796
rect 577492 697784 577516 697796
rect 577572 697784 577586 697796
rect 577266 697770 577276 697784
rect 577332 697770 577342 697784
rect 577074 697746 577086 697770
rect 577138 697746 577150 697770
rect 577202 697746 577214 697770
rect 577266 697746 577278 697770
rect 577330 697746 577342 697770
rect 577394 697746 577406 697770
rect 577458 697746 577470 697770
rect 577522 697746 577534 697770
rect 577266 697732 577276 697746
rect 577332 697732 577342 697746
rect 577022 697720 577036 697732
rect 577092 697720 577116 697732
rect 577172 697720 577196 697732
rect 577252 697720 577276 697732
rect 577332 697720 577356 697732
rect 577412 697720 577436 697732
rect 577492 697720 577516 697732
rect 577572 697720 577586 697732
rect 577266 697690 577276 697720
rect 577332 697690 577342 697720
rect 577074 697668 577086 697690
rect 577138 697668 577150 697690
rect 577202 697668 577214 697690
rect 577266 697668 577278 697690
rect 577330 697668 577342 697690
rect 577394 697668 577406 697690
rect 577458 697668 577470 697690
rect 577522 697668 577534 697690
rect 577022 697666 577586 697668
rect 577022 697656 577036 697666
rect 577092 697656 577116 697666
rect 577172 697656 577196 697666
rect 577252 697656 577276 697666
rect 577332 697656 577356 697666
rect 577412 697656 577436 697666
rect 577492 697656 577516 697666
rect 577572 697656 577586 697666
rect 577266 697610 577276 697656
rect 577332 697610 577342 697656
rect 577074 697604 577086 697610
rect 577138 697604 577150 697610
rect 577202 697604 577214 697610
rect 577266 697604 577278 697610
rect 577330 697604 577342 697610
rect 577394 697604 577406 697610
rect 577458 697604 577470 697610
rect 577522 697604 577534 697610
rect 577022 697598 577586 697604
rect 576605 697236 576661 697244
rect 576603 697235 576661 697236
rect 576603 697230 576605 697235
rect 576655 697178 576661 697179
rect 576603 697172 576661 697178
rect 576605 697170 576661 697172
rect 580906 697234 580962 697243
rect 580906 697169 580962 697178
rect 578262 697117 578826 697123
rect 578314 697111 578326 697117
rect 578378 697111 578390 697117
rect 578442 697111 578454 697117
rect 578506 697111 578518 697117
rect 578570 697111 578582 697117
rect 578634 697111 578646 697117
rect 578698 697111 578710 697117
rect 578762 697111 578774 697117
rect 578506 697065 578516 697111
rect 578572 697065 578582 697111
rect 578262 697055 578276 697065
rect 578332 697055 578356 697065
rect 578412 697055 578436 697065
rect 578492 697055 578516 697065
rect 578572 697055 578596 697065
rect 578652 697055 578676 697065
rect 578732 697055 578756 697065
rect 578812 697055 578826 697065
rect 578262 697053 578826 697055
rect 578314 697031 578326 697053
rect 578378 697031 578390 697053
rect 578442 697031 578454 697053
rect 578506 697031 578518 697053
rect 578570 697031 578582 697053
rect 578634 697031 578646 697053
rect 578698 697031 578710 697053
rect 578762 697031 578774 697053
rect 578506 697001 578516 697031
rect 578572 697001 578582 697031
rect 578262 696989 578276 697001
rect 578332 696989 578356 697001
rect 578412 696989 578436 697001
rect 578492 696989 578516 697001
rect 578572 696989 578596 697001
rect 578652 696989 578676 697001
rect 578732 696989 578756 697001
rect 578812 696989 578826 697001
rect 578506 696975 578516 696989
rect 578572 696975 578582 696989
rect 578314 696951 578326 696975
rect 578378 696951 578390 696975
rect 578442 696951 578454 696975
rect 578506 696951 578518 696975
rect 578570 696951 578582 696975
rect 578634 696951 578646 696975
rect 578698 696951 578710 696975
rect 578762 696951 578774 696975
rect 578506 696937 578516 696951
rect 578572 696937 578582 696951
rect 578262 696925 578276 696937
rect 578332 696925 578356 696937
rect 578412 696925 578436 696937
rect 578492 696925 578516 696937
rect 578572 696925 578596 696937
rect 578652 696925 578676 696937
rect 578732 696925 578756 696937
rect 578812 696925 578826 696937
rect 578506 696895 578516 696925
rect 578572 696895 578582 696925
rect 578314 696873 578326 696895
rect 578378 696873 578390 696895
rect 578442 696873 578454 696895
rect 578506 696873 578518 696895
rect 578570 696873 578582 696895
rect 578634 696873 578646 696895
rect 578698 696873 578710 696895
rect 578762 696873 578774 696895
rect 578262 696871 578826 696873
rect 578262 696861 578276 696871
rect 578332 696861 578356 696871
rect 578412 696861 578436 696871
rect 578492 696861 578516 696871
rect 578572 696861 578596 696871
rect 578652 696861 578676 696871
rect 578732 696861 578756 696871
rect 578812 696861 578826 696871
rect 578506 696815 578516 696861
rect 578572 696815 578582 696861
rect 578314 696809 578326 696815
rect 578378 696809 578390 696815
rect 578442 696809 578454 696815
rect 578506 696809 578518 696815
rect 578570 696809 578582 696815
rect 578634 696809 578646 696815
rect 578698 696809 578710 696815
rect 578762 696809 578774 696815
rect 578262 696803 578826 696809
rect 580262 670714 580318 670723
rect 580262 670649 580318 670658
rect 577022 644736 577586 644742
rect 577074 644730 577086 644736
rect 577138 644730 577150 644736
rect 577202 644730 577214 644736
rect 577266 644730 577278 644736
rect 577330 644730 577342 644736
rect 577394 644730 577406 644736
rect 577458 644730 577470 644736
rect 577522 644730 577534 644736
rect 577266 644684 577276 644730
rect 577332 644684 577342 644730
rect 577022 644674 577036 644684
rect 577092 644674 577116 644684
rect 577172 644674 577196 644684
rect 577252 644674 577276 644684
rect 577332 644674 577356 644684
rect 577412 644674 577436 644684
rect 577492 644674 577516 644684
rect 577572 644674 577586 644684
rect 577022 644672 577586 644674
rect 577074 644650 577086 644672
rect 577138 644650 577150 644672
rect 577202 644650 577214 644672
rect 577266 644650 577278 644672
rect 577330 644650 577342 644672
rect 577394 644650 577406 644672
rect 577458 644650 577470 644672
rect 577522 644650 577534 644672
rect 577266 644620 577276 644650
rect 577332 644620 577342 644650
rect 577022 644608 577036 644620
rect 577092 644608 577116 644620
rect 577172 644608 577196 644620
rect 577252 644608 577276 644620
rect 577332 644608 577356 644620
rect 577412 644608 577436 644620
rect 577492 644608 577516 644620
rect 577572 644608 577586 644620
rect 577266 644594 577276 644608
rect 577332 644594 577342 644608
rect 577074 644570 577086 644594
rect 577138 644570 577150 644594
rect 577202 644570 577214 644594
rect 577266 644570 577278 644594
rect 577330 644570 577342 644594
rect 577394 644570 577406 644594
rect 577458 644570 577470 644594
rect 577522 644570 577534 644594
rect 577266 644556 577276 644570
rect 577332 644556 577342 644570
rect 577022 644544 577036 644556
rect 577092 644544 577116 644556
rect 577172 644544 577196 644556
rect 577252 644544 577276 644556
rect 577332 644544 577356 644556
rect 577412 644544 577436 644556
rect 577492 644544 577516 644556
rect 577572 644544 577586 644556
rect 577266 644514 577276 644544
rect 577332 644514 577342 644544
rect 577074 644492 577086 644514
rect 577138 644492 577150 644514
rect 577202 644492 577214 644514
rect 577266 644492 577278 644514
rect 577330 644492 577342 644514
rect 577394 644492 577406 644514
rect 577458 644492 577470 644514
rect 577522 644492 577534 644514
rect 577022 644490 577586 644492
rect 577022 644480 577036 644490
rect 577092 644480 577116 644490
rect 577172 644480 577196 644490
rect 577252 644480 577276 644490
rect 577332 644480 577356 644490
rect 577412 644480 577436 644490
rect 577492 644480 577516 644490
rect 577572 644480 577586 644490
rect 577266 644434 577276 644480
rect 577332 644434 577342 644480
rect 577074 644428 577086 644434
rect 577138 644428 577150 644434
rect 577202 644428 577214 644434
rect 577266 644428 577278 644434
rect 577330 644428 577342 644434
rect 577394 644428 577406 644434
rect 577458 644428 577470 644434
rect 577522 644428 577534 644434
rect 577022 644422 577586 644428
rect 576605 644060 576661 644068
rect 576603 644059 576661 644060
rect 576603 644054 576605 644059
rect 576655 644002 576661 644003
rect 576603 643996 576661 644002
rect 576605 643994 576661 643996
rect 578262 643941 578826 643947
rect 578314 643935 578326 643941
rect 578378 643935 578390 643941
rect 578442 643935 578454 643941
rect 578506 643935 578518 643941
rect 578570 643935 578582 643941
rect 578634 643935 578646 643941
rect 578698 643935 578710 643941
rect 578762 643935 578774 643941
rect 578506 643889 578516 643935
rect 578572 643889 578582 643935
rect 578262 643879 578276 643889
rect 578332 643879 578356 643889
rect 578412 643879 578436 643889
rect 578492 643879 578516 643889
rect 578572 643879 578596 643889
rect 578652 643879 578676 643889
rect 578732 643879 578756 643889
rect 578812 643879 578826 643889
rect 578262 643877 578826 643879
rect 578314 643855 578326 643877
rect 578378 643855 578390 643877
rect 578442 643855 578454 643877
rect 578506 643855 578518 643877
rect 578570 643855 578582 643877
rect 578634 643855 578646 643877
rect 578698 643855 578710 643877
rect 578762 643855 578774 643877
rect 578506 643825 578516 643855
rect 578572 643825 578582 643855
rect 578262 643813 578276 643825
rect 578332 643813 578356 643825
rect 578412 643813 578436 643825
rect 578492 643813 578516 643825
rect 578572 643813 578596 643825
rect 578652 643813 578676 643825
rect 578732 643813 578756 643825
rect 578812 643813 578826 643825
rect 578506 643799 578516 643813
rect 578572 643799 578582 643813
rect 578314 643775 578326 643799
rect 578378 643775 578390 643799
rect 578442 643775 578454 643799
rect 578506 643775 578518 643799
rect 578570 643775 578582 643799
rect 578634 643775 578646 643799
rect 578698 643775 578710 643799
rect 578762 643775 578774 643799
rect 578506 643761 578516 643775
rect 578572 643761 578582 643775
rect 578262 643749 578276 643761
rect 578332 643749 578356 643761
rect 578412 643749 578436 643761
rect 578492 643749 578516 643761
rect 578572 643749 578596 643761
rect 578652 643749 578676 643761
rect 578732 643749 578756 643761
rect 578812 643749 578826 643761
rect 578506 643719 578516 643749
rect 578572 643719 578582 643749
rect 578314 643697 578326 643719
rect 578378 643697 578390 643719
rect 578442 643697 578454 643719
rect 578506 643697 578518 643719
rect 578570 643697 578582 643719
rect 578634 643697 578646 643719
rect 578698 643697 578710 643719
rect 578762 643697 578774 643719
rect 578262 643695 578826 643697
rect 578262 643685 578276 643695
rect 578332 643685 578356 643695
rect 578412 643685 578436 643695
rect 578492 643685 578516 643695
rect 578572 643685 578596 643695
rect 578652 643685 578676 643695
rect 578732 643685 578756 643695
rect 578812 643685 578826 643695
rect 578506 643639 578516 643685
rect 578572 643639 578582 643685
rect 578314 643633 578326 643639
rect 578378 643633 578390 643639
rect 578442 643633 578454 643639
rect 578506 643633 578518 643639
rect 578570 643633 578582 643639
rect 578634 643633 578646 643639
rect 578698 643633 578710 643639
rect 578762 643633 578774 643639
rect 578262 643627 578826 643633
rect 577022 591696 577586 591702
rect 577074 591690 577086 591696
rect 577138 591690 577150 591696
rect 577202 591690 577214 591696
rect 577266 591690 577278 591696
rect 577330 591690 577342 591696
rect 577394 591690 577406 591696
rect 577458 591690 577470 591696
rect 577522 591690 577534 591696
rect 577266 591644 577276 591690
rect 577332 591644 577342 591690
rect 577022 591634 577036 591644
rect 577092 591634 577116 591644
rect 577172 591634 577196 591644
rect 577252 591634 577276 591644
rect 577332 591634 577356 591644
rect 577412 591634 577436 591644
rect 577492 591634 577516 591644
rect 577572 591634 577586 591644
rect 577022 591632 577586 591634
rect 577074 591610 577086 591632
rect 577138 591610 577150 591632
rect 577202 591610 577214 591632
rect 577266 591610 577278 591632
rect 577330 591610 577342 591632
rect 577394 591610 577406 591632
rect 577458 591610 577470 591632
rect 577522 591610 577534 591632
rect 577266 591580 577276 591610
rect 577332 591580 577342 591610
rect 577022 591568 577036 591580
rect 577092 591568 577116 591580
rect 577172 591568 577196 591580
rect 577252 591568 577276 591580
rect 577332 591568 577356 591580
rect 577412 591568 577436 591580
rect 577492 591568 577516 591580
rect 577572 591568 577586 591580
rect 577266 591554 577276 591568
rect 577332 591554 577342 591568
rect 577074 591530 577086 591554
rect 577138 591530 577150 591554
rect 577202 591530 577214 591554
rect 577266 591530 577278 591554
rect 577330 591530 577342 591554
rect 577394 591530 577406 591554
rect 577458 591530 577470 591554
rect 577522 591530 577534 591554
rect 577266 591516 577276 591530
rect 577332 591516 577342 591530
rect 577022 591504 577036 591516
rect 577092 591504 577116 591516
rect 577172 591504 577196 591516
rect 577252 591504 577276 591516
rect 577332 591504 577356 591516
rect 577412 591504 577436 591516
rect 577492 591504 577516 591516
rect 577572 591504 577586 591516
rect 577266 591474 577276 591504
rect 577332 591474 577342 591504
rect 577074 591452 577086 591474
rect 577138 591452 577150 591474
rect 577202 591452 577214 591474
rect 577266 591452 577278 591474
rect 577330 591452 577342 591474
rect 577394 591452 577406 591474
rect 577458 591452 577470 591474
rect 577522 591452 577534 591474
rect 577022 591450 577586 591452
rect 577022 591440 577036 591450
rect 577092 591440 577116 591450
rect 577172 591440 577196 591450
rect 577252 591440 577276 591450
rect 577332 591440 577356 591450
rect 577412 591440 577436 591450
rect 577492 591440 577516 591450
rect 577572 591440 577586 591450
rect 577266 591394 577276 591440
rect 577332 591394 577342 591440
rect 577074 591388 577086 591394
rect 577138 591388 577150 591394
rect 577202 591388 577214 591394
rect 577266 591388 577278 591394
rect 577330 591388 577342 591394
rect 577394 591388 577406 591394
rect 577458 591388 577470 591394
rect 577522 591388 577534 591394
rect 577022 591382 577586 591388
rect 576605 591020 576661 591028
rect 576603 591019 576661 591020
rect 576603 591014 576605 591019
rect 576655 590962 576661 590963
rect 576603 590956 576661 590962
rect 576605 590954 576661 590956
rect 578262 590901 578826 590907
rect 578314 590895 578326 590901
rect 578378 590895 578390 590901
rect 578442 590895 578454 590901
rect 578506 590895 578518 590901
rect 578570 590895 578582 590901
rect 578634 590895 578646 590901
rect 578698 590895 578710 590901
rect 578762 590895 578774 590901
rect 578506 590849 578516 590895
rect 578572 590849 578582 590895
rect 578262 590839 578276 590849
rect 578332 590839 578356 590849
rect 578412 590839 578436 590849
rect 578492 590839 578516 590849
rect 578572 590839 578596 590849
rect 578652 590839 578676 590849
rect 578732 590839 578756 590849
rect 578812 590839 578826 590849
rect 578262 590837 578826 590839
rect 578314 590815 578326 590837
rect 578378 590815 578390 590837
rect 578442 590815 578454 590837
rect 578506 590815 578518 590837
rect 578570 590815 578582 590837
rect 578634 590815 578646 590837
rect 578698 590815 578710 590837
rect 578762 590815 578774 590837
rect 578506 590785 578516 590815
rect 578572 590785 578582 590815
rect 578262 590773 578276 590785
rect 578332 590773 578356 590785
rect 578412 590773 578436 590785
rect 578492 590773 578516 590785
rect 578572 590773 578596 590785
rect 578652 590773 578676 590785
rect 578732 590773 578756 590785
rect 578812 590773 578826 590785
rect 578506 590759 578516 590773
rect 578572 590759 578582 590773
rect 578314 590735 578326 590759
rect 578378 590735 578390 590759
rect 578442 590735 578454 590759
rect 578506 590735 578518 590759
rect 578570 590735 578582 590759
rect 578634 590735 578646 590759
rect 578698 590735 578710 590759
rect 578762 590735 578774 590759
rect 578506 590721 578516 590735
rect 578572 590721 578582 590735
rect 578262 590709 578276 590721
rect 578332 590709 578356 590721
rect 578412 590709 578436 590721
rect 578492 590709 578516 590721
rect 578572 590709 578596 590721
rect 578652 590709 578676 590721
rect 578732 590709 578756 590721
rect 578812 590709 578826 590721
rect 578506 590679 578516 590709
rect 578572 590679 578582 590709
rect 578314 590657 578326 590679
rect 578378 590657 578390 590679
rect 578442 590657 578454 590679
rect 578506 590657 578518 590679
rect 578570 590657 578582 590679
rect 578634 590657 578646 590679
rect 578698 590657 578710 590679
rect 578762 590657 578774 590679
rect 578262 590655 578826 590657
rect 578262 590645 578276 590655
rect 578332 590645 578356 590655
rect 578412 590645 578436 590655
rect 578492 590645 578516 590655
rect 578572 590645 578596 590655
rect 578652 590645 578676 590655
rect 578732 590645 578756 590655
rect 578812 590645 578826 590655
rect 578506 590599 578516 590645
rect 578572 590599 578582 590645
rect 578314 590593 578326 590599
rect 578378 590593 578390 590599
rect 578442 590593 578454 590599
rect 578506 590593 578518 590599
rect 578570 590593 578582 590599
rect 578634 590593 578646 590599
rect 578698 590593 578710 590599
rect 578762 590593 578774 590599
rect 578262 590587 578826 590593
rect 577022 538520 577586 538526
rect 577074 538514 577086 538520
rect 577138 538514 577150 538520
rect 577202 538514 577214 538520
rect 577266 538514 577278 538520
rect 577330 538514 577342 538520
rect 577394 538514 577406 538520
rect 577458 538514 577470 538520
rect 577522 538514 577534 538520
rect 577266 538468 577276 538514
rect 577332 538468 577342 538514
rect 577022 538458 577036 538468
rect 577092 538458 577116 538468
rect 577172 538458 577196 538468
rect 577252 538458 577276 538468
rect 577332 538458 577356 538468
rect 577412 538458 577436 538468
rect 577492 538458 577516 538468
rect 577572 538458 577586 538468
rect 577022 538456 577586 538458
rect 577074 538434 577086 538456
rect 577138 538434 577150 538456
rect 577202 538434 577214 538456
rect 577266 538434 577278 538456
rect 577330 538434 577342 538456
rect 577394 538434 577406 538456
rect 577458 538434 577470 538456
rect 577522 538434 577534 538456
rect 577266 538404 577276 538434
rect 577332 538404 577342 538434
rect 577022 538392 577036 538404
rect 577092 538392 577116 538404
rect 577172 538392 577196 538404
rect 577252 538392 577276 538404
rect 577332 538392 577356 538404
rect 577412 538392 577436 538404
rect 577492 538392 577516 538404
rect 577572 538392 577586 538404
rect 577266 538378 577276 538392
rect 577332 538378 577342 538392
rect 577074 538354 577086 538378
rect 577138 538354 577150 538378
rect 577202 538354 577214 538378
rect 577266 538354 577278 538378
rect 577330 538354 577342 538378
rect 577394 538354 577406 538378
rect 577458 538354 577470 538378
rect 577522 538354 577534 538378
rect 577266 538340 577276 538354
rect 577332 538340 577342 538354
rect 577022 538328 577036 538340
rect 577092 538328 577116 538340
rect 577172 538328 577196 538340
rect 577252 538328 577276 538340
rect 577332 538328 577356 538340
rect 577412 538328 577436 538340
rect 577492 538328 577516 538340
rect 577572 538328 577586 538340
rect 577266 538298 577276 538328
rect 577332 538298 577342 538328
rect 577074 538276 577086 538298
rect 577138 538276 577150 538298
rect 577202 538276 577214 538298
rect 577266 538276 577278 538298
rect 577330 538276 577342 538298
rect 577394 538276 577406 538298
rect 577458 538276 577470 538298
rect 577522 538276 577534 538298
rect 577022 538274 577586 538276
rect 577022 538264 577036 538274
rect 577092 538264 577116 538274
rect 577172 538264 577196 538274
rect 577252 538264 577276 538274
rect 577332 538264 577356 538274
rect 577412 538264 577436 538274
rect 577492 538264 577516 538274
rect 577572 538264 577586 538274
rect 577266 538218 577276 538264
rect 577332 538218 577342 538264
rect 577074 538212 577086 538218
rect 577138 538212 577150 538218
rect 577202 538212 577214 538218
rect 577266 538212 577278 538218
rect 577330 538212 577342 538218
rect 577394 538212 577406 538218
rect 577458 538212 577470 538218
rect 577522 538212 577534 538218
rect 577022 538206 577586 538212
rect 576605 537844 576661 537852
rect 576603 537843 576661 537844
rect 576603 537838 576605 537843
rect 576655 537786 576661 537787
rect 576603 537780 576661 537786
rect 576605 537778 576661 537780
rect 578262 537725 578826 537731
rect 578314 537719 578326 537725
rect 578378 537719 578390 537725
rect 578442 537719 578454 537725
rect 578506 537719 578518 537725
rect 578570 537719 578582 537725
rect 578634 537719 578646 537725
rect 578698 537719 578710 537725
rect 578762 537719 578774 537725
rect 578506 537673 578516 537719
rect 578572 537673 578582 537719
rect 578262 537663 578276 537673
rect 578332 537663 578356 537673
rect 578412 537663 578436 537673
rect 578492 537663 578516 537673
rect 578572 537663 578596 537673
rect 578652 537663 578676 537673
rect 578732 537663 578756 537673
rect 578812 537663 578826 537673
rect 578262 537661 578826 537663
rect 578314 537639 578326 537661
rect 578378 537639 578390 537661
rect 578442 537639 578454 537661
rect 578506 537639 578518 537661
rect 578570 537639 578582 537661
rect 578634 537639 578646 537661
rect 578698 537639 578710 537661
rect 578762 537639 578774 537661
rect 578506 537609 578516 537639
rect 578572 537609 578582 537639
rect 578262 537597 578276 537609
rect 578332 537597 578356 537609
rect 578412 537597 578436 537609
rect 578492 537597 578516 537609
rect 578572 537597 578596 537609
rect 578652 537597 578676 537609
rect 578732 537597 578756 537609
rect 578812 537597 578826 537609
rect 578506 537583 578516 537597
rect 578572 537583 578582 537597
rect 578314 537559 578326 537583
rect 578378 537559 578390 537583
rect 578442 537559 578454 537583
rect 578506 537559 578518 537583
rect 578570 537559 578582 537583
rect 578634 537559 578646 537583
rect 578698 537559 578710 537583
rect 578762 537559 578774 537583
rect 578506 537545 578516 537559
rect 578572 537545 578582 537559
rect 578262 537533 578276 537545
rect 578332 537533 578356 537545
rect 578412 537533 578436 537545
rect 578492 537533 578516 537545
rect 578572 537533 578596 537545
rect 578652 537533 578676 537545
rect 578732 537533 578756 537545
rect 578812 537533 578826 537545
rect 578506 537503 578516 537533
rect 578572 537503 578582 537533
rect 578314 537481 578326 537503
rect 578378 537481 578390 537503
rect 578442 537481 578454 537503
rect 578506 537481 578518 537503
rect 578570 537481 578582 537503
rect 578634 537481 578646 537503
rect 578698 537481 578710 537503
rect 578762 537481 578774 537503
rect 578262 537479 578826 537481
rect 578262 537469 578276 537479
rect 578332 537469 578356 537479
rect 578412 537469 578436 537479
rect 578492 537469 578516 537479
rect 578572 537469 578596 537479
rect 578652 537469 578676 537479
rect 578732 537469 578756 537479
rect 578812 537469 578826 537479
rect 578506 537423 578516 537469
rect 578572 537423 578582 537469
rect 578314 537417 578326 537423
rect 578378 537417 578390 537423
rect 578442 537417 578454 537423
rect 578506 537417 578518 537423
rect 578570 537417 578582 537423
rect 578634 537417 578646 537423
rect 578698 537417 578710 537423
rect 578762 537417 578774 537423
rect 578262 537411 578826 537417
rect 577022 485344 577586 485350
rect 577074 485338 577086 485344
rect 577138 485338 577150 485344
rect 577202 485338 577214 485344
rect 577266 485338 577278 485344
rect 577330 485338 577342 485344
rect 577394 485338 577406 485344
rect 577458 485338 577470 485344
rect 577522 485338 577534 485344
rect 577266 485292 577276 485338
rect 577332 485292 577342 485338
rect 577022 485282 577036 485292
rect 577092 485282 577116 485292
rect 577172 485282 577196 485292
rect 577252 485282 577276 485292
rect 577332 485282 577356 485292
rect 577412 485282 577436 485292
rect 577492 485282 577516 485292
rect 577572 485282 577586 485292
rect 577022 485280 577586 485282
rect 577074 485258 577086 485280
rect 577138 485258 577150 485280
rect 577202 485258 577214 485280
rect 577266 485258 577278 485280
rect 577330 485258 577342 485280
rect 577394 485258 577406 485280
rect 577458 485258 577470 485280
rect 577522 485258 577534 485280
rect 577266 485228 577276 485258
rect 577332 485228 577342 485258
rect 577022 485216 577036 485228
rect 577092 485216 577116 485228
rect 577172 485216 577196 485228
rect 577252 485216 577276 485228
rect 577332 485216 577356 485228
rect 577412 485216 577436 485228
rect 577492 485216 577516 485228
rect 577572 485216 577586 485228
rect 577266 485202 577276 485216
rect 577332 485202 577342 485216
rect 577074 485178 577086 485202
rect 577138 485178 577150 485202
rect 577202 485178 577214 485202
rect 577266 485178 577278 485202
rect 577330 485178 577342 485202
rect 577394 485178 577406 485202
rect 577458 485178 577470 485202
rect 577522 485178 577534 485202
rect 577266 485164 577276 485178
rect 577332 485164 577342 485178
rect 577022 485152 577036 485164
rect 577092 485152 577116 485164
rect 577172 485152 577196 485164
rect 577252 485152 577276 485164
rect 577332 485152 577356 485164
rect 577412 485152 577436 485164
rect 577492 485152 577516 485164
rect 577572 485152 577586 485164
rect 577266 485122 577276 485152
rect 577332 485122 577342 485152
rect 577074 485100 577086 485122
rect 577138 485100 577150 485122
rect 577202 485100 577214 485122
rect 577266 485100 577278 485122
rect 577330 485100 577342 485122
rect 577394 485100 577406 485122
rect 577458 485100 577470 485122
rect 577522 485100 577534 485122
rect 577022 485098 577586 485100
rect 577022 485088 577036 485098
rect 577092 485088 577116 485098
rect 577172 485088 577196 485098
rect 577252 485088 577276 485098
rect 577332 485088 577356 485098
rect 577412 485088 577436 485098
rect 577492 485088 577516 485098
rect 577572 485088 577586 485098
rect 577266 485042 577276 485088
rect 577332 485042 577342 485088
rect 577074 485036 577086 485042
rect 577138 485036 577150 485042
rect 577202 485036 577214 485042
rect 577266 485036 577278 485042
rect 577330 485036 577342 485042
rect 577394 485036 577406 485042
rect 577458 485036 577470 485042
rect 577522 485036 577534 485042
rect 577022 485030 577586 485036
rect 576605 484668 576661 484676
rect 576603 484667 576661 484668
rect 576603 484662 576605 484667
rect 576655 484610 576661 484611
rect 576603 484604 576661 484610
rect 576605 484602 576661 484604
rect 578262 484549 578826 484555
rect 578314 484543 578326 484549
rect 578378 484543 578390 484549
rect 578442 484543 578454 484549
rect 578506 484543 578518 484549
rect 578570 484543 578582 484549
rect 578634 484543 578646 484549
rect 578698 484543 578710 484549
rect 578762 484543 578774 484549
rect 578506 484497 578516 484543
rect 578572 484497 578582 484543
rect 578262 484487 578276 484497
rect 578332 484487 578356 484497
rect 578412 484487 578436 484497
rect 578492 484487 578516 484497
rect 578572 484487 578596 484497
rect 578652 484487 578676 484497
rect 578732 484487 578756 484497
rect 578812 484487 578826 484497
rect 578262 484485 578826 484487
rect 578314 484463 578326 484485
rect 578378 484463 578390 484485
rect 578442 484463 578454 484485
rect 578506 484463 578518 484485
rect 578570 484463 578582 484485
rect 578634 484463 578646 484485
rect 578698 484463 578710 484485
rect 578762 484463 578774 484485
rect 578506 484433 578516 484463
rect 578572 484433 578582 484463
rect 578262 484421 578276 484433
rect 578332 484421 578356 484433
rect 578412 484421 578436 484433
rect 578492 484421 578516 484433
rect 578572 484421 578596 484433
rect 578652 484421 578676 484433
rect 578732 484421 578756 484433
rect 578812 484421 578826 484433
rect 578506 484407 578516 484421
rect 578572 484407 578582 484421
rect 578314 484383 578326 484407
rect 578378 484383 578390 484407
rect 578442 484383 578454 484407
rect 578506 484383 578518 484407
rect 578570 484383 578582 484407
rect 578634 484383 578646 484407
rect 578698 484383 578710 484407
rect 578762 484383 578774 484407
rect 578506 484369 578516 484383
rect 578572 484369 578582 484383
rect 578262 484357 578276 484369
rect 578332 484357 578356 484369
rect 578412 484357 578436 484369
rect 578492 484357 578516 484369
rect 578572 484357 578596 484369
rect 578652 484357 578676 484369
rect 578732 484357 578756 484369
rect 578812 484357 578826 484369
rect 578506 484327 578516 484357
rect 578572 484327 578582 484357
rect 578314 484305 578326 484327
rect 578378 484305 578390 484327
rect 578442 484305 578454 484327
rect 578506 484305 578518 484327
rect 578570 484305 578582 484327
rect 578634 484305 578646 484327
rect 578698 484305 578710 484327
rect 578762 484305 578774 484327
rect 578262 484303 578826 484305
rect 578262 484293 578276 484303
rect 578332 484293 578356 484303
rect 578412 484293 578436 484303
rect 578492 484293 578516 484303
rect 578572 484293 578596 484303
rect 578652 484293 578676 484303
rect 578732 484293 578756 484303
rect 578812 484293 578826 484303
rect 578506 484247 578516 484293
rect 578572 484247 578582 484293
rect 578314 484241 578326 484247
rect 578378 484241 578390 484247
rect 578442 484241 578454 484247
rect 578506 484241 578518 484247
rect 578570 484241 578582 484247
rect 578634 484241 578646 484247
rect 578698 484241 578710 484247
rect 578762 484241 578774 484247
rect 578262 484235 578826 484241
rect 580170 458146 580226 458155
rect 580170 458081 580226 458090
rect 580184 453356 580212 458081
rect 580172 453350 580224 453356
rect 580172 453292 580224 453298
rect 580276 448091 580304 670649
rect 580906 644058 580962 644067
rect 580906 643993 580962 644002
rect 580446 617538 580502 617547
rect 580446 617473 580502 617482
rect 580262 448082 580318 448091
rect 580262 448017 580318 448026
rect 580460 447955 580488 617473
rect 580906 591018 580962 591027
rect 580906 590953 580962 590962
rect 580630 564362 580686 564371
rect 580630 564297 580686 564306
rect 580446 447946 580502 447955
rect 580446 447881 580502 447890
rect 580644 447275 580672 564297
rect 580906 537842 580962 537851
rect 580906 537777 580962 537786
rect 580814 511322 580870 511331
rect 580814 511257 580870 511266
rect 580828 447819 580856 511257
rect 580906 484666 580962 484675
rect 580906 484601 580962 484610
rect 580814 447810 580870 447819
rect 580814 447745 580870 447754
rect 580630 447266 580686 447275
rect 580630 447201 580686 447210
rect 548062 435434 548118 435443
rect 548062 435369 548118 435378
rect 577022 432304 577586 432310
rect 577074 432298 577086 432304
rect 577138 432298 577150 432304
rect 577202 432298 577214 432304
rect 577266 432298 577278 432304
rect 577330 432298 577342 432304
rect 577394 432298 577406 432304
rect 577458 432298 577470 432304
rect 577522 432298 577534 432304
rect 577266 432252 577276 432298
rect 577332 432252 577342 432298
rect 577022 432242 577036 432252
rect 577092 432242 577116 432252
rect 577172 432242 577196 432252
rect 577252 432242 577276 432252
rect 577332 432242 577356 432252
rect 577412 432242 577436 432252
rect 577492 432242 577516 432252
rect 577572 432242 577586 432252
rect 577022 432240 577586 432242
rect 577074 432218 577086 432240
rect 577138 432218 577150 432240
rect 577202 432218 577214 432240
rect 577266 432218 577278 432240
rect 577330 432218 577342 432240
rect 577394 432218 577406 432240
rect 577458 432218 577470 432240
rect 577522 432218 577534 432240
rect 577266 432188 577276 432218
rect 577332 432188 577342 432218
rect 577022 432176 577036 432188
rect 577092 432176 577116 432188
rect 577172 432176 577196 432188
rect 577252 432176 577276 432188
rect 577332 432176 577356 432188
rect 577412 432176 577436 432188
rect 577492 432176 577516 432188
rect 577572 432176 577586 432188
rect 577266 432162 577276 432176
rect 577332 432162 577342 432176
rect 577074 432138 577086 432162
rect 577138 432138 577150 432162
rect 577202 432138 577214 432162
rect 577266 432138 577278 432162
rect 577330 432138 577342 432162
rect 577394 432138 577406 432162
rect 577458 432138 577470 432162
rect 577522 432138 577534 432162
rect 577266 432124 577276 432138
rect 577332 432124 577342 432138
rect 577022 432112 577036 432124
rect 577092 432112 577116 432124
rect 577172 432112 577196 432124
rect 577252 432112 577276 432124
rect 577332 432112 577356 432124
rect 577412 432112 577436 432124
rect 577492 432112 577516 432124
rect 577572 432112 577586 432124
rect 577266 432082 577276 432112
rect 577332 432082 577342 432112
rect 577074 432060 577086 432082
rect 577138 432060 577150 432082
rect 577202 432060 577214 432082
rect 577266 432060 577278 432082
rect 577330 432060 577342 432082
rect 577394 432060 577406 432082
rect 577458 432060 577470 432082
rect 577522 432060 577534 432082
rect 577022 432058 577586 432060
rect 577022 432048 577036 432058
rect 577092 432048 577116 432058
rect 577172 432048 577196 432058
rect 577252 432048 577276 432058
rect 577332 432048 577356 432058
rect 577412 432048 577436 432058
rect 577492 432048 577516 432058
rect 577572 432048 577586 432058
rect 577266 432002 577276 432048
rect 577332 432002 577342 432048
rect 577074 431996 577086 432002
rect 577138 431996 577150 432002
rect 577202 431996 577214 432002
rect 577266 431996 577278 432002
rect 577330 431996 577342 432002
rect 577394 431996 577406 432002
rect 577458 431996 577470 432002
rect 577522 431996 577534 432002
rect 577022 431990 577586 431996
rect 576605 431628 576661 431636
rect 576603 431627 576661 431628
rect 576603 431622 576605 431627
rect 576655 431570 576661 431571
rect 576603 431564 576661 431570
rect 576605 431562 576661 431564
rect 580906 431626 580962 431635
rect 580906 431561 580962 431570
rect 578262 431509 578826 431515
rect 578314 431503 578326 431509
rect 578378 431503 578390 431509
rect 578442 431503 578454 431509
rect 578506 431503 578518 431509
rect 578570 431503 578582 431509
rect 578634 431503 578646 431509
rect 578698 431503 578710 431509
rect 578762 431503 578774 431509
rect 578506 431457 578516 431503
rect 578572 431457 578582 431503
rect 578262 431447 578276 431457
rect 578332 431447 578356 431457
rect 578412 431447 578436 431457
rect 578492 431447 578516 431457
rect 578572 431447 578596 431457
rect 578652 431447 578676 431457
rect 578732 431447 578756 431457
rect 578812 431447 578826 431457
rect 578262 431445 578826 431447
rect 578314 431423 578326 431445
rect 578378 431423 578390 431445
rect 578442 431423 578454 431445
rect 578506 431423 578518 431445
rect 578570 431423 578582 431445
rect 578634 431423 578646 431445
rect 578698 431423 578710 431445
rect 578762 431423 578774 431445
rect 578506 431393 578516 431423
rect 578572 431393 578582 431423
rect 578262 431381 578276 431393
rect 578332 431381 578356 431393
rect 578412 431381 578436 431393
rect 578492 431381 578516 431393
rect 578572 431381 578596 431393
rect 578652 431381 578676 431393
rect 578732 431381 578756 431393
rect 578812 431381 578826 431393
rect 578506 431367 578516 431381
rect 578572 431367 578582 431381
rect 578314 431343 578326 431367
rect 578378 431343 578390 431367
rect 578442 431343 578454 431367
rect 578506 431343 578518 431367
rect 578570 431343 578582 431367
rect 578634 431343 578646 431367
rect 578698 431343 578710 431367
rect 578762 431343 578774 431367
rect 578506 431329 578516 431343
rect 578572 431329 578582 431343
rect 578262 431317 578276 431329
rect 578332 431317 578356 431329
rect 578412 431317 578436 431329
rect 578492 431317 578516 431329
rect 578572 431317 578596 431329
rect 578652 431317 578676 431329
rect 578732 431317 578756 431329
rect 578812 431317 578826 431329
rect 578506 431287 578516 431317
rect 578572 431287 578582 431317
rect 578314 431265 578326 431287
rect 578378 431265 578390 431287
rect 578442 431265 578454 431287
rect 578506 431265 578518 431287
rect 578570 431265 578582 431287
rect 578634 431265 578646 431287
rect 578698 431265 578710 431287
rect 578762 431265 578774 431287
rect 578262 431263 578826 431265
rect 578262 431253 578276 431263
rect 578332 431253 578356 431263
rect 578412 431253 578436 431263
rect 578492 431253 578516 431263
rect 578572 431253 578596 431263
rect 578652 431253 578676 431263
rect 578732 431253 578756 431263
rect 578812 431253 578826 431263
rect 578506 431207 578516 431253
rect 578572 431207 578582 431253
rect 578314 431201 578326 431207
rect 578378 431201 578390 431207
rect 578442 431201 578454 431207
rect 578506 431201 578518 431207
rect 578570 431201 578582 431207
rect 578634 431201 578646 431207
rect 578698 431201 578710 431207
rect 578762 431201 578774 431207
rect 578262 431195 578826 431201
rect 580170 410002 580226 410011
rect 580170 409937 580226 409946
rect 580184 404979 580212 409937
rect 580170 404970 580226 404979
rect 580170 404905 580226 404914
rect 547970 398578 548026 398587
rect 547970 398513 548026 398522
rect 577022 379128 577586 379134
rect 577074 379122 577086 379128
rect 577138 379122 577150 379128
rect 577202 379122 577214 379128
rect 577266 379122 577278 379128
rect 577330 379122 577342 379128
rect 577394 379122 577406 379128
rect 577458 379122 577470 379128
rect 577522 379122 577534 379128
rect 577266 379076 577276 379122
rect 577332 379076 577342 379122
rect 577022 379066 577036 379076
rect 577092 379066 577116 379076
rect 577172 379066 577196 379076
rect 577252 379066 577276 379076
rect 577332 379066 577356 379076
rect 577412 379066 577436 379076
rect 577492 379066 577516 379076
rect 577572 379066 577586 379076
rect 577022 379064 577586 379066
rect 577074 379042 577086 379064
rect 577138 379042 577150 379064
rect 577202 379042 577214 379064
rect 577266 379042 577278 379064
rect 577330 379042 577342 379064
rect 577394 379042 577406 379064
rect 577458 379042 577470 379064
rect 577522 379042 577534 379064
rect 577266 379012 577276 379042
rect 577332 379012 577342 379042
rect 577022 379000 577036 379012
rect 577092 379000 577116 379012
rect 577172 379000 577196 379012
rect 577252 379000 577276 379012
rect 577332 379000 577356 379012
rect 577412 379000 577436 379012
rect 577492 379000 577516 379012
rect 577572 379000 577586 379012
rect 577266 378986 577276 379000
rect 577332 378986 577342 379000
rect 577074 378962 577086 378986
rect 577138 378962 577150 378986
rect 577202 378962 577214 378986
rect 577266 378962 577278 378986
rect 577330 378962 577342 378986
rect 577394 378962 577406 378986
rect 577458 378962 577470 378986
rect 577522 378962 577534 378986
rect 577266 378948 577276 378962
rect 577332 378948 577342 378962
rect 577022 378936 577036 378948
rect 577092 378936 577116 378948
rect 577172 378936 577196 378948
rect 577252 378936 577276 378948
rect 577332 378936 577356 378948
rect 577412 378936 577436 378948
rect 577492 378936 577516 378948
rect 577572 378936 577586 378948
rect 577266 378906 577276 378936
rect 577332 378906 577342 378936
rect 577074 378884 577086 378906
rect 577138 378884 577150 378906
rect 577202 378884 577214 378906
rect 577266 378884 577278 378906
rect 577330 378884 577342 378906
rect 577394 378884 577406 378906
rect 577458 378884 577470 378906
rect 577522 378884 577534 378906
rect 577022 378882 577586 378884
rect 577022 378872 577036 378882
rect 577092 378872 577116 378882
rect 577172 378872 577196 378882
rect 577252 378872 577276 378882
rect 577332 378872 577356 378882
rect 577412 378872 577436 378882
rect 577492 378872 577516 378882
rect 577572 378872 577586 378882
rect 577266 378826 577276 378872
rect 577332 378826 577342 378872
rect 577074 378820 577086 378826
rect 577138 378820 577150 378826
rect 577202 378820 577214 378826
rect 577266 378820 577278 378826
rect 577330 378820 577342 378826
rect 577394 378820 577406 378826
rect 577458 378820 577470 378826
rect 577522 378820 577534 378826
rect 577022 378814 577586 378820
rect 576605 378452 576661 378460
rect 576603 378451 576661 378452
rect 576603 378446 576605 378451
rect 576655 378394 576661 378395
rect 576603 378388 576661 378394
rect 576605 378386 576661 378388
rect 580906 378450 580962 378459
rect 580906 378385 580962 378394
rect 578262 378333 578826 378339
rect 578314 378327 578326 378333
rect 578378 378327 578390 378333
rect 578442 378327 578454 378333
rect 578506 378327 578518 378333
rect 578570 378327 578582 378333
rect 578634 378327 578646 378333
rect 578698 378327 578710 378333
rect 578762 378327 578774 378333
rect 578506 378281 578516 378327
rect 578572 378281 578582 378327
rect 578262 378271 578276 378281
rect 578332 378271 578356 378281
rect 578412 378271 578436 378281
rect 578492 378271 578516 378281
rect 578572 378271 578596 378281
rect 578652 378271 578676 378281
rect 578732 378271 578756 378281
rect 578812 378271 578826 378281
rect 578262 378269 578826 378271
rect 578314 378247 578326 378269
rect 578378 378247 578390 378269
rect 578442 378247 578454 378269
rect 578506 378247 578518 378269
rect 578570 378247 578582 378269
rect 578634 378247 578646 378269
rect 578698 378247 578710 378269
rect 578762 378247 578774 378269
rect 578506 378217 578516 378247
rect 578572 378217 578582 378247
rect 578262 378205 578276 378217
rect 578332 378205 578356 378217
rect 578412 378205 578436 378217
rect 578492 378205 578516 378217
rect 578572 378205 578596 378217
rect 578652 378205 578676 378217
rect 578732 378205 578756 378217
rect 578812 378205 578826 378217
rect 578506 378191 578516 378205
rect 578572 378191 578582 378205
rect 578314 378167 578326 378191
rect 578378 378167 578390 378191
rect 578442 378167 578454 378191
rect 578506 378167 578518 378191
rect 578570 378167 578582 378191
rect 578634 378167 578646 378191
rect 578698 378167 578710 378191
rect 578762 378167 578774 378191
rect 578506 378153 578516 378167
rect 578572 378153 578582 378167
rect 578262 378141 578276 378153
rect 578332 378141 578356 378153
rect 578412 378141 578436 378153
rect 578492 378141 578516 378153
rect 578572 378141 578596 378153
rect 578652 378141 578676 378153
rect 578732 378141 578756 378153
rect 578812 378141 578826 378153
rect 578506 378111 578516 378141
rect 578572 378111 578582 378141
rect 578314 378089 578326 378111
rect 578378 378089 578390 378111
rect 578442 378089 578454 378111
rect 578506 378089 578518 378111
rect 578570 378089 578582 378111
rect 578634 378089 578646 378111
rect 578698 378089 578710 378111
rect 578762 378089 578774 378111
rect 578262 378087 578826 378089
rect 578262 378077 578276 378087
rect 578332 378077 578356 378087
rect 578412 378077 578436 378087
rect 578492 378077 578516 378087
rect 578572 378077 578596 378087
rect 578652 378077 578676 378087
rect 578732 378077 578756 378087
rect 578812 378077 578826 378087
rect 578506 378031 578516 378077
rect 578572 378031 578582 378077
rect 578314 378025 578326 378031
rect 578378 378025 578390 378031
rect 578442 378025 578454 378031
rect 578506 378025 578518 378031
rect 578570 378025 578582 378031
rect 578634 378025 578646 378031
rect 578698 378025 578710 378031
rect 578762 378025 578774 378031
rect 578262 378019 578826 378025
rect 547878 362946 547934 362955
rect 547878 362881 547934 362890
rect 547512 345026 547564 345032
rect 547512 344968 547564 344974
rect 547512 337750 547564 337756
rect 547512 337692 547564 337698
rect 547418 327042 547474 327051
rect 547418 326977 547474 326986
rect 547524 303756 547552 337692
rect 577022 325952 577586 325958
rect 577074 325946 577086 325952
rect 577138 325946 577150 325952
rect 577202 325946 577214 325952
rect 577266 325946 577278 325952
rect 577330 325946 577342 325952
rect 577394 325946 577406 325952
rect 577458 325946 577470 325952
rect 577522 325946 577534 325952
rect 577266 325900 577276 325946
rect 577332 325900 577342 325946
rect 577022 325890 577036 325900
rect 577092 325890 577116 325900
rect 577172 325890 577196 325900
rect 577252 325890 577276 325900
rect 577332 325890 577356 325900
rect 577412 325890 577436 325900
rect 577492 325890 577516 325900
rect 577572 325890 577586 325900
rect 577022 325888 577586 325890
rect 577074 325866 577086 325888
rect 577138 325866 577150 325888
rect 577202 325866 577214 325888
rect 577266 325866 577278 325888
rect 577330 325866 577342 325888
rect 577394 325866 577406 325888
rect 577458 325866 577470 325888
rect 577522 325866 577534 325888
rect 577266 325836 577276 325866
rect 577332 325836 577342 325866
rect 577022 325824 577036 325836
rect 577092 325824 577116 325836
rect 577172 325824 577196 325836
rect 577252 325824 577276 325836
rect 577332 325824 577356 325836
rect 577412 325824 577436 325836
rect 577492 325824 577516 325836
rect 577572 325824 577586 325836
rect 577266 325810 577276 325824
rect 577332 325810 577342 325824
rect 577074 325786 577086 325810
rect 577138 325786 577150 325810
rect 577202 325786 577214 325810
rect 577266 325786 577278 325810
rect 577330 325786 577342 325810
rect 577394 325786 577406 325810
rect 577458 325786 577470 325810
rect 577522 325786 577534 325810
rect 577266 325772 577276 325786
rect 577332 325772 577342 325786
rect 577022 325760 577036 325772
rect 577092 325760 577116 325772
rect 577172 325760 577196 325772
rect 577252 325760 577276 325772
rect 577332 325760 577356 325772
rect 577412 325760 577436 325772
rect 577492 325760 577516 325772
rect 577572 325760 577586 325772
rect 577266 325730 577276 325760
rect 577332 325730 577342 325760
rect 577074 325708 577086 325730
rect 577138 325708 577150 325730
rect 577202 325708 577214 325730
rect 577266 325708 577278 325730
rect 577330 325708 577342 325730
rect 577394 325708 577406 325730
rect 577458 325708 577470 325730
rect 577522 325708 577534 325730
rect 577022 325706 577586 325708
rect 577022 325696 577036 325706
rect 577092 325696 577116 325706
rect 577172 325696 577196 325706
rect 577252 325696 577276 325706
rect 577332 325696 577356 325706
rect 577412 325696 577436 325706
rect 577492 325696 577516 325706
rect 577572 325696 577586 325706
rect 577266 325650 577276 325696
rect 577332 325650 577342 325696
rect 577074 325644 577086 325650
rect 577138 325644 577150 325650
rect 577202 325644 577214 325650
rect 577266 325644 577278 325650
rect 577330 325644 577342 325650
rect 577394 325644 577406 325650
rect 577458 325644 577470 325650
rect 577522 325644 577534 325650
rect 577022 325638 577586 325644
rect 576605 325276 576661 325284
rect 576603 325275 576661 325276
rect 576603 325270 576605 325275
rect 576655 325218 576661 325219
rect 576603 325212 576661 325218
rect 576605 325210 576661 325212
rect 580906 325274 580962 325283
rect 580906 325209 580962 325218
rect 578262 325157 578826 325163
rect 578314 325151 578326 325157
rect 578378 325151 578390 325157
rect 578442 325151 578454 325157
rect 578506 325151 578518 325157
rect 578570 325151 578582 325157
rect 578634 325151 578646 325157
rect 578698 325151 578710 325157
rect 578762 325151 578774 325157
rect 578506 325105 578516 325151
rect 578572 325105 578582 325151
rect 578262 325095 578276 325105
rect 578332 325095 578356 325105
rect 578412 325095 578436 325105
rect 578492 325095 578516 325105
rect 578572 325095 578596 325105
rect 578652 325095 578676 325105
rect 578732 325095 578756 325105
rect 578812 325095 578826 325105
rect 578262 325093 578826 325095
rect 578314 325071 578326 325093
rect 578378 325071 578390 325093
rect 578442 325071 578454 325093
rect 578506 325071 578518 325093
rect 578570 325071 578582 325093
rect 578634 325071 578646 325093
rect 578698 325071 578710 325093
rect 578762 325071 578774 325093
rect 578506 325041 578516 325071
rect 578572 325041 578582 325071
rect 578262 325029 578276 325041
rect 578332 325029 578356 325041
rect 578412 325029 578436 325041
rect 578492 325029 578516 325041
rect 578572 325029 578596 325041
rect 578652 325029 578676 325041
rect 578732 325029 578756 325041
rect 578812 325029 578826 325041
rect 578506 325015 578516 325029
rect 578572 325015 578582 325029
rect 578314 324991 578326 325015
rect 578378 324991 578390 325015
rect 578442 324991 578454 325015
rect 578506 324991 578518 325015
rect 578570 324991 578582 325015
rect 578634 324991 578646 325015
rect 578698 324991 578710 325015
rect 578762 324991 578774 325015
rect 578506 324977 578516 324991
rect 578572 324977 578582 324991
rect 578262 324965 578276 324977
rect 578332 324965 578356 324977
rect 578412 324965 578436 324977
rect 578492 324965 578516 324977
rect 578572 324965 578596 324977
rect 578652 324965 578676 324977
rect 578732 324965 578756 324977
rect 578812 324965 578826 324977
rect 578506 324935 578516 324965
rect 578572 324935 578582 324965
rect 578314 324913 578326 324935
rect 578378 324913 578390 324935
rect 578442 324913 578454 324935
rect 578506 324913 578518 324935
rect 578570 324913 578582 324935
rect 578634 324913 578646 324935
rect 578698 324913 578710 324935
rect 578762 324913 578774 324935
rect 578262 324911 578826 324913
rect 578262 324901 578276 324911
rect 578332 324901 578356 324911
rect 578412 324901 578436 324911
rect 578492 324901 578516 324911
rect 578572 324901 578596 324911
rect 578652 324901 578676 324911
rect 578732 324901 578756 324911
rect 578812 324901 578826 324911
rect 578506 324855 578516 324901
rect 578572 324855 578582 324901
rect 578314 324849 578326 324855
rect 578378 324849 578390 324855
rect 578442 324849 578454 324855
rect 578506 324849 578518 324855
rect 578570 324849 578582 324855
rect 578634 324849 578646 324855
rect 578698 324849 578710 324855
rect 578762 324849 578774 324855
rect 578262 324843 578826 324849
rect 547512 303750 547564 303756
rect 547512 303692 547564 303698
rect 580170 302290 580226 302299
rect 580170 302225 580226 302234
rect 580184 298763 580212 302225
rect 580170 298754 580226 298763
rect 580170 298689 580226 298698
rect 547326 291138 547382 291147
rect 547326 291073 547382 291082
rect 536746 287194 536802 287203
rect 536746 287129 536802 287138
rect 577022 272912 577586 272918
rect 577074 272906 577086 272912
rect 577138 272906 577150 272912
rect 577202 272906 577214 272912
rect 577266 272906 577278 272912
rect 577330 272906 577342 272912
rect 577394 272906 577406 272912
rect 577458 272906 577470 272912
rect 577522 272906 577534 272912
rect 577266 272860 577276 272906
rect 577332 272860 577342 272906
rect 577022 272850 577036 272860
rect 577092 272850 577116 272860
rect 577172 272850 577196 272860
rect 577252 272850 577276 272860
rect 577332 272850 577356 272860
rect 577412 272850 577436 272860
rect 577492 272850 577516 272860
rect 577572 272850 577586 272860
rect 577022 272848 577586 272850
rect 577074 272826 577086 272848
rect 577138 272826 577150 272848
rect 577202 272826 577214 272848
rect 577266 272826 577278 272848
rect 577330 272826 577342 272848
rect 577394 272826 577406 272848
rect 577458 272826 577470 272848
rect 577522 272826 577534 272848
rect 577266 272796 577276 272826
rect 577332 272796 577342 272826
rect 577022 272784 577036 272796
rect 577092 272784 577116 272796
rect 577172 272784 577196 272796
rect 577252 272784 577276 272796
rect 577332 272784 577356 272796
rect 577412 272784 577436 272796
rect 577492 272784 577516 272796
rect 577572 272784 577586 272796
rect 577266 272770 577276 272784
rect 577332 272770 577342 272784
rect 577074 272746 577086 272770
rect 577138 272746 577150 272770
rect 577202 272746 577214 272770
rect 577266 272746 577278 272770
rect 577330 272746 577342 272770
rect 577394 272746 577406 272770
rect 577458 272746 577470 272770
rect 577522 272746 577534 272770
rect 577266 272732 577276 272746
rect 577332 272732 577342 272746
rect 577022 272720 577036 272732
rect 577092 272720 577116 272732
rect 577172 272720 577196 272732
rect 577252 272720 577276 272732
rect 577332 272720 577356 272732
rect 577412 272720 577436 272732
rect 577492 272720 577516 272732
rect 577572 272720 577586 272732
rect 577266 272690 577276 272720
rect 577332 272690 577342 272720
rect 577074 272668 577086 272690
rect 577138 272668 577150 272690
rect 577202 272668 577214 272690
rect 577266 272668 577278 272690
rect 577330 272668 577342 272690
rect 577394 272668 577406 272690
rect 577458 272668 577470 272690
rect 577522 272668 577534 272690
rect 577022 272666 577586 272668
rect 577022 272656 577036 272666
rect 577092 272656 577116 272666
rect 577172 272656 577196 272666
rect 577252 272656 577276 272666
rect 577332 272656 577356 272666
rect 577412 272656 577436 272666
rect 577492 272656 577516 272666
rect 577572 272656 577586 272666
rect 577266 272610 577276 272656
rect 577332 272610 577342 272656
rect 577074 272604 577086 272610
rect 577138 272604 577150 272610
rect 577202 272604 577214 272610
rect 577266 272604 577278 272610
rect 577330 272604 577342 272610
rect 577394 272604 577406 272610
rect 577458 272604 577470 272610
rect 577522 272604 577534 272610
rect 577022 272598 577586 272604
rect 576605 272236 576661 272244
rect 576603 272235 576661 272236
rect 576603 272230 576605 272235
rect 576655 272178 576661 272179
rect 576603 272172 576661 272178
rect 576605 272170 576661 272172
rect 580906 272234 580962 272243
rect 580906 272169 580962 272178
rect 578262 272117 578826 272123
rect 578314 272111 578326 272117
rect 578378 272111 578390 272117
rect 578442 272111 578454 272117
rect 578506 272111 578518 272117
rect 578570 272111 578582 272117
rect 578634 272111 578646 272117
rect 578698 272111 578710 272117
rect 578762 272111 578774 272117
rect 578506 272065 578516 272111
rect 578572 272065 578582 272111
rect 578262 272055 578276 272065
rect 578332 272055 578356 272065
rect 578412 272055 578436 272065
rect 578492 272055 578516 272065
rect 578572 272055 578596 272065
rect 578652 272055 578676 272065
rect 578732 272055 578756 272065
rect 578812 272055 578826 272065
rect 578262 272053 578826 272055
rect 578314 272031 578326 272053
rect 578378 272031 578390 272053
rect 578442 272031 578454 272053
rect 578506 272031 578518 272053
rect 578570 272031 578582 272053
rect 578634 272031 578646 272053
rect 578698 272031 578710 272053
rect 578762 272031 578774 272053
rect 578506 272001 578516 272031
rect 578572 272001 578582 272031
rect 578262 271989 578276 272001
rect 578332 271989 578356 272001
rect 578412 271989 578436 272001
rect 578492 271989 578516 272001
rect 578572 271989 578596 272001
rect 578652 271989 578676 272001
rect 578732 271989 578756 272001
rect 578812 271989 578826 272001
rect 578506 271975 578516 271989
rect 578572 271975 578582 271989
rect 578314 271951 578326 271975
rect 578378 271951 578390 271975
rect 578442 271951 578454 271975
rect 578506 271951 578518 271975
rect 578570 271951 578582 271975
rect 578634 271951 578646 271975
rect 578698 271951 578710 271975
rect 578762 271951 578774 271975
rect 578506 271937 578516 271951
rect 578572 271937 578582 271951
rect 578262 271925 578276 271937
rect 578332 271925 578356 271937
rect 578412 271925 578436 271937
rect 578492 271925 578516 271937
rect 578572 271925 578596 271937
rect 578652 271925 578676 271937
rect 578732 271925 578756 271937
rect 578812 271925 578826 271937
rect 578506 271895 578516 271925
rect 578572 271895 578582 271925
rect 578314 271873 578326 271895
rect 578378 271873 578390 271895
rect 578442 271873 578454 271895
rect 578506 271873 578518 271895
rect 578570 271873 578582 271895
rect 578634 271873 578646 271895
rect 578698 271873 578710 271895
rect 578762 271873 578774 271895
rect 578262 271871 578826 271873
rect 578262 271861 578276 271871
rect 578332 271861 578356 271871
rect 578412 271861 578436 271871
rect 578492 271861 578516 271871
rect 578572 271861 578596 271871
rect 578652 271861 578676 271871
rect 578732 271861 578756 271871
rect 578812 271861 578826 271871
rect 578506 271815 578516 271861
rect 578572 271815 578582 271861
rect 578314 271809 578326 271815
rect 578378 271809 578390 271815
rect 578442 271809 578454 271815
rect 578506 271809 578518 271815
rect 578570 271809 578582 271815
rect 578634 271809 578646 271815
rect 578698 271809 578710 271815
rect 578762 271809 578774 271815
rect 578262 271803 578826 271809
rect 536380 263494 536432 263500
rect 536380 263436 536432 263442
rect 519544 263426 519596 263432
rect 519544 263368 519596 263374
rect 502984 263358 503036 263364
rect 502984 263300 503036 263306
rect 577022 233065 577586 233071
rect 577074 233059 577086 233065
rect 577138 233059 577150 233065
rect 577202 233059 577214 233065
rect 577266 233059 577278 233065
rect 577330 233059 577342 233065
rect 577394 233059 577406 233065
rect 577458 233059 577470 233065
rect 577522 233059 577534 233065
rect 577266 233013 577276 233059
rect 577332 233013 577342 233059
rect 577022 233003 577036 233013
rect 577092 233003 577116 233013
rect 577172 233003 577196 233013
rect 577252 233003 577276 233013
rect 577332 233003 577356 233013
rect 577412 233003 577436 233013
rect 577492 233003 577516 233013
rect 577572 233003 577586 233013
rect 577022 233001 577586 233003
rect 577074 232979 577086 233001
rect 577138 232979 577150 233001
rect 577202 232979 577214 233001
rect 577266 232979 577278 233001
rect 577330 232979 577342 233001
rect 577394 232979 577406 233001
rect 577458 232979 577470 233001
rect 577522 232979 577534 233001
rect 577266 232949 577276 232979
rect 577332 232949 577342 232979
rect 577022 232937 577036 232949
rect 577092 232937 577116 232949
rect 577172 232937 577196 232949
rect 577252 232937 577276 232949
rect 577332 232937 577356 232949
rect 577412 232937 577436 232949
rect 577492 232937 577516 232949
rect 577572 232937 577586 232949
rect 577266 232923 577276 232937
rect 577332 232923 577342 232937
rect 577074 232899 577086 232923
rect 577138 232899 577150 232923
rect 577202 232899 577214 232923
rect 577266 232899 577278 232923
rect 577330 232899 577342 232923
rect 577394 232899 577406 232923
rect 577458 232899 577470 232923
rect 577522 232899 577534 232923
rect 577266 232885 577276 232899
rect 577332 232885 577342 232899
rect 577022 232873 577036 232885
rect 577092 232873 577116 232885
rect 577172 232873 577196 232885
rect 577252 232873 577276 232885
rect 577332 232873 577356 232885
rect 577412 232873 577436 232885
rect 577492 232873 577516 232885
rect 577572 232873 577586 232885
rect 577266 232843 577276 232873
rect 577332 232843 577342 232873
rect 577074 232821 577086 232843
rect 577138 232821 577150 232843
rect 577202 232821 577214 232843
rect 577266 232821 577278 232843
rect 577330 232821 577342 232843
rect 577394 232821 577406 232843
rect 577458 232821 577470 232843
rect 577522 232821 577534 232843
rect 577022 232819 577586 232821
rect 577022 232809 577036 232819
rect 577092 232809 577116 232819
rect 577172 232809 577196 232819
rect 577252 232809 577276 232819
rect 577332 232809 577356 232819
rect 577412 232809 577436 232819
rect 577492 232809 577516 232819
rect 577572 232809 577586 232819
rect 577266 232763 577276 232809
rect 577332 232763 577342 232809
rect 577074 232757 577086 232763
rect 577138 232757 577150 232763
rect 577202 232757 577214 232763
rect 577266 232757 577278 232763
rect 577330 232757 577342 232763
rect 577394 232757 577406 232763
rect 577458 232757 577470 232763
rect 577522 232757 577534 232763
rect 577022 232751 577586 232757
rect 576605 232389 576661 232397
rect 576603 232388 576661 232389
rect 576603 232383 576605 232388
rect 576655 232331 576661 232332
rect 576603 232325 576661 232331
rect 576605 232323 576661 232325
rect 580906 232386 580962 232395
rect 580906 232321 580962 232330
rect 578262 232270 578826 232276
rect 578314 232264 578326 232270
rect 578378 232264 578390 232270
rect 578442 232264 578454 232270
rect 578506 232264 578518 232270
rect 578570 232264 578582 232270
rect 578634 232264 578646 232270
rect 578698 232264 578710 232270
rect 578762 232264 578774 232270
rect 578506 232218 578516 232264
rect 578572 232218 578582 232264
rect 578262 232208 578276 232218
rect 578332 232208 578356 232218
rect 578412 232208 578436 232218
rect 578492 232208 578516 232218
rect 578572 232208 578596 232218
rect 578652 232208 578676 232218
rect 578732 232208 578756 232218
rect 578812 232208 578826 232218
rect 578262 232206 578826 232208
rect 578314 232184 578326 232206
rect 578378 232184 578390 232206
rect 578442 232184 578454 232206
rect 578506 232184 578518 232206
rect 578570 232184 578582 232206
rect 578634 232184 578646 232206
rect 578698 232184 578710 232206
rect 578762 232184 578774 232206
rect 578506 232154 578516 232184
rect 578572 232154 578582 232184
rect 578262 232142 578276 232154
rect 578332 232142 578356 232154
rect 578412 232142 578436 232154
rect 578492 232142 578516 232154
rect 578572 232142 578596 232154
rect 578652 232142 578676 232154
rect 578732 232142 578756 232154
rect 578812 232142 578826 232154
rect 578506 232128 578516 232142
rect 578572 232128 578582 232142
rect 578314 232104 578326 232128
rect 578378 232104 578390 232128
rect 578442 232104 578454 232128
rect 578506 232104 578518 232128
rect 578570 232104 578582 232128
rect 578634 232104 578646 232128
rect 578698 232104 578710 232128
rect 578762 232104 578774 232128
rect 578506 232090 578516 232104
rect 578572 232090 578582 232104
rect 578262 232078 578276 232090
rect 578332 232078 578356 232090
rect 578412 232078 578436 232090
rect 578492 232078 578516 232090
rect 578572 232078 578596 232090
rect 578652 232078 578676 232090
rect 578732 232078 578756 232090
rect 578812 232078 578826 232090
rect 578506 232048 578516 232078
rect 578572 232048 578582 232078
rect 578314 232026 578326 232048
rect 578378 232026 578390 232048
rect 578442 232026 578454 232048
rect 578506 232026 578518 232048
rect 578570 232026 578582 232048
rect 578634 232026 578646 232048
rect 578698 232026 578710 232048
rect 578762 232026 578774 232048
rect 578262 232024 578826 232026
rect 578262 232014 578276 232024
rect 578332 232014 578356 232024
rect 578412 232014 578436 232024
rect 578492 232014 578516 232024
rect 578572 232014 578596 232024
rect 578652 232014 578676 232024
rect 578732 232014 578756 232024
rect 578812 232014 578826 232024
rect 578506 231968 578516 232014
rect 578572 231968 578582 232014
rect 578314 231962 578326 231968
rect 578378 231962 578390 231968
rect 578442 231962 578454 231968
rect 578506 231962 578518 231968
rect 578570 231962 578582 231968
rect 578634 231962 578646 231968
rect 578698 231962 578710 231968
rect 578762 231962 578774 231968
rect 578262 231956 578826 231962
rect 542 -958 654 482
rect 1646 -958 1758 482
rect 2842 -958 2954 482
rect 4038 -958 4150 482
rect 5234 -958 5346 482
rect 6430 -958 6542 482
rect 7626 -958 7738 482
rect 8730 -958 8842 482
rect 9926 -958 10038 482
rect 11122 -958 11234 482
rect 12318 -958 12430 482
rect 13514 -958 13626 482
rect 14710 -958 14822 482
rect 15906 -958 16018 482
rect 17010 -958 17122 482
rect 18206 -958 18318 482
rect 19402 -958 19514 482
rect 20598 -958 20710 482
rect 21794 -958 21906 482
rect 22990 -958 23102 482
rect 24186 -958 24298 482
rect 25290 -958 25402 482
rect 26486 -958 26598 482
rect 27682 -958 27794 482
rect 28878 -958 28990 482
rect 30074 -958 30186 482
rect 31270 -958 31382 482
rect 32374 -958 32486 482
rect 33570 -958 33682 482
rect 34766 -958 34878 482
rect 35962 -958 36074 482
rect 37158 -958 37270 482
rect 38354 -958 38466 482
rect 39550 -958 39662 482
rect 40654 -958 40766 482
rect 41850 -958 41962 482
rect 43046 -958 43158 482
rect 44242 -958 44354 482
rect 45438 -958 45550 482
rect 46634 -958 46746 482
rect 47830 -958 47942 482
rect 48934 -958 49046 482
rect 50130 -958 50242 482
rect 51326 -958 51438 482
rect 52522 -958 52634 482
rect 53718 -958 53830 482
rect 54914 -958 55026 482
rect 56018 -958 56130 482
rect 57214 -958 57326 482
rect 58410 -958 58522 482
rect 59606 -958 59718 482
rect 60802 -958 60914 482
rect 61998 -958 62110 482
rect 63194 -958 63306 482
rect 64298 -958 64410 482
rect 65494 -958 65606 482
rect 66690 -958 66802 482
rect 67886 -958 67998 482
rect 69082 -958 69194 482
rect 70278 -958 70390 482
rect 71474 -958 71586 482
rect 72578 -958 72690 482
rect 73774 -958 73886 482
rect 74970 -958 75082 482
rect 76166 -958 76278 482
rect 77362 -958 77474 482
rect 78558 -958 78670 482
rect 79662 -958 79774 482
rect 80858 -958 80970 482
rect 82054 -958 82166 482
rect 83250 -958 83362 482
rect 84446 -958 84558 482
rect 85642 -958 85754 482
rect 86838 -958 86950 482
rect 87942 -958 88054 482
rect 89138 -958 89250 482
rect 90334 -958 90446 482
rect 91530 -958 91642 482
rect 92726 -958 92838 482
rect 93922 -958 94034 482
rect 95118 -958 95230 482
rect 96222 -958 96334 482
rect 97418 -958 97530 482
rect 98614 -958 98726 482
rect 99810 -958 99922 482
rect 101006 -958 101118 482
rect 102202 -958 102314 482
rect 103306 -958 103418 482
rect 104502 -958 104614 482
rect 105698 -958 105810 482
rect 106894 -958 107006 482
rect 108090 -958 108202 482
rect 109286 -958 109398 482
rect 110482 -958 110594 482
rect 111586 -958 111698 482
rect 112782 -958 112894 482
rect 113978 -958 114090 482
rect 115174 -958 115286 482
rect 116370 -958 116482 482
rect 117566 -958 117678 482
rect 118762 -958 118874 482
rect 119866 -958 119978 482
rect 121062 -958 121174 482
rect 122258 -958 122370 482
rect 123454 -958 123566 482
rect 124650 -958 124762 482
rect 125846 -958 125958 482
rect 126950 -958 127062 482
rect 128146 -958 128258 482
rect 129342 -958 129454 482
rect 130538 -958 130650 482
rect 131734 -958 131846 482
rect 132930 -958 133042 482
rect 134126 -958 134238 482
rect 135230 -958 135342 482
rect 136426 -958 136538 482
rect 137622 -958 137734 482
rect 138818 -958 138930 482
rect 140014 -958 140126 482
rect 141210 -958 141322 482
rect 142406 -958 142518 482
rect 143510 -958 143622 482
rect 144706 -958 144818 482
rect 145902 -958 146014 482
rect 147098 -958 147210 482
rect 148294 -958 148406 482
rect 149490 -958 149602 482
rect 150594 -958 150706 482
rect 151790 -958 151902 482
rect 152986 -958 153098 482
rect 154182 -958 154294 482
rect 155378 -958 155490 482
rect 156574 -958 156686 482
rect 157770 -958 157882 482
rect 158874 -958 158986 482
rect 160070 -958 160182 482
rect 161266 -958 161378 482
rect 162462 -958 162574 482
rect 163658 -958 163770 482
rect 164854 -958 164966 482
rect 166050 -958 166162 482
rect 167154 -958 167266 482
rect 168350 -958 168462 482
rect 169546 -958 169658 482
rect 170742 -958 170854 482
rect 171938 -958 172050 482
rect 173134 -958 173246 482
rect 174238 -958 174350 482
rect 175434 -958 175546 482
rect 176630 -958 176742 482
rect 177826 -958 177938 482
rect 179022 -958 179134 482
rect 180218 -958 180330 482
rect 181414 -958 181526 482
rect 182518 -958 182630 482
rect 183714 -958 183826 482
rect 184910 -958 185022 482
rect 186106 -958 186218 482
rect 187302 -958 187414 482
rect 188498 -958 188610 482
rect 189694 -958 189806 482
rect 190798 -958 190910 482
rect 191994 -958 192106 482
rect 193190 -958 193302 482
rect 194386 -958 194498 482
rect 195582 -958 195694 482
rect 196778 -958 196890 482
rect 197882 -958 197994 482
rect 199078 -958 199190 482
rect 200274 -958 200386 482
rect 201470 -958 201582 482
rect 202666 -958 202778 482
rect 203862 -958 203974 482
rect 205058 -958 205170 482
rect 206162 -958 206274 482
rect 207358 -958 207470 482
rect 208554 -958 208666 482
rect 209750 -958 209862 482
rect 210946 -958 211058 482
rect 212142 -958 212254 482
rect 213338 -958 213450 482
rect 214442 -958 214554 482
rect 215638 -958 215750 482
rect 216834 -958 216946 482
rect 218030 -958 218142 482
rect 219226 -958 219338 482
rect 220422 -958 220534 482
rect 221526 -958 221638 482
rect 222722 -958 222834 482
rect 223918 -958 224030 482
rect 225114 -958 225226 482
rect 226310 -958 226422 482
rect 227506 -958 227618 482
rect 228702 -958 228814 482
rect 229806 -958 229918 482
rect 231002 -958 231114 482
rect 232198 -958 232310 482
rect 233394 -958 233506 482
rect 234590 -958 234702 482
rect 235786 -958 235898 482
rect 236982 -958 237094 482
rect 238086 -958 238198 482
rect 239282 -958 239394 482
rect 240478 -958 240590 482
rect 241674 -958 241786 482
rect 242870 -958 242982 482
rect 244066 -958 244178 482
rect 245170 -958 245282 482
rect 246366 -958 246478 482
rect 247562 -958 247674 482
rect 248758 -958 248870 482
rect 249954 -958 250066 482
rect 251150 -958 251262 482
rect 252346 -958 252458 482
rect 253450 -958 253562 482
rect 254646 -958 254758 482
rect 255842 -958 255954 482
rect 257038 -958 257150 482
rect 258234 -958 258346 482
rect 259430 -958 259542 482
rect 260626 -958 260738 482
rect 261730 -958 261842 482
rect 262926 -958 263038 482
rect 264122 -958 264234 482
rect 265318 -958 265430 482
rect 266514 -958 266626 482
rect 267710 -958 267822 482
rect 268814 -958 268926 482
rect 270010 -958 270122 482
rect 271206 -958 271318 482
rect 272402 -958 272514 482
rect 273598 -958 273710 482
rect 274794 -958 274906 482
rect 275990 -958 276102 482
rect 277094 -958 277206 482
rect 278290 -958 278402 482
rect 279486 -958 279598 482
rect 280682 -958 280794 482
rect 281878 -958 281990 482
rect 283074 -958 283186 482
rect 284270 -958 284382 482
rect 285374 -958 285486 482
rect 286570 -958 286682 482
rect 287766 -958 287878 482
rect 288962 -958 289074 482
rect 290158 -958 290270 482
rect 291354 -958 291466 482
rect 292550 -958 292662 482
rect 293654 -958 293766 482
rect 294850 -958 294962 482
rect 296046 -958 296158 482
rect 297242 -958 297354 482
rect 298438 -958 298550 482
rect 299634 -958 299746 482
rect 300738 -958 300850 482
rect 301934 -958 302046 482
rect 303130 -958 303242 482
rect 304326 -958 304438 482
rect 305522 -958 305634 482
rect 306718 -958 306830 482
rect 307914 -958 308026 482
rect 309018 -958 309130 482
rect 310214 -958 310326 482
rect 311410 -958 311522 482
rect 312606 -958 312718 482
rect 313802 -958 313914 482
rect 314998 -958 315110 482
rect 316194 -958 316306 482
rect 317298 -958 317410 482
rect 318494 -958 318606 482
rect 319690 -958 319802 482
rect 320886 -958 320998 482
rect 322082 -958 322194 482
rect 323278 -958 323390 482
rect 324382 -958 324494 482
rect 325578 -958 325690 482
rect 326774 -958 326886 482
rect 327970 -958 328082 482
rect 329166 -958 329278 482
rect 330362 -958 330474 482
rect 331558 -958 331670 482
rect 332662 -958 332774 482
rect 333858 -958 333970 482
rect 335054 -958 335166 482
rect 336250 -958 336362 482
rect 337446 -958 337558 482
rect 338642 -958 338754 482
rect 339838 -958 339950 482
rect 340942 -958 341054 482
rect 342138 -958 342250 482
rect 343334 -958 343446 482
rect 344530 -958 344642 482
rect 345726 -958 345838 482
rect 346922 -958 347034 482
rect 348026 -958 348138 482
rect 349222 -958 349334 482
rect 350418 -958 350530 482
rect 351614 -958 351726 482
rect 352810 -958 352922 482
rect 354006 -958 354118 482
rect 355202 -958 355314 482
rect 356306 -958 356418 482
rect 357502 -958 357614 482
rect 358698 -958 358810 482
rect 359894 -958 360006 482
rect 361090 -958 361202 482
rect 362286 -958 362398 482
rect 363482 -958 363594 482
rect 364586 -958 364698 482
rect 365782 -958 365894 482
rect 366978 -958 367090 482
rect 368174 -958 368286 482
rect 369370 -958 369482 482
rect 370566 -958 370678 482
rect 371670 -958 371782 482
rect 372866 -958 372978 482
rect 374062 -958 374174 482
rect 375258 -958 375370 482
rect 376454 -958 376566 482
rect 377650 -958 377762 482
rect 378846 -958 378958 482
rect 379950 -958 380062 482
rect 381146 -958 381258 482
rect 382342 -958 382454 482
rect 383538 -958 383650 482
rect 384734 -958 384846 482
rect 385930 -958 386042 482
rect 387126 -958 387238 482
rect 388230 -958 388342 482
rect 389426 -958 389538 482
rect 390622 -958 390734 482
rect 391818 -958 391930 482
rect 393014 -958 393126 482
rect 394210 -958 394322 482
rect 395314 -958 395426 482
rect 396510 -958 396622 482
rect 397706 -958 397818 482
rect 398902 -958 399014 482
rect 400098 -958 400210 482
rect 401294 -958 401406 482
rect 402490 -958 402602 482
rect 403594 -958 403706 482
rect 404790 -958 404902 482
rect 405986 -958 406098 482
rect 407182 -958 407294 482
rect 408378 -958 408490 482
rect 409574 -958 409686 482
rect 410770 -958 410882 482
rect 411874 -958 411986 482
rect 413070 -958 413182 482
rect 414266 -958 414378 482
rect 415462 -958 415574 482
rect 416658 -958 416770 482
rect 417854 -958 417966 482
rect 418958 -958 419070 482
rect 420154 -958 420266 482
rect 421350 -958 421462 482
rect 422546 -958 422658 482
rect 423742 -958 423854 482
rect 424938 -958 425050 482
rect 426134 -958 426246 482
rect 427238 -958 427350 482
rect 428434 -958 428546 482
rect 429630 -958 429742 482
rect 430826 -958 430938 482
rect 432022 -958 432134 482
rect 433218 -958 433330 482
rect 434414 -958 434526 482
rect 435518 -958 435630 482
rect 436714 -958 436826 482
rect 437910 -958 438022 482
rect 439106 -958 439218 482
rect 440302 -958 440414 482
rect 441498 -958 441610 482
rect 442602 -958 442714 482
rect 443798 -958 443910 482
rect 444994 -958 445106 482
rect 446190 -958 446302 482
rect 447386 -958 447498 482
rect 448582 -958 448694 482
rect 449778 -958 449890 482
rect 450882 -958 450994 482
rect 452078 -958 452190 482
rect 453274 -958 453386 482
rect 454470 -958 454582 482
rect 455666 -958 455778 482
rect 456862 -958 456974 482
rect 458058 -958 458170 482
rect 459162 -958 459274 482
rect 460358 -958 460470 482
rect 461554 -958 461666 482
rect 462750 -958 462862 482
rect 463946 -958 464058 482
rect 465142 -958 465254 482
rect 466246 -958 466358 482
rect 467442 -958 467554 482
rect 468638 -958 468750 482
rect 469834 -958 469946 482
rect 471030 -958 471142 482
rect 472226 -958 472338 482
rect 473422 -958 473534 482
rect 474526 -958 474638 482
rect 475722 -958 475834 482
rect 476918 -958 477030 482
rect 478114 -958 478226 482
rect 479310 -958 479422 482
rect 480506 -958 480618 482
rect 481702 -958 481814 482
rect 482806 -958 482918 482
rect 484002 -958 484114 482
rect 485198 -958 485310 482
rect 486394 -958 486506 482
rect 487590 -958 487702 482
rect 488786 -958 488898 482
rect 489890 -958 490002 482
rect 491086 -958 491198 482
rect 492282 -958 492394 482
rect 493478 -958 493590 482
rect 494674 -958 494786 482
rect 495870 -958 495982 482
rect 497066 -958 497178 482
rect 498170 -958 498282 482
rect 499366 -958 499478 482
rect 500562 -958 500674 482
rect 501758 -958 501870 482
rect 502954 -958 503066 482
rect 504150 -958 504262 482
rect 505346 -958 505458 482
rect 506450 -958 506562 482
rect 507646 -958 507758 482
rect 508842 -958 508954 482
rect 510038 -958 510150 482
rect 511234 -958 511346 482
rect 512430 -958 512542 482
rect 513534 -958 513646 482
rect 514730 -958 514842 482
rect 515926 -958 516038 482
rect 517122 -958 517234 482
rect 518318 -958 518430 482
rect 519514 -958 519626 482
rect 520710 -958 520822 482
rect 521814 -958 521926 482
rect 523010 -958 523122 482
rect 524206 -958 524318 482
rect 525402 -958 525514 482
rect 526598 -958 526710 482
rect 527794 -958 527906 482
rect 528990 -958 529102 482
rect 530094 -958 530206 482
rect 531290 -958 531402 482
rect 532486 -958 532598 482
rect 533682 -958 533794 482
rect 534878 -958 534990 482
rect 536074 -958 536186 482
rect 537178 -958 537290 482
rect 538374 -958 538486 482
rect 539570 -958 539682 482
rect 540766 -958 540878 482
rect 541962 -958 542074 482
rect 543158 -958 543270 482
rect 544354 -958 544466 482
rect 545458 -958 545570 482
rect 546654 -958 546766 482
rect 547850 -958 547962 482
rect 549046 -958 549158 482
rect 550242 -958 550354 482
rect 551438 -958 551550 482
rect 552634 -958 552746 482
rect 553738 -958 553850 482
rect 554934 -958 555046 482
rect 556130 -958 556242 482
rect 557326 -958 557438 482
rect 558522 -958 558634 482
rect 559718 -958 559830 482
rect 560822 -958 560934 482
rect 562018 -958 562130 482
rect 563214 -958 563326 482
rect 564410 -958 564522 482
rect 565606 -958 565718 482
rect 566802 -958 566914 482
rect 567998 -958 568110 482
rect 569102 -958 569214 482
rect 570298 -958 570410 482
rect 571494 -958 571606 482
rect 572690 -958 572802 482
rect 573886 -958 573998 482
rect 575082 -958 575194 482
rect 576278 -958 576390 482
rect 577382 -958 577494 482
rect 578578 -958 578690 482
rect 579774 -958 579886 482
rect 580970 -958 581082 482
rect 582166 -958 582278 482
rect 583362 -958 583474 482
<< via2 >>
rect 254276 703286 254314 703332
rect 254314 703286 254326 703332
rect 254326 703286 254332 703332
rect 254356 703286 254378 703332
rect 254378 703286 254390 703332
rect 254390 703286 254412 703332
rect 254436 703286 254442 703332
rect 254442 703286 254454 703332
rect 254454 703286 254492 703332
rect 254516 703286 254518 703332
rect 254518 703286 254570 703332
rect 254570 703286 254572 703332
rect 254596 703286 254634 703332
rect 254634 703286 254646 703332
rect 254646 703286 254652 703332
rect 254676 703286 254698 703332
rect 254698 703286 254710 703332
rect 254710 703286 254732 703332
rect 254756 703286 254762 703332
rect 254762 703286 254774 703332
rect 254774 703286 254812 703332
rect 254276 703276 254332 703286
rect 254356 703276 254412 703286
rect 254436 703276 254492 703286
rect 254516 703276 254572 703286
rect 254596 703276 254652 703286
rect 254676 703276 254732 703286
rect 254756 703276 254812 703286
rect 254276 703222 254314 703252
rect 254314 703222 254326 703252
rect 254326 703222 254332 703252
rect 254356 703222 254378 703252
rect 254378 703222 254390 703252
rect 254390 703222 254412 703252
rect 254436 703222 254442 703252
rect 254442 703222 254454 703252
rect 254454 703222 254492 703252
rect 254516 703222 254518 703252
rect 254518 703222 254570 703252
rect 254570 703222 254572 703252
rect 254596 703222 254634 703252
rect 254634 703222 254646 703252
rect 254646 703222 254652 703252
rect 254676 703222 254698 703252
rect 254698 703222 254710 703252
rect 254710 703222 254732 703252
rect 254756 703222 254762 703252
rect 254762 703222 254774 703252
rect 254774 703222 254812 703252
rect 254276 703210 254332 703222
rect 254356 703210 254412 703222
rect 254436 703210 254492 703222
rect 254516 703210 254572 703222
rect 254596 703210 254652 703222
rect 254676 703210 254732 703222
rect 254756 703210 254812 703222
rect 254276 703196 254314 703210
rect 254314 703196 254326 703210
rect 254326 703196 254332 703210
rect 254356 703196 254378 703210
rect 254378 703196 254390 703210
rect 254390 703196 254412 703210
rect 254436 703196 254442 703210
rect 254442 703196 254454 703210
rect 254454 703196 254492 703210
rect 254516 703196 254518 703210
rect 254518 703196 254570 703210
rect 254570 703196 254572 703210
rect 254596 703196 254634 703210
rect 254634 703196 254646 703210
rect 254646 703196 254652 703210
rect 254676 703196 254698 703210
rect 254698 703196 254710 703210
rect 254710 703196 254732 703210
rect 254756 703196 254762 703210
rect 254762 703196 254774 703210
rect 254774 703196 254812 703210
rect 254276 703158 254314 703172
rect 254314 703158 254326 703172
rect 254326 703158 254332 703172
rect 254356 703158 254378 703172
rect 254378 703158 254390 703172
rect 254390 703158 254412 703172
rect 254436 703158 254442 703172
rect 254442 703158 254454 703172
rect 254454 703158 254492 703172
rect 254516 703158 254518 703172
rect 254518 703158 254570 703172
rect 254570 703158 254572 703172
rect 254596 703158 254634 703172
rect 254634 703158 254646 703172
rect 254646 703158 254652 703172
rect 254676 703158 254698 703172
rect 254698 703158 254710 703172
rect 254710 703158 254732 703172
rect 254756 703158 254762 703172
rect 254762 703158 254774 703172
rect 254774 703158 254812 703172
rect 254276 703146 254332 703158
rect 254356 703146 254412 703158
rect 254436 703146 254492 703158
rect 254516 703146 254572 703158
rect 254596 703146 254652 703158
rect 254676 703146 254732 703158
rect 254756 703146 254812 703158
rect 254276 703116 254314 703146
rect 254314 703116 254326 703146
rect 254326 703116 254332 703146
rect 254356 703116 254378 703146
rect 254378 703116 254390 703146
rect 254390 703116 254412 703146
rect 254436 703116 254442 703146
rect 254442 703116 254454 703146
rect 254454 703116 254492 703146
rect 254516 703116 254518 703146
rect 254518 703116 254570 703146
rect 254570 703116 254572 703146
rect 254596 703116 254634 703146
rect 254634 703116 254646 703146
rect 254646 703116 254652 703146
rect 254676 703116 254698 703146
rect 254698 703116 254710 703146
rect 254710 703116 254732 703146
rect 254756 703116 254762 703146
rect 254762 703116 254774 703146
rect 254774 703116 254812 703146
rect 254276 703082 254332 703092
rect 254356 703082 254412 703092
rect 254436 703082 254492 703092
rect 254516 703082 254572 703092
rect 254596 703082 254652 703092
rect 254676 703082 254732 703092
rect 254756 703082 254812 703092
rect 254276 703036 254314 703082
rect 254314 703036 254326 703082
rect 254326 703036 254332 703082
rect 254356 703036 254378 703082
rect 254378 703036 254390 703082
rect 254390 703036 254412 703082
rect 254436 703036 254442 703082
rect 254442 703036 254454 703082
rect 254454 703036 254492 703082
rect 254516 703036 254518 703082
rect 254518 703036 254570 703082
rect 254570 703036 254572 703082
rect 254596 703036 254634 703082
rect 254634 703036 254646 703082
rect 254646 703036 254652 703082
rect 254676 703036 254698 703082
rect 254698 703036 254710 703082
rect 254710 703036 254732 703082
rect 254756 703036 254762 703082
rect 254762 703036 254774 703082
rect 254774 703036 254812 703082
rect 253036 702518 253074 702564
rect 253074 702518 253086 702564
rect 253086 702518 253092 702564
rect 253116 702518 253138 702564
rect 253138 702518 253150 702564
rect 253150 702518 253172 702564
rect 253196 702518 253202 702564
rect 253202 702518 253214 702564
rect 253214 702518 253252 702564
rect 253276 702518 253278 702564
rect 253278 702518 253330 702564
rect 253330 702518 253332 702564
rect 253356 702518 253394 702564
rect 253394 702518 253406 702564
rect 253406 702518 253412 702564
rect 253436 702518 253458 702564
rect 253458 702518 253470 702564
rect 253470 702518 253492 702564
rect 253516 702518 253522 702564
rect 253522 702518 253534 702564
rect 253534 702518 253572 702564
rect 253036 702508 253092 702518
rect 253116 702508 253172 702518
rect 253196 702508 253252 702518
rect 253276 702508 253332 702518
rect 253356 702508 253412 702518
rect 253436 702508 253492 702518
rect 253516 702508 253572 702518
rect 253036 702454 253074 702484
rect 253074 702454 253086 702484
rect 253086 702454 253092 702484
rect 253116 702454 253138 702484
rect 253138 702454 253150 702484
rect 253150 702454 253172 702484
rect 253196 702454 253202 702484
rect 253202 702454 253214 702484
rect 253214 702454 253252 702484
rect 253276 702454 253278 702484
rect 253278 702454 253330 702484
rect 253330 702454 253332 702484
rect 253356 702454 253394 702484
rect 253394 702454 253406 702484
rect 253406 702454 253412 702484
rect 253436 702454 253458 702484
rect 253458 702454 253470 702484
rect 253470 702454 253492 702484
rect 253516 702454 253522 702484
rect 253522 702454 253534 702484
rect 253534 702454 253572 702484
rect 253036 702442 253092 702454
rect 253116 702442 253172 702454
rect 253196 702442 253252 702454
rect 253276 702442 253332 702454
rect 253356 702442 253412 702454
rect 253436 702442 253492 702454
rect 253516 702442 253572 702454
rect 253036 702428 253074 702442
rect 253074 702428 253086 702442
rect 253086 702428 253092 702442
rect 253116 702428 253138 702442
rect 253138 702428 253150 702442
rect 253150 702428 253172 702442
rect 253196 702428 253202 702442
rect 253202 702428 253214 702442
rect 253214 702428 253252 702442
rect 253276 702428 253278 702442
rect 253278 702428 253330 702442
rect 253330 702428 253332 702442
rect 253356 702428 253394 702442
rect 253394 702428 253406 702442
rect 253406 702428 253412 702442
rect 253436 702428 253458 702442
rect 253458 702428 253470 702442
rect 253470 702428 253492 702442
rect 253516 702428 253522 702442
rect 253522 702428 253534 702442
rect 253534 702428 253572 702442
rect 253036 702390 253074 702404
rect 253074 702390 253086 702404
rect 253086 702390 253092 702404
rect 253116 702390 253138 702404
rect 253138 702390 253150 702404
rect 253150 702390 253172 702404
rect 253196 702390 253202 702404
rect 253202 702390 253214 702404
rect 253214 702390 253252 702404
rect 253276 702390 253278 702404
rect 253278 702390 253330 702404
rect 253330 702390 253332 702404
rect 253356 702390 253394 702404
rect 253394 702390 253406 702404
rect 253406 702390 253412 702404
rect 253436 702390 253458 702404
rect 253458 702390 253470 702404
rect 253470 702390 253492 702404
rect 253516 702390 253522 702404
rect 253522 702390 253534 702404
rect 253534 702390 253572 702404
rect 253036 702378 253092 702390
rect 253116 702378 253172 702390
rect 253196 702378 253252 702390
rect 253276 702378 253332 702390
rect 253356 702378 253412 702390
rect 253436 702378 253492 702390
rect 253516 702378 253572 702390
rect 253036 702348 253074 702378
rect 253074 702348 253086 702378
rect 253086 702348 253092 702378
rect 253116 702348 253138 702378
rect 253138 702348 253150 702378
rect 253150 702348 253172 702378
rect 253196 702348 253202 702378
rect 253202 702348 253214 702378
rect 253214 702348 253252 702378
rect 253276 702348 253278 702378
rect 253278 702348 253330 702378
rect 253330 702348 253332 702378
rect 253356 702348 253394 702378
rect 253394 702348 253406 702378
rect 253406 702348 253412 702378
rect 253436 702348 253458 702378
rect 253458 702348 253470 702378
rect 253470 702348 253492 702378
rect 253516 702348 253522 702378
rect 253522 702348 253534 702378
rect 253534 702348 253572 702378
rect 253036 702314 253092 702324
rect 253116 702314 253172 702324
rect 253196 702314 253252 702324
rect 253276 702314 253332 702324
rect 253356 702314 253412 702324
rect 253436 702314 253492 702324
rect 253516 702314 253572 702324
rect 253036 702268 253074 702314
rect 253074 702268 253086 702314
rect 253086 702268 253092 702314
rect 253116 702268 253138 702314
rect 253138 702268 253150 702314
rect 253150 702268 253172 702314
rect 253196 702268 253202 702314
rect 253202 702268 253214 702314
rect 253214 702268 253252 702314
rect 253276 702268 253278 702314
rect 253278 702268 253330 702314
rect 253330 702268 253332 702314
rect 253356 702268 253394 702314
rect 253394 702268 253406 702314
rect 253406 702268 253412 702314
rect 253436 702268 253458 702314
rect 253458 702268 253470 702314
rect 253470 702268 253492 702314
rect 253516 702268 253522 702314
rect 253522 702268 253534 702314
rect 253534 702268 253572 702314
rect 326276 703326 326314 703372
rect 326314 703326 326326 703372
rect 326326 703326 326332 703372
rect 326356 703326 326378 703372
rect 326378 703326 326390 703372
rect 326390 703326 326412 703372
rect 326436 703326 326442 703372
rect 326442 703326 326454 703372
rect 326454 703326 326492 703372
rect 326516 703326 326518 703372
rect 326518 703326 326570 703372
rect 326570 703326 326572 703372
rect 326596 703326 326634 703372
rect 326634 703326 326646 703372
rect 326646 703326 326652 703372
rect 326676 703326 326698 703372
rect 326698 703326 326710 703372
rect 326710 703326 326732 703372
rect 326756 703326 326762 703372
rect 326762 703326 326774 703372
rect 326774 703326 326812 703372
rect 326276 703316 326332 703326
rect 326356 703316 326412 703326
rect 326436 703316 326492 703326
rect 326516 703316 326572 703326
rect 326596 703316 326652 703326
rect 326676 703316 326732 703326
rect 326756 703316 326812 703326
rect 326276 703262 326314 703292
rect 326314 703262 326326 703292
rect 326326 703262 326332 703292
rect 326356 703262 326378 703292
rect 326378 703262 326390 703292
rect 326390 703262 326412 703292
rect 326436 703262 326442 703292
rect 326442 703262 326454 703292
rect 326454 703262 326492 703292
rect 326516 703262 326518 703292
rect 326518 703262 326570 703292
rect 326570 703262 326572 703292
rect 326596 703262 326634 703292
rect 326634 703262 326646 703292
rect 326646 703262 326652 703292
rect 326676 703262 326698 703292
rect 326698 703262 326710 703292
rect 326710 703262 326732 703292
rect 326756 703262 326762 703292
rect 326762 703262 326774 703292
rect 326774 703262 326812 703292
rect 326276 703250 326332 703262
rect 326356 703250 326412 703262
rect 326436 703250 326492 703262
rect 326516 703250 326572 703262
rect 326596 703250 326652 703262
rect 326676 703250 326732 703262
rect 326756 703250 326812 703262
rect 326276 703236 326314 703250
rect 326314 703236 326326 703250
rect 326326 703236 326332 703250
rect 326356 703236 326378 703250
rect 326378 703236 326390 703250
rect 326390 703236 326412 703250
rect 326436 703236 326442 703250
rect 326442 703236 326454 703250
rect 326454 703236 326492 703250
rect 326516 703236 326518 703250
rect 326518 703236 326570 703250
rect 326570 703236 326572 703250
rect 326596 703236 326634 703250
rect 326634 703236 326646 703250
rect 326646 703236 326652 703250
rect 326676 703236 326698 703250
rect 326698 703236 326710 703250
rect 326710 703236 326732 703250
rect 326756 703236 326762 703250
rect 326762 703236 326774 703250
rect 326774 703236 326812 703250
rect 326276 703198 326314 703212
rect 326314 703198 326326 703212
rect 326326 703198 326332 703212
rect 326356 703198 326378 703212
rect 326378 703198 326390 703212
rect 326390 703198 326412 703212
rect 326436 703198 326442 703212
rect 326442 703198 326454 703212
rect 326454 703198 326492 703212
rect 326516 703198 326518 703212
rect 326518 703198 326570 703212
rect 326570 703198 326572 703212
rect 326596 703198 326634 703212
rect 326634 703198 326646 703212
rect 326646 703198 326652 703212
rect 326676 703198 326698 703212
rect 326698 703198 326710 703212
rect 326710 703198 326732 703212
rect 326756 703198 326762 703212
rect 326762 703198 326774 703212
rect 326774 703198 326812 703212
rect 326276 703186 326332 703198
rect 326356 703186 326412 703198
rect 326436 703186 326492 703198
rect 326516 703186 326572 703198
rect 326596 703186 326652 703198
rect 326676 703186 326732 703198
rect 326756 703186 326812 703198
rect 326276 703156 326314 703186
rect 326314 703156 326326 703186
rect 326326 703156 326332 703186
rect 326356 703156 326378 703186
rect 326378 703156 326390 703186
rect 326390 703156 326412 703186
rect 326436 703156 326442 703186
rect 326442 703156 326454 703186
rect 326454 703156 326492 703186
rect 326516 703156 326518 703186
rect 326518 703156 326570 703186
rect 326570 703156 326572 703186
rect 326596 703156 326634 703186
rect 326634 703156 326646 703186
rect 326646 703156 326652 703186
rect 326676 703156 326698 703186
rect 326698 703156 326710 703186
rect 326710 703156 326732 703186
rect 326756 703156 326762 703186
rect 326762 703156 326774 703186
rect 326774 703156 326812 703186
rect 326276 703122 326332 703132
rect 326356 703122 326412 703132
rect 326436 703122 326492 703132
rect 326516 703122 326572 703132
rect 326596 703122 326652 703132
rect 326676 703122 326732 703132
rect 326756 703122 326812 703132
rect 326276 703076 326314 703122
rect 326314 703076 326326 703122
rect 326326 703076 326332 703122
rect 326356 703076 326378 703122
rect 326378 703076 326390 703122
rect 326390 703076 326412 703122
rect 326436 703076 326442 703122
rect 326442 703076 326454 703122
rect 326454 703076 326492 703122
rect 326516 703076 326518 703122
rect 326518 703076 326570 703122
rect 326570 703076 326572 703122
rect 326596 703076 326634 703122
rect 326634 703076 326646 703122
rect 326646 703076 326652 703122
rect 326676 703076 326698 703122
rect 326698 703076 326710 703122
rect 326710 703076 326732 703122
rect 326756 703076 326762 703122
rect 326762 703076 326774 703122
rect 326774 703076 326812 703122
rect 325036 702558 325074 702604
rect 325074 702558 325086 702604
rect 325086 702558 325092 702604
rect 325116 702558 325138 702604
rect 325138 702558 325150 702604
rect 325150 702558 325172 702604
rect 325196 702558 325202 702604
rect 325202 702558 325214 702604
rect 325214 702558 325252 702604
rect 325276 702558 325278 702604
rect 325278 702558 325330 702604
rect 325330 702558 325332 702604
rect 325356 702558 325394 702604
rect 325394 702558 325406 702604
rect 325406 702558 325412 702604
rect 325436 702558 325458 702604
rect 325458 702558 325470 702604
rect 325470 702558 325492 702604
rect 325516 702558 325522 702604
rect 325522 702558 325534 702604
rect 325534 702558 325572 702604
rect 325036 702548 325092 702558
rect 325116 702548 325172 702558
rect 325196 702548 325252 702558
rect 325276 702548 325332 702558
rect 325356 702548 325412 702558
rect 325436 702548 325492 702558
rect 325516 702548 325572 702558
rect 325036 702494 325074 702524
rect 325074 702494 325086 702524
rect 325086 702494 325092 702524
rect 325116 702494 325138 702524
rect 325138 702494 325150 702524
rect 325150 702494 325172 702524
rect 325196 702494 325202 702524
rect 325202 702494 325214 702524
rect 325214 702494 325252 702524
rect 325276 702494 325278 702524
rect 325278 702494 325330 702524
rect 325330 702494 325332 702524
rect 325356 702494 325394 702524
rect 325394 702494 325406 702524
rect 325406 702494 325412 702524
rect 325436 702494 325458 702524
rect 325458 702494 325470 702524
rect 325470 702494 325492 702524
rect 325516 702494 325522 702524
rect 325522 702494 325534 702524
rect 325534 702494 325572 702524
rect 325036 702482 325092 702494
rect 325116 702482 325172 702494
rect 325196 702482 325252 702494
rect 325276 702482 325332 702494
rect 325356 702482 325412 702494
rect 325436 702482 325492 702494
rect 325516 702482 325572 702494
rect 325036 702468 325074 702482
rect 325074 702468 325086 702482
rect 325086 702468 325092 702482
rect 325116 702468 325138 702482
rect 325138 702468 325150 702482
rect 325150 702468 325172 702482
rect 325196 702468 325202 702482
rect 325202 702468 325214 702482
rect 325214 702468 325252 702482
rect 325276 702468 325278 702482
rect 325278 702468 325330 702482
rect 325330 702468 325332 702482
rect 325356 702468 325394 702482
rect 325394 702468 325406 702482
rect 325406 702468 325412 702482
rect 325436 702468 325458 702482
rect 325458 702468 325470 702482
rect 325470 702468 325492 702482
rect 325516 702468 325522 702482
rect 325522 702468 325534 702482
rect 325534 702468 325572 702482
rect 325036 702430 325074 702444
rect 325074 702430 325086 702444
rect 325086 702430 325092 702444
rect 325116 702430 325138 702444
rect 325138 702430 325150 702444
rect 325150 702430 325172 702444
rect 325196 702430 325202 702444
rect 325202 702430 325214 702444
rect 325214 702430 325252 702444
rect 325276 702430 325278 702444
rect 325278 702430 325330 702444
rect 325330 702430 325332 702444
rect 325356 702430 325394 702444
rect 325394 702430 325406 702444
rect 325406 702430 325412 702444
rect 325436 702430 325458 702444
rect 325458 702430 325470 702444
rect 325470 702430 325492 702444
rect 325516 702430 325522 702444
rect 325522 702430 325534 702444
rect 325534 702430 325572 702444
rect 325036 702418 325092 702430
rect 325116 702418 325172 702430
rect 325196 702418 325252 702430
rect 325276 702418 325332 702430
rect 325356 702418 325412 702430
rect 325436 702418 325492 702430
rect 325516 702418 325572 702430
rect 325036 702388 325074 702418
rect 325074 702388 325086 702418
rect 325086 702388 325092 702418
rect 325116 702388 325138 702418
rect 325138 702388 325150 702418
rect 325150 702388 325172 702418
rect 325196 702388 325202 702418
rect 325202 702388 325214 702418
rect 325214 702388 325252 702418
rect 325276 702388 325278 702418
rect 325278 702388 325330 702418
rect 325330 702388 325332 702418
rect 325356 702388 325394 702418
rect 325394 702388 325406 702418
rect 325406 702388 325412 702418
rect 325436 702388 325458 702418
rect 325458 702388 325470 702418
rect 325470 702388 325492 702418
rect 325516 702388 325522 702418
rect 325522 702388 325534 702418
rect 325534 702388 325572 702418
rect 325036 702354 325092 702364
rect 325116 702354 325172 702364
rect 325196 702354 325252 702364
rect 325276 702354 325332 702364
rect 325356 702354 325412 702364
rect 325436 702354 325492 702364
rect 325516 702354 325572 702364
rect 325036 702308 325074 702354
rect 325074 702308 325086 702354
rect 325086 702308 325092 702354
rect 325116 702308 325138 702354
rect 325138 702308 325150 702354
rect 325150 702308 325172 702354
rect 325196 702308 325202 702354
rect 325202 702308 325214 702354
rect 325214 702308 325252 702354
rect 325276 702308 325278 702354
rect 325278 702308 325330 702354
rect 325330 702308 325332 702354
rect 325356 702308 325394 702354
rect 325394 702308 325406 702354
rect 325406 702308 325412 702354
rect 325436 702308 325458 702354
rect 325458 702308 325470 702354
rect 325470 702308 325492 702354
rect 325516 702308 325522 702354
rect 325522 702308 325534 702354
rect 325534 702308 325572 702354
rect 362276 702857 362314 702903
rect 362314 702857 362326 702903
rect 362326 702857 362332 702903
rect 362356 702857 362378 702903
rect 362378 702857 362390 702903
rect 362390 702857 362412 702903
rect 362436 702857 362442 702903
rect 362442 702857 362454 702903
rect 362454 702857 362492 702903
rect 362516 702857 362518 702903
rect 362518 702857 362570 702903
rect 362570 702857 362572 702903
rect 362596 702857 362634 702903
rect 362634 702857 362646 702903
rect 362646 702857 362652 702903
rect 362676 702857 362698 702903
rect 362698 702857 362710 702903
rect 362710 702857 362732 702903
rect 362756 702857 362762 702903
rect 362762 702857 362774 702903
rect 362774 702857 362812 702903
rect 362276 702847 362332 702857
rect 362356 702847 362412 702857
rect 362436 702847 362492 702857
rect 362516 702847 362572 702857
rect 362596 702847 362652 702857
rect 362676 702847 362732 702857
rect 362756 702847 362812 702857
rect 362276 702793 362314 702823
rect 362314 702793 362326 702823
rect 362326 702793 362332 702823
rect 362356 702793 362378 702823
rect 362378 702793 362390 702823
rect 362390 702793 362412 702823
rect 362436 702793 362442 702823
rect 362442 702793 362454 702823
rect 362454 702793 362492 702823
rect 362516 702793 362518 702823
rect 362518 702793 362570 702823
rect 362570 702793 362572 702823
rect 362596 702793 362634 702823
rect 362634 702793 362646 702823
rect 362646 702793 362652 702823
rect 362676 702793 362698 702823
rect 362698 702793 362710 702823
rect 362710 702793 362732 702823
rect 362756 702793 362762 702823
rect 362762 702793 362774 702823
rect 362774 702793 362812 702823
rect 362276 702781 362332 702793
rect 362356 702781 362412 702793
rect 362436 702781 362492 702793
rect 362516 702781 362572 702793
rect 362596 702781 362652 702793
rect 362676 702781 362732 702793
rect 362756 702781 362812 702793
rect 362276 702767 362314 702781
rect 362314 702767 362326 702781
rect 362326 702767 362332 702781
rect 362356 702767 362378 702781
rect 362378 702767 362390 702781
rect 362390 702767 362412 702781
rect 362436 702767 362442 702781
rect 362442 702767 362454 702781
rect 362454 702767 362492 702781
rect 362516 702767 362518 702781
rect 362518 702767 362570 702781
rect 362570 702767 362572 702781
rect 362596 702767 362634 702781
rect 362634 702767 362646 702781
rect 362646 702767 362652 702781
rect 362676 702767 362698 702781
rect 362698 702767 362710 702781
rect 362710 702767 362732 702781
rect 362756 702767 362762 702781
rect 362762 702767 362774 702781
rect 362774 702767 362812 702781
rect 362276 702729 362314 702743
rect 362314 702729 362326 702743
rect 362326 702729 362332 702743
rect 362356 702729 362378 702743
rect 362378 702729 362390 702743
rect 362390 702729 362412 702743
rect 362436 702729 362442 702743
rect 362442 702729 362454 702743
rect 362454 702729 362492 702743
rect 362516 702729 362518 702743
rect 362518 702729 362570 702743
rect 362570 702729 362572 702743
rect 362596 702729 362634 702743
rect 362634 702729 362646 702743
rect 362646 702729 362652 702743
rect 362676 702729 362698 702743
rect 362698 702729 362710 702743
rect 362710 702729 362732 702743
rect 362756 702729 362762 702743
rect 362762 702729 362774 702743
rect 362774 702729 362812 702743
rect 362276 702717 362332 702729
rect 362356 702717 362412 702729
rect 362436 702717 362492 702729
rect 362516 702717 362572 702729
rect 362596 702717 362652 702729
rect 362676 702717 362732 702729
rect 362756 702717 362812 702729
rect 362276 702687 362314 702717
rect 362314 702687 362326 702717
rect 362326 702687 362332 702717
rect 362356 702687 362378 702717
rect 362378 702687 362390 702717
rect 362390 702687 362412 702717
rect 362436 702687 362442 702717
rect 362442 702687 362454 702717
rect 362454 702687 362492 702717
rect 362516 702687 362518 702717
rect 362518 702687 362570 702717
rect 362570 702687 362572 702717
rect 362596 702687 362634 702717
rect 362634 702687 362646 702717
rect 362646 702687 362652 702717
rect 362676 702687 362698 702717
rect 362698 702687 362710 702717
rect 362710 702687 362732 702717
rect 362756 702687 362762 702717
rect 362762 702687 362774 702717
rect 362774 702687 362812 702717
rect 362276 702653 362332 702663
rect 362356 702653 362412 702663
rect 362436 702653 362492 702663
rect 362516 702653 362572 702663
rect 362596 702653 362652 702663
rect 362676 702653 362732 702663
rect 362756 702653 362812 702663
rect 362276 702607 362314 702653
rect 362314 702607 362326 702653
rect 362326 702607 362332 702653
rect 362356 702607 362378 702653
rect 362378 702607 362390 702653
rect 362390 702607 362412 702653
rect 362436 702607 362442 702653
rect 362442 702607 362454 702653
rect 362454 702607 362492 702653
rect 362516 702607 362518 702653
rect 362518 702607 362570 702653
rect 362570 702607 362572 702653
rect 362596 702607 362634 702653
rect 362634 702607 362646 702653
rect 362646 702607 362652 702653
rect 362676 702607 362698 702653
rect 362698 702607 362710 702653
rect 362710 702607 362732 702653
rect 362756 702607 362762 702653
rect 362762 702607 362774 702653
rect 362774 702607 362812 702653
rect 361036 702089 361074 702135
rect 361074 702089 361086 702135
rect 361086 702089 361092 702135
rect 361116 702089 361138 702135
rect 361138 702089 361150 702135
rect 361150 702089 361172 702135
rect 361196 702089 361202 702135
rect 361202 702089 361214 702135
rect 361214 702089 361252 702135
rect 361276 702089 361278 702135
rect 361278 702089 361330 702135
rect 361330 702089 361332 702135
rect 361356 702089 361394 702135
rect 361394 702089 361406 702135
rect 361406 702089 361412 702135
rect 361436 702089 361458 702135
rect 361458 702089 361470 702135
rect 361470 702089 361492 702135
rect 361516 702089 361522 702135
rect 361522 702089 361534 702135
rect 361534 702089 361572 702135
rect 361036 702079 361092 702089
rect 361116 702079 361172 702089
rect 361196 702079 361252 702089
rect 361276 702079 361332 702089
rect 361356 702079 361412 702089
rect 361436 702079 361492 702089
rect 361516 702079 361572 702089
rect 361036 702025 361074 702055
rect 361074 702025 361086 702055
rect 361086 702025 361092 702055
rect 361116 702025 361138 702055
rect 361138 702025 361150 702055
rect 361150 702025 361172 702055
rect 361196 702025 361202 702055
rect 361202 702025 361214 702055
rect 361214 702025 361252 702055
rect 361276 702025 361278 702055
rect 361278 702025 361330 702055
rect 361330 702025 361332 702055
rect 361356 702025 361394 702055
rect 361394 702025 361406 702055
rect 361406 702025 361412 702055
rect 361436 702025 361458 702055
rect 361458 702025 361470 702055
rect 361470 702025 361492 702055
rect 361516 702025 361522 702055
rect 361522 702025 361534 702055
rect 361534 702025 361572 702055
rect 361036 702013 361092 702025
rect 361116 702013 361172 702025
rect 361196 702013 361252 702025
rect 361276 702013 361332 702025
rect 361356 702013 361412 702025
rect 361436 702013 361492 702025
rect 361516 702013 361572 702025
rect 361036 701999 361074 702013
rect 361074 701999 361086 702013
rect 361086 701999 361092 702013
rect 361116 701999 361138 702013
rect 361138 701999 361150 702013
rect 361150 701999 361172 702013
rect 361196 701999 361202 702013
rect 361202 701999 361214 702013
rect 361214 701999 361252 702013
rect 361276 701999 361278 702013
rect 361278 701999 361330 702013
rect 361330 701999 361332 702013
rect 361356 701999 361394 702013
rect 361394 701999 361406 702013
rect 361406 701999 361412 702013
rect 361436 701999 361458 702013
rect 361458 701999 361470 702013
rect 361470 701999 361492 702013
rect 361516 701999 361522 702013
rect 361522 701999 361534 702013
rect 361534 701999 361572 702013
rect 361036 701961 361074 701975
rect 361074 701961 361086 701975
rect 361086 701961 361092 701975
rect 361116 701961 361138 701975
rect 361138 701961 361150 701975
rect 361150 701961 361172 701975
rect 361196 701961 361202 701975
rect 361202 701961 361214 701975
rect 361214 701961 361252 701975
rect 361276 701961 361278 701975
rect 361278 701961 361330 701975
rect 361330 701961 361332 701975
rect 361356 701961 361394 701975
rect 361394 701961 361406 701975
rect 361406 701961 361412 701975
rect 361436 701961 361458 701975
rect 361458 701961 361470 701975
rect 361470 701961 361492 701975
rect 361516 701961 361522 701975
rect 361522 701961 361534 701975
rect 361534 701961 361572 701975
rect 361036 701949 361092 701961
rect 361116 701949 361172 701961
rect 361196 701949 361252 701961
rect 361276 701949 361332 701961
rect 361356 701949 361412 701961
rect 361436 701949 361492 701961
rect 361516 701949 361572 701961
rect 361036 701919 361074 701949
rect 361074 701919 361086 701949
rect 361086 701919 361092 701949
rect 361116 701919 361138 701949
rect 361138 701919 361150 701949
rect 361150 701919 361172 701949
rect 361196 701919 361202 701949
rect 361202 701919 361214 701949
rect 361214 701919 361252 701949
rect 361276 701919 361278 701949
rect 361278 701919 361330 701949
rect 361330 701919 361332 701949
rect 361356 701919 361394 701949
rect 361394 701919 361406 701949
rect 361406 701919 361412 701949
rect 361436 701919 361458 701949
rect 361458 701919 361470 701949
rect 361470 701919 361492 701949
rect 361516 701919 361522 701949
rect 361522 701919 361534 701949
rect 361534 701919 361572 701949
rect 361036 701885 361092 701895
rect 361116 701885 361172 701895
rect 361196 701885 361252 701895
rect 361276 701885 361332 701895
rect 361356 701885 361412 701895
rect 361436 701885 361492 701895
rect 361516 701885 361572 701895
rect 361036 701839 361074 701885
rect 361074 701839 361086 701885
rect 361086 701839 361092 701885
rect 361116 701839 361138 701885
rect 361138 701839 361150 701885
rect 361150 701839 361172 701885
rect 361196 701839 361202 701885
rect 361202 701839 361214 701885
rect 361214 701839 361252 701885
rect 361276 701839 361278 701885
rect 361278 701839 361330 701885
rect 361330 701839 361332 701885
rect 361356 701839 361394 701885
rect 361394 701839 361406 701885
rect 361406 701839 361412 701885
rect 361436 701839 361458 701885
rect 361458 701839 361470 701885
rect 361470 701839 361492 701885
rect 361516 701839 361522 701885
rect 361522 701839 361534 701885
rect 361534 701839 361572 701885
rect 434276 702720 434314 702766
rect 434314 702720 434326 702766
rect 434326 702720 434332 702766
rect 434356 702720 434378 702766
rect 434378 702720 434390 702766
rect 434390 702720 434412 702766
rect 434436 702720 434442 702766
rect 434442 702720 434454 702766
rect 434454 702720 434492 702766
rect 434516 702720 434518 702766
rect 434518 702720 434570 702766
rect 434570 702720 434572 702766
rect 434596 702720 434634 702766
rect 434634 702720 434646 702766
rect 434646 702720 434652 702766
rect 434676 702720 434698 702766
rect 434698 702720 434710 702766
rect 434710 702720 434732 702766
rect 434756 702720 434762 702766
rect 434762 702720 434774 702766
rect 434774 702720 434812 702766
rect 434276 702710 434332 702720
rect 434356 702710 434412 702720
rect 434436 702710 434492 702720
rect 434516 702710 434572 702720
rect 434596 702710 434652 702720
rect 434676 702710 434732 702720
rect 434756 702710 434812 702720
rect 434276 702656 434314 702686
rect 434314 702656 434326 702686
rect 434326 702656 434332 702686
rect 434356 702656 434378 702686
rect 434378 702656 434390 702686
rect 434390 702656 434412 702686
rect 434436 702656 434442 702686
rect 434442 702656 434454 702686
rect 434454 702656 434492 702686
rect 434516 702656 434518 702686
rect 434518 702656 434570 702686
rect 434570 702656 434572 702686
rect 434596 702656 434634 702686
rect 434634 702656 434646 702686
rect 434646 702656 434652 702686
rect 434676 702656 434698 702686
rect 434698 702656 434710 702686
rect 434710 702656 434732 702686
rect 434756 702656 434762 702686
rect 434762 702656 434774 702686
rect 434774 702656 434812 702686
rect 434276 702644 434332 702656
rect 434356 702644 434412 702656
rect 434436 702644 434492 702656
rect 434516 702644 434572 702656
rect 434596 702644 434652 702656
rect 434676 702644 434732 702656
rect 434756 702644 434812 702656
rect 434276 702630 434314 702644
rect 434314 702630 434326 702644
rect 434326 702630 434332 702644
rect 434356 702630 434378 702644
rect 434378 702630 434390 702644
rect 434390 702630 434412 702644
rect 434436 702630 434442 702644
rect 434442 702630 434454 702644
rect 434454 702630 434492 702644
rect 434516 702630 434518 702644
rect 434518 702630 434570 702644
rect 434570 702630 434572 702644
rect 434596 702630 434634 702644
rect 434634 702630 434646 702644
rect 434646 702630 434652 702644
rect 434676 702630 434698 702644
rect 434698 702630 434710 702644
rect 434710 702630 434732 702644
rect 434756 702630 434762 702644
rect 434762 702630 434774 702644
rect 434774 702630 434812 702644
rect 434276 702592 434314 702606
rect 434314 702592 434326 702606
rect 434326 702592 434332 702606
rect 434356 702592 434378 702606
rect 434378 702592 434390 702606
rect 434390 702592 434412 702606
rect 434436 702592 434442 702606
rect 434442 702592 434454 702606
rect 434454 702592 434492 702606
rect 434516 702592 434518 702606
rect 434518 702592 434570 702606
rect 434570 702592 434572 702606
rect 434596 702592 434634 702606
rect 434634 702592 434646 702606
rect 434646 702592 434652 702606
rect 434676 702592 434698 702606
rect 434698 702592 434710 702606
rect 434710 702592 434732 702606
rect 434756 702592 434762 702606
rect 434762 702592 434774 702606
rect 434774 702592 434812 702606
rect 434276 702580 434332 702592
rect 434356 702580 434412 702592
rect 434436 702580 434492 702592
rect 434516 702580 434572 702592
rect 434596 702580 434652 702592
rect 434676 702580 434732 702592
rect 434756 702580 434812 702592
rect 434276 702550 434314 702580
rect 434314 702550 434326 702580
rect 434326 702550 434332 702580
rect 434356 702550 434378 702580
rect 434378 702550 434390 702580
rect 434390 702550 434412 702580
rect 434436 702550 434442 702580
rect 434442 702550 434454 702580
rect 434454 702550 434492 702580
rect 434516 702550 434518 702580
rect 434518 702550 434570 702580
rect 434570 702550 434572 702580
rect 434596 702550 434634 702580
rect 434634 702550 434646 702580
rect 434646 702550 434652 702580
rect 434676 702550 434698 702580
rect 434698 702550 434710 702580
rect 434710 702550 434732 702580
rect 434756 702550 434762 702580
rect 434762 702550 434774 702580
rect 434774 702550 434812 702580
rect 434276 702516 434332 702526
rect 434356 702516 434412 702526
rect 434436 702516 434492 702526
rect 434516 702516 434572 702526
rect 434596 702516 434652 702526
rect 434676 702516 434732 702526
rect 434756 702516 434812 702526
rect 434276 702470 434314 702516
rect 434314 702470 434326 702516
rect 434326 702470 434332 702516
rect 434356 702470 434378 702516
rect 434378 702470 434390 702516
rect 434390 702470 434412 702516
rect 434436 702470 434442 702516
rect 434442 702470 434454 702516
rect 434454 702470 434492 702516
rect 434516 702470 434518 702516
rect 434518 702470 434570 702516
rect 434570 702470 434572 702516
rect 434596 702470 434634 702516
rect 434634 702470 434646 702516
rect 434646 702470 434652 702516
rect 434676 702470 434698 702516
rect 434698 702470 434710 702516
rect 434710 702470 434732 702516
rect 434756 702470 434762 702516
rect 434762 702470 434774 702516
rect 434774 702470 434812 702516
rect 433036 701952 433074 701998
rect 433074 701952 433086 701998
rect 433086 701952 433092 701998
rect 433116 701952 433138 701998
rect 433138 701952 433150 701998
rect 433150 701952 433172 701998
rect 433196 701952 433202 701998
rect 433202 701952 433214 701998
rect 433214 701952 433252 701998
rect 433276 701952 433278 701998
rect 433278 701952 433330 701998
rect 433330 701952 433332 701998
rect 433356 701952 433394 701998
rect 433394 701952 433406 701998
rect 433406 701952 433412 701998
rect 433436 701952 433458 701998
rect 433458 701952 433470 701998
rect 433470 701952 433492 701998
rect 433516 701952 433522 701998
rect 433522 701952 433534 701998
rect 433534 701952 433572 701998
rect 433036 701942 433092 701952
rect 433116 701942 433172 701952
rect 433196 701942 433252 701952
rect 433276 701942 433332 701952
rect 433356 701942 433412 701952
rect 433436 701942 433492 701952
rect 433516 701942 433572 701952
rect 433036 701888 433074 701918
rect 433074 701888 433086 701918
rect 433086 701888 433092 701918
rect 433116 701888 433138 701918
rect 433138 701888 433150 701918
rect 433150 701888 433172 701918
rect 433196 701888 433202 701918
rect 433202 701888 433214 701918
rect 433214 701888 433252 701918
rect 433276 701888 433278 701918
rect 433278 701888 433330 701918
rect 433330 701888 433332 701918
rect 433356 701888 433394 701918
rect 433394 701888 433406 701918
rect 433406 701888 433412 701918
rect 433436 701888 433458 701918
rect 433458 701888 433470 701918
rect 433470 701888 433492 701918
rect 433516 701888 433522 701918
rect 433522 701888 433534 701918
rect 433534 701888 433572 701918
rect 433036 701876 433092 701888
rect 433116 701876 433172 701888
rect 433196 701876 433252 701888
rect 433276 701876 433332 701888
rect 433356 701876 433412 701888
rect 433436 701876 433492 701888
rect 433516 701876 433572 701888
rect 433036 701862 433074 701876
rect 433074 701862 433086 701876
rect 433086 701862 433092 701876
rect 433116 701862 433138 701876
rect 433138 701862 433150 701876
rect 433150 701862 433172 701876
rect 433196 701862 433202 701876
rect 433202 701862 433214 701876
rect 433214 701862 433252 701876
rect 433276 701862 433278 701876
rect 433278 701862 433330 701876
rect 433330 701862 433332 701876
rect 433356 701862 433394 701876
rect 433394 701862 433406 701876
rect 433406 701862 433412 701876
rect 433436 701862 433458 701876
rect 433458 701862 433470 701876
rect 433470 701862 433492 701876
rect 433516 701862 433522 701876
rect 433522 701862 433534 701876
rect 433534 701862 433572 701876
rect 433036 701824 433074 701838
rect 433074 701824 433086 701838
rect 433086 701824 433092 701838
rect 433116 701824 433138 701838
rect 433138 701824 433150 701838
rect 433150 701824 433172 701838
rect 433196 701824 433202 701838
rect 433202 701824 433214 701838
rect 433214 701824 433252 701838
rect 433276 701824 433278 701838
rect 433278 701824 433330 701838
rect 433330 701824 433332 701838
rect 433356 701824 433394 701838
rect 433394 701824 433406 701838
rect 433406 701824 433412 701838
rect 433436 701824 433458 701838
rect 433458 701824 433470 701838
rect 433470 701824 433492 701838
rect 433516 701824 433522 701838
rect 433522 701824 433534 701838
rect 433534 701824 433572 701838
rect 433036 701812 433092 701824
rect 433116 701812 433172 701824
rect 433196 701812 433252 701824
rect 433276 701812 433332 701824
rect 433356 701812 433412 701824
rect 433436 701812 433492 701824
rect 433516 701812 433572 701824
rect 433036 701782 433074 701812
rect 433074 701782 433086 701812
rect 433086 701782 433092 701812
rect 433116 701782 433138 701812
rect 433138 701782 433150 701812
rect 433150 701782 433172 701812
rect 433196 701782 433202 701812
rect 433202 701782 433214 701812
rect 433214 701782 433252 701812
rect 433276 701782 433278 701812
rect 433278 701782 433330 701812
rect 433330 701782 433332 701812
rect 433356 701782 433394 701812
rect 433394 701782 433406 701812
rect 433406 701782 433412 701812
rect 433436 701782 433458 701812
rect 433458 701782 433470 701812
rect 433470 701782 433492 701812
rect 433516 701782 433522 701812
rect 433522 701782 433534 701812
rect 433534 701782 433572 701812
rect 433036 701748 433092 701758
rect 433116 701748 433172 701758
rect 433196 701748 433252 701758
rect 433276 701748 433332 701758
rect 433356 701748 433412 701758
rect 433436 701748 433492 701758
rect 433516 701748 433572 701758
rect 433036 701702 433074 701748
rect 433074 701702 433086 701748
rect 433086 701702 433092 701748
rect 433116 701702 433138 701748
rect 433138 701702 433150 701748
rect 433150 701702 433172 701748
rect 433196 701702 433202 701748
rect 433202 701702 433214 701748
rect 433214 701702 433252 701748
rect 433276 701702 433278 701748
rect 433278 701702 433330 701748
rect 433330 701702 433332 701748
rect 433356 701702 433394 701748
rect 433394 701702 433406 701748
rect 433406 701702 433412 701748
rect 433436 701702 433458 701748
rect 433458 701702 433470 701748
rect 433470 701702 433492 701748
rect 433516 701702 433522 701748
rect 433522 701702 433534 701748
rect 433534 701702 433572 701748
rect 506276 702474 506314 702520
rect 506314 702474 506326 702520
rect 506326 702474 506332 702520
rect 506356 702474 506378 702520
rect 506378 702474 506390 702520
rect 506390 702474 506412 702520
rect 506436 702474 506442 702520
rect 506442 702474 506454 702520
rect 506454 702474 506492 702520
rect 506516 702474 506518 702520
rect 506518 702474 506570 702520
rect 506570 702474 506572 702520
rect 506596 702474 506634 702520
rect 506634 702474 506646 702520
rect 506646 702474 506652 702520
rect 506676 702474 506698 702520
rect 506698 702474 506710 702520
rect 506710 702474 506732 702520
rect 506756 702474 506762 702520
rect 506762 702474 506774 702520
rect 506774 702474 506812 702520
rect 506276 702464 506332 702474
rect 506356 702464 506412 702474
rect 506436 702464 506492 702474
rect 506516 702464 506572 702474
rect 506596 702464 506652 702474
rect 506676 702464 506732 702474
rect 506756 702464 506812 702474
rect 506276 702410 506314 702440
rect 506314 702410 506326 702440
rect 506326 702410 506332 702440
rect 506356 702410 506378 702440
rect 506378 702410 506390 702440
rect 506390 702410 506412 702440
rect 506436 702410 506442 702440
rect 506442 702410 506454 702440
rect 506454 702410 506492 702440
rect 506516 702410 506518 702440
rect 506518 702410 506570 702440
rect 506570 702410 506572 702440
rect 506596 702410 506634 702440
rect 506634 702410 506646 702440
rect 506646 702410 506652 702440
rect 506676 702410 506698 702440
rect 506698 702410 506710 702440
rect 506710 702410 506732 702440
rect 506756 702410 506762 702440
rect 506762 702410 506774 702440
rect 506774 702410 506812 702440
rect 506276 702398 506332 702410
rect 506356 702398 506412 702410
rect 506436 702398 506492 702410
rect 506516 702398 506572 702410
rect 506596 702398 506652 702410
rect 506676 702398 506732 702410
rect 506756 702398 506812 702410
rect 506276 702384 506314 702398
rect 506314 702384 506326 702398
rect 506326 702384 506332 702398
rect 506356 702384 506378 702398
rect 506378 702384 506390 702398
rect 506390 702384 506412 702398
rect 506436 702384 506442 702398
rect 506442 702384 506454 702398
rect 506454 702384 506492 702398
rect 506516 702384 506518 702398
rect 506518 702384 506570 702398
rect 506570 702384 506572 702398
rect 506596 702384 506634 702398
rect 506634 702384 506646 702398
rect 506646 702384 506652 702398
rect 506676 702384 506698 702398
rect 506698 702384 506710 702398
rect 506710 702384 506732 702398
rect 506756 702384 506762 702398
rect 506762 702384 506774 702398
rect 506774 702384 506812 702398
rect 506276 702346 506314 702360
rect 506314 702346 506326 702360
rect 506326 702346 506332 702360
rect 506356 702346 506378 702360
rect 506378 702346 506390 702360
rect 506390 702346 506412 702360
rect 506436 702346 506442 702360
rect 506442 702346 506454 702360
rect 506454 702346 506492 702360
rect 506516 702346 506518 702360
rect 506518 702346 506570 702360
rect 506570 702346 506572 702360
rect 506596 702346 506634 702360
rect 506634 702346 506646 702360
rect 506646 702346 506652 702360
rect 506676 702346 506698 702360
rect 506698 702346 506710 702360
rect 506710 702346 506732 702360
rect 506756 702346 506762 702360
rect 506762 702346 506774 702360
rect 506774 702346 506812 702360
rect 506276 702334 506332 702346
rect 506356 702334 506412 702346
rect 506436 702334 506492 702346
rect 506516 702334 506572 702346
rect 506596 702334 506652 702346
rect 506676 702334 506732 702346
rect 506756 702334 506812 702346
rect 506276 702304 506314 702334
rect 506314 702304 506326 702334
rect 506326 702304 506332 702334
rect 506356 702304 506378 702334
rect 506378 702304 506390 702334
rect 506390 702304 506412 702334
rect 506436 702304 506442 702334
rect 506442 702304 506454 702334
rect 506454 702304 506492 702334
rect 506516 702304 506518 702334
rect 506518 702304 506570 702334
rect 506570 702304 506572 702334
rect 506596 702304 506634 702334
rect 506634 702304 506646 702334
rect 506646 702304 506652 702334
rect 506676 702304 506698 702334
rect 506698 702304 506710 702334
rect 506710 702304 506732 702334
rect 506756 702304 506762 702334
rect 506762 702304 506774 702334
rect 506774 702304 506812 702334
rect 506276 702270 506332 702280
rect 506356 702270 506412 702280
rect 506436 702270 506492 702280
rect 506516 702270 506572 702280
rect 506596 702270 506652 702280
rect 506676 702270 506732 702280
rect 506756 702270 506812 702280
rect 506276 702224 506314 702270
rect 506314 702224 506326 702270
rect 506326 702224 506332 702270
rect 506356 702224 506378 702270
rect 506378 702224 506390 702270
rect 506390 702224 506412 702270
rect 506436 702224 506442 702270
rect 506442 702224 506454 702270
rect 506454 702224 506492 702270
rect 506516 702224 506518 702270
rect 506518 702224 506570 702270
rect 506570 702224 506572 702270
rect 506596 702224 506634 702270
rect 506634 702224 506646 702270
rect 506646 702224 506652 702270
rect 506676 702224 506698 702270
rect 506698 702224 506710 702270
rect 506710 702224 506732 702270
rect 506756 702224 506762 702270
rect 506762 702224 506774 702270
rect 506774 702224 506812 702270
rect 505036 701706 505074 701752
rect 505074 701706 505086 701752
rect 505086 701706 505092 701752
rect 505116 701706 505138 701752
rect 505138 701706 505150 701752
rect 505150 701706 505172 701752
rect 505196 701706 505202 701752
rect 505202 701706 505214 701752
rect 505214 701706 505252 701752
rect 505276 701706 505278 701752
rect 505278 701706 505330 701752
rect 505330 701706 505332 701752
rect 505356 701706 505394 701752
rect 505394 701706 505406 701752
rect 505406 701706 505412 701752
rect 505436 701706 505458 701752
rect 505458 701706 505470 701752
rect 505470 701706 505492 701752
rect 505516 701706 505522 701752
rect 505522 701706 505534 701752
rect 505534 701706 505572 701752
rect 505036 701696 505092 701706
rect 505116 701696 505172 701706
rect 505196 701696 505252 701706
rect 505276 701696 505332 701706
rect 505356 701696 505412 701706
rect 505436 701696 505492 701706
rect 505516 701696 505572 701706
rect 505036 701642 505074 701672
rect 505074 701642 505086 701672
rect 505086 701642 505092 701672
rect 505116 701642 505138 701672
rect 505138 701642 505150 701672
rect 505150 701642 505172 701672
rect 505196 701642 505202 701672
rect 505202 701642 505214 701672
rect 505214 701642 505252 701672
rect 505276 701642 505278 701672
rect 505278 701642 505330 701672
rect 505330 701642 505332 701672
rect 505356 701642 505394 701672
rect 505394 701642 505406 701672
rect 505406 701642 505412 701672
rect 505436 701642 505458 701672
rect 505458 701642 505470 701672
rect 505470 701642 505492 701672
rect 505516 701642 505522 701672
rect 505522 701642 505534 701672
rect 505534 701642 505572 701672
rect 505036 701630 505092 701642
rect 505116 701630 505172 701642
rect 505196 701630 505252 701642
rect 505276 701630 505332 701642
rect 505356 701630 505412 701642
rect 505436 701630 505492 701642
rect 505516 701630 505572 701642
rect 505036 701616 505074 701630
rect 505074 701616 505086 701630
rect 505086 701616 505092 701630
rect 505116 701616 505138 701630
rect 505138 701616 505150 701630
rect 505150 701616 505172 701630
rect 505196 701616 505202 701630
rect 505202 701616 505214 701630
rect 505214 701616 505252 701630
rect 505276 701616 505278 701630
rect 505278 701616 505330 701630
rect 505330 701616 505332 701630
rect 505356 701616 505394 701630
rect 505394 701616 505406 701630
rect 505406 701616 505412 701630
rect 505436 701616 505458 701630
rect 505458 701616 505470 701630
rect 505470 701616 505492 701630
rect 505516 701616 505522 701630
rect 505522 701616 505534 701630
rect 505534 701616 505572 701630
rect 505036 701578 505074 701592
rect 505074 701578 505086 701592
rect 505086 701578 505092 701592
rect 505116 701578 505138 701592
rect 505138 701578 505150 701592
rect 505150 701578 505172 701592
rect 505196 701578 505202 701592
rect 505202 701578 505214 701592
rect 505214 701578 505252 701592
rect 505276 701578 505278 701592
rect 505278 701578 505330 701592
rect 505330 701578 505332 701592
rect 505356 701578 505394 701592
rect 505394 701578 505406 701592
rect 505406 701578 505412 701592
rect 505436 701578 505458 701592
rect 505458 701578 505470 701592
rect 505470 701578 505492 701592
rect 505516 701578 505522 701592
rect 505522 701578 505534 701592
rect 505534 701578 505572 701592
rect 505036 701566 505092 701578
rect 505116 701566 505172 701578
rect 505196 701566 505252 701578
rect 505276 701566 505332 701578
rect 505356 701566 505412 701578
rect 505436 701566 505492 701578
rect 505516 701566 505572 701578
rect 505036 701536 505074 701566
rect 505074 701536 505086 701566
rect 505086 701536 505092 701566
rect 505116 701536 505138 701566
rect 505138 701536 505150 701566
rect 505150 701536 505172 701566
rect 505196 701536 505202 701566
rect 505202 701536 505214 701566
rect 505214 701536 505252 701566
rect 505276 701536 505278 701566
rect 505278 701536 505330 701566
rect 505330 701536 505332 701566
rect 505356 701536 505394 701566
rect 505394 701536 505406 701566
rect 505406 701536 505412 701566
rect 505436 701536 505458 701566
rect 505458 701536 505470 701566
rect 505470 701536 505492 701566
rect 505516 701536 505522 701566
rect 505522 701536 505534 701566
rect 505534 701536 505572 701566
rect 505036 701502 505092 701512
rect 505116 701502 505172 701512
rect 505196 701502 505252 701512
rect 505276 701502 505332 701512
rect 505356 701502 505412 701512
rect 505436 701502 505492 701512
rect 505516 701502 505572 701512
rect 505036 701456 505074 701502
rect 505074 701456 505086 701502
rect 505086 701456 505092 701502
rect 505116 701456 505138 701502
rect 505138 701456 505150 701502
rect 505150 701456 505172 701502
rect 505196 701456 505202 701502
rect 505202 701456 505214 701502
rect 505214 701456 505252 701502
rect 505276 701456 505278 701502
rect 505278 701456 505330 701502
rect 505330 701456 505332 701502
rect 505356 701456 505394 701502
rect 505394 701456 505406 701502
rect 505406 701456 505412 701502
rect 505436 701456 505458 701502
rect 505458 701456 505470 701502
rect 505470 701456 505492 701502
rect 505516 701456 505522 701502
rect 505522 701456 505534 701502
rect 505534 701456 505572 701502
rect 478510 700714 478566 700770
rect 413650 700578 413706 700634
rect 348790 700442 348846 700498
rect 283838 700306 283894 700362
rect 547970 700714 548026 700770
rect 547878 700578 547934 700634
rect 547418 700442 547474 700498
rect 547326 700306 547382 700362
rect 543462 699762 543518 699818
rect 505036 554552 505074 554598
rect 505074 554552 505086 554598
rect 505086 554552 505092 554598
rect 505116 554552 505138 554598
rect 505138 554552 505150 554598
rect 505150 554552 505172 554598
rect 505196 554552 505202 554598
rect 505202 554552 505214 554598
rect 505214 554552 505252 554598
rect 505276 554552 505278 554598
rect 505278 554552 505330 554598
rect 505330 554552 505332 554598
rect 505356 554552 505394 554598
rect 505394 554552 505406 554598
rect 505406 554552 505412 554598
rect 505436 554552 505458 554598
rect 505458 554552 505470 554598
rect 505470 554552 505492 554598
rect 505516 554552 505522 554598
rect 505522 554552 505534 554598
rect 505534 554552 505572 554598
rect 505036 554542 505092 554552
rect 505116 554542 505172 554552
rect 505196 554542 505252 554552
rect 505276 554542 505332 554552
rect 505356 554542 505412 554552
rect 505436 554542 505492 554552
rect 505516 554542 505572 554552
rect 505036 554488 505074 554518
rect 505074 554488 505086 554518
rect 505086 554488 505092 554518
rect 505116 554488 505138 554518
rect 505138 554488 505150 554518
rect 505150 554488 505172 554518
rect 505196 554488 505202 554518
rect 505202 554488 505214 554518
rect 505214 554488 505252 554518
rect 505276 554488 505278 554518
rect 505278 554488 505330 554518
rect 505330 554488 505332 554518
rect 505356 554488 505394 554518
rect 505394 554488 505406 554518
rect 505406 554488 505412 554518
rect 505436 554488 505458 554518
rect 505458 554488 505470 554518
rect 505470 554488 505492 554518
rect 505516 554488 505522 554518
rect 505522 554488 505534 554518
rect 505534 554488 505572 554518
rect 505036 554476 505092 554488
rect 505116 554476 505172 554488
rect 505196 554476 505252 554488
rect 505276 554476 505332 554488
rect 505356 554476 505412 554488
rect 505436 554476 505492 554488
rect 505516 554476 505572 554488
rect 505036 554462 505074 554476
rect 505074 554462 505086 554476
rect 505086 554462 505092 554476
rect 505116 554462 505138 554476
rect 505138 554462 505150 554476
rect 505150 554462 505172 554476
rect 505196 554462 505202 554476
rect 505202 554462 505214 554476
rect 505214 554462 505252 554476
rect 505276 554462 505278 554476
rect 505278 554462 505330 554476
rect 505330 554462 505332 554476
rect 505356 554462 505394 554476
rect 505394 554462 505406 554476
rect 505406 554462 505412 554476
rect 505436 554462 505458 554476
rect 505458 554462 505470 554476
rect 505470 554462 505492 554476
rect 505516 554462 505522 554476
rect 505522 554462 505534 554476
rect 505534 554462 505572 554476
rect 505036 554424 505074 554438
rect 505074 554424 505086 554438
rect 505086 554424 505092 554438
rect 505116 554424 505138 554438
rect 505138 554424 505150 554438
rect 505150 554424 505172 554438
rect 505196 554424 505202 554438
rect 505202 554424 505214 554438
rect 505214 554424 505252 554438
rect 505276 554424 505278 554438
rect 505278 554424 505330 554438
rect 505330 554424 505332 554438
rect 505356 554424 505394 554438
rect 505394 554424 505406 554438
rect 505406 554424 505412 554438
rect 505436 554424 505458 554438
rect 505458 554424 505470 554438
rect 505470 554424 505492 554438
rect 505516 554424 505522 554438
rect 505522 554424 505534 554438
rect 505534 554424 505572 554438
rect 505036 554412 505092 554424
rect 505116 554412 505172 554424
rect 505196 554412 505252 554424
rect 505276 554412 505332 554424
rect 505356 554412 505412 554424
rect 505436 554412 505492 554424
rect 505516 554412 505572 554424
rect 505036 554382 505074 554412
rect 505074 554382 505086 554412
rect 505086 554382 505092 554412
rect 505116 554382 505138 554412
rect 505138 554382 505150 554412
rect 505150 554382 505172 554412
rect 505196 554382 505202 554412
rect 505202 554382 505214 554412
rect 505214 554382 505252 554412
rect 505276 554382 505278 554412
rect 505278 554382 505330 554412
rect 505330 554382 505332 554412
rect 505356 554382 505394 554412
rect 505394 554382 505406 554412
rect 505406 554382 505412 554412
rect 505436 554382 505458 554412
rect 505458 554382 505470 554412
rect 505470 554382 505492 554412
rect 505516 554382 505522 554412
rect 505522 554382 505534 554412
rect 505534 554382 505572 554412
rect 505036 554348 505092 554358
rect 505116 554348 505172 554358
rect 505196 554348 505252 554358
rect 505276 554348 505332 554358
rect 505356 554348 505412 554358
rect 505436 554348 505492 554358
rect 505516 554348 505572 554358
rect 505036 554302 505074 554348
rect 505074 554302 505086 554348
rect 505086 554302 505092 554348
rect 505116 554302 505138 554348
rect 505138 554302 505150 554348
rect 505150 554302 505172 554348
rect 505196 554302 505202 554348
rect 505202 554302 505214 554348
rect 505214 554302 505252 554348
rect 505276 554302 505278 554348
rect 505278 554302 505330 554348
rect 505330 554302 505332 554348
rect 505356 554302 505394 554348
rect 505394 554302 505406 554348
rect 505406 554302 505412 554348
rect 505436 554302 505458 554348
rect 505458 554302 505470 554348
rect 505470 554302 505492 554348
rect 505516 554302 505522 554348
rect 505522 554302 505534 554348
rect 505534 554302 505572 554348
rect 506276 553757 506314 553803
rect 506314 553757 506326 553803
rect 506326 553757 506332 553803
rect 506356 553757 506378 553803
rect 506378 553757 506390 553803
rect 506390 553757 506412 553803
rect 506436 553757 506442 553803
rect 506442 553757 506454 553803
rect 506454 553757 506492 553803
rect 506516 553757 506518 553803
rect 506518 553757 506570 553803
rect 506570 553757 506572 553803
rect 506596 553757 506634 553803
rect 506634 553757 506646 553803
rect 506646 553757 506652 553803
rect 506676 553757 506698 553803
rect 506698 553757 506710 553803
rect 506710 553757 506732 553803
rect 506756 553757 506762 553803
rect 506762 553757 506774 553803
rect 506774 553757 506812 553803
rect 506276 553747 506332 553757
rect 506356 553747 506412 553757
rect 506436 553747 506492 553757
rect 506516 553747 506572 553757
rect 506596 553747 506652 553757
rect 506676 553747 506732 553757
rect 506756 553747 506812 553757
rect 506276 553693 506314 553723
rect 506314 553693 506326 553723
rect 506326 553693 506332 553723
rect 506356 553693 506378 553723
rect 506378 553693 506390 553723
rect 506390 553693 506412 553723
rect 506436 553693 506442 553723
rect 506442 553693 506454 553723
rect 506454 553693 506492 553723
rect 506516 553693 506518 553723
rect 506518 553693 506570 553723
rect 506570 553693 506572 553723
rect 506596 553693 506634 553723
rect 506634 553693 506646 553723
rect 506646 553693 506652 553723
rect 506676 553693 506698 553723
rect 506698 553693 506710 553723
rect 506710 553693 506732 553723
rect 506756 553693 506762 553723
rect 506762 553693 506774 553723
rect 506774 553693 506812 553723
rect 506276 553681 506332 553693
rect 506356 553681 506412 553693
rect 506436 553681 506492 553693
rect 506516 553681 506572 553693
rect 506596 553681 506652 553693
rect 506676 553681 506732 553693
rect 506756 553681 506812 553693
rect 506276 553667 506314 553681
rect 506314 553667 506326 553681
rect 506326 553667 506332 553681
rect 506356 553667 506378 553681
rect 506378 553667 506390 553681
rect 506390 553667 506412 553681
rect 506436 553667 506442 553681
rect 506442 553667 506454 553681
rect 506454 553667 506492 553681
rect 506516 553667 506518 553681
rect 506518 553667 506570 553681
rect 506570 553667 506572 553681
rect 506596 553667 506634 553681
rect 506634 553667 506646 553681
rect 506646 553667 506652 553681
rect 506676 553667 506698 553681
rect 506698 553667 506710 553681
rect 506710 553667 506732 553681
rect 506756 553667 506762 553681
rect 506762 553667 506774 553681
rect 506774 553667 506812 553681
rect 506276 553629 506314 553643
rect 506314 553629 506326 553643
rect 506326 553629 506332 553643
rect 506356 553629 506378 553643
rect 506378 553629 506390 553643
rect 506390 553629 506412 553643
rect 506436 553629 506442 553643
rect 506442 553629 506454 553643
rect 506454 553629 506492 553643
rect 506516 553629 506518 553643
rect 506518 553629 506570 553643
rect 506570 553629 506572 553643
rect 506596 553629 506634 553643
rect 506634 553629 506646 553643
rect 506646 553629 506652 553643
rect 506676 553629 506698 553643
rect 506698 553629 506710 553643
rect 506710 553629 506732 553643
rect 506756 553629 506762 553643
rect 506762 553629 506774 553643
rect 506774 553629 506812 553643
rect 506276 553617 506332 553629
rect 506356 553617 506412 553629
rect 506436 553617 506492 553629
rect 506516 553617 506572 553629
rect 506596 553617 506652 553629
rect 506676 553617 506732 553629
rect 506756 553617 506812 553629
rect 506276 553587 506314 553617
rect 506314 553587 506326 553617
rect 506326 553587 506332 553617
rect 506356 553587 506378 553617
rect 506378 553587 506390 553617
rect 506390 553587 506412 553617
rect 506436 553587 506442 553617
rect 506442 553587 506454 553617
rect 506454 553587 506492 553617
rect 506516 553587 506518 553617
rect 506518 553587 506570 553617
rect 506570 553587 506572 553617
rect 506596 553587 506634 553617
rect 506634 553587 506646 553617
rect 506646 553587 506652 553617
rect 506676 553587 506698 553617
rect 506698 553587 506710 553617
rect 506710 553587 506732 553617
rect 506756 553587 506762 553617
rect 506762 553587 506774 553617
rect 506774 553587 506812 553617
rect 506276 553553 506332 553563
rect 506356 553553 506412 553563
rect 506436 553553 506492 553563
rect 506516 553553 506572 553563
rect 506596 553553 506652 553563
rect 506676 553553 506732 553563
rect 506756 553553 506812 553563
rect 506276 553507 506314 553553
rect 506314 553507 506326 553553
rect 506326 553507 506332 553553
rect 506356 553507 506378 553553
rect 506378 553507 506390 553553
rect 506390 553507 506412 553553
rect 506436 553507 506442 553553
rect 506442 553507 506454 553553
rect 506454 553507 506492 553553
rect 506516 553507 506518 553553
rect 506518 553507 506570 553553
rect 506570 553507 506572 553553
rect 506596 553507 506634 553553
rect 506634 553507 506646 553553
rect 506646 553507 506652 553553
rect 506676 553507 506698 553553
rect 506698 553507 506710 553553
rect 506710 553507 506732 553553
rect 506756 553507 506762 553553
rect 506762 553507 506774 553553
rect 506774 553507 506812 553553
rect 470276 451435 470314 451481
rect 470314 451435 470326 451481
rect 470326 451435 470332 451481
rect 470356 451435 470378 451481
rect 470378 451435 470390 451481
rect 470390 451435 470412 451481
rect 470436 451435 470442 451481
rect 470442 451435 470454 451481
rect 470454 451435 470492 451481
rect 470516 451435 470518 451481
rect 470518 451435 470570 451481
rect 470570 451435 470572 451481
rect 470596 451435 470634 451481
rect 470634 451435 470646 451481
rect 470646 451435 470652 451481
rect 470676 451435 470698 451481
rect 470698 451435 470710 451481
rect 470710 451435 470732 451481
rect 470756 451435 470762 451481
rect 470762 451435 470774 451481
rect 470774 451435 470812 451481
rect 470276 451425 470332 451435
rect 470356 451425 470412 451435
rect 470436 451425 470492 451435
rect 470516 451425 470572 451435
rect 470596 451425 470652 451435
rect 470676 451425 470732 451435
rect 470756 451425 470812 451435
rect 470276 451371 470314 451401
rect 470314 451371 470326 451401
rect 470326 451371 470332 451401
rect 470356 451371 470378 451401
rect 470378 451371 470390 451401
rect 470390 451371 470412 451401
rect 470436 451371 470442 451401
rect 470442 451371 470454 451401
rect 470454 451371 470492 451401
rect 470516 451371 470518 451401
rect 470518 451371 470570 451401
rect 470570 451371 470572 451401
rect 470596 451371 470634 451401
rect 470634 451371 470646 451401
rect 470646 451371 470652 451401
rect 470676 451371 470698 451401
rect 470698 451371 470710 451401
rect 470710 451371 470732 451401
rect 470756 451371 470762 451401
rect 470762 451371 470774 451401
rect 470774 451371 470812 451401
rect 470276 451359 470332 451371
rect 470356 451359 470412 451371
rect 470436 451359 470492 451371
rect 470516 451359 470572 451371
rect 470596 451359 470652 451371
rect 470676 451359 470732 451371
rect 470756 451359 470812 451371
rect 470276 451345 470314 451359
rect 470314 451345 470326 451359
rect 470326 451345 470332 451359
rect 470356 451345 470378 451359
rect 470378 451345 470390 451359
rect 470390 451345 470412 451359
rect 470436 451345 470442 451359
rect 470442 451345 470454 451359
rect 470454 451345 470492 451359
rect 470516 451345 470518 451359
rect 470518 451345 470570 451359
rect 470570 451345 470572 451359
rect 470596 451345 470634 451359
rect 470634 451345 470646 451359
rect 470646 451345 470652 451359
rect 470676 451345 470698 451359
rect 470698 451345 470710 451359
rect 470710 451345 470732 451359
rect 470756 451345 470762 451359
rect 470762 451345 470774 451359
rect 470774 451345 470812 451359
rect 470276 451307 470314 451321
rect 470314 451307 470326 451321
rect 470326 451307 470332 451321
rect 470356 451307 470378 451321
rect 470378 451307 470390 451321
rect 470390 451307 470412 451321
rect 470436 451307 470442 451321
rect 470442 451307 470454 451321
rect 470454 451307 470492 451321
rect 470516 451307 470518 451321
rect 470518 451307 470570 451321
rect 470570 451307 470572 451321
rect 470596 451307 470634 451321
rect 470634 451307 470646 451321
rect 470646 451307 470652 451321
rect 470676 451307 470698 451321
rect 470698 451307 470710 451321
rect 470710 451307 470732 451321
rect 470756 451307 470762 451321
rect 470762 451307 470774 451321
rect 470774 451307 470812 451321
rect 470276 451295 470332 451307
rect 470356 451295 470412 451307
rect 470436 451295 470492 451307
rect 470516 451295 470572 451307
rect 470596 451295 470652 451307
rect 470676 451295 470732 451307
rect 470756 451295 470812 451307
rect 470276 451265 470314 451295
rect 470314 451265 470326 451295
rect 470326 451265 470332 451295
rect 470356 451265 470378 451295
rect 470378 451265 470390 451295
rect 470390 451265 470412 451295
rect 470436 451265 470442 451295
rect 470442 451265 470454 451295
rect 470454 451265 470492 451295
rect 470516 451265 470518 451295
rect 470518 451265 470570 451295
rect 470570 451265 470572 451295
rect 470596 451265 470634 451295
rect 470634 451265 470646 451295
rect 470646 451265 470652 451295
rect 470676 451265 470698 451295
rect 470698 451265 470710 451295
rect 470710 451265 470732 451295
rect 470756 451265 470762 451295
rect 470762 451265 470774 451295
rect 470774 451265 470812 451295
rect 470276 451231 470332 451241
rect 470356 451231 470412 451241
rect 470436 451231 470492 451241
rect 470516 451231 470572 451241
rect 470596 451231 470652 451241
rect 470676 451231 470732 451241
rect 470756 451231 470812 451241
rect 470276 451185 470314 451231
rect 470314 451185 470326 451231
rect 470326 451185 470332 451231
rect 470356 451185 470378 451231
rect 470378 451185 470390 451231
rect 470390 451185 470412 451231
rect 470436 451185 470442 451231
rect 470442 451185 470454 451231
rect 470454 451185 470492 451231
rect 470516 451185 470518 451231
rect 470518 451185 470570 451231
rect 470570 451185 470572 451231
rect 470596 451185 470634 451231
rect 470634 451185 470646 451231
rect 470646 451185 470652 451231
rect 470676 451185 470698 451231
rect 470698 451185 470710 451231
rect 470710 451185 470732 451231
rect 470756 451185 470762 451231
rect 470762 451185 470774 451231
rect 470774 451185 470812 451231
rect 469036 450349 469074 450395
rect 469074 450349 469086 450395
rect 469086 450349 469092 450395
rect 469116 450349 469138 450395
rect 469138 450349 469150 450395
rect 469150 450349 469172 450395
rect 469196 450349 469202 450395
rect 469202 450349 469214 450395
rect 469214 450349 469252 450395
rect 469276 450349 469278 450395
rect 469278 450349 469330 450395
rect 469330 450349 469332 450395
rect 469356 450349 469394 450395
rect 469394 450349 469406 450395
rect 469406 450349 469412 450395
rect 469436 450349 469458 450395
rect 469458 450349 469470 450395
rect 469470 450349 469492 450395
rect 469516 450349 469522 450395
rect 469522 450349 469534 450395
rect 469534 450349 469572 450395
rect 469036 450339 469092 450349
rect 469116 450339 469172 450349
rect 469196 450339 469252 450349
rect 469276 450339 469332 450349
rect 469356 450339 469412 450349
rect 469436 450339 469492 450349
rect 469516 450339 469572 450349
rect 469036 450285 469074 450315
rect 469074 450285 469086 450315
rect 469086 450285 469092 450315
rect 469116 450285 469138 450315
rect 469138 450285 469150 450315
rect 469150 450285 469172 450315
rect 469196 450285 469202 450315
rect 469202 450285 469214 450315
rect 469214 450285 469252 450315
rect 469276 450285 469278 450315
rect 469278 450285 469330 450315
rect 469330 450285 469332 450315
rect 469356 450285 469394 450315
rect 469394 450285 469406 450315
rect 469406 450285 469412 450315
rect 469436 450285 469458 450315
rect 469458 450285 469470 450315
rect 469470 450285 469492 450315
rect 469516 450285 469522 450315
rect 469522 450285 469534 450315
rect 469534 450285 469572 450315
rect 469036 450273 469092 450285
rect 469116 450273 469172 450285
rect 469196 450273 469252 450285
rect 469276 450273 469332 450285
rect 469356 450273 469412 450285
rect 469436 450273 469492 450285
rect 469516 450273 469572 450285
rect 469036 450259 469074 450273
rect 469074 450259 469086 450273
rect 469086 450259 469092 450273
rect 469116 450259 469138 450273
rect 469138 450259 469150 450273
rect 469150 450259 469172 450273
rect 469196 450259 469202 450273
rect 469202 450259 469214 450273
rect 469214 450259 469252 450273
rect 469276 450259 469278 450273
rect 469278 450259 469330 450273
rect 469330 450259 469332 450273
rect 469356 450259 469394 450273
rect 469394 450259 469406 450273
rect 469406 450259 469412 450273
rect 469436 450259 469458 450273
rect 469458 450259 469470 450273
rect 469470 450259 469492 450273
rect 469516 450259 469522 450273
rect 469522 450259 469534 450273
rect 469534 450259 469572 450273
rect 469036 450221 469074 450235
rect 469074 450221 469086 450235
rect 469086 450221 469092 450235
rect 469116 450221 469138 450235
rect 469138 450221 469150 450235
rect 469150 450221 469172 450235
rect 469196 450221 469202 450235
rect 469202 450221 469214 450235
rect 469214 450221 469252 450235
rect 469276 450221 469278 450235
rect 469278 450221 469330 450235
rect 469330 450221 469332 450235
rect 469356 450221 469394 450235
rect 469394 450221 469406 450235
rect 469406 450221 469412 450235
rect 469436 450221 469458 450235
rect 469458 450221 469470 450235
rect 469470 450221 469492 450235
rect 469516 450221 469522 450235
rect 469522 450221 469534 450235
rect 469534 450221 469572 450235
rect 469036 450209 469092 450221
rect 469116 450209 469172 450221
rect 469196 450209 469252 450221
rect 469276 450209 469332 450221
rect 469356 450209 469412 450221
rect 469436 450209 469492 450221
rect 469516 450209 469572 450221
rect 469036 450179 469074 450209
rect 469074 450179 469086 450209
rect 469086 450179 469092 450209
rect 469116 450179 469138 450209
rect 469138 450179 469150 450209
rect 469150 450179 469172 450209
rect 469196 450179 469202 450209
rect 469202 450179 469214 450209
rect 469214 450179 469252 450209
rect 469276 450179 469278 450209
rect 469278 450179 469330 450209
rect 469330 450179 469332 450209
rect 469356 450179 469394 450209
rect 469394 450179 469406 450209
rect 469406 450179 469412 450209
rect 469436 450179 469458 450209
rect 469458 450179 469470 450209
rect 469470 450179 469492 450209
rect 469516 450179 469522 450209
rect 469522 450179 469534 450209
rect 469534 450179 469572 450209
rect 469036 450145 469092 450155
rect 469116 450145 469172 450155
rect 469196 450145 469252 450155
rect 469276 450145 469332 450155
rect 469356 450145 469412 450155
rect 469436 450145 469492 450155
rect 469516 450145 469572 450155
rect 469036 450099 469074 450145
rect 469074 450099 469086 450145
rect 469086 450099 469092 450145
rect 469116 450099 469138 450145
rect 469138 450099 469150 450145
rect 469150 450099 469172 450145
rect 469196 450099 469202 450145
rect 469202 450099 469214 450145
rect 469214 450099 469252 450145
rect 469276 450099 469278 450145
rect 469278 450099 469330 450145
rect 469330 450099 469332 450145
rect 469356 450099 469394 450145
rect 469394 450099 469406 450145
rect 469406 450099 469412 450145
rect 469436 450099 469458 450145
rect 469458 450099 469470 450145
rect 469470 450099 469492 450145
rect 469516 450099 469522 450145
rect 469522 450099 469534 450145
rect 469534 450099 469572 450145
rect 470276 449264 470314 449310
rect 470314 449264 470326 449310
rect 470326 449264 470332 449310
rect 470356 449264 470378 449310
rect 470378 449264 470390 449310
rect 470390 449264 470412 449310
rect 470436 449264 470442 449310
rect 470442 449264 470454 449310
rect 470454 449264 470492 449310
rect 470516 449264 470518 449310
rect 470518 449264 470570 449310
rect 470570 449264 470572 449310
rect 470596 449264 470634 449310
rect 470634 449264 470646 449310
rect 470646 449264 470652 449310
rect 470676 449264 470698 449310
rect 470698 449264 470710 449310
rect 470710 449264 470732 449310
rect 470756 449264 470762 449310
rect 470762 449264 470774 449310
rect 470774 449264 470812 449310
rect 470276 449254 470332 449264
rect 470356 449254 470412 449264
rect 470436 449254 470492 449264
rect 470516 449254 470572 449264
rect 470596 449254 470652 449264
rect 470676 449254 470732 449264
rect 470756 449254 470812 449264
rect 470276 449200 470314 449230
rect 470314 449200 470326 449230
rect 470326 449200 470332 449230
rect 470356 449200 470378 449230
rect 470378 449200 470390 449230
rect 470390 449200 470412 449230
rect 470436 449200 470442 449230
rect 470442 449200 470454 449230
rect 470454 449200 470492 449230
rect 470516 449200 470518 449230
rect 470518 449200 470570 449230
rect 470570 449200 470572 449230
rect 470596 449200 470634 449230
rect 470634 449200 470646 449230
rect 470646 449200 470652 449230
rect 470676 449200 470698 449230
rect 470698 449200 470710 449230
rect 470710 449200 470732 449230
rect 470756 449200 470762 449230
rect 470762 449200 470774 449230
rect 470774 449200 470812 449230
rect 470276 449188 470332 449200
rect 470356 449188 470412 449200
rect 470436 449188 470492 449200
rect 470516 449188 470572 449200
rect 470596 449188 470652 449200
rect 470676 449188 470732 449200
rect 470756 449188 470812 449200
rect 470276 449174 470314 449188
rect 470314 449174 470326 449188
rect 470326 449174 470332 449188
rect 470356 449174 470378 449188
rect 470378 449174 470390 449188
rect 470390 449174 470412 449188
rect 470436 449174 470442 449188
rect 470442 449174 470454 449188
rect 470454 449174 470492 449188
rect 470516 449174 470518 449188
rect 470518 449174 470570 449188
rect 470570 449174 470572 449188
rect 470596 449174 470634 449188
rect 470634 449174 470646 449188
rect 470646 449174 470652 449188
rect 470676 449174 470698 449188
rect 470698 449174 470710 449188
rect 470710 449174 470732 449188
rect 470756 449174 470762 449188
rect 470762 449174 470774 449188
rect 470774 449174 470812 449188
rect 470276 449136 470314 449150
rect 470314 449136 470326 449150
rect 470326 449136 470332 449150
rect 470356 449136 470378 449150
rect 470378 449136 470390 449150
rect 470390 449136 470412 449150
rect 470436 449136 470442 449150
rect 470442 449136 470454 449150
rect 470454 449136 470492 449150
rect 470516 449136 470518 449150
rect 470518 449136 470570 449150
rect 470570 449136 470572 449150
rect 470596 449136 470634 449150
rect 470634 449136 470646 449150
rect 470646 449136 470652 449150
rect 470676 449136 470698 449150
rect 470698 449136 470710 449150
rect 470710 449136 470732 449150
rect 470756 449136 470762 449150
rect 470762 449136 470774 449150
rect 470774 449136 470812 449150
rect 470276 449124 470332 449136
rect 470356 449124 470412 449136
rect 470436 449124 470492 449136
rect 470516 449124 470572 449136
rect 470596 449124 470652 449136
rect 470676 449124 470732 449136
rect 470756 449124 470812 449136
rect 470276 449094 470314 449124
rect 470314 449094 470326 449124
rect 470326 449094 470332 449124
rect 470356 449094 470378 449124
rect 470378 449094 470390 449124
rect 470390 449094 470412 449124
rect 470436 449094 470442 449124
rect 470442 449094 470454 449124
rect 470454 449094 470492 449124
rect 470516 449094 470518 449124
rect 470518 449094 470570 449124
rect 470570 449094 470572 449124
rect 470596 449094 470634 449124
rect 470634 449094 470646 449124
rect 470646 449094 470652 449124
rect 470676 449094 470698 449124
rect 470698 449094 470710 449124
rect 470710 449094 470732 449124
rect 470756 449094 470762 449124
rect 470762 449094 470774 449124
rect 470774 449094 470812 449124
rect 470276 449060 470332 449070
rect 470356 449060 470412 449070
rect 470436 449060 470492 449070
rect 470516 449060 470572 449070
rect 470596 449060 470652 449070
rect 470676 449060 470732 449070
rect 470756 449060 470812 449070
rect 470276 449014 470314 449060
rect 470314 449014 470326 449060
rect 470326 449014 470332 449060
rect 470356 449014 470378 449060
rect 470378 449014 470390 449060
rect 470390 449014 470412 449060
rect 470436 449014 470442 449060
rect 470442 449014 470454 449060
rect 470454 449014 470492 449060
rect 470516 449014 470518 449060
rect 470518 449014 470570 449060
rect 470570 449014 470572 449060
rect 470596 449014 470634 449060
rect 470634 449014 470646 449060
rect 470646 449014 470652 449060
rect 470676 449014 470698 449060
rect 470698 449014 470710 449060
rect 470710 449014 470732 449060
rect 470756 449014 470762 449060
rect 470762 449014 470774 449060
rect 470774 449014 470812 449060
rect 477843 450202 477899 450258
rect 481160 450202 481216 450258
rect 487793 450202 487849 450258
rect 474094 449658 474150 449714
rect 470276 433036 470314 433082
rect 470314 433036 470326 433082
rect 470326 433036 470332 433082
rect 470356 433036 470378 433082
rect 470378 433036 470390 433082
rect 470390 433036 470412 433082
rect 470436 433036 470442 433082
rect 470442 433036 470454 433082
rect 470454 433036 470492 433082
rect 470516 433036 470518 433082
rect 470518 433036 470570 433082
rect 470570 433036 470572 433082
rect 470596 433036 470634 433082
rect 470634 433036 470646 433082
rect 470646 433036 470652 433082
rect 470676 433036 470698 433082
rect 470698 433036 470710 433082
rect 470710 433036 470732 433082
rect 470756 433036 470762 433082
rect 470762 433036 470774 433082
rect 470774 433036 470812 433082
rect 470276 433026 470332 433036
rect 470356 433026 470412 433036
rect 470436 433026 470492 433036
rect 470516 433026 470572 433036
rect 470596 433026 470652 433036
rect 470676 433026 470732 433036
rect 470756 433026 470812 433036
rect 470276 432972 470314 433002
rect 470314 432972 470326 433002
rect 470326 432972 470332 433002
rect 470356 432972 470378 433002
rect 470378 432972 470390 433002
rect 470390 432972 470412 433002
rect 470436 432972 470442 433002
rect 470442 432972 470454 433002
rect 470454 432972 470492 433002
rect 470516 432972 470518 433002
rect 470518 432972 470570 433002
rect 470570 432972 470572 433002
rect 470596 432972 470634 433002
rect 470634 432972 470646 433002
rect 470646 432972 470652 433002
rect 470676 432972 470698 433002
rect 470698 432972 470710 433002
rect 470710 432972 470732 433002
rect 470756 432972 470762 433002
rect 470762 432972 470774 433002
rect 470774 432972 470812 433002
rect 470276 432960 470332 432972
rect 470356 432960 470412 432972
rect 470436 432960 470492 432972
rect 470516 432960 470572 432972
rect 470596 432960 470652 432972
rect 470676 432960 470732 432972
rect 470756 432960 470812 432972
rect 470276 432946 470314 432960
rect 470314 432946 470326 432960
rect 470326 432946 470332 432960
rect 470356 432946 470378 432960
rect 470378 432946 470390 432960
rect 470390 432946 470412 432960
rect 470436 432946 470442 432960
rect 470442 432946 470454 432960
rect 470454 432946 470492 432960
rect 470516 432946 470518 432960
rect 470518 432946 470570 432960
rect 470570 432946 470572 432960
rect 470596 432946 470634 432960
rect 470634 432946 470646 432960
rect 470646 432946 470652 432960
rect 470676 432946 470698 432960
rect 470698 432946 470710 432960
rect 470710 432946 470732 432960
rect 470756 432946 470762 432960
rect 470762 432946 470774 432960
rect 470774 432946 470812 432960
rect 470276 432908 470314 432922
rect 470314 432908 470326 432922
rect 470326 432908 470332 432922
rect 470356 432908 470378 432922
rect 470378 432908 470390 432922
rect 470390 432908 470412 432922
rect 470436 432908 470442 432922
rect 470442 432908 470454 432922
rect 470454 432908 470492 432922
rect 470516 432908 470518 432922
rect 470518 432908 470570 432922
rect 470570 432908 470572 432922
rect 470596 432908 470634 432922
rect 470634 432908 470646 432922
rect 470646 432908 470652 432922
rect 470676 432908 470698 432922
rect 470698 432908 470710 432922
rect 470710 432908 470732 432922
rect 470756 432908 470762 432922
rect 470762 432908 470774 432922
rect 470774 432908 470812 432922
rect 470276 432896 470332 432908
rect 470356 432896 470412 432908
rect 470436 432896 470492 432908
rect 470516 432896 470572 432908
rect 470596 432896 470652 432908
rect 470676 432896 470732 432908
rect 470756 432896 470812 432908
rect 470276 432866 470314 432896
rect 470314 432866 470326 432896
rect 470326 432866 470332 432896
rect 470356 432866 470378 432896
rect 470378 432866 470390 432896
rect 470390 432866 470412 432896
rect 470436 432866 470442 432896
rect 470442 432866 470454 432896
rect 470454 432866 470492 432896
rect 470516 432866 470518 432896
rect 470518 432866 470570 432896
rect 470570 432866 470572 432896
rect 470596 432866 470634 432896
rect 470634 432866 470646 432896
rect 470646 432866 470652 432896
rect 470676 432866 470698 432896
rect 470698 432866 470710 432896
rect 470710 432866 470732 432896
rect 470756 432866 470762 432896
rect 470762 432866 470774 432896
rect 470774 432866 470812 432896
rect 470276 432832 470332 432842
rect 470356 432832 470412 432842
rect 470436 432832 470492 432842
rect 470516 432832 470572 432842
rect 470596 432832 470652 432842
rect 470676 432832 470732 432842
rect 470756 432832 470812 432842
rect 470276 432786 470314 432832
rect 470314 432786 470326 432832
rect 470326 432786 470332 432832
rect 470356 432786 470378 432832
rect 470378 432786 470390 432832
rect 470390 432786 470412 432832
rect 470436 432786 470442 432832
rect 470442 432786 470454 432832
rect 470454 432786 470492 432832
rect 470516 432786 470518 432832
rect 470518 432786 470570 432832
rect 470570 432786 470572 432832
rect 470596 432786 470634 432832
rect 470634 432786 470646 432832
rect 470646 432786 470652 432832
rect 470676 432786 470698 432832
rect 470698 432786 470710 432832
rect 470710 432786 470732 432832
rect 470756 432786 470762 432832
rect 470762 432786 470774 432832
rect 470774 432786 470812 432832
rect 483662 432794 483718 432850
rect 483570 432250 483626 432306
rect 469036 431949 469074 431995
rect 469074 431949 469086 431995
rect 469086 431949 469092 431995
rect 469116 431949 469138 431995
rect 469138 431949 469150 431995
rect 469150 431949 469172 431995
rect 469196 431949 469202 431995
rect 469202 431949 469214 431995
rect 469214 431949 469252 431995
rect 469276 431949 469278 431995
rect 469278 431949 469330 431995
rect 469330 431949 469332 431995
rect 469356 431949 469394 431995
rect 469394 431949 469406 431995
rect 469406 431949 469412 431995
rect 469436 431949 469458 431995
rect 469458 431949 469470 431995
rect 469470 431949 469492 431995
rect 469516 431949 469522 431995
rect 469522 431949 469534 431995
rect 469534 431949 469572 431995
rect 481270 432114 481326 432170
rect 469036 431939 469092 431949
rect 469116 431939 469172 431949
rect 469196 431939 469252 431949
rect 469276 431939 469332 431949
rect 469356 431939 469412 431949
rect 469436 431939 469492 431949
rect 469516 431939 469572 431949
rect 469036 431885 469074 431915
rect 469074 431885 469086 431915
rect 469086 431885 469092 431915
rect 469116 431885 469138 431915
rect 469138 431885 469150 431915
rect 469150 431885 469172 431915
rect 469196 431885 469202 431915
rect 469202 431885 469214 431915
rect 469214 431885 469252 431915
rect 469276 431885 469278 431915
rect 469278 431885 469330 431915
rect 469330 431885 469332 431915
rect 469356 431885 469394 431915
rect 469394 431885 469406 431915
rect 469406 431885 469412 431915
rect 469436 431885 469458 431915
rect 469458 431885 469470 431915
rect 469470 431885 469492 431915
rect 469516 431885 469522 431915
rect 469522 431885 469534 431915
rect 469534 431885 469572 431915
rect 469036 431873 469092 431885
rect 469116 431873 469172 431885
rect 469196 431873 469252 431885
rect 469276 431873 469332 431885
rect 469356 431873 469412 431885
rect 469436 431873 469492 431885
rect 469516 431873 469572 431885
rect 469036 431859 469074 431873
rect 469074 431859 469086 431873
rect 469086 431859 469092 431873
rect 469116 431859 469138 431873
rect 469138 431859 469150 431873
rect 469150 431859 469172 431873
rect 469196 431859 469202 431873
rect 469202 431859 469214 431873
rect 469214 431859 469252 431873
rect 469276 431859 469278 431873
rect 469278 431859 469330 431873
rect 469330 431859 469332 431873
rect 469356 431859 469394 431873
rect 469394 431859 469406 431873
rect 469406 431859 469412 431873
rect 469436 431859 469458 431873
rect 469458 431859 469470 431873
rect 469470 431859 469492 431873
rect 469516 431859 469522 431873
rect 469522 431859 469534 431873
rect 469534 431859 469572 431873
rect 469036 431821 469074 431835
rect 469074 431821 469086 431835
rect 469086 431821 469092 431835
rect 469116 431821 469138 431835
rect 469138 431821 469150 431835
rect 469150 431821 469172 431835
rect 469196 431821 469202 431835
rect 469202 431821 469214 431835
rect 469214 431821 469252 431835
rect 469276 431821 469278 431835
rect 469278 431821 469330 431835
rect 469330 431821 469332 431835
rect 469356 431821 469394 431835
rect 469394 431821 469406 431835
rect 469406 431821 469412 431835
rect 469436 431821 469458 431835
rect 469458 431821 469470 431835
rect 469470 431821 469492 431835
rect 469516 431821 469522 431835
rect 469522 431821 469534 431835
rect 469534 431821 469572 431835
rect 469036 431809 469092 431821
rect 469116 431809 469172 431821
rect 469196 431809 469252 431821
rect 469276 431809 469332 431821
rect 469356 431809 469412 431821
rect 469436 431809 469492 431821
rect 469516 431809 469572 431821
rect 469036 431779 469074 431809
rect 469074 431779 469086 431809
rect 469086 431779 469092 431809
rect 469116 431779 469138 431809
rect 469138 431779 469150 431809
rect 469150 431779 469172 431809
rect 469196 431779 469202 431809
rect 469202 431779 469214 431809
rect 469214 431779 469252 431809
rect 469276 431779 469278 431809
rect 469278 431779 469330 431809
rect 469330 431779 469332 431809
rect 469356 431779 469394 431809
rect 469394 431779 469406 431809
rect 469406 431779 469412 431809
rect 469436 431779 469458 431809
rect 469458 431779 469470 431809
rect 469470 431779 469492 431809
rect 469516 431779 469522 431809
rect 469522 431779 469534 431809
rect 469534 431779 469572 431809
rect 469036 431745 469092 431755
rect 469116 431745 469172 431755
rect 469196 431745 469252 431755
rect 469276 431745 469332 431755
rect 469356 431745 469412 431755
rect 469436 431745 469492 431755
rect 469516 431745 469572 431755
rect 469036 431699 469074 431745
rect 469074 431699 469086 431745
rect 469086 431699 469092 431745
rect 469116 431699 469138 431745
rect 469138 431699 469150 431745
rect 469150 431699 469172 431745
rect 469196 431699 469202 431745
rect 469202 431699 469214 431745
rect 469214 431699 469252 431745
rect 469276 431699 469278 431745
rect 469278 431699 469330 431745
rect 469330 431699 469332 431745
rect 469356 431699 469394 431745
rect 469394 431699 469406 431745
rect 469406 431699 469412 431745
rect 469436 431699 469458 431745
rect 469458 431699 469470 431745
rect 469470 431699 469492 431745
rect 469516 431699 469522 431745
rect 469522 431699 469534 431745
rect 469534 431699 469572 431745
rect 470276 430864 470314 430910
rect 470314 430864 470326 430910
rect 470326 430864 470332 430910
rect 470356 430864 470378 430910
rect 470378 430864 470390 430910
rect 470390 430864 470412 430910
rect 470436 430864 470442 430910
rect 470442 430864 470454 430910
rect 470454 430864 470492 430910
rect 470516 430864 470518 430910
rect 470518 430864 470570 430910
rect 470570 430864 470572 430910
rect 470596 430864 470634 430910
rect 470634 430864 470646 430910
rect 470646 430864 470652 430910
rect 470676 430864 470698 430910
rect 470698 430864 470710 430910
rect 470710 430864 470732 430910
rect 470756 430864 470762 430910
rect 470762 430864 470774 430910
rect 470774 430864 470812 430910
rect 470276 430854 470332 430864
rect 470356 430854 470412 430864
rect 470436 430854 470492 430864
rect 470516 430854 470572 430864
rect 470596 430854 470652 430864
rect 470676 430854 470732 430864
rect 470756 430854 470812 430864
rect 470276 430800 470314 430830
rect 470314 430800 470326 430830
rect 470326 430800 470332 430830
rect 470356 430800 470378 430830
rect 470378 430800 470390 430830
rect 470390 430800 470412 430830
rect 470436 430800 470442 430830
rect 470442 430800 470454 430830
rect 470454 430800 470492 430830
rect 470516 430800 470518 430830
rect 470518 430800 470570 430830
rect 470570 430800 470572 430830
rect 470596 430800 470634 430830
rect 470634 430800 470646 430830
rect 470646 430800 470652 430830
rect 470676 430800 470698 430830
rect 470698 430800 470710 430830
rect 470710 430800 470732 430830
rect 470756 430800 470762 430830
rect 470762 430800 470774 430830
rect 470774 430800 470812 430830
rect 470276 430788 470332 430800
rect 470356 430788 470412 430800
rect 470436 430788 470492 430800
rect 470516 430788 470572 430800
rect 470596 430788 470652 430800
rect 470676 430788 470732 430800
rect 470756 430788 470812 430800
rect 470276 430774 470314 430788
rect 470314 430774 470326 430788
rect 470326 430774 470332 430788
rect 470356 430774 470378 430788
rect 470378 430774 470390 430788
rect 470390 430774 470412 430788
rect 470436 430774 470442 430788
rect 470442 430774 470454 430788
rect 470454 430774 470492 430788
rect 470516 430774 470518 430788
rect 470518 430774 470570 430788
rect 470570 430774 470572 430788
rect 470596 430774 470634 430788
rect 470634 430774 470646 430788
rect 470646 430774 470652 430788
rect 470676 430774 470698 430788
rect 470698 430774 470710 430788
rect 470710 430774 470732 430788
rect 470756 430774 470762 430788
rect 470762 430774 470774 430788
rect 470774 430774 470812 430788
rect 470276 430736 470314 430750
rect 470314 430736 470326 430750
rect 470326 430736 470332 430750
rect 470356 430736 470378 430750
rect 470378 430736 470390 430750
rect 470390 430736 470412 430750
rect 470436 430736 470442 430750
rect 470442 430736 470454 430750
rect 470454 430736 470492 430750
rect 470516 430736 470518 430750
rect 470518 430736 470570 430750
rect 470570 430736 470572 430750
rect 470596 430736 470634 430750
rect 470634 430736 470646 430750
rect 470646 430736 470652 430750
rect 470676 430736 470698 430750
rect 470698 430736 470710 430750
rect 470710 430736 470732 430750
rect 470756 430736 470762 430750
rect 470762 430736 470774 430750
rect 470774 430736 470812 430750
rect 470276 430724 470332 430736
rect 470356 430724 470412 430736
rect 470436 430724 470492 430736
rect 470516 430724 470572 430736
rect 470596 430724 470652 430736
rect 470676 430724 470732 430736
rect 470756 430724 470812 430736
rect 470276 430694 470314 430724
rect 470314 430694 470326 430724
rect 470326 430694 470332 430724
rect 470356 430694 470378 430724
rect 470378 430694 470390 430724
rect 470390 430694 470412 430724
rect 470436 430694 470442 430724
rect 470442 430694 470454 430724
rect 470454 430694 470492 430724
rect 470516 430694 470518 430724
rect 470518 430694 470570 430724
rect 470570 430694 470572 430724
rect 470596 430694 470634 430724
rect 470634 430694 470646 430724
rect 470646 430694 470652 430724
rect 470676 430694 470698 430724
rect 470698 430694 470710 430724
rect 470710 430694 470732 430724
rect 470756 430694 470762 430724
rect 470762 430694 470774 430724
rect 470774 430694 470812 430724
rect 470276 430660 470332 430670
rect 470356 430660 470412 430670
rect 470436 430660 470492 430670
rect 470516 430660 470572 430670
rect 470596 430660 470652 430670
rect 470676 430660 470732 430670
rect 470756 430660 470812 430670
rect 470276 430614 470314 430660
rect 470314 430614 470326 430660
rect 470326 430614 470332 430660
rect 470356 430614 470378 430660
rect 470378 430614 470390 430660
rect 470390 430614 470412 430660
rect 470436 430614 470442 430660
rect 470442 430614 470454 430660
rect 470454 430614 470492 430660
rect 470516 430614 470518 430660
rect 470518 430614 470570 430660
rect 470570 430614 470572 430660
rect 470596 430614 470634 430660
rect 470634 430614 470646 430660
rect 470646 430614 470652 430660
rect 470676 430614 470698 430660
rect 470698 430614 470710 430660
rect 470710 430614 470732 430660
rect 470756 430614 470762 430660
rect 470762 430614 470774 430660
rect 470774 430614 470812 430660
rect 470276 412036 470314 412082
rect 470314 412036 470326 412082
rect 470326 412036 470332 412082
rect 470356 412036 470378 412082
rect 470378 412036 470390 412082
rect 470390 412036 470412 412082
rect 470436 412036 470442 412082
rect 470442 412036 470454 412082
rect 470454 412036 470492 412082
rect 470516 412036 470518 412082
rect 470518 412036 470570 412082
rect 470570 412036 470572 412082
rect 470596 412036 470634 412082
rect 470634 412036 470646 412082
rect 470646 412036 470652 412082
rect 470676 412036 470698 412082
rect 470698 412036 470710 412082
rect 470710 412036 470732 412082
rect 470756 412036 470762 412082
rect 470762 412036 470774 412082
rect 470774 412036 470812 412082
rect 470276 412026 470332 412036
rect 470356 412026 470412 412036
rect 470436 412026 470492 412036
rect 470516 412026 470572 412036
rect 470596 412026 470652 412036
rect 470676 412026 470732 412036
rect 470756 412026 470812 412036
rect 470276 411972 470314 412002
rect 470314 411972 470326 412002
rect 470326 411972 470332 412002
rect 470356 411972 470378 412002
rect 470378 411972 470390 412002
rect 470390 411972 470412 412002
rect 470436 411972 470442 412002
rect 470442 411972 470454 412002
rect 470454 411972 470492 412002
rect 470516 411972 470518 412002
rect 470518 411972 470570 412002
rect 470570 411972 470572 412002
rect 470596 411972 470634 412002
rect 470634 411972 470646 412002
rect 470646 411972 470652 412002
rect 470676 411972 470698 412002
rect 470698 411972 470710 412002
rect 470710 411972 470732 412002
rect 470756 411972 470762 412002
rect 470762 411972 470774 412002
rect 470774 411972 470812 412002
rect 470276 411960 470332 411972
rect 470356 411960 470412 411972
rect 470436 411960 470492 411972
rect 470516 411960 470572 411972
rect 470596 411960 470652 411972
rect 470676 411960 470732 411972
rect 470756 411960 470812 411972
rect 470276 411946 470314 411960
rect 470314 411946 470326 411960
rect 470326 411946 470332 411960
rect 470356 411946 470378 411960
rect 470378 411946 470390 411960
rect 470390 411946 470412 411960
rect 470436 411946 470442 411960
rect 470442 411946 470454 411960
rect 470454 411946 470492 411960
rect 470516 411946 470518 411960
rect 470518 411946 470570 411960
rect 470570 411946 470572 411960
rect 470596 411946 470634 411960
rect 470634 411946 470646 411960
rect 470646 411946 470652 411960
rect 470676 411946 470698 411960
rect 470698 411946 470710 411960
rect 470710 411946 470732 411960
rect 470756 411946 470762 411960
rect 470762 411946 470774 411960
rect 470774 411946 470812 411960
rect 470276 411908 470314 411922
rect 470314 411908 470326 411922
rect 470326 411908 470332 411922
rect 470356 411908 470378 411922
rect 470378 411908 470390 411922
rect 470390 411908 470412 411922
rect 470436 411908 470442 411922
rect 470442 411908 470454 411922
rect 470454 411908 470492 411922
rect 470516 411908 470518 411922
rect 470518 411908 470570 411922
rect 470570 411908 470572 411922
rect 470596 411908 470634 411922
rect 470634 411908 470646 411922
rect 470646 411908 470652 411922
rect 470676 411908 470698 411922
rect 470698 411908 470710 411922
rect 470710 411908 470732 411922
rect 470756 411908 470762 411922
rect 470762 411908 470774 411922
rect 470774 411908 470812 411922
rect 470276 411896 470332 411908
rect 470356 411896 470412 411908
rect 470436 411896 470492 411908
rect 470516 411896 470572 411908
rect 470596 411896 470652 411908
rect 470676 411896 470732 411908
rect 470756 411896 470812 411908
rect 470276 411866 470314 411896
rect 470314 411866 470326 411896
rect 470326 411866 470332 411896
rect 470356 411866 470378 411896
rect 470378 411866 470390 411896
rect 470390 411866 470412 411896
rect 470436 411866 470442 411896
rect 470442 411866 470454 411896
rect 470454 411866 470492 411896
rect 470516 411866 470518 411896
rect 470518 411866 470570 411896
rect 470570 411866 470572 411896
rect 470596 411866 470634 411896
rect 470634 411866 470646 411896
rect 470646 411866 470652 411896
rect 470676 411866 470698 411896
rect 470698 411866 470710 411896
rect 470710 411866 470732 411896
rect 470756 411866 470762 411896
rect 470762 411866 470774 411896
rect 470774 411866 470812 411896
rect 470276 411832 470332 411842
rect 470356 411832 470412 411842
rect 470436 411832 470492 411842
rect 470516 411832 470572 411842
rect 470596 411832 470652 411842
rect 470676 411832 470732 411842
rect 470756 411832 470812 411842
rect 470276 411786 470314 411832
rect 470314 411786 470326 411832
rect 470326 411786 470332 411832
rect 470356 411786 470378 411832
rect 470378 411786 470390 411832
rect 470390 411786 470412 411832
rect 470436 411786 470442 411832
rect 470442 411786 470454 411832
rect 470454 411786 470492 411832
rect 470516 411786 470518 411832
rect 470518 411786 470570 411832
rect 470570 411786 470572 411832
rect 470596 411786 470634 411832
rect 470634 411786 470646 411832
rect 470646 411786 470652 411832
rect 470676 411786 470698 411832
rect 470698 411786 470710 411832
rect 470710 411786 470732 411832
rect 470756 411786 470762 411832
rect 470762 411786 470774 411832
rect 470774 411786 470812 411832
rect 474278 431842 474334 431898
rect 478102 431570 478158 431626
rect 488433 431570 488489 431626
rect 478970 427898 479026 427954
rect 485778 427898 485834 427954
rect 488538 413890 488594 413946
rect 469036 410950 469074 410996
rect 469074 410950 469086 410996
rect 469086 410950 469092 410996
rect 469116 410950 469138 410996
rect 469138 410950 469150 410996
rect 469150 410950 469172 410996
rect 469196 410950 469202 410996
rect 469202 410950 469214 410996
rect 469214 410950 469252 410996
rect 469276 410950 469278 410996
rect 469278 410950 469330 410996
rect 469330 410950 469332 410996
rect 469356 410950 469394 410996
rect 469394 410950 469406 410996
rect 469406 410950 469412 410996
rect 469436 410950 469458 410996
rect 469458 410950 469470 410996
rect 469470 410950 469492 410996
rect 469516 410950 469522 410996
rect 469522 410950 469534 410996
rect 469534 410950 469572 410996
rect 469036 410940 469092 410950
rect 469116 410940 469172 410950
rect 469196 410940 469252 410950
rect 469276 410940 469332 410950
rect 469356 410940 469412 410950
rect 469436 410940 469492 410950
rect 469516 410940 469572 410950
rect 469036 410886 469074 410916
rect 469074 410886 469086 410916
rect 469086 410886 469092 410916
rect 469116 410886 469138 410916
rect 469138 410886 469150 410916
rect 469150 410886 469172 410916
rect 469196 410886 469202 410916
rect 469202 410886 469214 410916
rect 469214 410886 469252 410916
rect 469276 410886 469278 410916
rect 469278 410886 469330 410916
rect 469330 410886 469332 410916
rect 469356 410886 469394 410916
rect 469394 410886 469406 410916
rect 469406 410886 469412 410916
rect 469436 410886 469458 410916
rect 469458 410886 469470 410916
rect 469470 410886 469492 410916
rect 469516 410886 469522 410916
rect 469522 410886 469534 410916
rect 469534 410886 469572 410916
rect 469036 410874 469092 410886
rect 469116 410874 469172 410886
rect 469196 410874 469252 410886
rect 469276 410874 469332 410886
rect 469356 410874 469412 410886
rect 469436 410874 469492 410886
rect 469516 410874 469572 410886
rect 469036 410860 469074 410874
rect 469074 410860 469086 410874
rect 469086 410860 469092 410874
rect 469116 410860 469138 410874
rect 469138 410860 469150 410874
rect 469150 410860 469172 410874
rect 469196 410860 469202 410874
rect 469202 410860 469214 410874
rect 469214 410860 469252 410874
rect 469276 410860 469278 410874
rect 469278 410860 469330 410874
rect 469330 410860 469332 410874
rect 469356 410860 469394 410874
rect 469394 410860 469406 410874
rect 469406 410860 469412 410874
rect 469436 410860 469458 410874
rect 469458 410860 469470 410874
rect 469470 410860 469492 410874
rect 469516 410860 469522 410874
rect 469522 410860 469534 410874
rect 469534 410860 469572 410874
rect 469036 410822 469074 410836
rect 469074 410822 469086 410836
rect 469086 410822 469092 410836
rect 469116 410822 469138 410836
rect 469138 410822 469150 410836
rect 469150 410822 469172 410836
rect 469196 410822 469202 410836
rect 469202 410822 469214 410836
rect 469214 410822 469252 410836
rect 469276 410822 469278 410836
rect 469278 410822 469330 410836
rect 469330 410822 469332 410836
rect 469356 410822 469394 410836
rect 469394 410822 469406 410836
rect 469406 410822 469412 410836
rect 469436 410822 469458 410836
rect 469458 410822 469470 410836
rect 469470 410822 469492 410836
rect 469516 410822 469522 410836
rect 469522 410822 469534 410836
rect 469534 410822 469572 410836
rect 469036 410810 469092 410822
rect 469116 410810 469172 410822
rect 469196 410810 469252 410822
rect 469276 410810 469332 410822
rect 469356 410810 469412 410822
rect 469436 410810 469492 410822
rect 469516 410810 469572 410822
rect 469036 410780 469074 410810
rect 469074 410780 469086 410810
rect 469086 410780 469092 410810
rect 469116 410780 469138 410810
rect 469138 410780 469150 410810
rect 469150 410780 469172 410810
rect 469196 410780 469202 410810
rect 469202 410780 469214 410810
rect 469214 410780 469252 410810
rect 469276 410780 469278 410810
rect 469278 410780 469330 410810
rect 469330 410780 469332 410810
rect 469356 410780 469394 410810
rect 469394 410780 469406 410810
rect 469406 410780 469412 410810
rect 469436 410780 469458 410810
rect 469458 410780 469470 410810
rect 469470 410780 469492 410810
rect 469516 410780 469522 410810
rect 469522 410780 469534 410810
rect 469534 410780 469572 410810
rect 469036 410746 469092 410756
rect 469116 410746 469172 410756
rect 469196 410746 469252 410756
rect 469276 410746 469332 410756
rect 469356 410746 469412 410756
rect 469436 410746 469492 410756
rect 469516 410746 469572 410756
rect 469036 410700 469074 410746
rect 469074 410700 469086 410746
rect 469086 410700 469092 410746
rect 469116 410700 469138 410746
rect 469138 410700 469150 410746
rect 469150 410700 469172 410746
rect 469196 410700 469202 410746
rect 469202 410700 469214 410746
rect 469214 410700 469252 410746
rect 469276 410700 469278 410746
rect 469278 410700 469330 410746
rect 469330 410700 469332 410746
rect 469356 410700 469394 410746
rect 469394 410700 469406 410746
rect 469406 410700 469412 410746
rect 469436 410700 469458 410746
rect 469458 410700 469470 410746
rect 469470 410700 469492 410746
rect 469516 410700 469522 410746
rect 469522 410700 469534 410746
rect 469534 410700 469572 410746
rect 470276 409864 470314 409910
rect 470314 409864 470326 409910
rect 470326 409864 470332 409910
rect 470356 409864 470378 409910
rect 470378 409864 470390 409910
rect 470390 409864 470412 409910
rect 470436 409864 470442 409910
rect 470442 409864 470454 409910
rect 470454 409864 470492 409910
rect 470516 409864 470518 409910
rect 470518 409864 470570 409910
rect 470570 409864 470572 409910
rect 470596 409864 470634 409910
rect 470634 409864 470646 409910
rect 470646 409864 470652 409910
rect 470676 409864 470698 409910
rect 470698 409864 470710 409910
rect 470710 409864 470732 409910
rect 470756 409864 470762 409910
rect 470762 409864 470774 409910
rect 470774 409864 470812 409910
rect 470276 409854 470332 409864
rect 470356 409854 470412 409864
rect 470436 409854 470492 409864
rect 470516 409854 470572 409864
rect 470596 409854 470652 409864
rect 470676 409854 470732 409864
rect 470756 409854 470812 409864
rect 470276 409800 470314 409830
rect 470314 409800 470326 409830
rect 470326 409800 470332 409830
rect 470356 409800 470378 409830
rect 470378 409800 470390 409830
rect 470390 409800 470412 409830
rect 470436 409800 470442 409830
rect 470442 409800 470454 409830
rect 470454 409800 470492 409830
rect 470516 409800 470518 409830
rect 470518 409800 470570 409830
rect 470570 409800 470572 409830
rect 470596 409800 470634 409830
rect 470634 409800 470646 409830
rect 470646 409800 470652 409830
rect 470676 409800 470698 409830
rect 470698 409800 470710 409830
rect 470710 409800 470732 409830
rect 470756 409800 470762 409830
rect 470762 409800 470774 409830
rect 470774 409800 470812 409830
rect 470276 409788 470332 409800
rect 470356 409788 470412 409800
rect 470436 409788 470492 409800
rect 470516 409788 470572 409800
rect 470596 409788 470652 409800
rect 470676 409788 470732 409800
rect 470756 409788 470812 409800
rect 470276 409774 470314 409788
rect 470314 409774 470326 409788
rect 470326 409774 470332 409788
rect 470356 409774 470378 409788
rect 470378 409774 470390 409788
rect 470390 409774 470412 409788
rect 470436 409774 470442 409788
rect 470442 409774 470454 409788
rect 470454 409774 470492 409788
rect 470516 409774 470518 409788
rect 470518 409774 470570 409788
rect 470570 409774 470572 409788
rect 470596 409774 470634 409788
rect 470634 409774 470646 409788
rect 470646 409774 470652 409788
rect 470676 409774 470698 409788
rect 470698 409774 470710 409788
rect 470710 409774 470732 409788
rect 470756 409774 470762 409788
rect 470762 409774 470774 409788
rect 470774 409774 470812 409788
rect 470276 409736 470314 409750
rect 470314 409736 470326 409750
rect 470326 409736 470332 409750
rect 470356 409736 470378 409750
rect 470378 409736 470390 409750
rect 470390 409736 470412 409750
rect 470436 409736 470442 409750
rect 470442 409736 470454 409750
rect 470454 409736 470492 409750
rect 470516 409736 470518 409750
rect 470518 409736 470570 409750
rect 470570 409736 470572 409750
rect 470596 409736 470634 409750
rect 470634 409736 470646 409750
rect 470646 409736 470652 409750
rect 470676 409736 470698 409750
rect 470698 409736 470710 409750
rect 470710 409736 470732 409750
rect 470756 409736 470762 409750
rect 470762 409736 470774 409750
rect 470774 409736 470812 409750
rect 470276 409724 470332 409736
rect 470356 409724 470412 409736
rect 470436 409724 470492 409736
rect 470516 409724 470572 409736
rect 470596 409724 470652 409736
rect 470676 409724 470732 409736
rect 470756 409724 470812 409736
rect 470276 409694 470314 409724
rect 470314 409694 470326 409724
rect 470326 409694 470332 409724
rect 470356 409694 470378 409724
rect 470378 409694 470390 409724
rect 470390 409694 470412 409724
rect 470436 409694 470442 409724
rect 470442 409694 470454 409724
rect 470454 409694 470492 409724
rect 470516 409694 470518 409724
rect 470518 409694 470570 409724
rect 470570 409694 470572 409724
rect 470596 409694 470634 409724
rect 470634 409694 470646 409724
rect 470646 409694 470652 409724
rect 470676 409694 470698 409724
rect 470698 409694 470710 409724
rect 470710 409694 470732 409724
rect 470756 409694 470762 409724
rect 470762 409694 470774 409724
rect 470774 409694 470812 409724
rect 470276 409660 470332 409670
rect 470356 409660 470412 409670
rect 470436 409660 470492 409670
rect 470516 409660 470572 409670
rect 470596 409660 470652 409670
rect 470676 409660 470732 409670
rect 470756 409660 470812 409670
rect 470276 409614 470314 409660
rect 470314 409614 470326 409660
rect 470326 409614 470332 409660
rect 470356 409614 470378 409660
rect 470378 409614 470390 409660
rect 470390 409614 470412 409660
rect 470436 409614 470442 409660
rect 470442 409614 470454 409660
rect 470454 409614 470492 409660
rect 470516 409614 470518 409660
rect 470518 409614 470570 409660
rect 470570 409614 470572 409660
rect 470596 409614 470634 409660
rect 470634 409614 470646 409660
rect 470646 409614 470652 409660
rect 470676 409614 470698 409660
rect 470698 409614 470710 409660
rect 470710 409614 470732 409660
rect 470756 409614 470762 409660
rect 470762 409614 470774 409660
rect 470774 409614 470812 409660
rect 470276 391037 470314 391083
rect 470314 391037 470326 391083
rect 470326 391037 470332 391083
rect 470356 391037 470378 391083
rect 470378 391037 470390 391083
rect 470390 391037 470412 391083
rect 470436 391037 470442 391083
rect 470442 391037 470454 391083
rect 470454 391037 470492 391083
rect 470516 391037 470518 391083
rect 470518 391037 470570 391083
rect 470570 391037 470572 391083
rect 470596 391037 470634 391083
rect 470634 391037 470646 391083
rect 470646 391037 470652 391083
rect 470676 391037 470698 391083
rect 470698 391037 470710 391083
rect 470710 391037 470732 391083
rect 470756 391037 470762 391083
rect 470762 391037 470774 391083
rect 470774 391037 470812 391083
rect 470276 391027 470332 391037
rect 470356 391027 470412 391037
rect 470436 391027 470492 391037
rect 470516 391027 470572 391037
rect 470596 391027 470652 391037
rect 470676 391027 470732 391037
rect 470756 391027 470812 391037
rect 470276 390973 470314 391003
rect 470314 390973 470326 391003
rect 470326 390973 470332 391003
rect 470356 390973 470378 391003
rect 470378 390973 470390 391003
rect 470390 390973 470412 391003
rect 470436 390973 470442 391003
rect 470442 390973 470454 391003
rect 470454 390973 470492 391003
rect 470516 390973 470518 391003
rect 470518 390973 470570 391003
rect 470570 390973 470572 391003
rect 470596 390973 470634 391003
rect 470634 390973 470646 391003
rect 470646 390973 470652 391003
rect 470676 390973 470698 391003
rect 470698 390973 470710 391003
rect 470710 390973 470732 391003
rect 470756 390973 470762 391003
rect 470762 390973 470774 391003
rect 470774 390973 470812 391003
rect 470276 390961 470332 390973
rect 470356 390961 470412 390973
rect 470436 390961 470492 390973
rect 470516 390961 470572 390973
rect 470596 390961 470652 390973
rect 470676 390961 470732 390973
rect 470756 390961 470812 390973
rect 470276 390947 470314 390961
rect 470314 390947 470326 390961
rect 470326 390947 470332 390961
rect 470356 390947 470378 390961
rect 470378 390947 470390 390961
rect 470390 390947 470412 390961
rect 470436 390947 470442 390961
rect 470442 390947 470454 390961
rect 470454 390947 470492 390961
rect 470516 390947 470518 390961
rect 470518 390947 470570 390961
rect 470570 390947 470572 390961
rect 470596 390947 470634 390961
rect 470634 390947 470646 390961
rect 470646 390947 470652 390961
rect 470676 390947 470698 390961
rect 470698 390947 470710 390961
rect 470710 390947 470732 390961
rect 470756 390947 470762 390961
rect 470762 390947 470774 390961
rect 470774 390947 470812 390961
rect 470276 390909 470314 390923
rect 470314 390909 470326 390923
rect 470326 390909 470332 390923
rect 470356 390909 470378 390923
rect 470378 390909 470390 390923
rect 470390 390909 470412 390923
rect 470436 390909 470442 390923
rect 470442 390909 470454 390923
rect 470454 390909 470492 390923
rect 470516 390909 470518 390923
rect 470518 390909 470570 390923
rect 470570 390909 470572 390923
rect 470596 390909 470634 390923
rect 470634 390909 470646 390923
rect 470646 390909 470652 390923
rect 470676 390909 470698 390923
rect 470698 390909 470710 390923
rect 470710 390909 470732 390923
rect 470756 390909 470762 390923
rect 470762 390909 470774 390923
rect 470774 390909 470812 390923
rect 470276 390897 470332 390909
rect 470356 390897 470412 390909
rect 470436 390897 470492 390909
rect 470516 390897 470572 390909
rect 470596 390897 470652 390909
rect 470676 390897 470732 390909
rect 470756 390897 470812 390909
rect 470276 390867 470314 390897
rect 470314 390867 470326 390897
rect 470326 390867 470332 390897
rect 470356 390867 470378 390897
rect 470378 390867 470390 390897
rect 470390 390867 470412 390897
rect 470436 390867 470442 390897
rect 470442 390867 470454 390897
rect 470454 390867 470492 390897
rect 470516 390867 470518 390897
rect 470518 390867 470570 390897
rect 470570 390867 470572 390897
rect 470596 390867 470634 390897
rect 470634 390867 470646 390897
rect 470646 390867 470652 390897
rect 470676 390867 470698 390897
rect 470698 390867 470710 390897
rect 470710 390867 470732 390897
rect 470756 390867 470762 390897
rect 470762 390867 470774 390897
rect 470774 390867 470812 390897
rect 470276 390833 470332 390843
rect 470356 390833 470412 390843
rect 470436 390833 470492 390843
rect 470516 390833 470572 390843
rect 470596 390833 470652 390843
rect 470676 390833 470732 390843
rect 470756 390833 470812 390843
rect 470276 390787 470314 390833
rect 470314 390787 470326 390833
rect 470326 390787 470332 390833
rect 470356 390787 470378 390833
rect 470378 390787 470390 390833
rect 470390 390787 470412 390833
rect 470436 390787 470442 390833
rect 470442 390787 470454 390833
rect 470454 390787 470492 390833
rect 470516 390787 470518 390833
rect 470518 390787 470570 390833
rect 470570 390787 470572 390833
rect 470596 390787 470634 390833
rect 470634 390787 470646 390833
rect 470646 390787 470652 390833
rect 470676 390787 470698 390833
rect 470698 390787 470710 390833
rect 470710 390787 470732 390833
rect 470756 390787 470762 390833
rect 470762 390787 470774 390833
rect 470774 390787 470812 390833
rect 473726 410898 473782 410954
rect 478418 410082 478474 410138
rect 484122 410354 484178 410410
rect 481362 410082 481418 410138
rect 487618 409946 487674 410002
rect 488538 409946 488594 410002
rect 489826 409946 489882 410002
rect 481822 407090 481878 407146
rect 485134 407090 485190 407146
rect 489826 391994 489882 392050
rect 469036 389954 469074 390000
rect 469074 389954 469086 390000
rect 469086 389954 469092 390000
rect 469116 389954 469138 390000
rect 469138 389954 469150 390000
rect 469150 389954 469172 390000
rect 469196 389954 469202 390000
rect 469202 389954 469214 390000
rect 469214 389954 469252 390000
rect 469276 389954 469278 390000
rect 469278 389954 469330 390000
rect 469330 389954 469332 390000
rect 469356 389954 469394 390000
rect 469394 389954 469406 390000
rect 469406 389954 469412 390000
rect 469436 389954 469458 390000
rect 469458 389954 469470 390000
rect 469470 389954 469492 390000
rect 469516 389954 469522 390000
rect 469522 389954 469534 390000
rect 469534 389954 469572 390000
rect 469036 389944 469092 389954
rect 469116 389944 469172 389954
rect 469196 389944 469252 389954
rect 469276 389944 469332 389954
rect 469356 389944 469412 389954
rect 469436 389944 469492 389954
rect 469516 389944 469572 389954
rect 469036 389890 469074 389920
rect 469074 389890 469086 389920
rect 469086 389890 469092 389920
rect 469116 389890 469138 389920
rect 469138 389890 469150 389920
rect 469150 389890 469172 389920
rect 469196 389890 469202 389920
rect 469202 389890 469214 389920
rect 469214 389890 469252 389920
rect 469276 389890 469278 389920
rect 469278 389890 469330 389920
rect 469330 389890 469332 389920
rect 469356 389890 469394 389920
rect 469394 389890 469406 389920
rect 469406 389890 469412 389920
rect 469436 389890 469458 389920
rect 469458 389890 469470 389920
rect 469470 389890 469492 389920
rect 469516 389890 469522 389920
rect 469522 389890 469534 389920
rect 469534 389890 469572 389920
rect 469036 389878 469092 389890
rect 469116 389878 469172 389890
rect 469196 389878 469252 389890
rect 469276 389878 469332 389890
rect 469356 389878 469412 389890
rect 469436 389878 469492 389890
rect 469516 389878 469572 389890
rect 469036 389864 469074 389878
rect 469074 389864 469086 389878
rect 469086 389864 469092 389878
rect 469116 389864 469138 389878
rect 469138 389864 469150 389878
rect 469150 389864 469172 389878
rect 469196 389864 469202 389878
rect 469202 389864 469214 389878
rect 469214 389864 469252 389878
rect 469276 389864 469278 389878
rect 469278 389864 469330 389878
rect 469330 389864 469332 389878
rect 469356 389864 469394 389878
rect 469394 389864 469406 389878
rect 469406 389864 469412 389878
rect 469436 389864 469458 389878
rect 469458 389864 469470 389878
rect 469470 389864 469492 389878
rect 469516 389864 469522 389878
rect 469522 389864 469534 389878
rect 469534 389864 469572 389878
rect 469036 389826 469074 389840
rect 469074 389826 469086 389840
rect 469086 389826 469092 389840
rect 469116 389826 469138 389840
rect 469138 389826 469150 389840
rect 469150 389826 469172 389840
rect 469196 389826 469202 389840
rect 469202 389826 469214 389840
rect 469214 389826 469252 389840
rect 469276 389826 469278 389840
rect 469278 389826 469330 389840
rect 469330 389826 469332 389840
rect 469356 389826 469394 389840
rect 469394 389826 469406 389840
rect 469406 389826 469412 389840
rect 469436 389826 469458 389840
rect 469458 389826 469470 389840
rect 469470 389826 469492 389840
rect 469516 389826 469522 389840
rect 469522 389826 469534 389840
rect 469534 389826 469572 389840
rect 469036 389814 469092 389826
rect 469116 389814 469172 389826
rect 469196 389814 469252 389826
rect 469276 389814 469332 389826
rect 469356 389814 469412 389826
rect 469436 389814 469492 389826
rect 469516 389814 469572 389826
rect 469036 389784 469074 389814
rect 469074 389784 469086 389814
rect 469086 389784 469092 389814
rect 469116 389784 469138 389814
rect 469138 389784 469150 389814
rect 469150 389784 469172 389814
rect 469196 389784 469202 389814
rect 469202 389784 469214 389814
rect 469214 389784 469252 389814
rect 469276 389784 469278 389814
rect 469278 389784 469330 389814
rect 469330 389784 469332 389814
rect 469356 389784 469394 389814
rect 469394 389784 469406 389814
rect 469406 389784 469412 389814
rect 469436 389784 469458 389814
rect 469458 389784 469470 389814
rect 469470 389784 469492 389814
rect 469516 389784 469522 389814
rect 469522 389784 469534 389814
rect 469534 389784 469572 389814
rect 469036 389750 469092 389760
rect 469116 389750 469172 389760
rect 469196 389750 469252 389760
rect 469276 389750 469332 389760
rect 469356 389750 469412 389760
rect 469436 389750 469492 389760
rect 469516 389750 469572 389760
rect 469036 389704 469074 389750
rect 469074 389704 469086 389750
rect 469086 389704 469092 389750
rect 469116 389704 469138 389750
rect 469138 389704 469150 389750
rect 469150 389704 469172 389750
rect 469196 389704 469202 389750
rect 469202 389704 469214 389750
rect 469214 389704 469252 389750
rect 469276 389704 469278 389750
rect 469278 389704 469330 389750
rect 469330 389704 469332 389750
rect 469356 389704 469394 389750
rect 469394 389704 469406 389750
rect 469406 389704 469412 389750
rect 469436 389704 469458 389750
rect 469458 389704 469470 389750
rect 469470 389704 469492 389750
rect 469516 389704 469522 389750
rect 469522 389704 469534 389750
rect 469534 389704 469572 389750
rect 470276 388864 470314 388910
rect 470314 388864 470326 388910
rect 470326 388864 470332 388910
rect 470356 388864 470378 388910
rect 470378 388864 470390 388910
rect 470390 388864 470412 388910
rect 470436 388864 470442 388910
rect 470442 388864 470454 388910
rect 470454 388864 470492 388910
rect 470516 388864 470518 388910
rect 470518 388864 470570 388910
rect 470570 388864 470572 388910
rect 470596 388864 470634 388910
rect 470634 388864 470646 388910
rect 470646 388864 470652 388910
rect 470676 388864 470698 388910
rect 470698 388864 470710 388910
rect 470710 388864 470732 388910
rect 470756 388864 470762 388910
rect 470762 388864 470774 388910
rect 470774 388864 470812 388910
rect 470276 388854 470332 388864
rect 470356 388854 470412 388864
rect 470436 388854 470492 388864
rect 470516 388854 470572 388864
rect 470596 388854 470652 388864
rect 470676 388854 470732 388864
rect 470756 388854 470812 388864
rect 470276 388800 470314 388830
rect 470314 388800 470326 388830
rect 470326 388800 470332 388830
rect 470356 388800 470378 388830
rect 470378 388800 470390 388830
rect 470390 388800 470412 388830
rect 470436 388800 470442 388830
rect 470442 388800 470454 388830
rect 470454 388800 470492 388830
rect 470516 388800 470518 388830
rect 470518 388800 470570 388830
rect 470570 388800 470572 388830
rect 470596 388800 470634 388830
rect 470634 388800 470646 388830
rect 470646 388800 470652 388830
rect 470676 388800 470698 388830
rect 470698 388800 470710 388830
rect 470710 388800 470732 388830
rect 470756 388800 470762 388830
rect 470762 388800 470774 388830
rect 470774 388800 470812 388830
rect 470276 388788 470332 388800
rect 470356 388788 470412 388800
rect 470436 388788 470492 388800
rect 470516 388788 470572 388800
rect 470596 388788 470652 388800
rect 470676 388788 470732 388800
rect 470756 388788 470812 388800
rect 470276 388774 470314 388788
rect 470314 388774 470326 388788
rect 470326 388774 470332 388788
rect 470356 388774 470378 388788
rect 470378 388774 470390 388788
rect 470390 388774 470412 388788
rect 470436 388774 470442 388788
rect 470442 388774 470454 388788
rect 470454 388774 470492 388788
rect 470516 388774 470518 388788
rect 470518 388774 470570 388788
rect 470570 388774 470572 388788
rect 470596 388774 470634 388788
rect 470634 388774 470646 388788
rect 470646 388774 470652 388788
rect 470676 388774 470698 388788
rect 470698 388774 470710 388788
rect 470710 388774 470732 388788
rect 470756 388774 470762 388788
rect 470762 388774 470774 388788
rect 470774 388774 470812 388788
rect 470276 388736 470314 388750
rect 470314 388736 470326 388750
rect 470326 388736 470332 388750
rect 470356 388736 470378 388750
rect 470378 388736 470390 388750
rect 470390 388736 470412 388750
rect 470436 388736 470442 388750
rect 470442 388736 470454 388750
rect 470454 388736 470492 388750
rect 470516 388736 470518 388750
rect 470518 388736 470570 388750
rect 470570 388736 470572 388750
rect 470596 388736 470634 388750
rect 470634 388736 470646 388750
rect 470646 388736 470652 388750
rect 470676 388736 470698 388750
rect 470698 388736 470710 388750
rect 470710 388736 470732 388750
rect 470756 388736 470762 388750
rect 470762 388736 470774 388750
rect 470774 388736 470812 388750
rect 470276 388724 470332 388736
rect 470356 388724 470412 388736
rect 470436 388724 470492 388736
rect 470516 388724 470572 388736
rect 470596 388724 470652 388736
rect 470676 388724 470732 388736
rect 470756 388724 470812 388736
rect 470276 388694 470314 388724
rect 470314 388694 470326 388724
rect 470326 388694 470332 388724
rect 470356 388694 470378 388724
rect 470378 388694 470390 388724
rect 470390 388694 470412 388724
rect 470436 388694 470442 388724
rect 470442 388694 470454 388724
rect 470454 388694 470492 388724
rect 470516 388694 470518 388724
rect 470518 388694 470570 388724
rect 470570 388694 470572 388724
rect 470596 388694 470634 388724
rect 470634 388694 470646 388724
rect 470646 388694 470652 388724
rect 470676 388694 470698 388724
rect 470698 388694 470710 388724
rect 470710 388694 470732 388724
rect 470756 388694 470762 388724
rect 470762 388694 470774 388724
rect 470774 388694 470812 388724
rect 470276 388660 470332 388670
rect 470356 388660 470412 388670
rect 470436 388660 470492 388670
rect 470516 388660 470572 388670
rect 470596 388660 470652 388670
rect 470676 388660 470732 388670
rect 470756 388660 470812 388670
rect 470276 388614 470314 388660
rect 470314 388614 470326 388660
rect 470326 388614 470332 388660
rect 470356 388614 470378 388660
rect 470378 388614 470390 388660
rect 470390 388614 470412 388660
rect 470436 388614 470442 388660
rect 470442 388614 470454 388660
rect 470454 388614 470492 388660
rect 470516 388614 470518 388660
rect 470518 388614 470570 388660
rect 470570 388614 470572 388660
rect 470596 388614 470634 388660
rect 470634 388614 470646 388660
rect 470646 388614 470652 388660
rect 470676 388614 470698 388660
rect 470698 388614 470710 388660
rect 470710 388614 470732 388660
rect 470756 388614 470762 388660
rect 470762 388614 470774 388660
rect 470774 388614 470812 388660
rect 470276 358437 470314 358483
rect 470314 358437 470326 358483
rect 470326 358437 470332 358483
rect 470356 358437 470378 358483
rect 470378 358437 470390 358483
rect 470390 358437 470412 358483
rect 470436 358437 470442 358483
rect 470442 358437 470454 358483
rect 470454 358437 470492 358483
rect 470516 358437 470518 358483
rect 470518 358437 470570 358483
rect 470570 358437 470572 358483
rect 470596 358437 470634 358483
rect 470634 358437 470646 358483
rect 470646 358437 470652 358483
rect 470676 358437 470698 358483
rect 470698 358437 470710 358483
rect 470710 358437 470732 358483
rect 470756 358437 470762 358483
rect 470762 358437 470774 358483
rect 470774 358437 470812 358483
rect 470276 358427 470332 358437
rect 470356 358427 470412 358437
rect 470436 358427 470492 358437
rect 470516 358427 470572 358437
rect 470596 358427 470652 358437
rect 470676 358427 470732 358437
rect 470756 358427 470812 358437
rect 470276 358373 470314 358403
rect 470314 358373 470326 358403
rect 470326 358373 470332 358403
rect 470356 358373 470378 358403
rect 470378 358373 470390 358403
rect 470390 358373 470412 358403
rect 470436 358373 470442 358403
rect 470442 358373 470454 358403
rect 470454 358373 470492 358403
rect 470516 358373 470518 358403
rect 470518 358373 470570 358403
rect 470570 358373 470572 358403
rect 470596 358373 470634 358403
rect 470634 358373 470646 358403
rect 470646 358373 470652 358403
rect 470676 358373 470698 358403
rect 470698 358373 470710 358403
rect 470710 358373 470732 358403
rect 470756 358373 470762 358403
rect 470762 358373 470774 358403
rect 470774 358373 470812 358403
rect 470276 358361 470332 358373
rect 470356 358361 470412 358373
rect 470436 358361 470492 358373
rect 470516 358361 470572 358373
rect 470596 358361 470652 358373
rect 470676 358361 470732 358373
rect 470756 358361 470812 358373
rect 470276 358347 470314 358361
rect 470314 358347 470326 358361
rect 470326 358347 470332 358361
rect 470356 358347 470378 358361
rect 470378 358347 470390 358361
rect 470390 358347 470412 358361
rect 470436 358347 470442 358361
rect 470442 358347 470454 358361
rect 470454 358347 470492 358361
rect 470516 358347 470518 358361
rect 470518 358347 470570 358361
rect 470570 358347 470572 358361
rect 470596 358347 470634 358361
rect 470634 358347 470646 358361
rect 470646 358347 470652 358361
rect 470676 358347 470698 358361
rect 470698 358347 470710 358361
rect 470710 358347 470732 358361
rect 470756 358347 470762 358361
rect 470762 358347 470774 358361
rect 470774 358347 470812 358361
rect 470276 358309 470314 358323
rect 470314 358309 470326 358323
rect 470326 358309 470332 358323
rect 470356 358309 470378 358323
rect 470378 358309 470390 358323
rect 470390 358309 470412 358323
rect 470436 358309 470442 358323
rect 470442 358309 470454 358323
rect 470454 358309 470492 358323
rect 470516 358309 470518 358323
rect 470518 358309 470570 358323
rect 470570 358309 470572 358323
rect 470596 358309 470634 358323
rect 470634 358309 470646 358323
rect 470646 358309 470652 358323
rect 470676 358309 470698 358323
rect 470698 358309 470710 358323
rect 470710 358309 470732 358323
rect 470756 358309 470762 358323
rect 470762 358309 470774 358323
rect 470774 358309 470812 358323
rect 470276 358297 470332 358309
rect 470356 358297 470412 358309
rect 470436 358297 470492 358309
rect 470516 358297 470572 358309
rect 470596 358297 470652 358309
rect 470676 358297 470732 358309
rect 470756 358297 470812 358309
rect 470276 358267 470314 358297
rect 470314 358267 470326 358297
rect 470326 358267 470332 358297
rect 470356 358267 470378 358297
rect 470378 358267 470390 358297
rect 470390 358267 470412 358297
rect 470436 358267 470442 358297
rect 470442 358267 470454 358297
rect 470454 358267 470492 358297
rect 470516 358267 470518 358297
rect 470518 358267 470570 358297
rect 470570 358267 470572 358297
rect 470596 358267 470634 358297
rect 470634 358267 470646 358297
rect 470646 358267 470652 358297
rect 470676 358267 470698 358297
rect 470698 358267 470710 358297
rect 470710 358267 470732 358297
rect 470756 358267 470762 358297
rect 470762 358267 470774 358297
rect 470774 358267 470812 358297
rect 470276 358233 470332 358243
rect 470356 358233 470412 358243
rect 470436 358233 470492 358243
rect 470516 358233 470572 358243
rect 470596 358233 470652 358243
rect 470676 358233 470732 358243
rect 470756 358233 470812 358243
rect 470276 358187 470314 358233
rect 470314 358187 470326 358233
rect 470326 358187 470332 358233
rect 470356 358187 470378 358233
rect 470378 358187 470390 358233
rect 470390 358187 470412 358233
rect 470436 358187 470442 358233
rect 470442 358187 470454 358233
rect 470454 358187 470492 358233
rect 470516 358187 470518 358233
rect 470518 358187 470570 358233
rect 470570 358187 470572 358233
rect 470596 358187 470634 358233
rect 470634 358187 470646 358233
rect 470646 358187 470652 358233
rect 470676 358187 470698 358233
rect 470698 358187 470710 358233
rect 470710 358187 470732 358233
rect 470756 358187 470762 358233
rect 470762 358187 470774 358233
rect 470774 358187 470812 358233
rect 474922 389274 474978 389330
rect 478634 389274 478690 389330
rect 482098 389410 482154 389466
rect 489366 389410 489422 389466
rect 486882 386418 486938 386474
rect 478878 357994 478934 358050
rect 481822 357994 481878 358050
rect 484950 357994 485006 358050
rect 488446 357994 488502 358050
rect 469036 357351 469074 357397
rect 469074 357351 469086 357397
rect 469086 357351 469092 357397
rect 469116 357351 469138 357397
rect 469138 357351 469150 357397
rect 469150 357351 469172 357397
rect 469196 357351 469202 357397
rect 469202 357351 469214 357397
rect 469214 357351 469252 357397
rect 469276 357351 469278 357397
rect 469278 357351 469330 357397
rect 469330 357351 469332 357397
rect 469356 357351 469394 357397
rect 469394 357351 469406 357397
rect 469406 357351 469412 357397
rect 469436 357351 469458 357397
rect 469458 357351 469470 357397
rect 469470 357351 469492 357397
rect 469516 357351 469522 357397
rect 469522 357351 469534 357397
rect 469534 357351 469572 357397
rect 469036 357341 469092 357351
rect 469116 357341 469172 357351
rect 469196 357341 469252 357351
rect 469276 357341 469332 357351
rect 469356 357341 469412 357351
rect 469436 357341 469492 357351
rect 469516 357341 469572 357351
rect 469036 357287 469074 357317
rect 469074 357287 469086 357317
rect 469086 357287 469092 357317
rect 469116 357287 469138 357317
rect 469138 357287 469150 357317
rect 469150 357287 469172 357317
rect 469196 357287 469202 357317
rect 469202 357287 469214 357317
rect 469214 357287 469252 357317
rect 469276 357287 469278 357317
rect 469278 357287 469330 357317
rect 469330 357287 469332 357317
rect 469356 357287 469394 357317
rect 469394 357287 469406 357317
rect 469406 357287 469412 357317
rect 469436 357287 469458 357317
rect 469458 357287 469470 357317
rect 469470 357287 469492 357317
rect 469516 357287 469522 357317
rect 469522 357287 469534 357317
rect 469534 357287 469572 357317
rect 469036 357275 469092 357287
rect 469116 357275 469172 357287
rect 469196 357275 469252 357287
rect 469276 357275 469332 357287
rect 469356 357275 469412 357287
rect 469436 357275 469492 357287
rect 469516 357275 469572 357287
rect 469036 357261 469074 357275
rect 469074 357261 469086 357275
rect 469086 357261 469092 357275
rect 469116 357261 469138 357275
rect 469138 357261 469150 357275
rect 469150 357261 469172 357275
rect 469196 357261 469202 357275
rect 469202 357261 469214 357275
rect 469214 357261 469252 357275
rect 469276 357261 469278 357275
rect 469278 357261 469330 357275
rect 469330 357261 469332 357275
rect 469356 357261 469394 357275
rect 469394 357261 469406 357275
rect 469406 357261 469412 357275
rect 469436 357261 469458 357275
rect 469458 357261 469470 357275
rect 469470 357261 469492 357275
rect 469516 357261 469522 357275
rect 469522 357261 469534 357275
rect 469534 357261 469572 357275
rect 469036 357223 469074 357237
rect 469074 357223 469086 357237
rect 469086 357223 469092 357237
rect 469116 357223 469138 357237
rect 469138 357223 469150 357237
rect 469150 357223 469172 357237
rect 469196 357223 469202 357237
rect 469202 357223 469214 357237
rect 469214 357223 469252 357237
rect 469276 357223 469278 357237
rect 469278 357223 469330 357237
rect 469330 357223 469332 357237
rect 469356 357223 469394 357237
rect 469394 357223 469406 357237
rect 469406 357223 469412 357237
rect 469436 357223 469458 357237
rect 469458 357223 469470 357237
rect 469470 357223 469492 357237
rect 469516 357223 469522 357237
rect 469522 357223 469534 357237
rect 469534 357223 469572 357237
rect 469036 357211 469092 357223
rect 469116 357211 469172 357223
rect 469196 357211 469252 357223
rect 469276 357211 469332 357223
rect 469356 357211 469412 357223
rect 469436 357211 469492 357223
rect 469516 357211 469572 357223
rect 469036 357181 469074 357211
rect 469074 357181 469086 357211
rect 469086 357181 469092 357211
rect 469116 357181 469138 357211
rect 469138 357181 469150 357211
rect 469150 357181 469172 357211
rect 469196 357181 469202 357211
rect 469202 357181 469214 357211
rect 469214 357181 469252 357211
rect 469276 357181 469278 357211
rect 469278 357181 469330 357211
rect 469330 357181 469332 357211
rect 469356 357181 469394 357211
rect 469394 357181 469406 357211
rect 469406 357181 469412 357211
rect 469436 357181 469458 357211
rect 469458 357181 469470 357211
rect 469470 357181 469492 357211
rect 469516 357181 469522 357211
rect 469522 357181 469534 357211
rect 469534 357181 469572 357211
rect 469036 357147 469092 357157
rect 469116 357147 469172 357157
rect 469196 357147 469252 357157
rect 469276 357147 469332 357157
rect 469356 357147 469412 357157
rect 469436 357147 469492 357157
rect 469516 357147 469572 357157
rect 469036 357101 469074 357147
rect 469074 357101 469086 357147
rect 469086 357101 469092 357147
rect 469116 357101 469138 357147
rect 469138 357101 469150 357147
rect 469150 357101 469172 357147
rect 469196 357101 469202 357147
rect 469202 357101 469214 357147
rect 469214 357101 469252 357147
rect 469276 357101 469278 357147
rect 469278 357101 469330 357147
rect 469330 357101 469332 357147
rect 469356 357101 469394 357147
rect 469394 357101 469406 357147
rect 469406 357101 469412 357147
rect 469436 357101 469458 357147
rect 469458 357101 469470 357147
rect 469470 357101 469492 357147
rect 469516 357101 469522 357147
rect 469522 357101 469534 357147
rect 469534 357101 469572 357147
rect 470276 356264 470314 356310
rect 470314 356264 470326 356310
rect 470326 356264 470332 356310
rect 470356 356264 470378 356310
rect 470378 356264 470390 356310
rect 470390 356264 470412 356310
rect 470436 356264 470442 356310
rect 470442 356264 470454 356310
rect 470454 356264 470492 356310
rect 470516 356264 470518 356310
rect 470518 356264 470570 356310
rect 470570 356264 470572 356310
rect 470596 356264 470634 356310
rect 470634 356264 470646 356310
rect 470646 356264 470652 356310
rect 470676 356264 470698 356310
rect 470698 356264 470710 356310
rect 470710 356264 470732 356310
rect 470756 356264 470762 356310
rect 470762 356264 470774 356310
rect 470774 356264 470812 356310
rect 470276 356254 470332 356264
rect 470356 356254 470412 356264
rect 470436 356254 470492 356264
rect 470516 356254 470572 356264
rect 470596 356254 470652 356264
rect 470676 356254 470732 356264
rect 470756 356254 470812 356264
rect 470276 356200 470314 356230
rect 470314 356200 470326 356230
rect 470326 356200 470332 356230
rect 470356 356200 470378 356230
rect 470378 356200 470390 356230
rect 470390 356200 470412 356230
rect 470436 356200 470442 356230
rect 470442 356200 470454 356230
rect 470454 356200 470492 356230
rect 470516 356200 470518 356230
rect 470518 356200 470570 356230
rect 470570 356200 470572 356230
rect 470596 356200 470634 356230
rect 470634 356200 470646 356230
rect 470646 356200 470652 356230
rect 470676 356200 470698 356230
rect 470698 356200 470710 356230
rect 470710 356200 470732 356230
rect 470756 356200 470762 356230
rect 470762 356200 470774 356230
rect 470774 356200 470812 356230
rect 470276 356188 470332 356200
rect 470356 356188 470412 356200
rect 470436 356188 470492 356200
rect 470516 356188 470572 356200
rect 470596 356188 470652 356200
rect 470676 356188 470732 356200
rect 470756 356188 470812 356200
rect 470276 356174 470314 356188
rect 470314 356174 470326 356188
rect 470326 356174 470332 356188
rect 470356 356174 470378 356188
rect 470378 356174 470390 356188
rect 470390 356174 470412 356188
rect 470436 356174 470442 356188
rect 470442 356174 470454 356188
rect 470454 356174 470492 356188
rect 470516 356174 470518 356188
rect 470518 356174 470570 356188
rect 470570 356174 470572 356188
rect 470596 356174 470634 356188
rect 470634 356174 470646 356188
rect 470646 356174 470652 356188
rect 470676 356174 470698 356188
rect 470698 356174 470710 356188
rect 470710 356174 470732 356188
rect 470756 356174 470762 356188
rect 470762 356174 470774 356188
rect 470774 356174 470812 356188
rect 470276 356136 470314 356150
rect 470314 356136 470326 356150
rect 470326 356136 470332 356150
rect 470356 356136 470378 356150
rect 470378 356136 470390 356150
rect 470390 356136 470412 356150
rect 470436 356136 470442 356150
rect 470442 356136 470454 356150
rect 470454 356136 470492 356150
rect 470516 356136 470518 356150
rect 470518 356136 470570 356150
rect 470570 356136 470572 356150
rect 470596 356136 470634 356150
rect 470634 356136 470646 356150
rect 470646 356136 470652 356150
rect 470676 356136 470698 356150
rect 470698 356136 470710 356150
rect 470710 356136 470732 356150
rect 470756 356136 470762 356150
rect 470762 356136 470774 356150
rect 470774 356136 470812 356150
rect 470276 356124 470332 356136
rect 470356 356124 470412 356136
rect 470436 356124 470492 356136
rect 470516 356124 470572 356136
rect 470596 356124 470652 356136
rect 470676 356124 470732 356136
rect 470756 356124 470812 356136
rect 470276 356094 470314 356124
rect 470314 356094 470326 356124
rect 470326 356094 470332 356124
rect 470356 356094 470378 356124
rect 470378 356094 470390 356124
rect 470390 356094 470412 356124
rect 470436 356094 470442 356124
rect 470442 356094 470454 356124
rect 470454 356094 470492 356124
rect 470516 356094 470518 356124
rect 470518 356094 470570 356124
rect 470570 356094 470572 356124
rect 470596 356094 470634 356124
rect 470634 356094 470646 356124
rect 470646 356094 470652 356124
rect 470676 356094 470698 356124
rect 470698 356094 470710 356124
rect 470710 356094 470732 356124
rect 470756 356094 470762 356124
rect 470762 356094 470774 356124
rect 470774 356094 470812 356124
rect 470276 356060 470332 356070
rect 470356 356060 470412 356070
rect 470436 356060 470492 356070
rect 470516 356060 470572 356070
rect 470596 356060 470652 356070
rect 470676 356060 470732 356070
rect 470756 356060 470812 356070
rect 470276 356014 470314 356060
rect 470314 356014 470326 356060
rect 470326 356014 470332 356060
rect 470356 356014 470378 356060
rect 470378 356014 470390 356060
rect 470390 356014 470412 356060
rect 470436 356014 470442 356060
rect 470442 356014 470454 356060
rect 470454 356014 470492 356060
rect 470516 356014 470518 356060
rect 470518 356014 470570 356060
rect 470570 356014 470572 356060
rect 470596 356014 470634 356060
rect 470634 356014 470646 356060
rect 470646 356014 470652 356060
rect 470676 356014 470698 356060
rect 470698 356014 470710 356060
rect 470710 356014 470732 356060
rect 470756 356014 470762 356060
rect 470762 356014 470774 356060
rect 470774 356014 470812 356060
rect 475014 357450 475070 357506
rect 484582 351874 484638 351930
rect 470276 342436 470314 342482
rect 470314 342436 470326 342482
rect 470326 342436 470332 342482
rect 470356 342436 470378 342482
rect 470378 342436 470390 342482
rect 470390 342436 470412 342482
rect 470436 342436 470442 342482
rect 470442 342436 470454 342482
rect 470454 342436 470492 342482
rect 470516 342436 470518 342482
rect 470518 342436 470570 342482
rect 470570 342436 470572 342482
rect 470596 342436 470634 342482
rect 470634 342436 470646 342482
rect 470646 342436 470652 342482
rect 470676 342436 470698 342482
rect 470698 342436 470710 342482
rect 470710 342436 470732 342482
rect 470756 342436 470762 342482
rect 470762 342436 470774 342482
rect 470774 342436 470812 342482
rect 470276 342426 470332 342436
rect 470356 342426 470412 342436
rect 470436 342426 470492 342436
rect 470516 342426 470572 342436
rect 470596 342426 470652 342436
rect 470676 342426 470732 342436
rect 470756 342426 470812 342436
rect 470276 342372 470314 342402
rect 470314 342372 470326 342402
rect 470326 342372 470332 342402
rect 470356 342372 470378 342402
rect 470378 342372 470390 342402
rect 470390 342372 470412 342402
rect 470436 342372 470442 342402
rect 470442 342372 470454 342402
rect 470454 342372 470492 342402
rect 470516 342372 470518 342402
rect 470518 342372 470570 342402
rect 470570 342372 470572 342402
rect 470596 342372 470634 342402
rect 470634 342372 470646 342402
rect 470646 342372 470652 342402
rect 470676 342372 470698 342402
rect 470698 342372 470710 342402
rect 470710 342372 470732 342402
rect 470756 342372 470762 342402
rect 470762 342372 470774 342402
rect 470774 342372 470812 342402
rect 470276 342360 470332 342372
rect 470356 342360 470412 342372
rect 470436 342360 470492 342372
rect 470516 342360 470572 342372
rect 470596 342360 470652 342372
rect 470676 342360 470732 342372
rect 470756 342360 470812 342372
rect 470276 342346 470314 342360
rect 470314 342346 470326 342360
rect 470326 342346 470332 342360
rect 470356 342346 470378 342360
rect 470378 342346 470390 342360
rect 470390 342346 470412 342360
rect 470436 342346 470442 342360
rect 470442 342346 470454 342360
rect 470454 342346 470492 342360
rect 470516 342346 470518 342360
rect 470518 342346 470570 342360
rect 470570 342346 470572 342360
rect 470596 342346 470634 342360
rect 470634 342346 470646 342360
rect 470646 342346 470652 342360
rect 470676 342346 470698 342360
rect 470698 342346 470710 342360
rect 470710 342346 470732 342360
rect 470756 342346 470762 342360
rect 470762 342346 470774 342360
rect 470774 342346 470812 342360
rect 470276 342308 470314 342322
rect 470314 342308 470326 342322
rect 470326 342308 470332 342322
rect 470356 342308 470378 342322
rect 470378 342308 470390 342322
rect 470390 342308 470412 342322
rect 470436 342308 470442 342322
rect 470442 342308 470454 342322
rect 470454 342308 470492 342322
rect 470516 342308 470518 342322
rect 470518 342308 470570 342322
rect 470570 342308 470572 342322
rect 470596 342308 470634 342322
rect 470634 342308 470646 342322
rect 470646 342308 470652 342322
rect 470676 342308 470698 342322
rect 470698 342308 470710 342322
rect 470710 342308 470732 342322
rect 470756 342308 470762 342322
rect 470762 342308 470774 342322
rect 470774 342308 470812 342322
rect 470276 342296 470332 342308
rect 470356 342296 470412 342308
rect 470436 342296 470492 342308
rect 470516 342296 470572 342308
rect 470596 342296 470652 342308
rect 470676 342296 470732 342308
rect 470756 342296 470812 342308
rect 470276 342266 470314 342296
rect 470314 342266 470326 342296
rect 470326 342266 470332 342296
rect 470356 342266 470378 342296
rect 470378 342266 470390 342296
rect 470390 342266 470412 342296
rect 470436 342266 470442 342296
rect 470442 342266 470454 342296
rect 470454 342266 470492 342296
rect 470516 342266 470518 342296
rect 470518 342266 470570 342296
rect 470570 342266 470572 342296
rect 470596 342266 470634 342296
rect 470634 342266 470646 342296
rect 470646 342266 470652 342296
rect 470676 342266 470698 342296
rect 470698 342266 470710 342296
rect 470710 342266 470732 342296
rect 470756 342266 470762 342296
rect 470762 342266 470774 342296
rect 470774 342266 470812 342296
rect 470276 342232 470332 342242
rect 470356 342232 470412 342242
rect 470436 342232 470492 342242
rect 470516 342232 470572 342242
rect 470596 342232 470652 342242
rect 470676 342232 470732 342242
rect 470756 342232 470812 342242
rect 470276 342186 470314 342232
rect 470314 342186 470326 342232
rect 470326 342186 470332 342232
rect 470356 342186 470378 342232
rect 470378 342186 470390 342232
rect 470390 342186 470412 342232
rect 470436 342186 470442 342232
rect 470442 342186 470454 342232
rect 470454 342186 470492 342232
rect 470516 342186 470518 342232
rect 470518 342186 470570 342232
rect 470570 342186 470572 342232
rect 470596 342186 470634 342232
rect 470634 342186 470646 342232
rect 470646 342186 470652 342232
rect 470676 342186 470698 342232
rect 470698 342186 470710 342232
rect 470710 342186 470732 342232
rect 470756 342186 470762 342232
rect 470762 342186 470774 342232
rect 470774 342186 470812 342232
rect 484582 342218 484638 342274
rect 469036 341349 469074 341395
rect 469074 341349 469086 341395
rect 469086 341349 469092 341395
rect 469116 341349 469138 341395
rect 469138 341349 469150 341395
rect 469150 341349 469172 341395
rect 469196 341349 469202 341395
rect 469202 341349 469214 341395
rect 469214 341349 469252 341395
rect 469276 341349 469278 341395
rect 469278 341349 469330 341395
rect 469330 341349 469332 341395
rect 469356 341349 469394 341395
rect 469394 341349 469406 341395
rect 469406 341349 469412 341395
rect 469436 341349 469458 341395
rect 469458 341349 469470 341395
rect 469470 341349 469492 341395
rect 469516 341349 469522 341395
rect 469522 341349 469534 341395
rect 469534 341349 469572 341395
rect 469036 341339 469092 341349
rect 469116 341339 469172 341349
rect 469196 341339 469252 341349
rect 469276 341339 469332 341349
rect 469356 341339 469412 341349
rect 469436 341339 469492 341349
rect 469516 341339 469572 341349
rect 469036 341285 469074 341315
rect 469074 341285 469086 341315
rect 469086 341285 469092 341315
rect 469116 341285 469138 341315
rect 469138 341285 469150 341315
rect 469150 341285 469172 341315
rect 469196 341285 469202 341315
rect 469202 341285 469214 341315
rect 469214 341285 469252 341315
rect 469276 341285 469278 341315
rect 469278 341285 469330 341315
rect 469330 341285 469332 341315
rect 469356 341285 469394 341315
rect 469394 341285 469406 341315
rect 469406 341285 469412 341315
rect 469436 341285 469458 341315
rect 469458 341285 469470 341315
rect 469470 341285 469492 341315
rect 469516 341285 469522 341315
rect 469522 341285 469534 341315
rect 469534 341285 469572 341315
rect 469036 341273 469092 341285
rect 469116 341273 469172 341285
rect 469196 341273 469252 341285
rect 469276 341273 469332 341285
rect 469356 341273 469412 341285
rect 469436 341273 469492 341285
rect 469516 341273 469572 341285
rect 469036 341259 469074 341273
rect 469074 341259 469086 341273
rect 469086 341259 469092 341273
rect 469116 341259 469138 341273
rect 469138 341259 469150 341273
rect 469150 341259 469172 341273
rect 469196 341259 469202 341273
rect 469202 341259 469214 341273
rect 469214 341259 469252 341273
rect 469276 341259 469278 341273
rect 469278 341259 469330 341273
rect 469330 341259 469332 341273
rect 469356 341259 469394 341273
rect 469394 341259 469406 341273
rect 469406 341259 469412 341273
rect 469436 341259 469458 341273
rect 469458 341259 469470 341273
rect 469470 341259 469492 341273
rect 469516 341259 469522 341273
rect 469522 341259 469534 341273
rect 469534 341259 469572 341273
rect 469036 341221 469074 341235
rect 469074 341221 469086 341235
rect 469086 341221 469092 341235
rect 469116 341221 469138 341235
rect 469138 341221 469150 341235
rect 469150 341221 469172 341235
rect 469196 341221 469202 341235
rect 469202 341221 469214 341235
rect 469214 341221 469252 341235
rect 469276 341221 469278 341235
rect 469278 341221 469330 341235
rect 469330 341221 469332 341235
rect 469356 341221 469394 341235
rect 469394 341221 469406 341235
rect 469406 341221 469412 341235
rect 469436 341221 469458 341235
rect 469458 341221 469470 341235
rect 469470 341221 469492 341235
rect 469516 341221 469522 341235
rect 469522 341221 469534 341235
rect 469534 341221 469572 341235
rect 469036 341209 469092 341221
rect 469116 341209 469172 341221
rect 469196 341209 469252 341221
rect 469276 341209 469332 341221
rect 469356 341209 469412 341221
rect 469436 341209 469492 341221
rect 469516 341209 469572 341221
rect 469036 341179 469074 341209
rect 469074 341179 469086 341209
rect 469086 341179 469092 341209
rect 469116 341179 469138 341209
rect 469138 341179 469150 341209
rect 469150 341179 469172 341209
rect 469196 341179 469202 341209
rect 469202 341179 469214 341209
rect 469214 341179 469252 341209
rect 469276 341179 469278 341209
rect 469278 341179 469330 341209
rect 469330 341179 469332 341209
rect 469356 341179 469394 341209
rect 469394 341179 469406 341209
rect 469406 341179 469412 341209
rect 469436 341179 469458 341209
rect 469458 341179 469470 341209
rect 469470 341179 469492 341209
rect 469516 341179 469522 341209
rect 469522 341179 469534 341209
rect 469534 341179 469572 341209
rect 469036 341145 469092 341155
rect 469116 341145 469172 341155
rect 469196 341145 469252 341155
rect 469276 341145 469332 341155
rect 469356 341145 469412 341155
rect 469436 341145 469492 341155
rect 469516 341145 469572 341155
rect 469036 341099 469074 341145
rect 469074 341099 469086 341145
rect 469086 341099 469092 341145
rect 469116 341099 469138 341145
rect 469138 341099 469150 341145
rect 469150 341099 469172 341145
rect 469196 341099 469202 341145
rect 469202 341099 469214 341145
rect 469214 341099 469252 341145
rect 469276 341099 469278 341145
rect 469278 341099 469330 341145
rect 469330 341099 469332 341145
rect 469356 341099 469394 341145
rect 469394 341099 469406 341145
rect 469406 341099 469412 341145
rect 469436 341099 469458 341145
rect 469458 341099 469470 341145
rect 469470 341099 469492 341145
rect 469516 341099 469522 341145
rect 469522 341099 469534 341145
rect 469534 341099 469572 341145
rect 470276 340264 470314 340310
rect 470314 340264 470326 340310
rect 470326 340264 470332 340310
rect 470356 340264 470378 340310
rect 470378 340264 470390 340310
rect 470390 340264 470412 340310
rect 470436 340264 470442 340310
rect 470442 340264 470454 340310
rect 470454 340264 470492 340310
rect 470516 340264 470518 340310
rect 470518 340264 470570 340310
rect 470570 340264 470572 340310
rect 470596 340264 470634 340310
rect 470634 340264 470646 340310
rect 470646 340264 470652 340310
rect 470676 340264 470698 340310
rect 470698 340264 470710 340310
rect 470710 340264 470732 340310
rect 470756 340264 470762 340310
rect 470762 340264 470774 340310
rect 470774 340264 470812 340310
rect 470276 340254 470332 340264
rect 470356 340254 470412 340264
rect 470436 340254 470492 340264
rect 470516 340254 470572 340264
rect 470596 340254 470652 340264
rect 470676 340254 470732 340264
rect 470756 340254 470812 340264
rect 470276 340200 470314 340230
rect 470314 340200 470326 340230
rect 470326 340200 470332 340230
rect 470356 340200 470378 340230
rect 470378 340200 470390 340230
rect 470390 340200 470412 340230
rect 470436 340200 470442 340230
rect 470442 340200 470454 340230
rect 470454 340200 470492 340230
rect 470516 340200 470518 340230
rect 470518 340200 470570 340230
rect 470570 340200 470572 340230
rect 470596 340200 470634 340230
rect 470634 340200 470646 340230
rect 470646 340200 470652 340230
rect 470676 340200 470698 340230
rect 470698 340200 470710 340230
rect 470710 340200 470732 340230
rect 470756 340200 470762 340230
rect 470762 340200 470774 340230
rect 470774 340200 470812 340230
rect 470276 340188 470332 340200
rect 470356 340188 470412 340200
rect 470436 340188 470492 340200
rect 470516 340188 470572 340200
rect 470596 340188 470652 340200
rect 470676 340188 470732 340200
rect 470756 340188 470812 340200
rect 470276 340174 470314 340188
rect 470314 340174 470326 340188
rect 470326 340174 470332 340188
rect 470356 340174 470378 340188
rect 470378 340174 470390 340188
rect 470390 340174 470412 340188
rect 470436 340174 470442 340188
rect 470442 340174 470454 340188
rect 470454 340174 470492 340188
rect 470516 340174 470518 340188
rect 470518 340174 470570 340188
rect 470570 340174 470572 340188
rect 470596 340174 470634 340188
rect 470634 340174 470646 340188
rect 470646 340174 470652 340188
rect 470676 340174 470698 340188
rect 470698 340174 470710 340188
rect 470710 340174 470732 340188
rect 470756 340174 470762 340188
rect 470762 340174 470774 340188
rect 470774 340174 470812 340188
rect 470276 340136 470314 340150
rect 470314 340136 470326 340150
rect 470326 340136 470332 340150
rect 470356 340136 470378 340150
rect 470378 340136 470390 340150
rect 470390 340136 470412 340150
rect 470436 340136 470442 340150
rect 470442 340136 470454 340150
rect 470454 340136 470492 340150
rect 470516 340136 470518 340150
rect 470518 340136 470570 340150
rect 470570 340136 470572 340150
rect 470596 340136 470634 340150
rect 470634 340136 470646 340150
rect 470646 340136 470652 340150
rect 470676 340136 470698 340150
rect 470698 340136 470710 340150
rect 470710 340136 470732 340150
rect 470756 340136 470762 340150
rect 470762 340136 470774 340150
rect 470774 340136 470812 340150
rect 470276 340124 470332 340136
rect 470356 340124 470412 340136
rect 470436 340124 470492 340136
rect 470516 340124 470572 340136
rect 470596 340124 470652 340136
rect 470676 340124 470732 340136
rect 470756 340124 470812 340136
rect 470276 340094 470314 340124
rect 470314 340094 470326 340124
rect 470326 340094 470332 340124
rect 470356 340094 470378 340124
rect 470378 340094 470390 340124
rect 470390 340094 470412 340124
rect 470436 340094 470442 340124
rect 470442 340094 470454 340124
rect 470454 340094 470492 340124
rect 470516 340094 470518 340124
rect 470518 340094 470570 340124
rect 470570 340094 470572 340124
rect 470596 340094 470634 340124
rect 470634 340094 470646 340124
rect 470646 340094 470652 340124
rect 470676 340094 470698 340124
rect 470698 340094 470710 340124
rect 470710 340094 470732 340124
rect 470756 340094 470762 340124
rect 470762 340094 470774 340124
rect 470774 340094 470812 340124
rect 470276 340060 470332 340070
rect 470356 340060 470412 340070
rect 470436 340060 470492 340070
rect 470516 340060 470572 340070
rect 470596 340060 470652 340070
rect 470676 340060 470732 340070
rect 470756 340060 470812 340070
rect 470276 340014 470314 340060
rect 470314 340014 470326 340060
rect 470326 340014 470332 340060
rect 470356 340014 470378 340060
rect 470378 340014 470390 340060
rect 470390 340014 470412 340060
rect 470436 340014 470442 340060
rect 470442 340014 470454 340060
rect 470454 340014 470492 340060
rect 470516 340014 470518 340060
rect 470518 340014 470570 340060
rect 470570 340014 470572 340060
rect 470596 340014 470634 340060
rect 470634 340014 470646 340060
rect 470646 340014 470652 340060
rect 470676 340014 470698 340060
rect 470698 340014 470710 340060
rect 470710 340014 470732 340060
rect 470756 340014 470762 340060
rect 470762 340014 470774 340060
rect 470774 340014 470812 340060
rect 470276 322436 470314 322482
rect 470314 322436 470326 322482
rect 470326 322436 470332 322482
rect 470356 322436 470378 322482
rect 470378 322436 470390 322482
rect 470390 322436 470412 322482
rect 470436 322436 470442 322482
rect 470442 322436 470454 322482
rect 470454 322436 470492 322482
rect 470516 322436 470518 322482
rect 470518 322436 470570 322482
rect 470570 322436 470572 322482
rect 470596 322436 470634 322482
rect 470634 322436 470646 322482
rect 470646 322436 470652 322482
rect 470676 322436 470698 322482
rect 470698 322436 470710 322482
rect 470710 322436 470732 322482
rect 470756 322436 470762 322482
rect 470762 322436 470774 322482
rect 470774 322436 470812 322482
rect 470276 322426 470332 322436
rect 470356 322426 470412 322436
rect 470436 322426 470492 322436
rect 470516 322426 470572 322436
rect 470596 322426 470652 322436
rect 470676 322426 470732 322436
rect 470756 322426 470812 322436
rect 470276 322372 470314 322402
rect 470314 322372 470326 322402
rect 470326 322372 470332 322402
rect 470356 322372 470378 322402
rect 470378 322372 470390 322402
rect 470390 322372 470412 322402
rect 470436 322372 470442 322402
rect 470442 322372 470454 322402
rect 470454 322372 470492 322402
rect 470516 322372 470518 322402
rect 470518 322372 470570 322402
rect 470570 322372 470572 322402
rect 470596 322372 470634 322402
rect 470634 322372 470646 322402
rect 470646 322372 470652 322402
rect 470676 322372 470698 322402
rect 470698 322372 470710 322402
rect 470710 322372 470732 322402
rect 470756 322372 470762 322402
rect 470762 322372 470774 322402
rect 470774 322372 470812 322402
rect 470276 322360 470332 322372
rect 470356 322360 470412 322372
rect 470436 322360 470492 322372
rect 470516 322360 470572 322372
rect 470596 322360 470652 322372
rect 470676 322360 470732 322372
rect 470756 322360 470812 322372
rect 470276 322346 470314 322360
rect 470314 322346 470326 322360
rect 470326 322346 470332 322360
rect 470356 322346 470378 322360
rect 470378 322346 470390 322360
rect 470390 322346 470412 322360
rect 470436 322346 470442 322360
rect 470442 322346 470454 322360
rect 470454 322346 470492 322360
rect 470516 322346 470518 322360
rect 470518 322346 470570 322360
rect 470570 322346 470572 322360
rect 470596 322346 470634 322360
rect 470634 322346 470646 322360
rect 470646 322346 470652 322360
rect 470676 322346 470698 322360
rect 470698 322346 470710 322360
rect 470710 322346 470732 322360
rect 470756 322346 470762 322360
rect 470762 322346 470774 322360
rect 470774 322346 470812 322360
rect 470276 322308 470314 322322
rect 470314 322308 470326 322322
rect 470326 322308 470332 322322
rect 470356 322308 470378 322322
rect 470378 322308 470390 322322
rect 470390 322308 470412 322322
rect 470436 322308 470442 322322
rect 470442 322308 470454 322322
rect 470454 322308 470492 322322
rect 470516 322308 470518 322322
rect 470518 322308 470570 322322
rect 470570 322308 470572 322322
rect 470596 322308 470634 322322
rect 470634 322308 470646 322322
rect 470646 322308 470652 322322
rect 470676 322308 470698 322322
rect 470698 322308 470710 322322
rect 470710 322308 470732 322322
rect 470756 322308 470762 322322
rect 470762 322308 470774 322322
rect 470774 322308 470812 322322
rect 470276 322296 470332 322308
rect 470356 322296 470412 322308
rect 470436 322296 470492 322308
rect 470516 322296 470572 322308
rect 470596 322296 470652 322308
rect 470676 322296 470732 322308
rect 470756 322296 470812 322308
rect 470276 322266 470314 322296
rect 470314 322266 470326 322296
rect 470326 322266 470332 322296
rect 470356 322266 470378 322296
rect 470378 322266 470390 322296
rect 470390 322266 470412 322296
rect 470436 322266 470442 322296
rect 470442 322266 470454 322296
rect 470454 322266 470492 322296
rect 470516 322266 470518 322296
rect 470518 322266 470570 322296
rect 470570 322266 470572 322296
rect 470596 322266 470634 322296
rect 470634 322266 470646 322296
rect 470646 322266 470652 322296
rect 470676 322266 470698 322296
rect 470698 322266 470710 322296
rect 470710 322266 470732 322296
rect 470756 322266 470762 322296
rect 470762 322266 470774 322296
rect 470774 322266 470812 322296
rect 470276 322232 470332 322242
rect 470356 322232 470412 322242
rect 470436 322232 470492 322242
rect 470516 322232 470572 322242
rect 470596 322232 470652 322242
rect 470676 322232 470732 322242
rect 470756 322232 470812 322242
rect 470276 322186 470314 322232
rect 470314 322186 470326 322232
rect 470326 322186 470332 322232
rect 470356 322186 470378 322232
rect 470378 322186 470390 322232
rect 470390 322186 470412 322232
rect 470436 322186 470442 322232
rect 470442 322186 470454 322232
rect 470454 322186 470492 322232
rect 470516 322186 470518 322232
rect 470518 322186 470570 322232
rect 470570 322186 470572 322232
rect 470596 322186 470634 322232
rect 470634 322186 470646 322232
rect 470646 322186 470652 322232
rect 470676 322186 470698 322232
rect 470698 322186 470710 322232
rect 470710 322186 470732 322232
rect 470756 322186 470762 322232
rect 470762 322186 470774 322232
rect 470774 322186 470812 322232
rect 484398 341674 484454 341730
rect 477915 340994 477971 341050
rect 481232 340994 481288 341050
rect 487894 340994 487950 341050
rect 474554 340450 474610 340506
rect 484306 322090 484362 322146
rect 469036 321349 469074 321395
rect 469074 321349 469086 321395
rect 469086 321349 469092 321395
rect 469116 321349 469138 321395
rect 469138 321349 469150 321395
rect 469150 321349 469172 321395
rect 469196 321349 469202 321395
rect 469202 321349 469214 321395
rect 469214 321349 469252 321395
rect 469276 321349 469278 321395
rect 469278 321349 469330 321395
rect 469330 321349 469332 321395
rect 469356 321349 469394 321395
rect 469394 321349 469406 321395
rect 469406 321349 469412 321395
rect 469436 321349 469458 321395
rect 469458 321349 469470 321395
rect 469470 321349 469492 321395
rect 469516 321349 469522 321395
rect 469522 321349 469534 321395
rect 469534 321349 469572 321395
rect 469036 321339 469092 321349
rect 469116 321339 469172 321349
rect 469196 321339 469252 321349
rect 469276 321339 469332 321349
rect 469356 321339 469412 321349
rect 469436 321339 469492 321349
rect 469516 321339 469572 321349
rect 469036 321285 469074 321315
rect 469074 321285 469086 321315
rect 469086 321285 469092 321315
rect 469116 321285 469138 321315
rect 469138 321285 469150 321315
rect 469150 321285 469172 321315
rect 469196 321285 469202 321315
rect 469202 321285 469214 321315
rect 469214 321285 469252 321315
rect 469276 321285 469278 321315
rect 469278 321285 469330 321315
rect 469330 321285 469332 321315
rect 469356 321285 469394 321315
rect 469394 321285 469406 321315
rect 469406 321285 469412 321315
rect 469436 321285 469458 321315
rect 469458 321285 469470 321315
rect 469470 321285 469492 321315
rect 469516 321285 469522 321315
rect 469522 321285 469534 321315
rect 469534 321285 469572 321315
rect 469036 321273 469092 321285
rect 469116 321273 469172 321285
rect 469196 321273 469252 321285
rect 469276 321273 469332 321285
rect 469356 321273 469412 321285
rect 469436 321273 469492 321285
rect 469516 321273 469572 321285
rect 469036 321259 469074 321273
rect 469074 321259 469086 321273
rect 469086 321259 469092 321273
rect 469116 321259 469138 321273
rect 469138 321259 469150 321273
rect 469150 321259 469172 321273
rect 469196 321259 469202 321273
rect 469202 321259 469214 321273
rect 469214 321259 469252 321273
rect 469276 321259 469278 321273
rect 469278 321259 469330 321273
rect 469330 321259 469332 321273
rect 469356 321259 469394 321273
rect 469394 321259 469406 321273
rect 469406 321259 469412 321273
rect 469436 321259 469458 321273
rect 469458 321259 469470 321273
rect 469470 321259 469492 321273
rect 469516 321259 469522 321273
rect 469522 321259 469534 321273
rect 469534 321259 469572 321273
rect 469036 321221 469074 321235
rect 469074 321221 469086 321235
rect 469086 321221 469092 321235
rect 469116 321221 469138 321235
rect 469138 321221 469150 321235
rect 469150 321221 469172 321235
rect 469196 321221 469202 321235
rect 469202 321221 469214 321235
rect 469214 321221 469252 321235
rect 469276 321221 469278 321235
rect 469278 321221 469330 321235
rect 469330 321221 469332 321235
rect 469356 321221 469394 321235
rect 469394 321221 469406 321235
rect 469406 321221 469412 321235
rect 469436 321221 469458 321235
rect 469458 321221 469470 321235
rect 469470 321221 469492 321235
rect 469516 321221 469522 321235
rect 469522 321221 469534 321235
rect 469534 321221 469572 321235
rect 469036 321209 469092 321221
rect 469116 321209 469172 321221
rect 469196 321209 469252 321221
rect 469276 321209 469332 321221
rect 469356 321209 469412 321221
rect 469436 321209 469492 321221
rect 469516 321209 469572 321221
rect 469036 321179 469074 321209
rect 469074 321179 469086 321209
rect 469086 321179 469092 321209
rect 469116 321179 469138 321209
rect 469138 321179 469150 321209
rect 469150 321179 469172 321209
rect 469196 321179 469202 321209
rect 469202 321179 469214 321209
rect 469214 321179 469252 321209
rect 469276 321179 469278 321209
rect 469278 321179 469330 321209
rect 469330 321179 469332 321209
rect 469356 321179 469394 321209
rect 469394 321179 469406 321209
rect 469406 321179 469412 321209
rect 469436 321179 469458 321209
rect 469458 321179 469470 321209
rect 469470 321179 469492 321209
rect 469516 321179 469522 321209
rect 469522 321179 469534 321209
rect 469534 321179 469572 321209
rect 469036 321145 469092 321155
rect 469116 321145 469172 321155
rect 469196 321145 469252 321155
rect 469276 321145 469332 321155
rect 469356 321145 469412 321155
rect 469436 321145 469492 321155
rect 469516 321145 469572 321155
rect 469036 321099 469074 321145
rect 469074 321099 469086 321145
rect 469086 321099 469092 321145
rect 469116 321099 469138 321145
rect 469138 321099 469150 321145
rect 469150 321099 469172 321145
rect 469196 321099 469202 321145
rect 469202 321099 469214 321145
rect 469214 321099 469252 321145
rect 469276 321099 469278 321145
rect 469278 321099 469330 321145
rect 469330 321099 469332 321145
rect 469356 321099 469394 321145
rect 469394 321099 469406 321145
rect 469406 321099 469412 321145
rect 469436 321099 469458 321145
rect 469458 321099 469470 321145
rect 469470 321099 469492 321145
rect 469516 321099 469522 321145
rect 469522 321099 469534 321145
rect 469534 321099 469572 321145
rect 470276 320264 470314 320310
rect 470314 320264 470326 320310
rect 470326 320264 470332 320310
rect 470356 320264 470378 320310
rect 470378 320264 470390 320310
rect 470390 320264 470412 320310
rect 470436 320264 470442 320310
rect 470442 320264 470454 320310
rect 470454 320264 470492 320310
rect 470516 320264 470518 320310
rect 470518 320264 470570 320310
rect 470570 320264 470572 320310
rect 470596 320264 470634 320310
rect 470634 320264 470646 320310
rect 470646 320264 470652 320310
rect 470676 320264 470698 320310
rect 470698 320264 470710 320310
rect 470710 320264 470732 320310
rect 470756 320264 470762 320310
rect 470762 320264 470774 320310
rect 470774 320264 470812 320310
rect 470276 320254 470332 320264
rect 470356 320254 470412 320264
rect 470436 320254 470492 320264
rect 470516 320254 470572 320264
rect 470596 320254 470652 320264
rect 470676 320254 470732 320264
rect 470756 320254 470812 320264
rect 470276 320200 470314 320230
rect 470314 320200 470326 320230
rect 470326 320200 470332 320230
rect 470356 320200 470378 320230
rect 470378 320200 470390 320230
rect 470390 320200 470412 320230
rect 470436 320200 470442 320230
rect 470442 320200 470454 320230
rect 470454 320200 470492 320230
rect 470516 320200 470518 320230
rect 470518 320200 470570 320230
rect 470570 320200 470572 320230
rect 470596 320200 470634 320230
rect 470634 320200 470646 320230
rect 470646 320200 470652 320230
rect 470676 320200 470698 320230
rect 470698 320200 470710 320230
rect 470710 320200 470732 320230
rect 470756 320200 470762 320230
rect 470762 320200 470774 320230
rect 470774 320200 470812 320230
rect 470276 320188 470332 320200
rect 470356 320188 470412 320200
rect 470436 320188 470492 320200
rect 470516 320188 470572 320200
rect 470596 320188 470652 320200
rect 470676 320188 470732 320200
rect 470756 320188 470812 320200
rect 470276 320174 470314 320188
rect 470314 320174 470326 320188
rect 470326 320174 470332 320188
rect 470356 320174 470378 320188
rect 470378 320174 470390 320188
rect 470390 320174 470412 320188
rect 470436 320174 470442 320188
rect 470442 320174 470454 320188
rect 470454 320174 470492 320188
rect 470516 320174 470518 320188
rect 470518 320174 470570 320188
rect 470570 320174 470572 320188
rect 470596 320174 470634 320188
rect 470634 320174 470646 320188
rect 470646 320174 470652 320188
rect 470676 320174 470698 320188
rect 470698 320174 470710 320188
rect 470710 320174 470732 320188
rect 470756 320174 470762 320188
rect 470762 320174 470774 320188
rect 470774 320174 470812 320188
rect 470276 320136 470314 320150
rect 470314 320136 470326 320150
rect 470326 320136 470332 320150
rect 470356 320136 470378 320150
rect 470378 320136 470390 320150
rect 470390 320136 470412 320150
rect 470436 320136 470442 320150
rect 470442 320136 470454 320150
rect 470454 320136 470492 320150
rect 470516 320136 470518 320150
rect 470518 320136 470570 320150
rect 470570 320136 470572 320150
rect 470596 320136 470634 320150
rect 470634 320136 470646 320150
rect 470646 320136 470652 320150
rect 470676 320136 470698 320150
rect 470698 320136 470710 320150
rect 470710 320136 470732 320150
rect 470756 320136 470762 320150
rect 470762 320136 470774 320150
rect 470774 320136 470812 320150
rect 470276 320124 470332 320136
rect 470356 320124 470412 320136
rect 470436 320124 470492 320136
rect 470516 320124 470572 320136
rect 470596 320124 470652 320136
rect 470676 320124 470732 320136
rect 470756 320124 470812 320136
rect 470276 320094 470314 320124
rect 470314 320094 470326 320124
rect 470326 320094 470332 320124
rect 470356 320094 470378 320124
rect 470378 320094 470390 320124
rect 470390 320094 470412 320124
rect 470436 320094 470442 320124
rect 470442 320094 470454 320124
rect 470454 320094 470492 320124
rect 470516 320094 470518 320124
rect 470518 320094 470570 320124
rect 470570 320094 470572 320124
rect 470596 320094 470634 320124
rect 470634 320094 470646 320124
rect 470646 320094 470652 320124
rect 470676 320094 470698 320124
rect 470698 320094 470710 320124
rect 470710 320094 470732 320124
rect 470756 320094 470762 320124
rect 470762 320094 470774 320124
rect 470774 320094 470812 320124
rect 470276 320060 470332 320070
rect 470356 320060 470412 320070
rect 470436 320060 470492 320070
rect 470516 320060 470572 320070
rect 470596 320060 470652 320070
rect 470676 320060 470732 320070
rect 470756 320060 470812 320070
rect 470276 320014 470314 320060
rect 470314 320014 470326 320060
rect 470326 320014 470332 320060
rect 470356 320014 470378 320060
rect 470378 320014 470390 320060
rect 470390 320014 470412 320060
rect 470436 320014 470442 320060
rect 470442 320014 470454 320060
rect 470454 320014 470492 320060
rect 470516 320014 470518 320060
rect 470518 320014 470570 320060
rect 470570 320014 470572 320060
rect 470596 320014 470634 320060
rect 470634 320014 470646 320060
rect 470646 320014 470652 320060
rect 470676 320014 470698 320060
rect 470698 320014 470710 320060
rect 470710 320014 470732 320060
rect 470756 320014 470762 320060
rect 470762 320014 470774 320060
rect 470774 320014 470812 320060
rect 470276 307036 470314 307082
rect 470314 307036 470326 307082
rect 470326 307036 470332 307082
rect 470356 307036 470378 307082
rect 470378 307036 470390 307082
rect 470390 307036 470412 307082
rect 470436 307036 470442 307082
rect 470442 307036 470454 307082
rect 470454 307036 470492 307082
rect 470516 307036 470518 307082
rect 470518 307036 470570 307082
rect 470570 307036 470572 307082
rect 470596 307036 470634 307082
rect 470634 307036 470646 307082
rect 470646 307036 470652 307082
rect 470676 307036 470698 307082
rect 470698 307036 470710 307082
rect 470710 307036 470732 307082
rect 470756 307036 470762 307082
rect 470762 307036 470774 307082
rect 470774 307036 470812 307082
rect 470276 307026 470332 307036
rect 470356 307026 470412 307036
rect 470436 307026 470492 307036
rect 470516 307026 470572 307036
rect 470596 307026 470652 307036
rect 470676 307026 470732 307036
rect 470756 307026 470812 307036
rect 470276 306972 470314 307002
rect 470314 306972 470326 307002
rect 470326 306972 470332 307002
rect 470356 306972 470378 307002
rect 470378 306972 470390 307002
rect 470390 306972 470412 307002
rect 470436 306972 470442 307002
rect 470442 306972 470454 307002
rect 470454 306972 470492 307002
rect 470516 306972 470518 307002
rect 470518 306972 470570 307002
rect 470570 306972 470572 307002
rect 470596 306972 470634 307002
rect 470634 306972 470646 307002
rect 470646 306972 470652 307002
rect 470676 306972 470698 307002
rect 470698 306972 470710 307002
rect 470710 306972 470732 307002
rect 470756 306972 470762 307002
rect 470762 306972 470774 307002
rect 470774 306972 470812 307002
rect 470276 306960 470332 306972
rect 470356 306960 470412 306972
rect 470436 306960 470492 306972
rect 470516 306960 470572 306972
rect 470596 306960 470652 306972
rect 470676 306960 470732 306972
rect 470756 306960 470812 306972
rect 470276 306946 470314 306960
rect 470314 306946 470326 306960
rect 470326 306946 470332 306960
rect 470356 306946 470378 306960
rect 470378 306946 470390 306960
rect 470390 306946 470412 306960
rect 470436 306946 470442 306960
rect 470442 306946 470454 306960
rect 470454 306946 470492 306960
rect 470516 306946 470518 306960
rect 470518 306946 470570 306960
rect 470570 306946 470572 306960
rect 470596 306946 470634 306960
rect 470634 306946 470646 306960
rect 470646 306946 470652 306960
rect 470676 306946 470698 306960
rect 470698 306946 470710 306960
rect 470710 306946 470732 306960
rect 470756 306946 470762 306960
rect 470762 306946 470774 306960
rect 470774 306946 470812 306960
rect 470276 306908 470314 306922
rect 470314 306908 470326 306922
rect 470326 306908 470332 306922
rect 470356 306908 470378 306922
rect 470378 306908 470390 306922
rect 470390 306908 470412 306922
rect 470436 306908 470442 306922
rect 470442 306908 470454 306922
rect 470454 306908 470492 306922
rect 470516 306908 470518 306922
rect 470518 306908 470570 306922
rect 470570 306908 470572 306922
rect 470596 306908 470634 306922
rect 470634 306908 470646 306922
rect 470646 306908 470652 306922
rect 470676 306908 470698 306922
rect 470698 306908 470710 306922
rect 470710 306908 470732 306922
rect 470756 306908 470762 306922
rect 470762 306908 470774 306922
rect 470774 306908 470812 306922
rect 470276 306896 470332 306908
rect 470356 306896 470412 306908
rect 470436 306896 470492 306908
rect 470516 306896 470572 306908
rect 470596 306896 470652 306908
rect 470676 306896 470732 306908
rect 470756 306896 470812 306908
rect 470276 306866 470314 306896
rect 470314 306866 470326 306896
rect 470326 306866 470332 306896
rect 470356 306866 470378 306896
rect 470378 306866 470390 306896
rect 470390 306866 470412 306896
rect 470436 306866 470442 306896
rect 470442 306866 470454 306896
rect 470454 306866 470492 306896
rect 470516 306866 470518 306896
rect 470518 306866 470570 306896
rect 470570 306866 470572 306896
rect 470596 306866 470634 306896
rect 470634 306866 470646 306896
rect 470646 306866 470652 306896
rect 470676 306866 470698 306896
rect 470698 306866 470710 306896
rect 470710 306866 470732 306896
rect 470756 306866 470762 306896
rect 470762 306866 470774 306896
rect 470774 306866 470812 306896
rect 470276 306832 470332 306842
rect 470356 306832 470412 306842
rect 470436 306832 470492 306842
rect 470516 306832 470572 306842
rect 470596 306832 470652 306842
rect 470676 306832 470732 306842
rect 470756 306832 470812 306842
rect 470276 306786 470314 306832
rect 470314 306786 470326 306832
rect 470326 306786 470332 306832
rect 470356 306786 470378 306832
rect 470378 306786 470390 306832
rect 470390 306786 470412 306832
rect 470436 306786 470442 306832
rect 470442 306786 470454 306832
rect 470454 306786 470492 306832
rect 470516 306786 470518 306832
rect 470518 306786 470570 306832
rect 470570 306786 470572 306832
rect 470596 306786 470634 306832
rect 470634 306786 470646 306832
rect 470646 306786 470652 306832
rect 470676 306786 470698 306832
rect 470698 306786 470710 306832
rect 470710 306786 470732 306832
rect 470756 306786 470762 306832
rect 470762 306786 470774 306832
rect 470774 306786 470812 306832
rect 483478 321546 483534 321602
rect 474278 321274 474334 321330
rect 481178 321002 481234 321058
rect 488170 321002 488226 321058
rect 478142 320866 478198 320922
rect 480902 306450 480958 306506
rect 469036 305951 469074 305997
rect 469074 305951 469086 305997
rect 469086 305951 469092 305997
rect 469116 305951 469138 305997
rect 469138 305951 469150 305997
rect 469150 305951 469172 305997
rect 469196 305951 469202 305997
rect 469202 305951 469214 305997
rect 469214 305951 469252 305997
rect 469276 305951 469278 305997
rect 469278 305951 469330 305997
rect 469330 305951 469332 305997
rect 469356 305951 469394 305997
rect 469394 305951 469406 305997
rect 469406 305951 469412 305997
rect 469436 305951 469458 305997
rect 469458 305951 469470 305997
rect 469470 305951 469492 305997
rect 469516 305951 469522 305997
rect 469522 305951 469534 305997
rect 469534 305951 469572 305997
rect 469036 305941 469092 305951
rect 469116 305941 469172 305951
rect 469196 305941 469252 305951
rect 469276 305941 469332 305951
rect 469356 305941 469412 305951
rect 469436 305941 469492 305951
rect 469516 305941 469572 305951
rect 469036 305887 469074 305917
rect 469074 305887 469086 305917
rect 469086 305887 469092 305917
rect 469116 305887 469138 305917
rect 469138 305887 469150 305917
rect 469150 305887 469172 305917
rect 469196 305887 469202 305917
rect 469202 305887 469214 305917
rect 469214 305887 469252 305917
rect 469276 305887 469278 305917
rect 469278 305887 469330 305917
rect 469330 305887 469332 305917
rect 469356 305887 469394 305917
rect 469394 305887 469406 305917
rect 469406 305887 469412 305917
rect 469436 305887 469458 305917
rect 469458 305887 469470 305917
rect 469470 305887 469492 305917
rect 469516 305887 469522 305917
rect 469522 305887 469534 305917
rect 469534 305887 469572 305917
rect 469036 305875 469092 305887
rect 469116 305875 469172 305887
rect 469196 305875 469252 305887
rect 469276 305875 469332 305887
rect 469356 305875 469412 305887
rect 469436 305875 469492 305887
rect 469516 305875 469572 305887
rect 469036 305861 469074 305875
rect 469074 305861 469086 305875
rect 469086 305861 469092 305875
rect 469116 305861 469138 305875
rect 469138 305861 469150 305875
rect 469150 305861 469172 305875
rect 469196 305861 469202 305875
rect 469202 305861 469214 305875
rect 469214 305861 469252 305875
rect 469276 305861 469278 305875
rect 469278 305861 469330 305875
rect 469330 305861 469332 305875
rect 469356 305861 469394 305875
rect 469394 305861 469406 305875
rect 469406 305861 469412 305875
rect 469436 305861 469458 305875
rect 469458 305861 469470 305875
rect 469470 305861 469492 305875
rect 469516 305861 469522 305875
rect 469522 305861 469534 305875
rect 469534 305861 469572 305875
rect 469036 305823 469074 305837
rect 469074 305823 469086 305837
rect 469086 305823 469092 305837
rect 469116 305823 469138 305837
rect 469138 305823 469150 305837
rect 469150 305823 469172 305837
rect 469196 305823 469202 305837
rect 469202 305823 469214 305837
rect 469214 305823 469252 305837
rect 469276 305823 469278 305837
rect 469278 305823 469330 305837
rect 469330 305823 469332 305837
rect 469356 305823 469394 305837
rect 469394 305823 469406 305837
rect 469406 305823 469412 305837
rect 469436 305823 469458 305837
rect 469458 305823 469470 305837
rect 469470 305823 469492 305837
rect 469516 305823 469522 305837
rect 469522 305823 469534 305837
rect 469534 305823 469572 305837
rect 469036 305811 469092 305823
rect 469116 305811 469172 305823
rect 469196 305811 469252 305823
rect 469276 305811 469332 305823
rect 469356 305811 469412 305823
rect 469436 305811 469492 305823
rect 469516 305811 469572 305823
rect 469036 305781 469074 305811
rect 469074 305781 469086 305811
rect 469086 305781 469092 305811
rect 469116 305781 469138 305811
rect 469138 305781 469150 305811
rect 469150 305781 469172 305811
rect 469196 305781 469202 305811
rect 469202 305781 469214 305811
rect 469214 305781 469252 305811
rect 469276 305781 469278 305811
rect 469278 305781 469330 305811
rect 469330 305781 469332 305811
rect 469356 305781 469394 305811
rect 469394 305781 469406 305811
rect 469406 305781 469412 305811
rect 469436 305781 469458 305811
rect 469458 305781 469470 305811
rect 469470 305781 469492 305811
rect 469516 305781 469522 305811
rect 469522 305781 469534 305811
rect 469534 305781 469572 305811
rect 469036 305747 469092 305757
rect 469116 305747 469172 305757
rect 469196 305747 469252 305757
rect 469276 305747 469332 305757
rect 469356 305747 469412 305757
rect 469436 305747 469492 305757
rect 469516 305747 469572 305757
rect 469036 305701 469074 305747
rect 469074 305701 469086 305747
rect 469086 305701 469092 305747
rect 469116 305701 469138 305747
rect 469138 305701 469150 305747
rect 469150 305701 469172 305747
rect 469196 305701 469202 305747
rect 469202 305701 469214 305747
rect 469214 305701 469252 305747
rect 469276 305701 469278 305747
rect 469278 305701 469330 305747
rect 469330 305701 469332 305747
rect 469356 305701 469394 305747
rect 469394 305701 469406 305747
rect 469406 305701 469412 305747
rect 469436 305701 469458 305747
rect 469458 305701 469470 305747
rect 469470 305701 469492 305747
rect 469516 305701 469522 305747
rect 469522 305701 469534 305747
rect 469534 305701 469572 305747
rect 470276 304864 470314 304910
rect 470314 304864 470326 304910
rect 470326 304864 470332 304910
rect 470356 304864 470378 304910
rect 470378 304864 470390 304910
rect 470390 304864 470412 304910
rect 470436 304864 470442 304910
rect 470442 304864 470454 304910
rect 470454 304864 470492 304910
rect 470516 304864 470518 304910
rect 470518 304864 470570 304910
rect 470570 304864 470572 304910
rect 470596 304864 470634 304910
rect 470634 304864 470646 304910
rect 470646 304864 470652 304910
rect 470676 304864 470698 304910
rect 470698 304864 470710 304910
rect 470710 304864 470732 304910
rect 470756 304864 470762 304910
rect 470762 304864 470774 304910
rect 470774 304864 470812 304910
rect 470276 304854 470332 304864
rect 470356 304854 470412 304864
rect 470436 304854 470492 304864
rect 470516 304854 470572 304864
rect 470596 304854 470652 304864
rect 470676 304854 470732 304864
rect 470756 304854 470812 304864
rect 470276 304800 470314 304830
rect 470314 304800 470326 304830
rect 470326 304800 470332 304830
rect 470356 304800 470378 304830
rect 470378 304800 470390 304830
rect 470390 304800 470412 304830
rect 470436 304800 470442 304830
rect 470442 304800 470454 304830
rect 470454 304800 470492 304830
rect 470516 304800 470518 304830
rect 470518 304800 470570 304830
rect 470570 304800 470572 304830
rect 470596 304800 470634 304830
rect 470634 304800 470646 304830
rect 470646 304800 470652 304830
rect 470676 304800 470698 304830
rect 470698 304800 470710 304830
rect 470710 304800 470732 304830
rect 470756 304800 470762 304830
rect 470762 304800 470774 304830
rect 470774 304800 470812 304830
rect 470276 304788 470332 304800
rect 470356 304788 470412 304800
rect 470436 304788 470492 304800
rect 470516 304788 470572 304800
rect 470596 304788 470652 304800
rect 470676 304788 470732 304800
rect 470756 304788 470812 304800
rect 470276 304774 470314 304788
rect 470314 304774 470326 304788
rect 470326 304774 470332 304788
rect 470356 304774 470378 304788
rect 470378 304774 470390 304788
rect 470390 304774 470412 304788
rect 470436 304774 470442 304788
rect 470442 304774 470454 304788
rect 470454 304774 470492 304788
rect 470516 304774 470518 304788
rect 470518 304774 470570 304788
rect 470570 304774 470572 304788
rect 470596 304774 470634 304788
rect 470634 304774 470646 304788
rect 470646 304774 470652 304788
rect 470676 304774 470698 304788
rect 470698 304774 470710 304788
rect 470710 304774 470732 304788
rect 470756 304774 470762 304788
rect 470762 304774 470774 304788
rect 470774 304774 470812 304788
rect 470276 304736 470314 304750
rect 470314 304736 470326 304750
rect 470326 304736 470332 304750
rect 470356 304736 470378 304750
rect 470378 304736 470390 304750
rect 470390 304736 470412 304750
rect 470436 304736 470442 304750
rect 470442 304736 470454 304750
rect 470454 304736 470492 304750
rect 470516 304736 470518 304750
rect 470518 304736 470570 304750
rect 470570 304736 470572 304750
rect 470596 304736 470634 304750
rect 470634 304736 470646 304750
rect 470646 304736 470652 304750
rect 470676 304736 470698 304750
rect 470698 304736 470710 304750
rect 470710 304736 470732 304750
rect 470756 304736 470762 304750
rect 470762 304736 470774 304750
rect 470774 304736 470812 304750
rect 470276 304724 470332 304736
rect 470356 304724 470412 304736
rect 470436 304724 470492 304736
rect 470516 304724 470572 304736
rect 470596 304724 470652 304736
rect 470676 304724 470732 304736
rect 470756 304724 470812 304736
rect 470276 304694 470314 304724
rect 470314 304694 470326 304724
rect 470326 304694 470332 304724
rect 470356 304694 470378 304724
rect 470378 304694 470390 304724
rect 470390 304694 470412 304724
rect 470436 304694 470442 304724
rect 470442 304694 470454 304724
rect 470454 304694 470492 304724
rect 470516 304694 470518 304724
rect 470518 304694 470570 304724
rect 470570 304694 470572 304724
rect 470596 304694 470634 304724
rect 470634 304694 470646 304724
rect 470646 304694 470652 304724
rect 470676 304694 470698 304724
rect 470698 304694 470710 304724
rect 470710 304694 470732 304724
rect 470756 304694 470762 304724
rect 470762 304694 470774 304724
rect 470774 304694 470812 304724
rect 470276 304660 470332 304670
rect 470356 304660 470412 304670
rect 470436 304660 470492 304670
rect 470516 304660 470572 304670
rect 470596 304660 470652 304670
rect 470676 304660 470732 304670
rect 470756 304660 470812 304670
rect 470276 304614 470314 304660
rect 470314 304614 470326 304660
rect 470326 304614 470332 304660
rect 470356 304614 470378 304660
rect 470378 304614 470390 304660
rect 470390 304614 470412 304660
rect 470436 304614 470442 304660
rect 470442 304614 470454 304660
rect 470454 304614 470492 304660
rect 470516 304614 470518 304660
rect 470518 304614 470570 304660
rect 470570 304614 470572 304660
rect 470596 304614 470634 304660
rect 470634 304614 470646 304660
rect 470646 304614 470652 304660
rect 470676 304614 470698 304660
rect 470698 304614 470710 304660
rect 470710 304614 470732 304660
rect 470756 304614 470762 304660
rect 470762 304614 470774 304660
rect 470774 304614 470812 304660
rect 470276 287437 470314 287483
rect 470314 287437 470326 287483
rect 470326 287437 470332 287483
rect 470356 287437 470378 287483
rect 470378 287437 470390 287483
rect 470390 287437 470412 287483
rect 470436 287437 470442 287483
rect 470442 287437 470454 287483
rect 470454 287437 470492 287483
rect 470516 287437 470518 287483
rect 470518 287437 470570 287483
rect 470570 287437 470572 287483
rect 470596 287437 470634 287483
rect 470634 287437 470646 287483
rect 470646 287437 470652 287483
rect 470676 287437 470698 287483
rect 470698 287437 470710 287483
rect 470710 287437 470732 287483
rect 470756 287437 470762 287483
rect 470762 287437 470774 287483
rect 470774 287437 470812 287483
rect 470276 287427 470332 287437
rect 470356 287427 470412 287437
rect 470436 287427 470492 287437
rect 470516 287427 470572 287437
rect 470596 287427 470652 287437
rect 470676 287427 470732 287437
rect 470756 287427 470812 287437
rect 470276 287373 470314 287403
rect 470314 287373 470326 287403
rect 470326 287373 470332 287403
rect 470356 287373 470378 287403
rect 470378 287373 470390 287403
rect 470390 287373 470412 287403
rect 470436 287373 470442 287403
rect 470442 287373 470454 287403
rect 470454 287373 470492 287403
rect 470516 287373 470518 287403
rect 470518 287373 470570 287403
rect 470570 287373 470572 287403
rect 470596 287373 470634 287403
rect 470634 287373 470646 287403
rect 470646 287373 470652 287403
rect 470676 287373 470698 287403
rect 470698 287373 470710 287403
rect 470710 287373 470732 287403
rect 470756 287373 470762 287403
rect 470762 287373 470774 287403
rect 470774 287373 470812 287403
rect 470276 287361 470332 287373
rect 470356 287361 470412 287373
rect 470436 287361 470492 287373
rect 470516 287361 470572 287373
rect 470596 287361 470652 287373
rect 470676 287361 470732 287373
rect 470756 287361 470812 287373
rect 470276 287347 470314 287361
rect 470314 287347 470326 287361
rect 470326 287347 470332 287361
rect 470356 287347 470378 287361
rect 470378 287347 470390 287361
rect 470390 287347 470412 287361
rect 470436 287347 470442 287361
rect 470442 287347 470454 287361
rect 470454 287347 470492 287361
rect 470516 287347 470518 287361
rect 470518 287347 470570 287361
rect 470570 287347 470572 287361
rect 470596 287347 470634 287361
rect 470634 287347 470646 287361
rect 470646 287347 470652 287361
rect 470676 287347 470698 287361
rect 470698 287347 470710 287361
rect 470710 287347 470732 287361
rect 470756 287347 470762 287361
rect 470762 287347 470774 287361
rect 470774 287347 470812 287361
rect 470276 287309 470314 287323
rect 470314 287309 470326 287323
rect 470326 287309 470332 287323
rect 470356 287309 470378 287323
rect 470378 287309 470390 287323
rect 470390 287309 470412 287323
rect 470436 287309 470442 287323
rect 470442 287309 470454 287323
rect 470454 287309 470492 287323
rect 470516 287309 470518 287323
rect 470518 287309 470570 287323
rect 470570 287309 470572 287323
rect 470596 287309 470634 287323
rect 470634 287309 470646 287323
rect 470646 287309 470652 287323
rect 470676 287309 470698 287323
rect 470698 287309 470710 287323
rect 470710 287309 470732 287323
rect 470756 287309 470762 287323
rect 470762 287309 470774 287323
rect 470774 287309 470812 287323
rect 470276 287297 470332 287309
rect 470356 287297 470412 287309
rect 470436 287297 470492 287309
rect 470516 287297 470572 287309
rect 470596 287297 470652 287309
rect 470676 287297 470732 287309
rect 470756 287297 470812 287309
rect 470276 287267 470314 287297
rect 470314 287267 470326 287297
rect 470326 287267 470332 287297
rect 470356 287267 470378 287297
rect 470378 287267 470390 287297
rect 470390 287267 470412 287297
rect 470436 287267 470442 287297
rect 470442 287267 470454 287297
rect 470454 287267 470492 287297
rect 470516 287267 470518 287297
rect 470518 287267 470570 287297
rect 470570 287267 470572 287297
rect 470596 287267 470634 287297
rect 470634 287267 470646 287297
rect 470646 287267 470652 287297
rect 470676 287267 470698 287297
rect 470698 287267 470710 287297
rect 470710 287267 470732 287297
rect 470756 287267 470762 287297
rect 470762 287267 470774 287297
rect 470774 287267 470812 287297
rect 470276 287233 470332 287243
rect 470356 287233 470412 287243
rect 470436 287233 470492 287243
rect 470516 287233 470572 287243
rect 470596 287233 470652 287243
rect 470676 287233 470732 287243
rect 470756 287233 470812 287243
rect 470276 287187 470314 287233
rect 470314 287187 470326 287233
rect 470326 287187 470332 287233
rect 470356 287187 470378 287233
rect 470378 287187 470390 287233
rect 470390 287187 470412 287233
rect 470436 287187 470442 287233
rect 470442 287187 470454 287233
rect 470454 287187 470492 287233
rect 470516 287187 470518 287233
rect 470518 287187 470570 287233
rect 470570 287187 470572 287233
rect 470596 287187 470634 287233
rect 470634 287187 470646 287233
rect 470646 287187 470652 287233
rect 470676 287187 470698 287233
rect 470698 287187 470710 287233
rect 470710 287187 470732 287233
rect 470756 287187 470762 287233
rect 470762 287187 470774 287233
rect 470774 287187 470812 287233
rect 487534 306178 487590 306234
rect 473726 305906 473782 305962
rect 477739 305634 477795 305690
rect 484122 305498 484178 305554
rect 482282 302234 482338 302290
rect 482282 288362 482338 288418
rect 478633 286866 478689 286922
rect 474921 286594 474977 286650
rect 484766 286594 484822 286650
rect 488538 286594 488594 286650
rect 469036 286352 469074 286398
rect 469074 286352 469086 286398
rect 469086 286352 469092 286398
rect 469116 286352 469138 286398
rect 469138 286352 469150 286398
rect 469150 286352 469172 286398
rect 469196 286352 469202 286398
rect 469202 286352 469214 286398
rect 469214 286352 469252 286398
rect 469276 286352 469278 286398
rect 469278 286352 469330 286398
rect 469330 286352 469332 286398
rect 469356 286352 469394 286398
rect 469394 286352 469406 286398
rect 469406 286352 469412 286398
rect 469436 286352 469458 286398
rect 469458 286352 469470 286398
rect 469470 286352 469492 286398
rect 469516 286352 469522 286398
rect 469522 286352 469534 286398
rect 469534 286352 469572 286398
rect 469036 286342 469092 286352
rect 469116 286342 469172 286352
rect 469196 286342 469252 286352
rect 469276 286342 469332 286352
rect 469356 286342 469412 286352
rect 469436 286342 469492 286352
rect 469516 286342 469572 286352
rect 469036 286288 469074 286318
rect 469074 286288 469086 286318
rect 469086 286288 469092 286318
rect 469116 286288 469138 286318
rect 469138 286288 469150 286318
rect 469150 286288 469172 286318
rect 469196 286288 469202 286318
rect 469202 286288 469214 286318
rect 469214 286288 469252 286318
rect 469276 286288 469278 286318
rect 469278 286288 469330 286318
rect 469330 286288 469332 286318
rect 469356 286288 469394 286318
rect 469394 286288 469406 286318
rect 469406 286288 469412 286318
rect 469436 286288 469458 286318
rect 469458 286288 469470 286318
rect 469470 286288 469492 286318
rect 469516 286288 469522 286318
rect 469522 286288 469534 286318
rect 469534 286288 469572 286318
rect 469036 286276 469092 286288
rect 469116 286276 469172 286288
rect 469196 286276 469252 286288
rect 469276 286276 469332 286288
rect 469356 286276 469412 286288
rect 469436 286276 469492 286288
rect 469516 286276 469572 286288
rect 469036 286262 469074 286276
rect 469074 286262 469086 286276
rect 469086 286262 469092 286276
rect 469116 286262 469138 286276
rect 469138 286262 469150 286276
rect 469150 286262 469172 286276
rect 469196 286262 469202 286276
rect 469202 286262 469214 286276
rect 469214 286262 469252 286276
rect 469276 286262 469278 286276
rect 469278 286262 469330 286276
rect 469330 286262 469332 286276
rect 469356 286262 469394 286276
rect 469394 286262 469406 286276
rect 469406 286262 469412 286276
rect 469436 286262 469458 286276
rect 469458 286262 469470 286276
rect 469470 286262 469492 286276
rect 469516 286262 469522 286276
rect 469522 286262 469534 286276
rect 469534 286262 469572 286276
rect 469036 286224 469074 286238
rect 469074 286224 469086 286238
rect 469086 286224 469092 286238
rect 469116 286224 469138 286238
rect 469138 286224 469150 286238
rect 469150 286224 469172 286238
rect 469196 286224 469202 286238
rect 469202 286224 469214 286238
rect 469214 286224 469252 286238
rect 469276 286224 469278 286238
rect 469278 286224 469330 286238
rect 469330 286224 469332 286238
rect 469356 286224 469394 286238
rect 469394 286224 469406 286238
rect 469406 286224 469412 286238
rect 469436 286224 469458 286238
rect 469458 286224 469470 286238
rect 469470 286224 469492 286238
rect 469516 286224 469522 286238
rect 469522 286224 469534 286238
rect 469534 286224 469572 286238
rect 469036 286212 469092 286224
rect 469116 286212 469172 286224
rect 469196 286212 469252 286224
rect 469276 286212 469332 286224
rect 469356 286212 469412 286224
rect 469436 286212 469492 286224
rect 469516 286212 469572 286224
rect 469036 286182 469074 286212
rect 469074 286182 469086 286212
rect 469086 286182 469092 286212
rect 469116 286182 469138 286212
rect 469138 286182 469150 286212
rect 469150 286182 469172 286212
rect 469196 286182 469202 286212
rect 469202 286182 469214 286212
rect 469214 286182 469252 286212
rect 469276 286182 469278 286212
rect 469278 286182 469330 286212
rect 469330 286182 469332 286212
rect 469356 286182 469394 286212
rect 469394 286182 469406 286212
rect 469406 286182 469412 286212
rect 469436 286182 469458 286212
rect 469458 286182 469470 286212
rect 469470 286182 469492 286212
rect 469516 286182 469522 286212
rect 469522 286182 469534 286212
rect 469534 286182 469572 286212
rect 469036 286148 469092 286158
rect 469116 286148 469172 286158
rect 469196 286148 469252 286158
rect 469276 286148 469332 286158
rect 469356 286148 469412 286158
rect 469436 286148 469492 286158
rect 469516 286148 469572 286158
rect 469036 286102 469074 286148
rect 469074 286102 469086 286148
rect 469086 286102 469092 286148
rect 469116 286102 469138 286148
rect 469138 286102 469150 286148
rect 469150 286102 469172 286148
rect 469196 286102 469202 286148
rect 469202 286102 469214 286148
rect 469214 286102 469252 286148
rect 469276 286102 469278 286148
rect 469278 286102 469330 286148
rect 469330 286102 469332 286148
rect 469356 286102 469394 286148
rect 469394 286102 469406 286148
rect 469406 286102 469412 286148
rect 469436 286102 469458 286148
rect 469458 286102 469470 286148
rect 469470 286102 469492 286148
rect 469516 286102 469522 286148
rect 469522 286102 469534 286148
rect 469534 286102 469572 286148
rect 470276 285264 470314 285310
rect 470314 285264 470326 285310
rect 470326 285264 470332 285310
rect 470356 285264 470378 285310
rect 470378 285264 470390 285310
rect 470390 285264 470412 285310
rect 470436 285264 470442 285310
rect 470442 285264 470454 285310
rect 470454 285264 470492 285310
rect 470516 285264 470518 285310
rect 470518 285264 470570 285310
rect 470570 285264 470572 285310
rect 470596 285264 470634 285310
rect 470634 285264 470646 285310
rect 470646 285264 470652 285310
rect 470676 285264 470698 285310
rect 470698 285264 470710 285310
rect 470710 285264 470732 285310
rect 470756 285264 470762 285310
rect 470762 285264 470774 285310
rect 470774 285264 470812 285310
rect 470276 285254 470332 285264
rect 470356 285254 470412 285264
rect 470436 285254 470492 285264
rect 470516 285254 470572 285264
rect 470596 285254 470652 285264
rect 470676 285254 470732 285264
rect 470756 285254 470812 285264
rect 470276 285200 470314 285230
rect 470314 285200 470326 285230
rect 470326 285200 470332 285230
rect 470356 285200 470378 285230
rect 470378 285200 470390 285230
rect 470390 285200 470412 285230
rect 470436 285200 470442 285230
rect 470442 285200 470454 285230
rect 470454 285200 470492 285230
rect 470516 285200 470518 285230
rect 470518 285200 470570 285230
rect 470570 285200 470572 285230
rect 470596 285200 470634 285230
rect 470634 285200 470646 285230
rect 470646 285200 470652 285230
rect 470676 285200 470698 285230
rect 470698 285200 470710 285230
rect 470710 285200 470732 285230
rect 470756 285200 470762 285230
rect 470762 285200 470774 285230
rect 470774 285200 470812 285230
rect 470276 285188 470332 285200
rect 470356 285188 470412 285200
rect 470436 285188 470492 285200
rect 470516 285188 470572 285200
rect 470596 285188 470652 285200
rect 470676 285188 470732 285200
rect 470756 285188 470812 285200
rect 470276 285174 470314 285188
rect 470314 285174 470326 285188
rect 470326 285174 470332 285188
rect 470356 285174 470378 285188
rect 470378 285174 470390 285188
rect 470390 285174 470412 285188
rect 470436 285174 470442 285188
rect 470442 285174 470454 285188
rect 470454 285174 470492 285188
rect 470516 285174 470518 285188
rect 470518 285174 470570 285188
rect 470570 285174 470572 285188
rect 470596 285174 470634 285188
rect 470634 285174 470646 285188
rect 470646 285174 470652 285188
rect 470676 285174 470698 285188
rect 470698 285174 470710 285188
rect 470710 285174 470732 285188
rect 470756 285174 470762 285188
rect 470762 285174 470774 285188
rect 470774 285174 470812 285188
rect 470276 285136 470314 285150
rect 470314 285136 470326 285150
rect 470326 285136 470332 285150
rect 470356 285136 470378 285150
rect 470378 285136 470390 285150
rect 470390 285136 470412 285150
rect 470436 285136 470442 285150
rect 470442 285136 470454 285150
rect 470454 285136 470492 285150
rect 470516 285136 470518 285150
rect 470518 285136 470570 285150
rect 470570 285136 470572 285150
rect 470596 285136 470634 285150
rect 470634 285136 470646 285150
rect 470646 285136 470652 285150
rect 470676 285136 470698 285150
rect 470698 285136 470710 285150
rect 470710 285136 470732 285150
rect 470756 285136 470762 285150
rect 470762 285136 470774 285150
rect 470774 285136 470812 285150
rect 470276 285124 470332 285136
rect 470356 285124 470412 285136
rect 470436 285124 470492 285136
rect 470516 285124 470572 285136
rect 470596 285124 470652 285136
rect 470676 285124 470732 285136
rect 470756 285124 470812 285136
rect 470276 285094 470314 285124
rect 470314 285094 470326 285124
rect 470326 285094 470332 285124
rect 470356 285094 470378 285124
rect 470378 285094 470390 285124
rect 470390 285094 470412 285124
rect 470436 285094 470442 285124
rect 470442 285094 470454 285124
rect 470454 285094 470492 285124
rect 470516 285094 470518 285124
rect 470518 285094 470570 285124
rect 470570 285094 470572 285124
rect 470596 285094 470634 285124
rect 470634 285094 470646 285124
rect 470646 285094 470652 285124
rect 470676 285094 470698 285124
rect 470698 285094 470710 285124
rect 470710 285094 470732 285124
rect 470756 285094 470762 285124
rect 470762 285094 470774 285124
rect 470774 285094 470812 285124
rect 470276 285060 470332 285070
rect 470356 285060 470412 285070
rect 470436 285060 470492 285070
rect 470516 285060 470572 285070
rect 470596 285060 470652 285070
rect 470676 285060 470732 285070
rect 470756 285060 470812 285070
rect 470276 285014 470314 285060
rect 470314 285014 470326 285060
rect 470326 285014 470332 285060
rect 470356 285014 470378 285060
rect 470378 285014 470390 285060
rect 470390 285014 470412 285060
rect 470436 285014 470442 285060
rect 470442 285014 470454 285060
rect 470454 285014 470492 285060
rect 470516 285014 470518 285060
rect 470518 285014 470570 285060
rect 470570 285014 470572 285060
rect 470596 285014 470634 285060
rect 470634 285014 470646 285060
rect 470646 285014 470652 285060
rect 470676 285014 470698 285060
rect 470698 285014 470710 285060
rect 470710 285014 470732 285060
rect 470756 285014 470762 285060
rect 470762 285014 470774 285060
rect 470774 285014 470812 285060
rect 482190 285642 482246 285698
rect 482374 273266 482430 273322
rect 470276 267437 470314 267483
rect 470314 267437 470326 267483
rect 470326 267437 470332 267483
rect 470356 267437 470378 267483
rect 470378 267437 470390 267483
rect 470390 267437 470412 267483
rect 470436 267437 470442 267483
rect 470442 267437 470454 267483
rect 470454 267437 470492 267483
rect 470516 267437 470518 267483
rect 470518 267437 470570 267483
rect 470570 267437 470572 267483
rect 470596 267437 470634 267483
rect 470634 267437 470646 267483
rect 470646 267437 470652 267483
rect 470676 267437 470698 267483
rect 470698 267437 470710 267483
rect 470710 267437 470732 267483
rect 470756 267437 470762 267483
rect 470762 267437 470774 267483
rect 470774 267437 470812 267483
rect 470276 267427 470332 267437
rect 470356 267427 470412 267437
rect 470436 267427 470492 267437
rect 470516 267427 470572 267437
rect 470596 267427 470652 267437
rect 470676 267427 470732 267437
rect 470756 267427 470812 267437
rect 470276 267373 470314 267403
rect 470314 267373 470326 267403
rect 470326 267373 470332 267403
rect 470356 267373 470378 267403
rect 470378 267373 470390 267403
rect 470390 267373 470412 267403
rect 470436 267373 470442 267403
rect 470442 267373 470454 267403
rect 470454 267373 470492 267403
rect 470516 267373 470518 267403
rect 470518 267373 470570 267403
rect 470570 267373 470572 267403
rect 470596 267373 470634 267403
rect 470634 267373 470646 267403
rect 470646 267373 470652 267403
rect 470676 267373 470698 267403
rect 470698 267373 470710 267403
rect 470710 267373 470732 267403
rect 470756 267373 470762 267403
rect 470762 267373 470774 267403
rect 470774 267373 470812 267403
rect 470276 267361 470332 267373
rect 470356 267361 470412 267373
rect 470436 267361 470492 267373
rect 470516 267361 470572 267373
rect 470596 267361 470652 267373
rect 470676 267361 470732 267373
rect 470756 267361 470812 267373
rect 470276 267347 470314 267361
rect 470314 267347 470326 267361
rect 470326 267347 470332 267361
rect 470356 267347 470378 267361
rect 470378 267347 470390 267361
rect 470390 267347 470412 267361
rect 470436 267347 470442 267361
rect 470442 267347 470454 267361
rect 470454 267347 470492 267361
rect 470516 267347 470518 267361
rect 470518 267347 470570 267361
rect 470570 267347 470572 267361
rect 470596 267347 470634 267361
rect 470634 267347 470646 267361
rect 470646 267347 470652 267361
rect 470676 267347 470698 267361
rect 470698 267347 470710 267361
rect 470710 267347 470732 267361
rect 470756 267347 470762 267361
rect 470762 267347 470774 267361
rect 470774 267347 470812 267361
rect 470276 267309 470314 267323
rect 470314 267309 470326 267323
rect 470326 267309 470332 267323
rect 470356 267309 470378 267323
rect 470378 267309 470390 267323
rect 470390 267309 470412 267323
rect 470436 267309 470442 267323
rect 470442 267309 470454 267323
rect 470454 267309 470492 267323
rect 470516 267309 470518 267323
rect 470518 267309 470570 267323
rect 470570 267309 470572 267323
rect 470596 267309 470634 267323
rect 470634 267309 470646 267323
rect 470646 267309 470652 267323
rect 470676 267309 470698 267323
rect 470698 267309 470710 267323
rect 470710 267309 470732 267323
rect 470756 267309 470762 267323
rect 470762 267309 470774 267323
rect 470774 267309 470812 267323
rect 470276 267297 470332 267309
rect 470356 267297 470412 267309
rect 470436 267297 470492 267309
rect 470516 267297 470572 267309
rect 470596 267297 470652 267309
rect 470676 267297 470732 267309
rect 470756 267297 470812 267309
rect 470276 267267 470314 267297
rect 470314 267267 470326 267297
rect 470326 267267 470332 267297
rect 470356 267267 470378 267297
rect 470378 267267 470390 267297
rect 470390 267267 470412 267297
rect 470436 267267 470442 267297
rect 470442 267267 470454 267297
rect 470454 267267 470492 267297
rect 470516 267267 470518 267297
rect 470518 267267 470570 267297
rect 470570 267267 470572 267297
rect 470596 267267 470634 267297
rect 470634 267267 470646 267297
rect 470646 267267 470652 267297
rect 470676 267267 470698 267297
rect 470698 267267 470710 267297
rect 470710 267267 470732 267297
rect 470756 267267 470762 267297
rect 470762 267267 470774 267297
rect 470774 267267 470812 267297
rect 470276 267233 470332 267243
rect 470356 267233 470412 267243
rect 470436 267233 470492 267243
rect 470516 267233 470572 267243
rect 470596 267233 470652 267243
rect 470676 267233 470732 267243
rect 470756 267233 470812 267243
rect 470276 267187 470314 267233
rect 470314 267187 470326 267233
rect 470326 267187 470332 267233
rect 470356 267187 470378 267233
rect 470378 267187 470390 267233
rect 470390 267187 470412 267233
rect 470436 267187 470442 267233
rect 470442 267187 470454 267233
rect 470454 267187 470492 267233
rect 470516 267187 470518 267233
rect 470518 267187 470570 267233
rect 470570 267187 470572 267233
rect 470596 267187 470634 267233
rect 470634 267187 470646 267233
rect 470646 267187 470652 267233
rect 470676 267187 470698 267233
rect 470698 267187 470710 267233
rect 470710 267187 470732 267233
rect 470756 267187 470762 267233
rect 470762 267187 470774 267233
rect 470774 267187 470812 267233
rect 485502 272586 485558 272642
rect 482374 267282 482430 267338
rect 485502 267282 485558 267338
rect 482374 267010 482430 267066
rect 485410 267010 485466 267066
rect 488446 267010 488502 267066
rect 469036 266351 469074 266397
rect 469074 266351 469086 266397
rect 469086 266351 469092 266397
rect 469116 266351 469138 266397
rect 469138 266351 469150 266397
rect 469150 266351 469172 266397
rect 469196 266351 469202 266397
rect 469202 266351 469214 266397
rect 469214 266351 469252 266397
rect 469276 266351 469278 266397
rect 469278 266351 469330 266397
rect 469330 266351 469332 266397
rect 469356 266351 469394 266397
rect 469394 266351 469406 266397
rect 469406 266351 469412 266397
rect 469436 266351 469458 266397
rect 469458 266351 469470 266397
rect 469470 266351 469492 266397
rect 469516 266351 469522 266397
rect 469522 266351 469534 266397
rect 469534 266351 469572 266397
rect 469036 266341 469092 266351
rect 469116 266341 469172 266351
rect 469196 266341 469252 266351
rect 469276 266341 469332 266351
rect 469356 266341 469412 266351
rect 469436 266341 469492 266351
rect 469516 266341 469572 266351
rect 469036 266287 469074 266317
rect 469074 266287 469086 266317
rect 469086 266287 469092 266317
rect 469116 266287 469138 266317
rect 469138 266287 469150 266317
rect 469150 266287 469172 266317
rect 469196 266287 469202 266317
rect 469202 266287 469214 266317
rect 469214 266287 469252 266317
rect 469276 266287 469278 266317
rect 469278 266287 469330 266317
rect 469330 266287 469332 266317
rect 469356 266287 469394 266317
rect 469394 266287 469406 266317
rect 469406 266287 469412 266317
rect 469436 266287 469458 266317
rect 469458 266287 469470 266317
rect 469470 266287 469492 266317
rect 469516 266287 469522 266317
rect 469522 266287 469534 266317
rect 469534 266287 469572 266317
rect 469036 266275 469092 266287
rect 469116 266275 469172 266287
rect 469196 266275 469252 266287
rect 469276 266275 469332 266287
rect 469356 266275 469412 266287
rect 469436 266275 469492 266287
rect 469516 266275 469572 266287
rect 469036 266261 469074 266275
rect 469074 266261 469086 266275
rect 469086 266261 469092 266275
rect 469116 266261 469138 266275
rect 469138 266261 469150 266275
rect 469150 266261 469172 266275
rect 469196 266261 469202 266275
rect 469202 266261 469214 266275
rect 469214 266261 469252 266275
rect 469276 266261 469278 266275
rect 469278 266261 469330 266275
rect 469330 266261 469332 266275
rect 469356 266261 469394 266275
rect 469394 266261 469406 266275
rect 469406 266261 469412 266275
rect 469436 266261 469458 266275
rect 469458 266261 469470 266275
rect 469470 266261 469492 266275
rect 469516 266261 469522 266275
rect 469522 266261 469534 266275
rect 469534 266261 469572 266275
rect 469036 266223 469074 266237
rect 469074 266223 469086 266237
rect 469086 266223 469092 266237
rect 469116 266223 469138 266237
rect 469138 266223 469150 266237
rect 469150 266223 469172 266237
rect 469196 266223 469202 266237
rect 469202 266223 469214 266237
rect 469214 266223 469252 266237
rect 469276 266223 469278 266237
rect 469278 266223 469330 266237
rect 469330 266223 469332 266237
rect 469356 266223 469394 266237
rect 469394 266223 469406 266237
rect 469406 266223 469412 266237
rect 469436 266223 469458 266237
rect 469458 266223 469470 266237
rect 469470 266223 469492 266237
rect 469516 266223 469522 266237
rect 469522 266223 469534 266237
rect 469534 266223 469572 266237
rect 469036 266211 469092 266223
rect 469116 266211 469172 266223
rect 469196 266211 469252 266223
rect 469276 266211 469332 266223
rect 469356 266211 469412 266223
rect 469436 266211 469492 266223
rect 469516 266211 469572 266223
rect 469036 266181 469074 266211
rect 469074 266181 469086 266211
rect 469086 266181 469092 266211
rect 469116 266181 469138 266211
rect 469138 266181 469150 266211
rect 469150 266181 469172 266211
rect 469196 266181 469202 266211
rect 469202 266181 469214 266211
rect 469214 266181 469252 266211
rect 469276 266181 469278 266211
rect 469278 266181 469330 266211
rect 469330 266181 469332 266211
rect 469356 266181 469394 266211
rect 469394 266181 469406 266211
rect 469406 266181 469412 266211
rect 469436 266181 469458 266211
rect 469458 266181 469470 266211
rect 469470 266181 469492 266211
rect 469516 266181 469522 266211
rect 469522 266181 469534 266211
rect 469534 266181 469572 266211
rect 469036 266147 469092 266157
rect 469116 266147 469172 266157
rect 469196 266147 469252 266157
rect 469276 266147 469332 266157
rect 469356 266147 469412 266157
rect 469436 266147 469492 266157
rect 469516 266147 469572 266157
rect 469036 266101 469074 266147
rect 469074 266101 469086 266147
rect 469086 266101 469092 266147
rect 469116 266101 469138 266147
rect 469138 266101 469150 266147
rect 469150 266101 469172 266147
rect 469196 266101 469202 266147
rect 469202 266101 469214 266147
rect 469214 266101 469252 266147
rect 469276 266101 469278 266147
rect 469278 266101 469330 266147
rect 469330 266101 469332 266147
rect 469356 266101 469394 266147
rect 469394 266101 469406 266147
rect 469406 266101 469412 266147
rect 469436 266101 469458 266147
rect 469458 266101 469470 266147
rect 469470 266101 469492 266147
rect 469516 266101 469522 266147
rect 469522 266101 469534 266147
rect 469534 266101 469572 266147
rect 479062 265922 479118 265978
rect 470276 265264 470314 265310
rect 470314 265264 470326 265310
rect 470326 265264 470332 265310
rect 470356 265264 470378 265310
rect 470378 265264 470390 265310
rect 470390 265264 470412 265310
rect 470436 265264 470442 265310
rect 470442 265264 470454 265310
rect 470454 265264 470492 265310
rect 470516 265264 470518 265310
rect 470518 265264 470570 265310
rect 470570 265264 470572 265310
rect 470596 265264 470634 265310
rect 470634 265264 470646 265310
rect 470646 265264 470652 265310
rect 470676 265264 470698 265310
rect 470698 265264 470710 265310
rect 470710 265264 470732 265310
rect 470756 265264 470762 265310
rect 470762 265264 470774 265310
rect 470774 265264 470812 265310
rect 470276 265254 470332 265264
rect 470356 265254 470412 265264
rect 470436 265254 470492 265264
rect 470516 265254 470572 265264
rect 470596 265254 470652 265264
rect 470676 265254 470732 265264
rect 470756 265254 470812 265264
rect 470276 265200 470314 265230
rect 470314 265200 470326 265230
rect 470326 265200 470332 265230
rect 470356 265200 470378 265230
rect 470378 265200 470390 265230
rect 470390 265200 470412 265230
rect 470436 265200 470442 265230
rect 470442 265200 470454 265230
rect 470454 265200 470492 265230
rect 470516 265200 470518 265230
rect 470518 265200 470570 265230
rect 470570 265200 470572 265230
rect 470596 265200 470634 265230
rect 470634 265200 470646 265230
rect 470646 265200 470652 265230
rect 470676 265200 470698 265230
rect 470698 265200 470710 265230
rect 470710 265200 470732 265230
rect 470756 265200 470762 265230
rect 470762 265200 470774 265230
rect 470774 265200 470812 265230
rect 470276 265188 470332 265200
rect 470356 265188 470412 265200
rect 470436 265188 470492 265200
rect 470516 265188 470572 265200
rect 470596 265188 470652 265200
rect 470676 265188 470732 265200
rect 470756 265188 470812 265200
rect 470276 265174 470314 265188
rect 470314 265174 470326 265188
rect 470326 265174 470332 265188
rect 470356 265174 470378 265188
rect 470378 265174 470390 265188
rect 470390 265174 470412 265188
rect 470436 265174 470442 265188
rect 470442 265174 470454 265188
rect 470454 265174 470492 265188
rect 470516 265174 470518 265188
rect 470518 265174 470570 265188
rect 470570 265174 470572 265188
rect 470596 265174 470634 265188
rect 470634 265174 470646 265188
rect 470646 265174 470652 265188
rect 470676 265174 470698 265188
rect 470698 265174 470710 265188
rect 470710 265174 470732 265188
rect 470756 265174 470762 265188
rect 470762 265174 470774 265188
rect 470774 265174 470812 265188
rect 470276 265136 470314 265150
rect 470314 265136 470326 265150
rect 470326 265136 470332 265150
rect 470356 265136 470378 265150
rect 470378 265136 470390 265150
rect 470390 265136 470412 265150
rect 470436 265136 470442 265150
rect 470442 265136 470454 265150
rect 470454 265136 470492 265150
rect 470516 265136 470518 265150
rect 470518 265136 470570 265150
rect 470570 265136 470572 265150
rect 470596 265136 470634 265150
rect 470634 265136 470646 265150
rect 470646 265136 470652 265150
rect 470676 265136 470698 265150
rect 470698 265136 470710 265150
rect 470710 265136 470732 265150
rect 470756 265136 470762 265150
rect 470762 265136 470774 265150
rect 470774 265136 470812 265150
rect 470276 265124 470332 265136
rect 470356 265124 470412 265136
rect 470436 265124 470492 265136
rect 470516 265124 470572 265136
rect 470596 265124 470652 265136
rect 470676 265124 470732 265136
rect 470756 265124 470812 265136
rect 470276 265094 470314 265124
rect 470314 265094 470326 265124
rect 470326 265094 470332 265124
rect 470356 265094 470378 265124
rect 470378 265094 470390 265124
rect 470390 265094 470412 265124
rect 470436 265094 470442 265124
rect 470442 265094 470454 265124
rect 470454 265094 470492 265124
rect 470516 265094 470518 265124
rect 470518 265094 470570 265124
rect 470570 265094 470572 265124
rect 470596 265094 470634 265124
rect 470634 265094 470646 265124
rect 470646 265094 470652 265124
rect 470676 265094 470698 265124
rect 470698 265094 470710 265124
rect 470710 265094 470732 265124
rect 470756 265094 470762 265124
rect 470762 265094 470774 265124
rect 470774 265094 470812 265124
rect 470276 265060 470332 265070
rect 470356 265060 470412 265070
rect 470436 265060 470492 265070
rect 470516 265060 470572 265070
rect 470596 265060 470652 265070
rect 470676 265060 470732 265070
rect 470756 265060 470812 265070
rect 470276 265014 470314 265060
rect 470314 265014 470326 265060
rect 470326 265014 470332 265060
rect 470356 265014 470378 265060
rect 470378 265014 470390 265060
rect 470390 265014 470412 265060
rect 470436 265014 470442 265060
rect 470442 265014 470454 265060
rect 470454 265014 470492 265060
rect 470516 265014 470518 265060
rect 470518 265014 470570 265060
rect 470570 265014 470572 265060
rect 470596 265014 470634 265060
rect 470634 265014 470646 265060
rect 470646 265014 470652 265060
rect 470676 265014 470698 265060
rect 470698 265014 470710 265060
rect 470710 265014 470732 265060
rect 470756 265014 470762 265060
rect 470762 265014 470774 265060
rect 470774 265014 470812 265060
rect 476486 264970 476542 265026
rect 479522 264970 479578 265026
rect 535458 444762 535514 444818
rect 535458 443402 535514 443458
rect 535458 442042 535514 442098
rect 535458 440682 535514 440738
rect 535458 439322 535514 439378
rect 535458 437962 535514 438018
rect 535458 436602 535514 436658
rect 535458 435242 535514 435298
rect 535458 433882 535514 433938
rect 535458 432522 535514 432578
rect 546682 448026 546738 448082
rect 544198 447890 544254 447946
rect 539230 447754 539286 447810
rect 541714 447210 541770 447266
rect 536102 431162 536158 431218
rect 536746 424362 536802 424418
rect 535458 409266 535514 409322
rect 535458 406546 535514 406602
rect 535458 404506 535514 404562
rect 535458 403146 535514 403202
rect 536378 401650 536434 401706
rect 536286 400290 536342 400346
rect 535458 399066 535514 399122
rect 536102 397434 536158 397490
rect 535458 396346 535514 396402
rect 535458 372818 535514 372874
rect 535458 371458 535514 371514
rect 535458 368738 535514 368794
rect 535458 367378 535514 367434
rect 535458 366018 535514 366074
rect 535458 361938 535514 361994
rect 535458 336778 535514 336834
rect 535458 331338 535514 331394
rect 535458 329978 535514 330034
rect 536010 328618 536066 328674
rect 535458 325898 535514 325954
rect 535458 300774 535460 300794
rect 535460 300774 535512 300794
rect 535512 300774 535514 300794
rect 535458 300738 535514 300774
rect 535458 299414 535460 299434
rect 535460 299414 535512 299434
rect 535512 299414 535514 299434
rect 535458 299378 535514 299414
rect 535458 298054 535460 298074
rect 535460 298054 535512 298074
rect 535512 298054 535514 298074
rect 535458 298018 535514 298054
rect 535458 296658 535514 296714
rect 535550 295298 535606 295354
rect 535458 293938 535514 293994
rect 535550 292578 535606 292634
rect 535458 291218 535514 291274
rect 535458 289878 535514 289914
rect 535458 289858 535460 289878
rect 535460 289858 535512 289878
rect 535512 289858 535514 289878
rect 535458 288498 535514 288554
rect 536194 360578 536250 360634
rect 544198 445714 544254 445770
rect 541714 445306 541770 445362
rect 541714 409266 541770 409322
rect 544290 409266 544346 409322
rect 536746 395938 536802 395994
rect 536746 388322 536802 388378
rect 536562 364658 536618 364714
rect 536470 363298 536526 363354
rect 536378 324538 536434 324594
rect 536746 359218 536802 359274
rect 541714 373090 541770 373146
rect 544198 373090 544254 373146
rect 536746 352418 536802 352474
rect 536654 327258 536710 327314
rect 541714 339498 541770 339554
rect 544198 339498 544254 339554
rect 536746 323178 536802 323234
rect 536746 316378 536802 316434
rect 541714 303730 541770 303786
rect 544198 303730 544254 303786
rect 548062 699762 548118 699818
rect 577036 697860 577074 697906
rect 577074 697860 577086 697906
rect 577086 697860 577092 697906
rect 577116 697860 577138 697906
rect 577138 697860 577150 697906
rect 577150 697860 577172 697906
rect 577196 697860 577202 697906
rect 577202 697860 577214 697906
rect 577214 697860 577252 697906
rect 577276 697860 577278 697906
rect 577278 697860 577330 697906
rect 577330 697860 577332 697906
rect 577356 697860 577394 697906
rect 577394 697860 577406 697906
rect 577406 697860 577412 697906
rect 577436 697860 577458 697906
rect 577458 697860 577470 697906
rect 577470 697860 577492 697906
rect 577516 697860 577522 697906
rect 577522 697860 577534 697906
rect 577534 697860 577572 697906
rect 577036 697850 577092 697860
rect 577116 697850 577172 697860
rect 577196 697850 577252 697860
rect 577276 697850 577332 697860
rect 577356 697850 577412 697860
rect 577436 697850 577492 697860
rect 577516 697850 577572 697860
rect 577036 697796 577074 697826
rect 577074 697796 577086 697826
rect 577086 697796 577092 697826
rect 577116 697796 577138 697826
rect 577138 697796 577150 697826
rect 577150 697796 577172 697826
rect 577196 697796 577202 697826
rect 577202 697796 577214 697826
rect 577214 697796 577252 697826
rect 577276 697796 577278 697826
rect 577278 697796 577330 697826
rect 577330 697796 577332 697826
rect 577356 697796 577394 697826
rect 577394 697796 577406 697826
rect 577406 697796 577412 697826
rect 577436 697796 577458 697826
rect 577458 697796 577470 697826
rect 577470 697796 577492 697826
rect 577516 697796 577522 697826
rect 577522 697796 577534 697826
rect 577534 697796 577572 697826
rect 577036 697784 577092 697796
rect 577116 697784 577172 697796
rect 577196 697784 577252 697796
rect 577276 697784 577332 697796
rect 577356 697784 577412 697796
rect 577436 697784 577492 697796
rect 577516 697784 577572 697796
rect 577036 697770 577074 697784
rect 577074 697770 577086 697784
rect 577086 697770 577092 697784
rect 577116 697770 577138 697784
rect 577138 697770 577150 697784
rect 577150 697770 577172 697784
rect 577196 697770 577202 697784
rect 577202 697770 577214 697784
rect 577214 697770 577252 697784
rect 577276 697770 577278 697784
rect 577278 697770 577330 697784
rect 577330 697770 577332 697784
rect 577356 697770 577394 697784
rect 577394 697770 577406 697784
rect 577406 697770 577412 697784
rect 577436 697770 577458 697784
rect 577458 697770 577470 697784
rect 577470 697770 577492 697784
rect 577516 697770 577522 697784
rect 577522 697770 577534 697784
rect 577534 697770 577572 697784
rect 577036 697732 577074 697746
rect 577074 697732 577086 697746
rect 577086 697732 577092 697746
rect 577116 697732 577138 697746
rect 577138 697732 577150 697746
rect 577150 697732 577172 697746
rect 577196 697732 577202 697746
rect 577202 697732 577214 697746
rect 577214 697732 577252 697746
rect 577276 697732 577278 697746
rect 577278 697732 577330 697746
rect 577330 697732 577332 697746
rect 577356 697732 577394 697746
rect 577394 697732 577406 697746
rect 577406 697732 577412 697746
rect 577436 697732 577458 697746
rect 577458 697732 577470 697746
rect 577470 697732 577492 697746
rect 577516 697732 577522 697746
rect 577522 697732 577534 697746
rect 577534 697732 577572 697746
rect 577036 697720 577092 697732
rect 577116 697720 577172 697732
rect 577196 697720 577252 697732
rect 577276 697720 577332 697732
rect 577356 697720 577412 697732
rect 577436 697720 577492 697732
rect 577516 697720 577572 697732
rect 577036 697690 577074 697720
rect 577074 697690 577086 697720
rect 577086 697690 577092 697720
rect 577116 697690 577138 697720
rect 577138 697690 577150 697720
rect 577150 697690 577172 697720
rect 577196 697690 577202 697720
rect 577202 697690 577214 697720
rect 577214 697690 577252 697720
rect 577276 697690 577278 697720
rect 577278 697690 577330 697720
rect 577330 697690 577332 697720
rect 577356 697690 577394 697720
rect 577394 697690 577406 697720
rect 577406 697690 577412 697720
rect 577436 697690 577458 697720
rect 577458 697690 577470 697720
rect 577470 697690 577492 697720
rect 577516 697690 577522 697720
rect 577522 697690 577534 697720
rect 577534 697690 577572 697720
rect 577036 697656 577092 697666
rect 577116 697656 577172 697666
rect 577196 697656 577252 697666
rect 577276 697656 577332 697666
rect 577356 697656 577412 697666
rect 577436 697656 577492 697666
rect 577516 697656 577572 697666
rect 577036 697610 577074 697656
rect 577074 697610 577086 697656
rect 577086 697610 577092 697656
rect 577116 697610 577138 697656
rect 577138 697610 577150 697656
rect 577150 697610 577172 697656
rect 577196 697610 577202 697656
rect 577202 697610 577214 697656
rect 577214 697610 577252 697656
rect 577276 697610 577278 697656
rect 577278 697610 577330 697656
rect 577330 697610 577332 697656
rect 577356 697610 577394 697656
rect 577394 697610 577406 697656
rect 577406 697610 577412 697656
rect 577436 697610 577458 697656
rect 577458 697610 577470 697656
rect 577470 697610 577492 697656
rect 577516 697610 577522 697656
rect 577522 697610 577534 697656
rect 577534 697610 577572 697656
rect 576605 697230 576661 697235
rect 576605 697179 576655 697230
rect 576655 697179 576661 697230
rect 580906 697178 580962 697234
rect 578276 697065 578314 697111
rect 578314 697065 578326 697111
rect 578326 697065 578332 697111
rect 578356 697065 578378 697111
rect 578378 697065 578390 697111
rect 578390 697065 578412 697111
rect 578436 697065 578442 697111
rect 578442 697065 578454 697111
rect 578454 697065 578492 697111
rect 578516 697065 578518 697111
rect 578518 697065 578570 697111
rect 578570 697065 578572 697111
rect 578596 697065 578634 697111
rect 578634 697065 578646 697111
rect 578646 697065 578652 697111
rect 578676 697065 578698 697111
rect 578698 697065 578710 697111
rect 578710 697065 578732 697111
rect 578756 697065 578762 697111
rect 578762 697065 578774 697111
rect 578774 697065 578812 697111
rect 578276 697055 578332 697065
rect 578356 697055 578412 697065
rect 578436 697055 578492 697065
rect 578516 697055 578572 697065
rect 578596 697055 578652 697065
rect 578676 697055 578732 697065
rect 578756 697055 578812 697065
rect 578276 697001 578314 697031
rect 578314 697001 578326 697031
rect 578326 697001 578332 697031
rect 578356 697001 578378 697031
rect 578378 697001 578390 697031
rect 578390 697001 578412 697031
rect 578436 697001 578442 697031
rect 578442 697001 578454 697031
rect 578454 697001 578492 697031
rect 578516 697001 578518 697031
rect 578518 697001 578570 697031
rect 578570 697001 578572 697031
rect 578596 697001 578634 697031
rect 578634 697001 578646 697031
rect 578646 697001 578652 697031
rect 578676 697001 578698 697031
rect 578698 697001 578710 697031
rect 578710 697001 578732 697031
rect 578756 697001 578762 697031
rect 578762 697001 578774 697031
rect 578774 697001 578812 697031
rect 578276 696989 578332 697001
rect 578356 696989 578412 697001
rect 578436 696989 578492 697001
rect 578516 696989 578572 697001
rect 578596 696989 578652 697001
rect 578676 696989 578732 697001
rect 578756 696989 578812 697001
rect 578276 696975 578314 696989
rect 578314 696975 578326 696989
rect 578326 696975 578332 696989
rect 578356 696975 578378 696989
rect 578378 696975 578390 696989
rect 578390 696975 578412 696989
rect 578436 696975 578442 696989
rect 578442 696975 578454 696989
rect 578454 696975 578492 696989
rect 578516 696975 578518 696989
rect 578518 696975 578570 696989
rect 578570 696975 578572 696989
rect 578596 696975 578634 696989
rect 578634 696975 578646 696989
rect 578646 696975 578652 696989
rect 578676 696975 578698 696989
rect 578698 696975 578710 696989
rect 578710 696975 578732 696989
rect 578756 696975 578762 696989
rect 578762 696975 578774 696989
rect 578774 696975 578812 696989
rect 578276 696937 578314 696951
rect 578314 696937 578326 696951
rect 578326 696937 578332 696951
rect 578356 696937 578378 696951
rect 578378 696937 578390 696951
rect 578390 696937 578412 696951
rect 578436 696937 578442 696951
rect 578442 696937 578454 696951
rect 578454 696937 578492 696951
rect 578516 696937 578518 696951
rect 578518 696937 578570 696951
rect 578570 696937 578572 696951
rect 578596 696937 578634 696951
rect 578634 696937 578646 696951
rect 578646 696937 578652 696951
rect 578676 696937 578698 696951
rect 578698 696937 578710 696951
rect 578710 696937 578732 696951
rect 578756 696937 578762 696951
rect 578762 696937 578774 696951
rect 578774 696937 578812 696951
rect 578276 696925 578332 696937
rect 578356 696925 578412 696937
rect 578436 696925 578492 696937
rect 578516 696925 578572 696937
rect 578596 696925 578652 696937
rect 578676 696925 578732 696937
rect 578756 696925 578812 696937
rect 578276 696895 578314 696925
rect 578314 696895 578326 696925
rect 578326 696895 578332 696925
rect 578356 696895 578378 696925
rect 578378 696895 578390 696925
rect 578390 696895 578412 696925
rect 578436 696895 578442 696925
rect 578442 696895 578454 696925
rect 578454 696895 578492 696925
rect 578516 696895 578518 696925
rect 578518 696895 578570 696925
rect 578570 696895 578572 696925
rect 578596 696895 578634 696925
rect 578634 696895 578646 696925
rect 578646 696895 578652 696925
rect 578676 696895 578698 696925
rect 578698 696895 578710 696925
rect 578710 696895 578732 696925
rect 578756 696895 578762 696925
rect 578762 696895 578774 696925
rect 578774 696895 578812 696925
rect 578276 696861 578332 696871
rect 578356 696861 578412 696871
rect 578436 696861 578492 696871
rect 578516 696861 578572 696871
rect 578596 696861 578652 696871
rect 578676 696861 578732 696871
rect 578756 696861 578812 696871
rect 578276 696815 578314 696861
rect 578314 696815 578326 696861
rect 578326 696815 578332 696861
rect 578356 696815 578378 696861
rect 578378 696815 578390 696861
rect 578390 696815 578412 696861
rect 578436 696815 578442 696861
rect 578442 696815 578454 696861
rect 578454 696815 578492 696861
rect 578516 696815 578518 696861
rect 578518 696815 578570 696861
rect 578570 696815 578572 696861
rect 578596 696815 578634 696861
rect 578634 696815 578646 696861
rect 578646 696815 578652 696861
rect 578676 696815 578698 696861
rect 578698 696815 578710 696861
rect 578710 696815 578732 696861
rect 578756 696815 578762 696861
rect 578762 696815 578774 696861
rect 578774 696815 578812 696861
rect 580262 670658 580318 670714
rect 577036 644684 577074 644730
rect 577074 644684 577086 644730
rect 577086 644684 577092 644730
rect 577116 644684 577138 644730
rect 577138 644684 577150 644730
rect 577150 644684 577172 644730
rect 577196 644684 577202 644730
rect 577202 644684 577214 644730
rect 577214 644684 577252 644730
rect 577276 644684 577278 644730
rect 577278 644684 577330 644730
rect 577330 644684 577332 644730
rect 577356 644684 577394 644730
rect 577394 644684 577406 644730
rect 577406 644684 577412 644730
rect 577436 644684 577458 644730
rect 577458 644684 577470 644730
rect 577470 644684 577492 644730
rect 577516 644684 577522 644730
rect 577522 644684 577534 644730
rect 577534 644684 577572 644730
rect 577036 644674 577092 644684
rect 577116 644674 577172 644684
rect 577196 644674 577252 644684
rect 577276 644674 577332 644684
rect 577356 644674 577412 644684
rect 577436 644674 577492 644684
rect 577516 644674 577572 644684
rect 577036 644620 577074 644650
rect 577074 644620 577086 644650
rect 577086 644620 577092 644650
rect 577116 644620 577138 644650
rect 577138 644620 577150 644650
rect 577150 644620 577172 644650
rect 577196 644620 577202 644650
rect 577202 644620 577214 644650
rect 577214 644620 577252 644650
rect 577276 644620 577278 644650
rect 577278 644620 577330 644650
rect 577330 644620 577332 644650
rect 577356 644620 577394 644650
rect 577394 644620 577406 644650
rect 577406 644620 577412 644650
rect 577436 644620 577458 644650
rect 577458 644620 577470 644650
rect 577470 644620 577492 644650
rect 577516 644620 577522 644650
rect 577522 644620 577534 644650
rect 577534 644620 577572 644650
rect 577036 644608 577092 644620
rect 577116 644608 577172 644620
rect 577196 644608 577252 644620
rect 577276 644608 577332 644620
rect 577356 644608 577412 644620
rect 577436 644608 577492 644620
rect 577516 644608 577572 644620
rect 577036 644594 577074 644608
rect 577074 644594 577086 644608
rect 577086 644594 577092 644608
rect 577116 644594 577138 644608
rect 577138 644594 577150 644608
rect 577150 644594 577172 644608
rect 577196 644594 577202 644608
rect 577202 644594 577214 644608
rect 577214 644594 577252 644608
rect 577276 644594 577278 644608
rect 577278 644594 577330 644608
rect 577330 644594 577332 644608
rect 577356 644594 577394 644608
rect 577394 644594 577406 644608
rect 577406 644594 577412 644608
rect 577436 644594 577458 644608
rect 577458 644594 577470 644608
rect 577470 644594 577492 644608
rect 577516 644594 577522 644608
rect 577522 644594 577534 644608
rect 577534 644594 577572 644608
rect 577036 644556 577074 644570
rect 577074 644556 577086 644570
rect 577086 644556 577092 644570
rect 577116 644556 577138 644570
rect 577138 644556 577150 644570
rect 577150 644556 577172 644570
rect 577196 644556 577202 644570
rect 577202 644556 577214 644570
rect 577214 644556 577252 644570
rect 577276 644556 577278 644570
rect 577278 644556 577330 644570
rect 577330 644556 577332 644570
rect 577356 644556 577394 644570
rect 577394 644556 577406 644570
rect 577406 644556 577412 644570
rect 577436 644556 577458 644570
rect 577458 644556 577470 644570
rect 577470 644556 577492 644570
rect 577516 644556 577522 644570
rect 577522 644556 577534 644570
rect 577534 644556 577572 644570
rect 577036 644544 577092 644556
rect 577116 644544 577172 644556
rect 577196 644544 577252 644556
rect 577276 644544 577332 644556
rect 577356 644544 577412 644556
rect 577436 644544 577492 644556
rect 577516 644544 577572 644556
rect 577036 644514 577074 644544
rect 577074 644514 577086 644544
rect 577086 644514 577092 644544
rect 577116 644514 577138 644544
rect 577138 644514 577150 644544
rect 577150 644514 577172 644544
rect 577196 644514 577202 644544
rect 577202 644514 577214 644544
rect 577214 644514 577252 644544
rect 577276 644514 577278 644544
rect 577278 644514 577330 644544
rect 577330 644514 577332 644544
rect 577356 644514 577394 644544
rect 577394 644514 577406 644544
rect 577406 644514 577412 644544
rect 577436 644514 577458 644544
rect 577458 644514 577470 644544
rect 577470 644514 577492 644544
rect 577516 644514 577522 644544
rect 577522 644514 577534 644544
rect 577534 644514 577572 644544
rect 577036 644480 577092 644490
rect 577116 644480 577172 644490
rect 577196 644480 577252 644490
rect 577276 644480 577332 644490
rect 577356 644480 577412 644490
rect 577436 644480 577492 644490
rect 577516 644480 577572 644490
rect 577036 644434 577074 644480
rect 577074 644434 577086 644480
rect 577086 644434 577092 644480
rect 577116 644434 577138 644480
rect 577138 644434 577150 644480
rect 577150 644434 577172 644480
rect 577196 644434 577202 644480
rect 577202 644434 577214 644480
rect 577214 644434 577252 644480
rect 577276 644434 577278 644480
rect 577278 644434 577330 644480
rect 577330 644434 577332 644480
rect 577356 644434 577394 644480
rect 577394 644434 577406 644480
rect 577406 644434 577412 644480
rect 577436 644434 577458 644480
rect 577458 644434 577470 644480
rect 577470 644434 577492 644480
rect 577516 644434 577522 644480
rect 577522 644434 577534 644480
rect 577534 644434 577572 644480
rect 576605 644054 576661 644059
rect 576605 644003 576655 644054
rect 576655 644003 576661 644054
rect 578276 643889 578314 643935
rect 578314 643889 578326 643935
rect 578326 643889 578332 643935
rect 578356 643889 578378 643935
rect 578378 643889 578390 643935
rect 578390 643889 578412 643935
rect 578436 643889 578442 643935
rect 578442 643889 578454 643935
rect 578454 643889 578492 643935
rect 578516 643889 578518 643935
rect 578518 643889 578570 643935
rect 578570 643889 578572 643935
rect 578596 643889 578634 643935
rect 578634 643889 578646 643935
rect 578646 643889 578652 643935
rect 578676 643889 578698 643935
rect 578698 643889 578710 643935
rect 578710 643889 578732 643935
rect 578756 643889 578762 643935
rect 578762 643889 578774 643935
rect 578774 643889 578812 643935
rect 578276 643879 578332 643889
rect 578356 643879 578412 643889
rect 578436 643879 578492 643889
rect 578516 643879 578572 643889
rect 578596 643879 578652 643889
rect 578676 643879 578732 643889
rect 578756 643879 578812 643889
rect 578276 643825 578314 643855
rect 578314 643825 578326 643855
rect 578326 643825 578332 643855
rect 578356 643825 578378 643855
rect 578378 643825 578390 643855
rect 578390 643825 578412 643855
rect 578436 643825 578442 643855
rect 578442 643825 578454 643855
rect 578454 643825 578492 643855
rect 578516 643825 578518 643855
rect 578518 643825 578570 643855
rect 578570 643825 578572 643855
rect 578596 643825 578634 643855
rect 578634 643825 578646 643855
rect 578646 643825 578652 643855
rect 578676 643825 578698 643855
rect 578698 643825 578710 643855
rect 578710 643825 578732 643855
rect 578756 643825 578762 643855
rect 578762 643825 578774 643855
rect 578774 643825 578812 643855
rect 578276 643813 578332 643825
rect 578356 643813 578412 643825
rect 578436 643813 578492 643825
rect 578516 643813 578572 643825
rect 578596 643813 578652 643825
rect 578676 643813 578732 643825
rect 578756 643813 578812 643825
rect 578276 643799 578314 643813
rect 578314 643799 578326 643813
rect 578326 643799 578332 643813
rect 578356 643799 578378 643813
rect 578378 643799 578390 643813
rect 578390 643799 578412 643813
rect 578436 643799 578442 643813
rect 578442 643799 578454 643813
rect 578454 643799 578492 643813
rect 578516 643799 578518 643813
rect 578518 643799 578570 643813
rect 578570 643799 578572 643813
rect 578596 643799 578634 643813
rect 578634 643799 578646 643813
rect 578646 643799 578652 643813
rect 578676 643799 578698 643813
rect 578698 643799 578710 643813
rect 578710 643799 578732 643813
rect 578756 643799 578762 643813
rect 578762 643799 578774 643813
rect 578774 643799 578812 643813
rect 578276 643761 578314 643775
rect 578314 643761 578326 643775
rect 578326 643761 578332 643775
rect 578356 643761 578378 643775
rect 578378 643761 578390 643775
rect 578390 643761 578412 643775
rect 578436 643761 578442 643775
rect 578442 643761 578454 643775
rect 578454 643761 578492 643775
rect 578516 643761 578518 643775
rect 578518 643761 578570 643775
rect 578570 643761 578572 643775
rect 578596 643761 578634 643775
rect 578634 643761 578646 643775
rect 578646 643761 578652 643775
rect 578676 643761 578698 643775
rect 578698 643761 578710 643775
rect 578710 643761 578732 643775
rect 578756 643761 578762 643775
rect 578762 643761 578774 643775
rect 578774 643761 578812 643775
rect 578276 643749 578332 643761
rect 578356 643749 578412 643761
rect 578436 643749 578492 643761
rect 578516 643749 578572 643761
rect 578596 643749 578652 643761
rect 578676 643749 578732 643761
rect 578756 643749 578812 643761
rect 578276 643719 578314 643749
rect 578314 643719 578326 643749
rect 578326 643719 578332 643749
rect 578356 643719 578378 643749
rect 578378 643719 578390 643749
rect 578390 643719 578412 643749
rect 578436 643719 578442 643749
rect 578442 643719 578454 643749
rect 578454 643719 578492 643749
rect 578516 643719 578518 643749
rect 578518 643719 578570 643749
rect 578570 643719 578572 643749
rect 578596 643719 578634 643749
rect 578634 643719 578646 643749
rect 578646 643719 578652 643749
rect 578676 643719 578698 643749
rect 578698 643719 578710 643749
rect 578710 643719 578732 643749
rect 578756 643719 578762 643749
rect 578762 643719 578774 643749
rect 578774 643719 578812 643749
rect 578276 643685 578332 643695
rect 578356 643685 578412 643695
rect 578436 643685 578492 643695
rect 578516 643685 578572 643695
rect 578596 643685 578652 643695
rect 578676 643685 578732 643695
rect 578756 643685 578812 643695
rect 578276 643639 578314 643685
rect 578314 643639 578326 643685
rect 578326 643639 578332 643685
rect 578356 643639 578378 643685
rect 578378 643639 578390 643685
rect 578390 643639 578412 643685
rect 578436 643639 578442 643685
rect 578442 643639 578454 643685
rect 578454 643639 578492 643685
rect 578516 643639 578518 643685
rect 578518 643639 578570 643685
rect 578570 643639 578572 643685
rect 578596 643639 578634 643685
rect 578634 643639 578646 643685
rect 578646 643639 578652 643685
rect 578676 643639 578698 643685
rect 578698 643639 578710 643685
rect 578710 643639 578732 643685
rect 578756 643639 578762 643685
rect 578762 643639 578774 643685
rect 578774 643639 578812 643685
rect 577036 591644 577074 591690
rect 577074 591644 577086 591690
rect 577086 591644 577092 591690
rect 577116 591644 577138 591690
rect 577138 591644 577150 591690
rect 577150 591644 577172 591690
rect 577196 591644 577202 591690
rect 577202 591644 577214 591690
rect 577214 591644 577252 591690
rect 577276 591644 577278 591690
rect 577278 591644 577330 591690
rect 577330 591644 577332 591690
rect 577356 591644 577394 591690
rect 577394 591644 577406 591690
rect 577406 591644 577412 591690
rect 577436 591644 577458 591690
rect 577458 591644 577470 591690
rect 577470 591644 577492 591690
rect 577516 591644 577522 591690
rect 577522 591644 577534 591690
rect 577534 591644 577572 591690
rect 577036 591634 577092 591644
rect 577116 591634 577172 591644
rect 577196 591634 577252 591644
rect 577276 591634 577332 591644
rect 577356 591634 577412 591644
rect 577436 591634 577492 591644
rect 577516 591634 577572 591644
rect 577036 591580 577074 591610
rect 577074 591580 577086 591610
rect 577086 591580 577092 591610
rect 577116 591580 577138 591610
rect 577138 591580 577150 591610
rect 577150 591580 577172 591610
rect 577196 591580 577202 591610
rect 577202 591580 577214 591610
rect 577214 591580 577252 591610
rect 577276 591580 577278 591610
rect 577278 591580 577330 591610
rect 577330 591580 577332 591610
rect 577356 591580 577394 591610
rect 577394 591580 577406 591610
rect 577406 591580 577412 591610
rect 577436 591580 577458 591610
rect 577458 591580 577470 591610
rect 577470 591580 577492 591610
rect 577516 591580 577522 591610
rect 577522 591580 577534 591610
rect 577534 591580 577572 591610
rect 577036 591568 577092 591580
rect 577116 591568 577172 591580
rect 577196 591568 577252 591580
rect 577276 591568 577332 591580
rect 577356 591568 577412 591580
rect 577436 591568 577492 591580
rect 577516 591568 577572 591580
rect 577036 591554 577074 591568
rect 577074 591554 577086 591568
rect 577086 591554 577092 591568
rect 577116 591554 577138 591568
rect 577138 591554 577150 591568
rect 577150 591554 577172 591568
rect 577196 591554 577202 591568
rect 577202 591554 577214 591568
rect 577214 591554 577252 591568
rect 577276 591554 577278 591568
rect 577278 591554 577330 591568
rect 577330 591554 577332 591568
rect 577356 591554 577394 591568
rect 577394 591554 577406 591568
rect 577406 591554 577412 591568
rect 577436 591554 577458 591568
rect 577458 591554 577470 591568
rect 577470 591554 577492 591568
rect 577516 591554 577522 591568
rect 577522 591554 577534 591568
rect 577534 591554 577572 591568
rect 577036 591516 577074 591530
rect 577074 591516 577086 591530
rect 577086 591516 577092 591530
rect 577116 591516 577138 591530
rect 577138 591516 577150 591530
rect 577150 591516 577172 591530
rect 577196 591516 577202 591530
rect 577202 591516 577214 591530
rect 577214 591516 577252 591530
rect 577276 591516 577278 591530
rect 577278 591516 577330 591530
rect 577330 591516 577332 591530
rect 577356 591516 577394 591530
rect 577394 591516 577406 591530
rect 577406 591516 577412 591530
rect 577436 591516 577458 591530
rect 577458 591516 577470 591530
rect 577470 591516 577492 591530
rect 577516 591516 577522 591530
rect 577522 591516 577534 591530
rect 577534 591516 577572 591530
rect 577036 591504 577092 591516
rect 577116 591504 577172 591516
rect 577196 591504 577252 591516
rect 577276 591504 577332 591516
rect 577356 591504 577412 591516
rect 577436 591504 577492 591516
rect 577516 591504 577572 591516
rect 577036 591474 577074 591504
rect 577074 591474 577086 591504
rect 577086 591474 577092 591504
rect 577116 591474 577138 591504
rect 577138 591474 577150 591504
rect 577150 591474 577172 591504
rect 577196 591474 577202 591504
rect 577202 591474 577214 591504
rect 577214 591474 577252 591504
rect 577276 591474 577278 591504
rect 577278 591474 577330 591504
rect 577330 591474 577332 591504
rect 577356 591474 577394 591504
rect 577394 591474 577406 591504
rect 577406 591474 577412 591504
rect 577436 591474 577458 591504
rect 577458 591474 577470 591504
rect 577470 591474 577492 591504
rect 577516 591474 577522 591504
rect 577522 591474 577534 591504
rect 577534 591474 577572 591504
rect 577036 591440 577092 591450
rect 577116 591440 577172 591450
rect 577196 591440 577252 591450
rect 577276 591440 577332 591450
rect 577356 591440 577412 591450
rect 577436 591440 577492 591450
rect 577516 591440 577572 591450
rect 577036 591394 577074 591440
rect 577074 591394 577086 591440
rect 577086 591394 577092 591440
rect 577116 591394 577138 591440
rect 577138 591394 577150 591440
rect 577150 591394 577172 591440
rect 577196 591394 577202 591440
rect 577202 591394 577214 591440
rect 577214 591394 577252 591440
rect 577276 591394 577278 591440
rect 577278 591394 577330 591440
rect 577330 591394 577332 591440
rect 577356 591394 577394 591440
rect 577394 591394 577406 591440
rect 577406 591394 577412 591440
rect 577436 591394 577458 591440
rect 577458 591394 577470 591440
rect 577470 591394 577492 591440
rect 577516 591394 577522 591440
rect 577522 591394 577534 591440
rect 577534 591394 577572 591440
rect 576605 591014 576661 591019
rect 576605 590963 576655 591014
rect 576655 590963 576661 591014
rect 578276 590849 578314 590895
rect 578314 590849 578326 590895
rect 578326 590849 578332 590895
rect 578356 590849 578378 590895
rect 578378 590849 578390 590895
rect 578390 590849 578412 590895
rect 578436 590849 578442 590895
rect 578442 590849 578454 590895
rect 578454 590849 578492 590895
rect 578516 590849 578518 590895
rect 578518 590849 578570 590895
rect 578570 590849 578572 590895
rect 578596 590849 578634 590895
rect 578634 590849 578646 590895
rect 578646 590849 578652 590895
rect 578676 590849 578698 590895
rect 578698 590849 578710 590895
rect 578710 590849 578732 590895
rect 578756 590849 578762 590895
rect 578762 590849 578774 590895
rect 578774 590849 578812 590895
rect 578276 590839 578332 590849
rect 578356 590839 578412 590849
rect 578436 590839 578492 590849
rect 578516 590839 578572 590849
rect 578596 590839 578652 590849
rect 578676 590839 578732 590849
rect 578756 590839 578812 590849
rect 578276 590785 578314 590815
rect 578314 590785 578326 590815
rect 578326 590785 578332 590815
rect 578356 590785 578378 590815
rect 578378 590785 578390 590815
rect 578390 590785 578412 590815
rect 578436 590785 578442 590815
rect 578442 590785 578454 590815
rect 578454 590785 578492 590815
rect 578516 590785 578518 590815
rect 578518 590785 578570 590815
rect 578570 590785 578572 590815
rect 578596 590785 578634 590815
rect 578634 590785 578646 590815
rect 578646 590785 578652 590815
rect 578676 590785 578698 590815
rect 578698 590785 578710 590815
rect 578710 590785 578732 590815
rect 578756 590785 578762 590815
rect 578762 590785 578774 590815
rect 578774 590785 578812 590815
rect 578276 590773 578332 590785
rect 578356 590773 578412 590785
rect 578436 590773 578492 590785
rect 578516 590773 578572 590785
rect 578596 590773 578652 590785
rect 578676 590773 578732 590785
rect 578756 590773 578812 590785
rect 578276 590759 578314 590773
rect 578314 590759 578326 590773
rect 578326 590759 578332 590773
rect 578356 590759 578378 590773
rect 578378 590759 578390 590773
rect 578390 590759 578412 590773
rect 578436 590759 578442 590773
rect 578442 590759 578454 590773
rect 578454 590759 578492 590773
rect 578516 590759 578518 590773
rect 578518 590759 578570 590773
rect 578570 590759 578572 590773
rect 578596 590759 578634 590773
rect 578634 590759 578646 590773
rect 578646 590759 578652 590773
rect 578676 590759 578698 590773
rect 578698 590759 578710 590773
rect 578710 590759 578732 590773
rect 578756 590759 578762 590773
rect 578762 590759 578774 590773
rect 578774 590759 578812 590773
rect 578276 590721 578314 590735
rect 578314 590721 578326 590735
rect 578326 590721 578332 590735
rect 578356 590721 578378 590735
rect 578378 590721 578390 590735
rect 578390 590721 578412 590735
rect 578436 590721 578442 590735
rect 578442 590721 578454 590735
rect 578454 590721 578492 590735
rect 578516 590721 578518 590735
rect 578518 590721 578570 590735
rect 578570 590721 578572 590735
rect 578596 590721 578634 590735
rect 578634 590721 578646 590735
rect 578646 590721 578652 590735
rect 578676 590721 578698 590735
rect 578698 590721 578710 590735
rect 578710 590721 578732 590735
rect 578756 590721 578762 590735
rect 578762 590721 578774 590735
rect 578774 590721 578812 590735
rect 578276 590709 578332 590721
rect 578356 590709 578412 590721
rect 578436 590709 578492 590721
rect 578516 590709 578572 590721
rect 578596 590709 578652 590721
rect 578676 590709 578732 590721
rect 578756 590709 578812 590721
rect 578276 590679 578314 590709
rect 578314 590679 578326 590709
rect 578326 590679 578332 590709
rect 578356 590679 578378 590709
rect 578378 590679 578390 590709
rect 578390 590679 578412 590709
rect 578436 590679 578442 590709
rect 578442 590679 578454 590709
rect 578454 590679 578492 590709
rect 578516 590679 578518 590709
rect 578518 590679 578570 590709
rect 578570 590679 578572 590709
rect 578596 590679 578634 590709
rect 578634 590679 578646 590709
rect 578646 590679 578652 590709
rect 578676 590679 578698 590709
rect 578698 590679 578710 590709
rect 578710 590679 578732 590709
rect 578756 590679 578762 590709
rect 578762 590679 578774 590709
rect 578774 590679 578812 590709
rect 578276 590645 578332 590655
rect 578356 590645 578412 590655
rect 578436 590645 578492 590655
rect 578516 590645 578572 590655
rect 578596 590645 578652 590655
rect 578676 590645 578732 590655
rect 578756 590645 578812 590655
rect 578276 590599 578314 590645
rect 578314 590599 578326 590645
rect 578326 590599 578332 590645
rect 578356 590599 578378 590645
rect 578378 590599 578390 590645
rect 578390 590599 578412 590645
rect 578436 590599 578442 590645
rect 578442 590599 578454 590645
rect 578454 590599 578492 590645
rect 578516 590599 578518 590645
rect 578518 590599 578570 590645
rect 578570 590599 578572 590645
rect 578596 590599 578634 590645
rect 578634 590599 578646 590645
rect 578646 590599 578652 590645
rect 578676 590599 578698 590645
rect 578698 590599 578710 590645
rect 578710 590599 578732 590645
rect 578756 590599 578762 590645
rect 578762 590599 578774 590645
rect 578774 590599 578812 590645
rect 577036 538468 577074 538514
rect 577074 538468 577086 538514
rect 577086 538468 577092 538514
rect 577116 538468 577138 538514
rect 577138 538468 577150 538514
rect 577150 538468 577172 538514
rect 577196 538468 577202 538514
rect 577202 538468 577214 538514
rect 577214 538468 577252 538514
rect 577276 538468 577278 538514
rect 577278 538468 577330 538514
rect 577330 538468 577332 538514
rect 577356 538468 577394 538514
rect 577394 538468 577406 538514
rect 577406 538468 577412 538514
rect 577436 538468 577458 538514
rect 577458 538468 577470 538514
rect 577470 538468 577492 538514
rect 577516 538468 577522 538514
rect 577522 538468 577534 538514
rect 577534 538468 577572 538514
rect 577036 538458 577092 538468
rect 577116 538458 577172 538468
rect 577196 538458 577252 538468
rect 577276 538458 577332 538468
rect 577356 538458 577412 538468
rect 577436 538458 577492 538468
rect 577516 538458 577572 538468
rect 577036 538404 577074 538434
rect 577074 538404 577086 538434
rect 577086 538404 577092 538434
rect 577116 538404 577138 538434
rect 577138 538404 577150 538434
rect 577150 538404 577172 538434
rect 577196 538404 577202 538434
rect 577202 538404 577214 538434
rect 577214 538404 577252 538434
rect 577276 538404 577278 538434
rect 577278 538404 577330 538434
rect 577330 538404 577332 538434
rect 577356 538404 577394 538434
rect 577394 538404 577406 538434
rect 577406 538404 577412 538434
rect 577436 538404 577458 538434
rect 577458 538404 577470 538434
rect 577470 538404 577492 538434
rect 577516 538404 577522 538434
rect 577522 538404 577534 538434
rect 577534 538404 577572 538434
rect 577036 538392 577092 538404
rect 577116 538392 577172 538404
rect 577196 538392 577252 538404
rect 577276 538392 577332 538404
rect 577356 538392 577412 538404
rect 577436 538392 577492 538404
rect 577516 538392 577572 538404
rect 577036 538378 577074 538392
rect 577074 538378 577086 538392
rect 577086 538378 577092 538392
rect 577116 538378 577138 538392
rect 577138 538378 577150 538392
rect 577150 538378 577172 538392
rect 577196 538378 577202 538392
rect 577202 538378 577214 538392
rect 577214 538378 577252 538392
rect 577276 538378 577278 538392
rect 577278 538378 577330 538392
rect 577330 538378 577332 538392
rect 577356 538378 577394 538392
rect 577394 538378 577406 538392
rect 577406 538378 577412 538392
rect 577436 538378 577458 538392
rect 577458 538378 577470 538392
rect 577470 538378 577492 538392
rect 577516 538378 577522 538392
rect 577522 538378 577534 538392
rect 577534 538378 577572 538392
rect 577036 538340 577074 538354
rect 577074 538340 577086 538354
rect 577086 538340 577092 538354
rect 577116 538340 577138 538354
rect 577138 538340 577150 538354
rect 577150 538340 577172 538354
rect 577196 538340 577202 538354
rect 577202 538340 577214 538354
rect 577214 538340 577252 538354
rect 577276 538340 577278 538354
rect 577278 538340 577330 538354
rect 577330 538340 577332 538354
rect 577356 538340 577394 538354
rect 577394 538340 577406 538354
rect 577406 538340 577412 538354
rect 577436 538340 577458 538354
rect 577458 538340 577470 538354
rect 577470 538340 577492 538354
rect 577516 538340 577522 538354
rect 577522 538340 577534 538354
rect 577534 538340 577572 538354
rect 577036 538328 577092 538340
rect 577116 538328 577172 538340
rect 577196 538328 577252 538340
rect 577276 538328 577332 538340
rect 577356 538328 577412 538340
rect 577436 538328 577492 538340
rect 577516 538328 577572 538340
rect 577036 538298 577074 538328
rect 577074 538298 577086 538328
rect 577086 538298 577092 538328
rect 577116 538298 577138 538328
rect 577138 538298 577150 538328
rect 577150 538298 577172 538328
rect 577196 538298 577202 538328
rect 577202 538298 577214 538328
rect 577214 538298 577252 538328
rect 577276 538298 577278 538328
rect 577278 538298 577330 538328
rect 577330 538298 577332 538328
rect 577356 538298 577394 538328
rect 577394 538298 577406 538328
rect 577406 538298 577412 538328
rect 577436 538298 577458 538328
rect 577458 538298 577470 538328
rect 577470 538298 577492 538328
rect 577516 538298 577522 538328
rect 577522 538298 577534 538328
rect 577534 538298 577572 538328
rect 577036 538264 577092 538274
rect 577116 538264 577172 538274
rect 577196 538264 577252 538274
rect 577276 538264 577332 538274
rect 577356 538264 577412 538274
rect 577436 538264 577492 538274
rect 577516 538264 577572 538274
rect 577036 538218 577074 538264
rect 577074 538218 577086 538264
rect 577086 538218 577092 538264
rect 577116 538218 577138 538264
rect 577138 538218 577150 538264
rect 577150 538218 577172 538264
rect 577196 538218 577202 538264
rect 577202 538218 577214 538264
rect 577214 538218 577252 538264
rect 577276 538218 577278 538264
rect 577278 538218 577330 538264
rect 577330 538218 577332 538264
rect 577356 538218 577394 538264
rect 577394 538218 577406 538264
rect 577406 538218 577412 538264
rect 577436 538218 577458 538264
rect 577458 538218 577470 538264
rect 577470 538218 577492 538264
rect 577516 538218 577522 538264
rect 577522 538218 577534 538264
rect 577534 538218 577572 538264
rect 576605 537838 576661 537843
rect 576605 537787 576655 537838
rect 576655 537787 576661 537838
rect 578276 537673 578314 537719
rect 578314 537673 578326 537719
rect 578326 537673 578332 537719
rect 578356 537673 578378 537719
rect 578378 537673 578390 537719
rect 578390 537673 578412 537719
rect 578436 537673 578442 537719
rect 578442 537673 578454 537719
rect 578454 537673 578492 537719
rect 578516 537673 578518 537719
rect 578518 537673 578570 537719
rect 578570 537673 578572 537719
rect 578596 537673 578634 537719
rect 578634 537673 578646 537719
rect 578646 537673 578652 537719
rect 578676 537673 578698 537719
rect 578698 537673 578710 537719
rect 578710 537673 578732 537719
rect 578756 537673 578762 537719
rect 578762 537673 578774 537719
rect 578774 537673 578812 537719
rect 578276 537663 578332 537673
rect 578356 537663 578412 537673
rect 578436 537663 578492 537673
rect 578516 537663 578572 537673
rect 578596 537663 578652 537673
rect 578676 537663 578732 537673
rect 578756 537663 578812 537673
rect 578276 537609 578314 537639
rect 578314 537609 578326 537639
rect 578326 537609 578332 537639
rect 578356 537609 578378 537639
rect 578378 537609 578390 537639
rect 578390 537609 578412 537639
rect 578436 537609 578442 537639
rect 578442 537609 578454 537639
rect 578454 537609 578492 537639
rect 578516 537609 578518 537639
rect 578518 537609 578570 537639
rect 578570 537609 578572 537639
rect 578596 537609 578634 537639
rect 578634 537609 578646 537639
rect 578646 537609 578652 537639
rect 578676 537609 578698 537639
rect 578698 537609 578710 537639
rect 578710 537609 578732 537639
rect 578756 537609 578762 537639
rect 578762 537609 578774 537639
rect 578774 537609 578812 537639
rect 578276 537597 578332 537609
rect 578356 537597 578412 537609
rect 578436 537597 578492 537609
rect 578516 537597 578572 537609
rect 578596 537597 578652 537609
rect 578676 537597 578732 537609
rect 578756 537597 578812 537609
rect 578276 537583 578314 537597
rect 578314 537583 578326 537597
rect 578326 537583 578332 537597
rect 578356 537583 578378 537597
rect 578378 537583 578390 537597
rect 578390 537583 578412 537597
rect 578436 537583 578442 537597
rect 578442 537583 578454 537597
rect 578454 537583 578492 537597
rect 578516 537583 578518 537597
rect 578518 537583 578570 537597
rect 578570 537583 578572 537597
rect 578596 537583 578634 537597
rect 578634 537583 578646 537597
rect 578646 537583 578652 537597
rect 578676 537583 578698 537597
rect 578698 537583 578710 537597
rect 578710 537583 578732 537597
rect 578756 537583 578762 537597
rect 578762 537583 578774 537597
rect 578774 537583 578812 537597
rect 578276 537545 578314 537559
rect 578314 537545 578326 537559
rect 578326 537545 578332 537559
rect 578356 537545 578378 537559
rect 578378 537545 578390 537559
rect 578390 537545 578412 537559
rect 578436 537545 578442 537559
rect 578442 537545 578454 537559
rect 578454 537545 578492 537559
rect 578516 537545 578518 537559
rect 578518 537545 578570 537559
rect 578570 537545 578572 537559
rect 578596 537545 578634 537559
rect 578634 537545 578646 537559
rect 578646 537545 578652 537559
rect 578676 537545 578698 537559
rect 578698 537545 578710 537559
rect 578710 537545 578732 537559
rect 578756 537545 578762 537559
rect 578762 537545 578774 537559
rect 578774 537545 578812 537559
rect 578276 537533 578332 537545
rect 578356 537533 578412 537545
rect 578436 537533 578492 537545
rect 578516 537533 578572 537545
rect 578596 537533 578652 537545
rect 578676 537533 578732 537545
rect 578756 537533 578812 537545
rect 578276 537503 578314 537533
rect 578314 537503 578326 537533
rect 578326 537503 578332 537533
rect 578356 537503 578378 537533
rect 578378 537503 578390 537533
rect 578390 537503 578412 537533
rect 578436 537503 578442 537533
rect 578442 537503 578454 537533
rect 578454 537503 578492 537533
rect 578516 537503 578518 537533
rect 578518 537503 578570 537533
rect 578570 537503 578572 537533
rect 578596 537503 578634 537533
rect 578634 537503 578646 537533
rect 578646 537503 578652 537533
rect 578676 537503 578698 537533
rect 578698 537503 578710 537533
rect 578710 537503 578732 537533
rect 578756 537503 578762 537533
rect 578762 537503 578774 537533
rect 578774 537503 578812 537533
rect 578276 537469 578332 537479
rect 578356 537469 578412 537479
rect 578436 537469 578492 537479
rect 578516 537469 578572 537479
rect 578596 537469 578652 537479
rect 578676 537469 578732 537479
rect 578756 537469 578812 537479
rect 578276 537423 578314 537469
rect 578314 537423 578326 537469
rect 578326 537423 578332 537469
rect 578356 537423 578378 537469
rect 578378 537423 578390 537469
rect 578390 537423 578412 537469
rect 578436 537423 578442 537469
rect 578442 537423 578454 537469
rect 578454 537423 578492 537469
rect 578516 537423 578518 537469
rect 578518 537423 578570 537469
rect 578570 537423 578572 537469
rect 578596 537423 578634 537469
rect 578634 537423 578646 537469
rect 578646 537423 578652 537469
rect 578676 537423 578698 537469
rect 578698 537423 578710 537469
rect 578710 537423 578732 537469
rect 578756 537423 578762 537469
rect 578762 537423 578774 537469
rect 578774 537423 578812 537469
rect 577036 485292 577074 485338
rect 577074 485292 577086 485338
rect 577086 485292 577092 485338
rect 577116 485292 577138 485338
rect 577138 485292 577150 485338
rect 577150 485292 577172 485338
rect 577196 485292 577202 485338
rect 577202 485292 577214 485338
rect 577214 485292 577252 485338
rect 577276 485292 577278 485338
rect 577278 485292 577330 485338
rect 577330 485292 577332 485338
rect 577356 485292 577394 485338
rect 577394 485292 577406 485338
rect 577406 485292 577412 485338
rect 577436 485292 577458 485338
rect 577458 485292 577470 485338
rect 577470 485292 577492 485338
rect 577516 485292 577522 485338
rect 577522 485292 577534 485338
rect 577534 485292 577572 485338
rect 577036 485282 577092 485292
rect 577116 485282 577172 485292
rect 577196 485282 577252 485292
rect 577276 485282 577332 485292
rect 577356 485282 577412 485292
rect 577436 485282 577492 485292
rect 577516 485282 577572 485292
rect 577036 485228 577074 485258
rect 577074 485228 577086 485258
rect 577086 485228 577092 485258
rect 577116 485228 577138 485258
rect 577138 485228 577150 485258
rect 577150 485228 577172 485258
rect 577196 485228 577202 485258
rect 577202 485228 577214 485258
rect 577214 485228 577252 485258
rect 577276 485228 577278 485258
rect 577278 485228 577330 485258
rect 577330 485228 577332 485258
rect 577356 485228 577394 485258
rect 577394 485228 577406 485258
rect 577406 485228 577412 485258
rect 577436 485228 577458 485258
rect 577458 485228 577470 485258
rect 577470 485228 577492 485258
rect 577516 485228 577522 485258
rect 577522 485228 577534 485258
rect 577534 485228 577572 485258
rect 577036 485216 577092 485228
rect 577116 485216 577172 485228
rect 577196 485216 577252 485228
rect 577276 485216 577332 485228
rect 577356 485216 577412 485228
rect 577436 485216 577492 485228
rect 577516 485216 577572 485228
rect 577036 485202 577074 485216
rect 577074 485202 577086 485216
rect 577086 485202 577092 485216
rect 577116 485202 577138 485216
rect 577138 485202 577150 485216
rect 577150 485202 577172 485216
rect 577196 485202 577202 485216
rect 577202 485202 577214 485216
rect 577214 485202 577252 485216
rect 577276 485202 577278 485216
rect 577278 485202 577330 485216
rect 577330 485202 577332 485216
rect 577356 485202 577394 485216
rect 577394 485202 577406 485216
rect 577406 485202 577412 485216
rect 577436 485202 577458 485216
rect 577458 485202 577470 485216
rect 577470 485202 577492 485216
rect 577516 485202 577522 485216
rect 577522 485202 577534 485216
rect 577534 485202 577572 485216
rect 577036 485164 577074 485178
rect 577074 485164 577086 485178
rect 577086 485164 577092 485178
rect 577116 485164 577138 485178
rect 577138 485164 577150 485178
rect 577150 485164 577172 485178
rect 577196 485164 577202 485178
rect 577202 485164 577214 485178
rect 577214 485164 577252 485178
rect 577276 485164 577278 485178
rect 577278 485164 577330 485178
rect 577330 485164 577332 485178
rect 577356 485164 577394 485178
rect 577394 485164 577406 485178
rect 577406 485164 577412 485178
rect 577436 485164 577458 485178
rect 577458 485164 577470 485178
rect 577470 485164 577492 485178
rect 577516 485164 577522 485178
rect 577522 485164 577534 485178
rect 577534 485164 577572 485178
rect 577036 485152 577092 485164
rect 577116 485152 577172 485164
rect 577196 485152 577252 485164
rect 577276 485152 577332 485164
rect 577356 485152 577412 485164
rect 577436 485152 577492 485164
rect 577516 485152 577572 485164
rect 577036 485122 577074 485152
rect 577074 485122 577086 485152
rect 577086 485122 577092 485152
rect 577116 485122 577138 485152
rect 577138 485122 577150 485152
rect 577150 485122 577172 485152
rect 577196 485122 577202 485152
rect 577202 485122 577214 485152
rect 577214 485122 577252 485152
rect 577276 485122 577278 485152
rect 577278 485122 577330 485152
rect 577330 485122 577332 485152
rect 577356 485122 577394 485152
rect 577394 485122 577406 485152
rect 577406 485122 577412 485152
rect 577436 485122 577458 485152
rect 577458 485122 577470 485152
rect 577470 485122 577492 485152
rect 577516 485122 577522 485152
rect 577522 485122 577534 485152
rect 577534 485122 577572 485152
rect 577036 485088 577092 485098
rect 577116 485088 577172 485098
rect 577196 485088 577252 485098
rect 577276 485088 577332 485098
rect 577356 485088 577412 485098
rect 577436 485088 577492 485098
rect 577516 485088 577572 485098
rect 577036 485042 577074 485088
rect 577074 485042 577086 485088
rect 577086 485042 577092 485088
rect 577116 485042 577138 485088
rect 577138 485042 577150 485088
rect 577150 485042 577172 485088
rect 577196 485042 577202 485088
rect 577202 485042 577214 485088
rect 577214 485042 577252 485088
rect 577276 485042 577278 485088
rect 577278 485042 577330 485088
rect 577330 485042 577332 485088
rect 577356 485042 577394 485088
rect 577394 485042 577406 485088
rect 577406 485042 577412 485088
rect 577436 485042 577458 485088
rect 577458 485042 577470 485088
rect 577470 485042 577492 485088
rect 577516 485042 577522 485088
rect 577522 485042 577534 485088
rect 577534 485042 577572 485088
rect 576605 484662 576661 484667
rect 576605 484611 576655 484662
rect 576655 484611 576661 484662
rect 578276 484497 578314 484543
rect 578314 484497 578326 484543
rect 578326 484497 578332 484543
rect 578356 484497 578378 484543
rect 578378 484497 578390 484543
rect 578390 484497 578412 484543
rect 578436 484497 578442 484543
rect 578442 484497 578454 484543
rect 578454 484497 578492 484543
rect 578516 484497 578518 484543
rect 578518 484497 578570 484543
rect 578570 484497 578572 484543
rect 578596 484497 578634 484543
rect 578634 484497 578646 484543
rect 578646 484497 578652 484543
rect 578676 484497 578698 484543
rect 578698 484497 578710 484543
rect 578710 484497 578732 484543
rect 578756 484497 578762 484543
rect 578762 484497 578774 484543
rect 578774 484497 578812 484543
rect 578276 484487 578332 484497
rect 578356 484487 578412 484497
rect 578436 484487 578492 484497
rect 578516 484487 578572 484497
rect 578596 484487 578652 484497
rect 578676 484487 578732 484497
rect 578756 484487 578812 484497
rect 578276 484433 578314 484463
rect 578314 484433 578326 484463
rect 578326 484433 578332 484463
rect 578356 484433 578378 484463
rect 578378 484433 578390 484463
rect 578390 484433 578412 484463
rect 578436 484433 578442 484463
rect 578442 484433 578454 484463
rect 578454 484433 578492 484463
rect 578516 484433 578518 484463
rect 578518 484433 578570 484463
rect 578570 484433 578572 484463
rect 578596 484433 578634 484463
rect 578634 484433 578646 484463
rect 578646 484433 578652 484463
rect 578676 484433 578698 484463
rect 578698 484433 578710 484463
rect 578710 484433 578732 484463
rect 578756 484433 578762 484463
rect 578762 484433 578774 484463
rect 578774 484433 578812 484463
rect 578276 484421 578332 484433
rect 578356 484421 578412 484433
rect 578436 484421 578492 484433
rect 578516 484421 578572 484433
rect 578596 484421 578652 484433
rect 578676 484421 578732 484433
rect 578756 484421 578812 484433
rect 578276 484407 578314 484421
rect 578314 484407 578326 484421
rect 578326 484407 578332 484421
rect 578356 484407 578378 484421
rect 578378 484407 578390 484421
rect 578390 484407 578412 484421
rect 578436 484407 578442 484421
rect 578442 484407 578454 484421
rect 578454 484407 578492 484421
rect 578516 484407 578518 484421
rect 578518 484407 578570 484421
rect 578570 484407 578572 484421
rect 578596 484407 578634 484421
rect 578634 484407 578646 484421
rect 578646 484407 578652 484421
rect 578676 484407 578698 484421
rect 578698 484407 578710 484421
rect 578710 484407 578732 484421
rect 578756 484407 578762 484421
rect 578762 484407 578774 484421
rect 578774 484407 578812 484421
rect 578276 484369 578314 484383
rect 578314 484369 578326 484383
rect 578326 484369 578332 484383
rect 578356 484369 578378 484383
rect 578378 484369 578390 484383
rect 578390 484369 578412 484383
rect 578436 484369 578442 484383
rect 578442 484369 578454 484383
rect 578454 484369 578492 484383
rect 578516 484369 578518 484383
rect 578518 484369 578570 484383
rect 578570 484369 578572 484383
rect 578596 484369 578634 484383
rect 578634 484369 578646 484383
rect 578646 484369 578652 484383
rect 578676 484369 578698 484383
rect 578698 484369 578710 484383
rect 578710 484369 578732 484383
rect 578756 484369 578762 484383
rect 578762 484369 578774 484383
rect 578774 484369 578812 484383
rect 578276 484357 578332 484369
rect 578356 484357 578412 484369
rect 578436 484357 578492 484369
rect 578516 484357 578572 484369
rect 578596 484357 578652 484369
rect 578676 484357 578732 484369
rect 578756 484357 578812 484369
rect 578276 484327 578314 484357
rect 578314 484327 578326 484357
rect 578326 484327 578332 484357
rect 578356 484327 578378 484357
rect 578378 484327 578390 484357
rect 578390 484327 578412 484357
rect 578436 484327 578442 484357
rect 578442 484327 578454 484357
rect 578454 484327 578492 484357
rect 578516 484327 578518 484357
rect 578518 484327 578570 484357
rect 578570 484327 578572 484357
rect 578596 484327 578634 484357
rect 578634 484327 578646 484357
rect 578646 484327 578652 484357
rect 578676 484327 578698 484357
rect 578698 484327 578710 484357
rect 578710 484327 578732 484357
rect 578756 484327 578762 484357
rect 578762 484327 578774 484357
rect 578774 484327 578812 484357
rect 578276 484293 578332 484303
rect 578356 484293 578412 484303
rect 578436 484293 578492 484303
rect 578516 484293 578572 484303
rect 578596 484293 578652 484303
rect 578676 484293 578732 484303
rect 578756 484293 578812 484303
rect 578276 484247 578314 484293
rect 578314 484247 578326 484293
rect 578326 484247 578332 484293
rect 578356 484247 578378 484293
rect 578378 484247 578390 484293
rect 578390 484247 578412 484293
rect 578436 484247 578442 484293
rect 578442 484247 578454 484293
rect 578454 484247 578492 484293
rect 578516 484247 578518 484293
rect 578518 484247 578570 484293
rect 578570 484247 578572 484293
rect 578596 484247 578634 484293
rect 578634 484247 578646 484293
rect 578646 484247 578652 484293
rect 578676 484247 578698 484293
rect 578698 484247 578710 484293
rect 578710 484247 578732 484293
rect 578756 484247 578762 484293
rect 578762 484247 578774 484293
rect 578774 484247 578812 484293
rect 580170 458090 580226 458146
rect 580906 644002 580962 644058
rect 580446 617482 580502 617538
rect 580262 448026 580318 448082
rect 580906 590962 580962 591018
rect 580630 564306 580686 564362
rect 580446 447890 580502 447946
rect 580906 537786 580962 537842
rect 580814 511266 580870 511322
rect 580906 484610 580962 484666
rect 580814 447754 580870 447810
rect 580630 447210 580686 447266
rect 548062 435378 548118 435434
rect 577036 432252 577074 432298
rect 577074 432252 577086 432298
rect 577086 432252 577092 432298
rect 577116 432252 577138 432298
rect 577138 432252 577150 432298
rect 577150 432252 577172 432298
rect 577196 432252 577202 432298
rect 577202 432252 577214 432298
rect 577214 432252 577252 432298
rect 577276 432252 577278 432298
rect 577278 432252 577330 432298
rect 577330 432252 577332 432298
rect 577356 432252 577394 432298
rect 577394 432252 577406 432298
rect 577406 432252 577412 432298
rect 577436 432252 577458 432298
rect 577458 432252 577470 432298
rect 577470 432252 577492 432298
rect 577516 432252 577522 432298
rect 577522 432252 577534 432298
rect 577534 432252 577572 432298
rect 577036 432242 577092 432252
rect 577116 432242 577172 432252
rect 577196 432242 577252 432252
rect 577276 432242 577332 432252
rect 577356 432242 577412 432252
rect 577436 432242 577492 432252
rect 577516 432242 577572 432252
rect 577036 432188 577074 432218
rect 577074 432188 577086 432218
rect 577086 432188 577092 432218
rect 577116 432188 577138 432218
rect 577138 432188 577150 432218
rect 577150 432188 577172 432218
rect 577196 432188 577202 432218
rect 577202 432188 577214 432218
rect 577214 432188 577252 432218
rect 577276 432188 577278 432218
rect 577278 432188 577330 432218
rect 577330 432188 577332 432218
rect 577356 432188 577394 432218
rect 577394 432188 577406 432218
rect 577406 432188 577412 432218
rect 577436 432188 577458 432218
rect 577458 432188 577470 432218
rect 577470 432188 577492 432218
rect 577516 432188 577522 432218
rect 577522 432188 577534 432218
rect 577534 432188 577572 432218
rect 577036 432176 577092 432188
rect 577116 432176 577172 432188
rect 577196 432176 577252 432188
rect 577276 432176 577332 432188
rect 577356 432176 577412 432188
rect 577436 432176 577492 432188
rect 577516 432176 577572 432188
rect 577036 432162 577074 432176
rect 577074 432162 577086 432176
rect 577086 432162 577092 432176
rect 577116 432162 577138 432176
rect 577138 432162 577150 432176
rect 577150 432162 577172 432176
rect 577196 432162 577202 432176
rect 577202 432162 577214 432176
rect 577214 432162 577252 432176
rect 577276 432162 577278 432176
rect 577278 432162 577330 432176
rect 577330 432162 577332 432176
rect 577356 432162 577394 432176
rect 577394 432162 577406 432176
rect 577406 432162 577412 432176
rect 577436 432162 577458 432176
rect 577458 432162 577470 432176
rect 577470 432162 577492 432176
rect 577516 432162 577522 432176
rect 577522 432162 577534 432176
rect 577534 432162 577572 432176
rect 577036 432124 577074 432138
rect 577074 432124 577086 432138
rect 577086 432124 577092 432138
rect 577116 432124 577138 432138
rect 577138 432124 577150 432138
rect 577150 432124 577172 432138
rect 577196 432124 577202 432138
rect 577202 432124 577214 432138
rect 577214 432124 577252 432138
rect 577276 432124 577278 432138
rect 577278 432124 577330 432138
rect 577330 432124 577332 432138
rect 577356 432124 577394 432138
rect 577394 432124 577406 432138
rect 577406 432124 577412 432138
rect 577436 432124 577458 432138
rect 577458 432124 577470 432138
rect 577470 432124 577492 432138
rect 577516 432124 577522 432138
rect 577522 432124 577534 432138
rect 577534 432124 577572 432138
rect 577036 432112 577092 432124
rect 577116 432112 577172 432124
rect 577196 432112 577252 432124
rect 577276 432112 577332 432124
rect 577356 432112 577412 432124
rect 577436 432112 577492 432124
rect 577516 432112 577572 432124
rect 577036 432082 577074 432112
rect 577074 432082 577086 432112
rect 577086 432082 577092 432112
rect 577116 432082 577138 432112
rect 577138 432082 577150 432112
rect 577150 432082 577172 432112
rect 577196 432082 577202 432112
rect 577202 432082 577214 432112
rect 577214 432082 577252 432112
rect 577276 432082 577278 432112
rect 577278 432082 577330 432112
rect 577330 432082 577332 432112
rect 577356 432082 577394 432112
rect 577394 432082 577406 432112
rect 577406 432082 577412 432112
rect 577436 432082 577458 432112
rect 577458 432082 577470 432112
rect 577470 432082 577492 432112
rect 577516 432082 577522 432112
rect 577522 432082 577534 432112
rect 577534 432082 577572 432112
rect 577036 432048 577092 432058
rect 577116 432048 577172 432058
rect 577196 432048 577252 432058
rect 577276 432048 577332 432058
rect 577356 432048 577412 432058
rect 577436 432048 577492 432058
rect 577516 432048 577572 432058
rect 577036 432002 577074 432048
rect 577074 432002 577086 432048
rect 577086 432002 577092 432048
rect 577116 432002 577138 432048
rect 577138 432002 577150 432048
rect 577150 432002 577172 432048
rect 577196 432002 577202 432048
rect 577202 432002 577214 432048
rect 577214 432002 577252 432048
rect 577276 432002 577278 432048
rect 577278 432002 577330 432048
rect 577330 432002 577332 432048
rect 577356 432002 577394 432048
rect 577394 432002 577406 432048
rect 577406 432002 577412 432048
rect 577436 432002 577458 432048
rect 577458 432002 577470 432048
rect 577470 432002 577492 432048
rect 577516 432002 577522 432048
rect 577522 432002 577534 432048
rect 577534 432002 577572 432048
rect 576605 431622 576661 431627
rect 576605 431571 576655 431622
rect 576655 431571 576661 431622
rect 580906 431570 580962 431626
rect 578276 431457 578314 431503
rect 578314 431457 578326 431503
rect 578326 431457 578332 431503
rect 578356 431457 578378 431503
rect 578378 431457 578390 431503
rect 578390 431457 578412 431503
rect 578436 431457 578442 431503
rect 578442 431457 578454 431503
rect 578454 431457 578492 431503
rect 578516 431457 578518 431503
rect 578518 431457 578570 431503
rect 578570 431457 578572 431503
rect 578596 431457 578634 431503
rect 578634 431457 578646 431503
rect 578646 431457 578652 431503
rect 578676 431457 578698 431503
rect 578698 431457 578710 431503
rect 578710 431457 578732 431503
rect 578756 431457 578762 431503
rect 578762 431457 578774 431503
rect 578774 431457 578812 431503
rect 578276 431447 578332 431457
rect 578356 431447 578412 431457
rect 578436 431447 578492 431457
rect 578516 431447 578572 431457
rect 578596 431447 578652 431457
rect 578676 431447 578732 431457
rect 578756 431447 578812 431457
rect 578276 431393 578314 431423
rect 578314 431393 578326 431423
rect 578326 431393 578332 431423
rect 578356 431393 578378 431423
rect 578378 431393 578390 431423
rect 578390 431393 578412 431423
rect 578436 431393 578442 431423
rect 578442 431393 578454 431423
rect 578454 431393 578492 431423
rect 578516 431393 578518 431423
rect 578518 431393 578570 431423
rect 578570 431393 578572 431423
rect 578596 431393 578634 431423
rect 578634 431393 578646 431423
rect 578646 431393 578652 431423
rect 578676 431393 578698 431423
rect 578698 431393 578710 431423
rect 578710 431393 578732 431423
rect 578756 431393 578762 431423
rect 578762 431393 578774 431423
rect 578774 431393 578812 431423
rect 578276 431381 578332 431393
rect 578356 431381 578412 431393
rect 578436 431381 578492 431393
rect 578516 431381 578572 431393
rect 578596 431381 578652 431393
rect 578676 431381 578732 431393
rect 578756 431381 578812 431393
rect 578276 431367 578314 431381
rect 578314 431367 578326 431381
rect 578326 431367 578332 431381
rect 578356 431367 578378 431381
rect 578378 431367 578390 431381
rect 578390 431367 578412 431381
rect 578436 431367 578442 431381
rect 578442 431367 578454 431381
rect 578454 431367 578492 431381
rect 578516 431367 578518 431381
rect 578518 431367 578570 431381
rect 578570 431367 578572 431381
rect 578596 431367 578634 431381
rect 578634 431367 578646 431381
rect 578646 431367 578652 431381
rect 578676 431367 578698 431381
rect 578698 431367 578710 431381
rect 578710 431367 578732 431381
rect 578756 431367 578762 431381
rect 578762 431367 578774 431381
rect 578774 431367 578812 431381
rect 578276 431329 578314 431343
rect 578314 431329 578326 431343
rect 578326 431329 578332 431343
rect 578356 431329 578378 431343
rect 578378 431329 578390 431343
rect 578390 431329 578412 431343
rect 578436 431329 578442 431343
rect 578442 431329 578454 431343
rect 578454 431329 578492 431343
rect 578516 431329 578518 431343
rect 578518 431329 578570 431343
rect 578570 431329 578572 431343
rect 578596 431329 578634 431343
rect 578634 431329 578646 431343
rect 578646 431329 578652 431343
rect 578676 431329 578698 431343
rect 578698 431329 578710 431343
rect 578710 431329 578732 431343
rect 578756 431329 578762 431343
rect 578762 431329 578774 431343
rect 578774 431329 578812 431343
rect 578276 431317 578332 431329
rect 578356 431317 578412 431329
rect 578436 431317 578492 431329
rect 578516 431317 578572 431329
rect 578596 431317 578652 431329
rect 578676 431317 578732 431329
rect 578756 431317 578812 431329
rect 578276 431287 578314 431317
rect 578314 431287 578326 431317
rect 578326 431287 578332 431317
rect 578356 431287 578378 431317
rect 578378 431287 578390 431317
rect 578390 431287 578412 431317
rect 578436 431287 578442 431317
rect 578442 431287 578454 431317
rect 578454 431287 578492 431317
rect 578516 431287 578518 431317
rect 578518 431287 578570 431317
rect 578570 431287 578572 431317
rect 578596 431287 578634 431317
rect 578634 431287 578646 431317
rect 578646 431287 578652 431317
rect 578676 431287 578698 431317
rect 578698 431287 578710 431317
rect 578710 431287 578732 431317
rect 578756 431287 578762 431317
rect 578762 431287 578774 431317
rect 578774 431287 578812 431317
rect 578276 431253 578332 431263
rect 578356 431253 578412 431263
rect 578436 431253 578492 431263
rect 578516 431253 578572 431263
rect 578596 431253 578652 431263
rect 578676 431253 578732 431263
rect 578756 431253 578812 431263
rect 578276 431207 578314 431253
rect 578314 431207 578326 431253
rect 578326 431207 578332 431253
rect 578356 431207 578378 431253
rect 578378 431207 578390 431253
rect 578390 431207 578412 431253
rect 578436 431207 578442 431253
rect 578442 431207 578454 431253
rect 578454 431207 578492 431253
rect 578516 431207 578518 431253
rect 578518 431207 578570 431253
rect 578570 431207 578572 431253
rect 578596 431207 578634 431253
rect 578634 431207 578646 431253
rect 578646 431207 578652 431253
rect 578676 431207 578698 431253
rect 578698 431207 578710 431253
rect 578710 431207 578732 431253
rect 578756 431207 578762 431253
rect 578762 431207 578774 431253
rect 578774 431207 578812 431253
rect 580170 409946 580226 410002
rect 580170 404914 580226 404970
rect 547970 398522 548026 398578
rect 577036 379076 577074 379122
rect 577074 379076 577086 379122
rect 577086 379076 577092 379122
rect 577116 379076 577138 379122
rect 577138 379076 577150 379122
rect 577150 379076 577172 379122
rect 577196 379076 577202 379122
rect 577202 379076 577214 379122
rect 577214 379076 577252 379122
rect 577276 379076 577278 379122
rect 577278 379076 577330 379122
rect 577330 379076 577332 379122
rect 577356 379076 577394 379122
rect 577394 379076 577406 379122
rect 577406 379076 577412 379122
rect 577436 379076 577458 379122
rect 577458 379076 577470 379122
rect 577470 379076 577492 379122
rect 577516 379076 577522 379122
rect 577522 379076 577534 379122
rect 577534 379076 577572 379122
rect 577036 379066 577092 379076
rect 577116 379066 577172 379076
rect 577196 379066 577252 379076
rect 577276 379066 577332 379076
rect 577356 379066 577412 379076
rect 577436 379066 577492 379076
rect 577516 379066 577572 379076
rect 577036 379012 577074 379042
rect 577074 379012 577086 379042
rect 577086 379012 577092 379042
rect 577116 379012 577138 379042
rect 577138 379012 577150 379042
rect 577150 379012 577172 379042
rect 577196 379012 577202 379042
rect 577202 379012 577214 379042
rect 577214 379012 577252 379042
rect 577276 379012 577278 379042
rect 577278 379012 577330 379042
rect 577330 379012 577332 379042
rect 577356 379012 577394 379042
rect 577394 379012 577406 379042
rect 577406 379012 577412 379042
rect 577436 379012 577458 379042
rect 577458 379012 577470 379042
rect 577470 379012 577492 379042
rect 577516 379012 577522 379042
rect 577522 379012 577534 379042
rect 577534 379012 577572 379042
rect 577036 379000 577092 379012
rect 577116 379000 577172 379012
rect 577196 379000 577252 379012
rect 577276 379000 577332 379012
rect 577356 379000 577412 379012
rect 577436 379000 577492 379012
rect 577516 379000 577572 379012
rect 577036 378986 577074 379000
rect 577074 378986 577086 379000
rect 577086 378986 577092 379000
rect 577116 378986 577138 379000
rect 577138 378986 577150 379000
rect 577150 378986 577172 379000
rect 577196 378986 577202 379000
rect 577202 378986 577214 379000
rect 577214 378986 577252 379000
rect 577276 378986 577278 379000
rect 577278 378986 577330 379000
rect 577330 378986 577332 379000
rect 577356 378986 577394 379000
rect 577394 378986 577406 379000
rect 577406 378986 577412 379000
rect 577436 378986 577458 379000
rect 577458 378986 577470 379000
rect 577470 378986 577492 379000
rect 577516 378986 577522 379000
rect 577522 378986 577534 379000
rect 577534 378986 577572 379000
rect 577036 378948 577074 378962
rect 577074 378948 577086 378962
rect 577086 378948 577092 378962
rect 577116 378948 577138 378962
rect 577138 378948 577150 378962
rect 577150 378948 577172 378962
rect 577196 378948 577202 378962
rect 577202 378948 577214 378962
rect 577214 378948 577252 378962
rect 577276 378948 577278 378962
rect 577278 378948 577330 378962
rect 577330 378948 577332 378962
rect 577356 378948 577394 378962
rect 577394 378948 577406 378962
rect 577406 378948 577412 378962
rect 577436 378948 577458 378962
rect 577458 378948 577470 378962
rect 577470 378948 577492 378962
rect 577516 378948 577522 378962
rect 577522 378948 577534 378962
rect 577534 378948 577572 378962
rect 577036 378936 577092 378948
rect 577116 378936 577172 378948
rect 577196 378936 577252 378948
rect 577276 378936 577332 378948
rect 577356 378936 577412 378948
rect 577436 378936 577492 378948
rect 577516 378936 577572 378948
rect 577036 378906 577074 378936
rect 577074 378906 577086 378936
rect 577086 378906 577092 378936
rect 577116 378906 577138 378936
rect 577138 378906 577150 378936
rect 577150 378906 577172 378936
rect 577196 378906 577202 378936
rect 577202 378906 577214 378936
rect 577214 378906 577252 378936
rect 577276 378906 577278 378936
rect 577278 378906 577330 378936
rect 577330 378906 577332 378936
rect 577356 378906 577394 378936
rect 577394 378906 577406 378936
rect 577406 378906 577412 378936
rect 577436 378906 577458 378936
rect 577458 378906 577470 378936
rect 577470 378906 577492 378936
rect 577516 378906 577522 378936
rect 577522 378906 577534 378936
rect 577534 378906 577572 378936
rect 577036 378872 577092 378882
rect 577116 378872 577172 378882
rect 577196 378872 577252 378882
rect 577276 378872 577332 378882
rect 577356 378872 577412 378882
rect 577436 378872 577492 378882
rect 577516 378872 577572 378882
rect 577036 378826 577074 378872
rect 577074 378826 577086 378872
rect 577086 378826 577092 378872
rect 577116 378826 577138 378872
rect 577138 378826 577150 378872
rect 577150 378826 577172 378872
rect 577196 378826 577202 378872
rect 577202 378826 577214 378872
rect 577214 378826 577252 378872
rect 577276 378826 577278 378872
rect 577278 378826 577330 378872
rect 577330 378826 577332 378872
rect 577356 378826 577394 378872
rect 577394 378826 577406 378872
rect 577406 378826 577412 378872
rect 577436 378826 577458 378872
rect 577458 378826 577470 378872
rect 577470 378826 577492 378872
rect 577516 378826 577522 378872
rect 577522 378826 577534 378872
rect 577534 378826 577572 378872
rect 576605 378446 576661 378451
rect 576605 378395 576655 378446
rect 576655 378395 576661 378446
rect 580906 378394 580962 378450
rect 578276 378281 578314 378327
rect 578314 378281 578326 378327
rect 578326 378281 578332 378327
rect 578356 378281 578378 378327
rect 578378 378281 578390 378327
rect 578390 378281 578412 378327
rect 578436 378281 578442 378327
rect 578442 378281 578454 378327
rect 578454 378281 578492 378327
rect 578516 378281 578518 378327
rect 578518 378281 578570 378327
rect 578570 378281 578572 378327
rect 578596 378281 578634 378327
rect 578634 378281 578646 378327
rect 578646 378281 578652 378327
rect 578676 378281 578698 378327
rect 578698 378281 578710 378327
rect 578710 378281 578732 378327
rect 578756 378281 578762 378327
rect 578762 378281 578774 378327
rect 578774 378281 578812 378327
rect 578276 378271 578332 378281
rect 578356 378271 578412 378281
rect 578436 378271 578492 378281
rect 578516 378271 578572 378281
rect 578596 378271 578652 378281
rect 578676 378271 578732 378281
rect 578756 378271 578812 378281
rect 578276 378217 578314 378247
rect 578314 378217 578326 378247
rect 578326 378217 578332 378247
rect 578356 378217 578378 378247
rect 578378 378217 578390 378247
rect 578390 378217 578412 378247
rect 578436 378217 578442 378247
rect 578442 378217 578454 378247
rect 578454 378217 578492 378247
rect 578516 378217 578518 378247
rect 578518 378217 578570 378247
rect 578570 378217 578572 378247
rect 578596 378217 578634 378247
rect 578634 378217 578646 378247
rect 578646 378217 578652 378247
rect 578676 378217 578698 378247
rect 578698 378217 578710 378247
rect 578710 378217 578732 378247
rect 578756 378217 578762 378247
rect 578762 378217 578774 378247
rect 578774 378217 578812 378247
rect 578276 378205 578332 378217
rect 578356 378205 578412 378217
rect 578436 378205 578492 378217
rect 578516 378205 578572 378217
rect 578596 378205 578652 378217
rect 578676 378205 578732 378217
rect 578756 378205 578812 378217
rect 578276 378191 578314 378205
rect 578314 378191 578326 378205
rect 578326 378191 578332 378205
rect 578356 378191 578378 378205
rect 578378 378191 578390 378205
rect 578390 378191 578412 378205
rect 578436 378191 578442 378205
rect 578442 378191 578454 378205
rect 578454 378191 578492 378205
rect 578516 378191 578518 378205
rect 578518 378191 578570 378205
rect 578570 378191 578572 378205
rect 578596 378191 578634 378205
rect 578634 378191 578646 378205
rect 578646 378191 578652 378205
rect 578676 378191 578698 378205
rect 578698 378191 578710 378205
rect 578710 378191 578732 378205
rect 578756 378191 578762 378205
rect 578762 378191 578774 378205
rect 578774 378191 578812 378205
rect 578276 378153 578314 378167
rect 578314 378153 578326 378167
rect 578326 378153 578332 378167
rect 578356 378153 578378 378167
rect 578378 378153 578390 378167
rect 578390 378153 578412 378167
rect 578436 378153 578442 378167
rect 578442 378153 578454 378167
rect 578454 378153 578492 378167
rect 578516 378153 578518 378167
rect 578518 378153 578570 378167
rect 578570 378153 578572 378167
rect 578596 378153 578634 378167
rect 578634 378153 578646 378167
rect 578646 378153 578652 378167
rect 578676 378153 578698 378167
rect 578698 378153 578710 378167
rect 578710 378153 578732 378167
rect 578756 378153 578762 378167
rect 578762 378153 578774 378167
rect 578774 378153 578812 378167
rect 578276 378141 578332 378153
rect 578356 378141 578412 378153
rect 578436 378141 578492 378153
rect 578516 378141 578572 378153
rect 578596 378141 578652 378153
rect 578676 378141 578732 378153
rect 578756 378141 578812 378153
rect 578276 378111 578314 378141
rect 578314 378111 578326 378141
rect 578326 378111 578332 378141
rect 578356 378111 578378 378141
rect 578378 378111 578390 378141
rect 578390 378111 578412 378141
rect 578436 378111 578442 378141
rect 578442 378111 578454 378141
rect 578454 378111 578492 378141
rect 578516 378111 578518 378141
rect 578518 378111 578570 378141
rect 578570 378111 578572 378141
rect 578596 378111 578634 378141
rect 578634 378111 578646 378141
rect 578646 378111 578652 378141
rect 578676 378111 578698 378141
rect 578698 378111 578710 378141
rect 578710 378111 578732 378141
rect 578756 378111 578762 378141
rect 578762 378111 578774 378141
rect 578774 378111 578812 378141
rect 578276 378077 578332 378087
rect 578356 378077 578412 378087
rect 578436 378077 578492 378087
rect 578516 378077 578572 378087
rect 578596 378077 578652 378087
rect 578676 378077 578732 378087
rect 578756 378077 578812 378087
rect 578276 378031 578314 378077
rect 578314 378031 578326 378077
rect 578326 378031 578332 378077
rect 578356 378031 578378 378077
rect 578378 378031 578390 378077
rect 578390 378031 578412 378077
rect 578436 378031 578442 378077
rect 578442 378031 578454 378077
rect 578454 378031 578492 378077
rect 578516 378031 578518 378077
rect 578518 378031 578570 378077
rect 578570 378031 578572 378077
rect 578596 378031 578634 378077
rect 578634 378031 578646 378077
rect 578646 378031 578652 378077
rect 578676 378031 578698 378077
rect 578698 378031 578710 378077
rect 578710 378031 578732 378077
rect 578756 378031 578762 378077
rect 578762 378031 578774 378077
rect 578774 378031 578812 378077
rect 547878 362890 547934 362946
rect 547418 326986 547474 327042
rect 577036 325900 577074 325946
rect 577074 325900 577086 325946
rect 577086 325900 577092 325946
rect 577116 325900 577138 325946
rect 577138 325900 577150 325946
rect 577150 325900 577172 325946
rect 577196 325900 577202 325946
rect 577202 325900 577214 325946
rect 577214 325900 577252 325946
rect 577276 325900 577278 325946
rect 577278 325900 577330 325946
rect 577330 325900 577332 325946
rect 577356 325900 577394 325946
rect 577394 325900 577406 325946
rect 577406 325900 577412 325946
rect 577436 325900 577458 325946
rect 577458 325900 577470 325946
rect 577470 325900 577492 325946
rect 577516 325900 577522 325946
rect 577522 325900 577534 325946
rect 577534 325900 577572 325946
rect 577036 325890 577092 325900
rect 577116 325890 577172 325900
rect 577196 325890 577252 325900
rect 577276 325890 577332 325900
rect 577356 325890 577412 325900
rect 577436 325890 577492 325900
rect 577516 325890 577572 325900
rect 577036 325836 577074 325866
rect 577074 325836 577086 325866
rect 577086 325836 577092 325866
rect 577116 325836 577138 325866
rect 577138 325836 577150 325866
rect 577150 325836 577172 325866
rect 577196 325836 577202 325866
rect 577202 325836 577214 325866
rect 577214 325836 577252 325866
rect 577276 325836 577278 325866
rect 577278 325836 577330 325866
rect 577330 325836 577332 325866
rect 577356 325836 577394 325866
rect 577394 325836 577406 325866
rect 577406 325836 577412 325866
rect 577436 325836 577458 325866
rect 577458 325836 577470 325866
rect 577470 325836 577492 325866
rect 577516 325836 577522 325866
rect 577522 325836 577534 325866
rect 577534 325836 577572 325866
rect 577036 325824 577092 325836
rect 577116 325824 577172 325836
rect 577196 325824 577252 325836
rect 577276 325824 577332 325836
rect 577356 325824 577412 325836
rect 577436 325824 577492 325836
rect 577516 325824 577572 325836
rect 577036 325810 577074 325824
rect 577074 325810 577086 325824
rect 577086 325810 577092 325824
rect 577116 325810 577138 325824
rect 577138 325810 577150 325824
rect 577150 325810 577172 325824
rect 577196 325810 577202 325824
rect 577202 325810 577214 325824
rect 577214 325810 577252 325824
rect 577276 325810 577278 325824
rect 577278 325810 577330 325824
rect 577330 325810 577332 325824
rect 577356 325810 577394 325824
rect 577394 325810 577406 325824
rect 577406 325810 577412 325824
rect 577436 325810 577458 325824
rect 577458 325810 577470 325824
rect 577470 325810 577492 325824
rect 577516 325810 577522 325824
rect 577522 325810 577534 325824
rect 577534 325810 577572 325824
rect 577036 325772 577074 325786
rect 577074 325772 577086 325786
rect 577086 325772 577092 325786
rect 577116 325772 577138 325786
rect 577138 325772 577150 325786
rect 577150 325772 577172 325786
rect 577196 325772 577202 325786
rect 577202 325772 577214 325786
rect 577214 325772 577252 325786
rect 577276 325772 577278 325786
rect 577278 325772 577330 325786
rect 577330 325772 577332 325786
rect 577356 325772 577394 325786
rect 577394 325772 577406 325786
rect 577406 325772 577412 325786
rect 577436 325772 577458 325786
rect 577458 325772 577470 325786
rect 577470 325772 577492 325786
rect 577516 325772 577522 325786
rect 577522 325772 577534 325786
rect 577534 325772 577572 325786
rect 577036 325760 577092 325772
rect 577116 325760 577172 325772
rect 577196 325760 577252 325772
rect 577276 325760 577332 325772
rect 577356 325760 577412 325772
rect 577436 325760 577492 325772
rect 577516 325760 577572 325772
rect 577036 325730 577074 325760
rect 577074 325730 577086 325760
rect 577086 325730 577092 325760
rect 577116 325730 577138 325760
rect 577138 325730 577150 325760
rect 577150 325730 577172 325760
rect 577196 325730 577202 325760
rect 577202 325730 577214 325760
rect 577214 325730 577252 325760
rect 577276 325730 577278 325760
rect 577278 325730 577330 325760
rect 577330 325730 577332 325760
rect 577356 325730 577394 325760
rect 577394 325730 577406 325760
rect 577406 325730 577412 325760
rect 577436 325730 577458 325760
rect 577458 325730 577470 325760
rect 577470 325730 577492 325760
rect 577516 325730 577522 325760
rect 577522 325730 577534 325760
rect 577534 325730 577572 325760
rect 577036 325696 577092 325706
rect 577116 325696 577172 325706
rect 577196 325696 577252 325706
rect 577276 325696 577332 325706
rect 577356 325696 577412 325706
rect 577436 325696 577492 325706
rect 577516 325696 577572 325706
rect 577036 325650 577074 325696
rect 577074 325650 577086 325696
rect 577086 325650 577092 325696
rect 577116 325650 577138 325696
rect 577138 325650 577150 325696
rect 577150 325650 577172 325696
rect 577196 325650 577202 325696
rect 577202 325650 577214 325696
rect 577214 325650 577252 325696
rect 577276 325650 577278 325696
rect 577278 325650 577330 325696
rect 577330 325650 577332 325696
rect 577356 325650 577394 325696
rect 577394 325650 577406 325696
rect 577406 325650 577412 325696
rect 577436 325650 577458 325696
rect 577458 325650 577470 325696
rect 577470 325650 577492 325696
rect 577516 325650 577522 325696
rect 577522 325650 577534 325696
rect 577534 325650 577572 325696
rect 576605 325270 576661 325275
rect 576605 325219 576655 325270
rect 576655 325219 576661 325270
rect 580906 325218 580962 325274
rect 578276 325105 578314 325151
rect 578314 325105 578326 325151
rect 578326 325105 578332 325151
rect 578356 325105 578378 325151
rect 578378 325105 578390 325151
rect 578390 325105 578412 325151
rect 578436 325105 578442 325151
rect 578442 325105 578454 325151
rect 578454 325105 578492 325151
rect 578516 325105 578518 325151
rect 578518 325105 578570 325151
rect 578570 325105 578572 325151
rect 578596 325105 578634 325151
rect 578634 325105 578646 325151
rect 578646 325105 578652 325151
rect 578676 325105 578698 325151
rect 578698 325105 578710 325151
rect 578710 325105 578732 325151
rect 578756 325105 578762 325151
rect 578762 325105 578774 325151
rect 578774 325105 578812 325151
rect 578276 325095 578332 325105
rect 578356 325095 578412 325105
rect 578436 325095 578492 325105
rect 578516 325095 578572 325105
rect 578596 325095 578652 325105
rect 578676 325095 578732 325105
rect 578756 325095 578812 325105
rect 578276 325041 578314 325071
rect 578314 325041 578326 325071
rect 578326 325041 578332 325071
rect 578356 325041 578378 325071
rect 578378 325041 578390 325071
rect 578390 325041 578412 325071
rect 578436 325041 578442 325071
rect 578442 325041 578454 325071
rect 578454 325041 578492 325071
rect 578516 325041 578518 325071
rect 578518 325041 578570 325071
rect 578570 325041 578572 325071
rect 578596 325041 578634 325071
rect 578634 325041 578646 325071
rect 578646 325041 578652 325071
rect 578676 325041 578698 325071
rect 578698 325041 578710 325071
rect 578710 325041 578732 325071
rect 578756 325041 578762 325071
rect 578762 325041 578774 325071
rect 578774 325041 578812 325071
rect 578276 325029 578332 325041
rect 578356 325029 578412 325041
rect 578436 325029 578492 325041
rect 578516 325029 578572 325041
rect 578596 325029 578652 325041
rect 578676 325029 578732 325041
rect 578756 325029 578812 325041
rect 578276 325015 578314 325029
rect 578314 325015 578326 325029
rect 578326 325015 578332 325029
rect 578356 325015 578378 325029
rect 578378 325015 578390 325029
rect 578390 325015 578412 325029
rect 578436 325015 578442 325029
rect 578442 325015 578454 325029
rect 578454 325015 578492 325029
rect 578516 325015 578518 325029
rect 578518 325015 578570 325029
rect 578570 325015 578572 325029
rect 578596 325015 578634 325029
rect 578634 325015 578646 325029
rect 578646 325015 578652 325029
rect 578676 325015 578698 325029
rect 578698 325015 578710 325029
rect 578710 325015 578732 325029
rect 578756 325015 578762 325029
rect 578762 325015 578774 325029
rect 578774 325015 578812 325029
rect 578276 324977 578314 324991
rect 578314 324977 578326 324991
rect 578326 324977 578332 324991
rect 578356 324977 578378 324991
rect 578378 324977 578390 324991
rect 578390 324977 578412 324991
rect 578436 324977 578442 324991
rect 578442 324977 578454 324991
rect 578454 324977 578492 324991
rect 578516 324977 578518 324991
rect 578518 324977 578570 324991
rect 578570 324977 578572 324991
rect 578596 324977 578634 324991
rect 578634 324977 578646 324991
rect 578646 324977 578652 324991
rect 578676 324977 578698 324991
rect 578698 324977 578710 324991
rect 578710 324977 578732 324991
rect 578756 324977 578762 324991
rect 578762 324977 578774 324991
rect 578774 324977 578812 324991
rect 578276 324965 578332 324977
rect 578356 324965 578412 324977
rect 578436 324965 578492 324977
rect 578516 324965 578572 324977
rect 578596 324965 578652 324977
rect 578676 324965 578732 324977
rect 578756 324965 578812 324977
rect 578276 324935 578314 324965
rect 578314 324935 578326 324965
rect 578326 324935 578332 324965
rect 578356 324935 578378 324965
rect 578378 324935 578390 324965
rect 578390 324935 578412 324965
rect 578436 324935 578442 324965
rect 578442 324935 578454 324965
rect 578454 324935 578492 324965
rect 578516 324935 578518 324965
rect 578518 324935 578570 324965
rect 578570 324935 578572 324965
rect 578596 324935 578634 324965
rect 578634 324935 578646 324965
rect 578646 324935 578652 324965
rect 578676 324935 578698 324965
rect 578698 324935 578710 324965
rect 578710 324935 578732 324965
rect 578756 324935 578762 324965
rect 578762 324935 578774 324965
rect 578774 324935 578812 324965
rect 578276 324901 578332 324911
rect 578356 324901 578412 324911
rect 578436 324901 578492 324911
rect 578516 324901 578572 324911
rect 578596 324901 578652 324911
rect 578676 324901 578732 324911
rect 578756 324901 578812 324911
rect 578276 324855 578314 324901
rect 578314 324855 578326 324901
rect 578326 324855 578332 324901
rect 578356 324855 578378 324901
rect 578378 324855 578390 324901
rect 578390 324855 578412 324901
rect 578436 324855 578442 324901
rect 578442 324855 578454 324901
rect 578454 324855 578492 324901
rect 578516 324855 578518 324901
rect 578518 324855 578570 324901
rect 578570 324855 578572 324901
rect 578596 324855 578634 324901
rect 578634 324855 578646 324901
rect 578646 324855 578652 324901
rect 578676 324855 578698 324901
rect 578698 324855 578710 324901
rect 578710 324855 578732 324901
rect 578756 324855 578762 324901
rect 578762 324855 578774 324901
rect 578774 324855 578812 324901
rect 580170 302234 580226 302290
rect 580170 298698 580226 298754
rect 547326 291082 547382 291138
rect 536746 287138 536802 287194
rect 577036 272860 577074 272906
rect 577074 272860 577086 272906
rect 577086 272860 577092 272906
rect 577116 272860 577138 272906
rect 577138 272860 577150 272906
rect 577150 272860 577172 272906
rect 577196 272860 577202 272906
rect 577202 272860 577214 272906
rect 577214 272860 577252 272906
rect 577276 272860 577278 272906
rect 577278 272860 577330 272906
rect 577330 272860 577332 272906
rect 577356 272860 577394 272906
rect 577394 272860 577406 272906
rect 577406 272860 577412 272906
rect 577436 272860 577458 272906
rect 577458 272860 577470 272906
rect 577470 272860 577492 272906
rect 577516 272860 577522 272906
rect 577522 272860 577534 272906
rect 577534 272860 577572 272906
rect 577036 272850 577092 272860
rect 577116 272850 577172 272860
rect 577196 272850 577252 272860
rect 577276 272850 577332 272860
rect 577356 272850 577412 272860
rect 577436 272850 577492 272860
rect 577516 272850 577572 272860
rect 577036 272796 577074 272826
rect 577074 272796 577086 272826
rect 577086 272796 577092 272826
rect 577116 272796 577138 272826
rect 577138 272796 577150 272826
rect 577150 272796 577172 272826
rect 577196 272796 577202 272826
rect 577202 272796 577214 272826
rect 577214 272796 577252 272826
rect 577276 272796 577278 272826
rect 577278 272796 577330 272826
rect 577330 272796 577332 272826
rect 577356 272796 577394 272826
rect 577394 272796 577406 272826
rect 577406 272796 577412 272826
rect 577436 272796 577458 272826
rect 577458 272796 577470 272826
rect 577470 272796 577492 272826
rect 577516 272796 577522 272826
rect 577522 272796 577534 272826
rect 577534 272796 577572 272826
rect 577036 272784 577092 272796
rect 577116 272784 577172 272796
rect 577196 272784 577252 272796
rect 577276 272784 577332 272796
rect 577356 272784 577412 272796
rect 577436 272784 577492 272796
rect 577516 272784 577572 272796
rect 577036 272770 577074 272784
rect 577074 272770 577086 272784
rect 577086 272770 577092 272784
rect 577116 272770 577138 272784
rect 577138 272770 577150 272784
rect 577150 272770 577172 272784
rect 577196 272770 577202 272784
rect 577202 272770 577214 272784
rect 577214 272770 577252 272784
rect 577276 272770 577278 272784
rect 577278 272770 577330 272784
rect 577330 272770 577332 272784
rect 577356 272770 577394 272784
rect 577394 272770 577406 272784
rect 577406 272770 577412 272784
rect 577436 272770 577458 272784
rect 577458 272770 577470 272784
rect 577470 272770 577492 272784
rect 577516 272770 577522 272784
rect 577522 272770 577534 272784
rect 577534 272770 577572 272784
rect 577036 272732 577074 272746
rect 577074 272732 577086 272746
rect 577086 272732 577092 272746
rect 577116 272732 577138 272746
rect 577138 272732 577150 272746
rect 577150 272732 577172 272746
rect 577196 272732 577202 272746
rect 577202 272732 577214 272746
rect 577214 272732 577252 272746
rect 577276 272732 577278 272746
rect 577278 272732 577330 272746
rect 577330 272732 577332 272746
rect 577356 272732 577394 272746
rect 577394 272732 577406 272746
rect 577406 272732 577412 272746
rect 577436 272732 577458 272746
rect 577458 272732 577470 272746
rect 577470 272732 577492 272746
rect 577516 272732 577522 272746
rect 577522 272732 577534 272746
rect 577534 272732 577572 272746
rect 577036 272720 577092 272732
rect 577116 272720 577172 272732
rect 577196 272720 577252 272732
rect 577276 272720 577332 272732
rect 577356 272720 577412 272732
rect 577436 272720 577492 272732
rect 577516 272720 577572 272732
rect 577036 272690 577074 272720
rect 577074 272690 577086 272720
rect 577086 272690 577092 272720
rect 577116 272690 577138 272720
rect 577138 272690 577150 272720
rect 577150 272690 577172 272720
rect 577196 272690 577202 272720
rect 577202 272690 577214 272720
rect 577214 272690 577252 272720
rect 577276 272690 577278 272720
rect 577278 272690 577330 272720
rect 577330 272690 577332 272720
rect 577356 272690 577394 272720
rect 577394 272690 577406 272720
rect 577406 272690 577412 272720
rect 577436 272690 577458 272720
rect 577458 272690 577470 272720
rect 577470 272690 577492 272720
rect 577516 272690 577522 272720
rect 577522 272690 577534 272720
rect 577534 272690 577572 272720
rect 577036 272656 577092 272666
rect 577116 272656 577172 272666
rect 577196 272656 577252 272666
rect 577276 272656 577332 272666
rect 577356 272656 577412 272666
rect 577436 272656 577492 272666
rect 577516 272656 577572 272666
rect 577036 272610 577074 272656
rect 577074 272610 577086 272656
rect 577086 272610 577092 272656
rect 577116 272610 577138 272656
rect 577138 272610 577150 272656
rect 577150 272610 577172 272656
rect 577196 272610 577202 272656
rect 577202 272610 577214 272656
rect 577214 272610 577252 272656
rect 577276 272610 577278 272656
rect 577278 272610 577330 272656
rect 577330 272610 577332 272656
rect 577356 272610 577394 272656
rect 577394 272610 577406 272656
rect 577406 272610 577412 272656
rect 577436 272610 577458 272656
rect 577458 272610 577470 272656
rect 577470 272610 577492 272656
rect 577516 272610 577522 272656
rect 577522 272610 577534 272656
rect 577534 272610 577572 272656
rect 576605 272230 576661 272235
rect 576605 272179 576655 272230
rect 576655 272179 576661 272230
rect 580906 272178 580962 272234
rect 578276 272065 578314 272111
rect 578314 272065 578326 272111
rect 578326 272065 578332 272111
rect 578356 272065 578378 272111
rect 578378 272065 578390 272111
rect 578390 272065 578412 272111
rect 578436 272065 578442 272111
rect 578442 272065 578454 272111
rect 578454 272065 578492 272111
rect 578516 272065 578518 272111
rect 578518 272065 578570 272111
rect 578570 272065 578572 272111
rect 578596 272065 578634 272111
rect 578634 272065 578646 272111
rect 578646 272065 578652 272111
rect 578676 272065 578698 272111
rect 578698 272065 578710 272111
rect 578710 272065 578732 272111
rect 578756 272065 578762 272111
rect 578762 272065 578774 272111
rect 578774 272065 578812 272111
rect 578276 272055 578332 272065
rect 578356 272055 578412 272065
rect 578436 272055 578492 272065
rect 578516 272055 578572 272065
rect 578596 272055 578652 272065
rect 578676 272055 578732 272065
rect 578756 272055 578812 272065
rect 578276 272001 578314 272031
rect 578314 272001 578326 272031
rect 578326 272001 578332 272031
rect 578356 272001 578378 272031
rect 578378 272001 578390 272031
rect 578390 272001 578412 272031
rect 578436 272001 578442 272031
rect 578442 272001 578454 272031
rect 578454 272001 578492 272031
rect 578516 272001 578518 272031
rect 578518 272001 578570 272031
rect 578570 272001 578572 272031
rect 578596 272001 578634 272031
rect 578634 272001 578646 272031
rect 578646 272001 578652 272031
rect 578676 272001 578698 272031
rect 578698 272001 578710 272031
rect 578710 272001 578732 272031
rect 578756 272001 578762 272031
rect 578762 272001 578774 272031
rect 578774 272001 578812 272031
rect 578276 271989 578332 272001
rect 578356 271989 578412 272001
rect 578436 271989 578492 272001
rect 578516 271989 578572 272001
rect 578596 271989 578652 272001
rect 578676 271989 578732 272001
rect 578756 271989 578812 272001
rect 578276 271975 578314 271989
rect 578314 271975 578326 271989
rect 578326 271975 578332 271989
rect 578356 271975 578378 271989
rect 578378 271975 578390 271989
rect 578390 271975 578412 271989
rect 578436 271975 578442 271989
rect 578442 271975 578454 271989
rect 578454 271975 578492 271989
rect 578516 271975 578518 271989
rect 578518 271975 578570 271989
rect 578570 271975 578572 271989
rect 578596 271975 578634 271989
rect 578634 271975 578646 271989
rect 578646 271975 578652 271989
rect 578676 271975 578698 271989
rect 578698 271975 578710 271989
rect 578710 271975 578732 271989
rect 578756 271975 578762 271989
rect 578762 271975 578774 271989
rect 578774 271975 578812 271989
rect 578276 271937 578314 271951
rect 578314 271937 578326 271951
rect 578326 271937 578332 271951
rect 578356 271937 578378 271951
rect 578378 271937 578390 271951
rect 578390 271937 578412 271951
rect 578436 271937 578442 271951
rect 578442 271937 578454 271951
rect 578454 271937 578492 271951
rect 578516 271937 578518 271951
rect 578518 271937 578570 271951
rect 578570 271937 578572 271951
rect 578596 271937 578634 271951
rect 578634 271937 578646 271951
rect 578646 271937 578652 271951
rect 578676 271937 578698 271951
rect 578698 271937 578710 271951
rect 578710 271937 578732 271951
rect 578756 271937 578762 271951
rect 578762 271937 578774 271951
rect 578774 271937 578812 271951
rect 578276 271925 578332 271937
rect 578356 271925 578412 271937
rect 578436 271925 578492 271937
rect 578516 271925 578572 271937
rect 578596 271925 578652 271937
rect 578676 271925 578732 271937
rect 578756 271925 578812 271937
rect 578276 271895 578314 271925
rect 578314 271895 578326 271925
rect 578326 271895 578332 271925
rect 578356 271895 578378 271925
rect 578378 271895 578390 271925
rect 578390 271895 578412 271925
rect 578436 271895 578442 271925
rect 578442 271895 578454 271925
rect 578454 271895 578492 271925
rect 578516 271895 578518 271925
rect 578518 271895 578570 271925
rect 578570 271895 578572 271925
rect 578596 271895 578634 271925
rect 578634 271895 578646 271925
rect 578646 271895 578652 271925
rect 578676 271895 578698 271925
rect 578698 271895 578710 271925
rect 578710 271895 578732 271925
rect 578756 271895 578762 271925
rect 578762 271895 578774 271925
rect 578774 271895 578812 271925
rect 578276 271861 578332 271871
rect 578356 271861 578412 271871
rect 578436 271861 578492 271871
rect 578516 271861 578572 271871
rect 578596 271861 578652 271871
rect 578676 271861 578732 271871
rect 578756 271861 578812 271871
rect 578276 271815 578314 271861
rect 578314 271815 578326 271861
rect 578326 271815 578332 271861
rect 578356 271815 578378 271861
rect 578378 271815 578390 271861
rect 578390 271815 578412 271861
rect 578436 271815 578442 271861
rect 578442 271815 578454 271861
rect 578454 271815 578492 271861
rect 578516 271815 578518 271861
rect 578518 271815 578570 271861
rect 578570 271815 578572 271861
rect 578596 271815 578634 271861
rect 578634 271815 578646 271861
rect 578646 271815 578652 271861
rect 578676 271815 578698 271861
rect 578698 271815 578710 271861
rect 578710 271815 578732 271861
rect 578756 271815 578762 271861
rect 578762 271815 578774 271861
rect 578774 271815 578812 271861
rect 577036 233013 577074 233059
rect 577074 233013 577086 233059
rect 577086 233013 577092 233059
rect 577116 233013 577138 233059
rect 577138 233013 577150 233059
rect 577150 233013 577172 233059
rect 577196 233013 577202 233059
rect 577202 233013 577214 233059
rect 577214 233013 577252 233059
rect 577276 233013 577278 233059
rect 577278 233013 577330 233059
rect 577330 233013 577332 233059
rect 577356 233013 577394 233059
rect 577394 233013 577406 233059
rect 577406 233013 577412 233059
rect 577436 233013 577458 233059
rect 577458 233013 577470 233059
rect 577470 233013 577492 233059
rect 577516 233013 577522 233059
rect 577522 233013 577534 233059
rect 577534 233013 577572 233059
rect 577036 233003 577092 233013
rect 577116 233003 577172 233013
rect 577196 233003 577252 233013
rect 577276 233003 577332 233013
rect 577356 233003 577412 233013
rect 577436 233003 577492 233013
rect 577516 233003 577572 233013
rect 577036 232949 577074 232979
rect 577074 232949 577086 232979
rect 577086 232949 577092 232979
rect 577116 232949 577138 232979
rect 577138 232949 577150 232979
rect 577150 232949 577172 232979
rect 577196 232949 577202 232979
rect 577202 232949 577214 232979
rect 577214 232949 577252 232979
rect 577276 232949 577278 232979
rect 577278 232949 577330 232979
rect 577330 232949 577332 232979
rect 577356 232949 577394 232979
rect 577394 232949 577406 232979
rect 577406 232949 577412 232979
rect 577436 232949 577458 232979
rect 577458 232949 577470 232979
rect 577470 232949 577492 232979
rect 577516 232949 577522 232979
rect 577522 232949 577534 232979
rect 577534 232949 577572 232979
rect 577036 232937 577092 232949
rect 577116 232937 577172 232949
rect 577196 232937 577252 232949
rect 577276 232937 577332 232949
rect 577356 232937 577412 232949
rect 577436 232937 577492 232949
rect 577516 232937 577572 232949
rect 577036 232923 577074 232937
rect 577074 232923 577086 232937
rect 577086 232923 577092 232937
rect 577116 232923 577138 232937
rect 577138 232923 577150 232937
rect 577150 232923 577172 232937
rect 577196 232923 577202 232937
rect 577202 232923 577214 232937
rect 577214 232923 577252 232937
rect 577276 232923 577278 232937
rect 577278 232923 577330 232937
rect 577330 232923 577332 232937
rect 577356 232923 577394 232937
rect 577394 232923 577406 232937
rect 577406 232923 577412 232937
rect 577436 232923 577458 232937
rect 577458 232923 577470 232937
rect 577470 232923 577492 232937
rect 577516 232923 577522 232937
rect 577522 232923 577534 232937
rect 577534 232923 577572 232937
rect 577036 232885 577074 232899
rect 577074 232885 577086 232899
rect 577086 232885 577092 232899
rect 577116 232885 577138 232899
rect 577138 232885 577150 232899
rect 577150 232885 577172 232899
rect 577196 232885 577202 232899
rect 577202 232885 577214 232899
rect 577214 232885 577252 232899
rect 577276 232885 577278 232899
rect 577278 232885 577330 232899
rect 577330 232885 577332 232899
rect 577356 232885 577394 232899
rect 577394 232885 577406 232899
rect 577406 232885 577412 232899
rect 577436 232885 577458 232899
rect 577458 232885 577470 232899
rect 577470 232885 577492 232899
rect 577516 232885 577522 232899
rect 577522 232885 577534 232899
rect 577534 232885 577572 232899
rect 577036 232873 577092 232885
rect 577116 232873 577172 232885
rect 577196 232873 577252 232885
rect 577276 232873 577332 232885
rect 577356 232873 577412 232885
rect 577436 232873 577492 232885
rect 577516 232873 577572 232885
rect 577036 232843 577074 232873
rect 577074 232843 577086 232873
rect 577086 232843 577092 232873
rect 577116 232843 577138 232873
rect 577138 232843 577150 232873
rect 577150 232843 577172 232873
rect 577196 232843 577202 232873
rect 577202 232843 577214 232873
rect 577214 232843 577252 232873
rect 577276 232843 577278 232873
rect 577278 232843 577330 232873
rect 577330 232843 577332 232873
rect 577356 232843 577394 232873
rect 577394 232843 577406 232873
rect 577406 232843 577412 232873
rect 577436 232843 577458 232873
rect 577458 232843 577470 232873
rect 577470 232843 577492 232873
rect 577516 232843 577522 232873
rect 577522 232843 577534 232873
rect 577534 232843 577572 232873
rect 577036 232809 577092 232819
rect 577116 232809 577172 232819
rect 577196 232809 577252 232819
rect 577276 232809 577332 232819
rect 577356 232809 577412 232819
rect 577436 232809 577492 232819
rect 577516 232809 577572 232819
rect 577036 232763 577074 232809
rect 577074 232763 577086 232809
rect 577086 232763 577092 232809
rect 577116 232763 577138 232809
rect 577138 232763 577150 232809
rect 577150 232763 577172 232809
rect 577196 232763 577202 232809
rect 577202 232763 577214 232809
rect 577214 232763 577252 232809
rect 577276 232763 577278 232809
rect 577278 232763 577330 232809
rect 577330 232763 577332 232809
rect 577356 232763 577394 232809
rect 577394 232763 577406 232809
rect 577406 232763 577412 232809
rect 577436 232763 577458 232809
rect 577458 232763 577470 232809
rect 577470 232763 577492 232809
rect 577516 232763 577522 232809
rect 577522 232763 577534 232809
rect 577534 232763 577572 232809
rect 576605 232383 576661 232388
rect 576605 232332 576655 232383
rect 576655 232332 576661 232383
rect 580906 232330 580962 232386
rect 578276 232218 578314 232264
rect 578314 232218 578326 232264
rect 578326 232218 578332 232264
rect 578356 232218 578378 232264
rect 578378 232218 578390 232264
rect 578390 232218 578412 232264
rect 578436 232218 578442 232264
rect 578442 232218 578454 232264
rect 578454 232218 578492 232264
rect 578516 232218 578518 232264
rect 578518 232218 578570 232264
rect 578570 232218 578572 232264
rect 578596 232218 578634 232264
rect 578634 232218 578646 232264
rect 578646 232218 578652 232264
rect 578676 232218 578698 232264
rect 578698 232218 578710 232264
rect 578710 232218 578732 232264
rect 578756 232218 578762 232264
rect 578762 232218 578774 232264
rect 578774 232218 578812 232264
rect 578276 232208 578332 232218
rect 578356 232208 578412 232218
rect 578436 232208 578492 232218
rect 578516 232208 578572 232218
rect 578596 232208 578652 232218
rect 578676 232208 578732 232218
rect 578756 232208 578812 232218
rect 578276 232154 578314 232184
rect 578314 232154 578326 232184
rect 578326 232154 578332 232184
rect 578356 232154 578378 232184
rect 578378 232154 578390 232184
rect 578390 232154 578412 232184
rect 578436 232154 578442 232184
rect 578442 232154 578454 232184
rect 578454 232154 578492 232184
rect 578516 232154 578518 232184
rect 578518 232154 578570 232184
rect 578570 232154 578572 232184
rect 578596 232154 578634 232184
rect 578634 232154 578646 232184
rect 578646 232154 578652 232184
rect 578676 232154 578698 232184
rect 578698 232154 578710 232184
rect 578710 232154 578732 232184
rect 578756 232154 578762 232184
rect 578762 232154 578774 232184
rect 578774 232154 578812 232184
rect 578276 232142 578332 232154
rect 578356 232142 578412 232154
rect 578436 232142 578492 232154
rect 578516 232142 578572 232154
rect 578596 232142 578652 232154
rect 578676 232142 578732 232154
rect 578756 232142 578812 232154
rect 578276 232128 578314 232142
rect 578314 232128 578326 232142
rect 578326 232128 578332 232142
rect 578356 232128 578378 232142
rect 578378 232128 578390 232142
rect 578390 232128 578412 232142
rect 578436 232128 578442 232142
rect 578442 232128 578454 232142
rect 578454 232128 578492 232142
rect 578516 232128 578518 232142
rect 578518 232128 578570 232142
rect 578570 232128 578572 232142
rect 578596 232128 578634 232142
rect 578634 232128 578646 232142
rect 578646 232128 578652 232142
rect 578676 232128 578698 232142
rect 578698 232128 578710 232142
rect 578710 232128 578732 232142
rect 578756 232128 578762 232142
rect 578762 232128 578774 232142
rect 578774 232128 578812 232142
rect 578276 232090 578314 232104
rect 578314 232090 578326 232104
rect 578326 232090 578332 232104
rect 578356 232090 578378 232104
rect 578378 232090 578390 232104
rect 578390 232090 578412 232104
rect 578436 232090 578442 232104
rect 578442 232090 578454 232104
rect 578454 232090 578492 232104
rect 578516 232090 578518 232104
rect 578518 232090 578570 232104
rect 578570 232090 578572 232104
rect 578596 232090 578634 232104
rect 578634 232090 578646 232104
rect 578646 232090 578652 232104
rect 578676 232090 578698 232104
rect 578698 232090 578710 232104
rect 578710 232090 578732 232104
rect 578756 232090 578762 232104
rect 578762 232090 578774 232104
rect 578774 232090 578812 232104
rect 578276 232078 578332 232090
rect 578356 232078 578412 232090
rect 578436 232078 578492 232090
rect 578516 232078 578572 232090
rect 578596 232078 578652 232090
rect 578676 232078 578732 232090
rect 578756 232078 578812 232090
rect 578276 232048 578314 232078
rect 578314 232048 578326 232078
rect 578326 232048 578332 232078
rect 578356 232048 578378 232078
rect 578378 232048 578390 232078
rect 578390 232048 578412 232078
rect 578436 232048 578442 232078
rect 578442 232048 578454 232078
rect 578454 232048 578492 232078
rect 578516 232048 578518 232078
rect 578518 232048 578570 232078
rect 578570 232048 578572 232078
rect 578596 232048 578634 232078
rect 578634 232048 578646 232078
rect 578646 232048 578652 232078
rect 578676 232048 578698 232078
rect 578698 232048 578710 232078
rect 578710 232048 578732 232078
rect 578756 232048 578762 232078
rect 578762 232048 578774 232078
rect 578774 232048 578812 232078
rect 578276 232014 578332 232024
rect 578356 232014 578412 232024
rect 578436 232014 578492 232024
rect 578516 232014 578572 232024
rect 578596 232014 578652 232024
rect 578676 232014 578732 232024
rect 578756 232014 578812 232024
rect 578276 231968 578314 232014
rect 578314 231968 578326 232014
rect 578326 231968 578332 232014
rect 578356 231968 578378 232014
rect 578378 231968 578390 232014
rect 578390 231968 578412 232014
rect 578436 231968 578442 232014
rect 578442 231968 578454 232014
rect 578454 231968 578492 232014
rect 578516 231968 578518 232014
rect 578518 231968 578570 232014
rect 578570 231968 578572 232014
rect 578596 231968 578634 232014
rect 578634 231968 578646 232014
rect 578646 231968 578652 232014
rect 578676 231968 578698 232014
rect 578698 231968 578710 232014
rect 578710 231968 578732 232014
rect 578756 231968 578762 232014
rect 578762 231968 578774 232014
rect 578774 231968 578812 232014
<< metal3 >>
rect 326266 703376 326822 703377
rect 254266 703336 254822 703337
rect 254266 703272 254272 703336
rect 254336 703272 254352 703336
rect 254416 703272 254432 703336
rect 254496 703272 254512 703336
rect 254576 703272 254592 703336
rect 254656 703272 254672 703336
rect 254736 703272 254752 703336
rect 254816 703272 254822 703336
rect 254266 703256 254822 703272
rect 254266 703192 254272 703256
rect 254336 703192 254352 703256
rect 254416 703192 254432 703256
rect 254496 703192 254512 703256
rect 254576 703192 254592 703256
rect 254656 703192 254672 703256
rect 254736 703192 254752 703256
rect 254816 703192 254822 703256
rect 254266 703176 254822 703192
rect 254266 703112 254272 703176
rect 254336 703112 254352 703176
rect 254416 703112 254432 703176
rect 254496 703112 254512 703176
rect 254576 703112 254592 703176
rect 254656 703112 254672 703176
rect 254736 703112 254752 703176
rect 254816 703112 254822 703176
rect 254266 703096 254822 703112
rect 254266 703032 254272 703096
rect 254336 703032 254352 703096
rect 254416 703032 254432 703096
rect 254496 703032 254512 703096
rect 254576 703032 254592 703096
rect 254656 703032 254672 703096
rect 254736 703032 254752 703096
rect 254816 703032 254822 703096
rect 326266 703312 326272 703376
rect 326336 703312 326352 703376
rect 326416 703312 326432 703376
rect 326496 703312 326512 703376
rect 326576 703312 326592 703376
rect 326656 703312 326672 703376
rect 326736 703312 326752 703376
rect 326816 703312 326822 703376
rect 326266 703296 326822 703312
rect 326266 703232 326272 703296
rect 326336 703232 326352 703296
rect 326416 703232 326432 703296
rect 326496 703232 326512 703296
rect 326576 703232 326592 703296
rect 326656 703232 326672 703296
rect 326736 703232 326752 703296
rect 326816 703232 326822 703296
rect 326266 703216 326822 703232
rect 326266 703152 326272 703216
rect 326336 703152 326352 703216
rect 326416 703152 326432 703216
rect 326496 703152 326512 703216
rect 326576 703152 326592 703216
rect 326656 703152 326672 703216
rect 326736 703152 326752 703216
rect 326816 703152 326822 703216
rect 326266 703136 326822 703152
rect 326266 703072 326272 703136
rect 326336 703072 326352 703136
rect 326416 703072 326432 703136
rect 326496 703072 326512 703136
rect 326576 703072 326592 703136
rect 326656 703072 326672 703136
rect 326736 703072 326752 703136
rect 326816 703072 326822 703136
rect 326266 703071 326822 703072
rect 254266 703031 254822 703032
rect 362266 702907 362822 702908
rect 362266 702843 362272 702907
rect 362336 702843 362352 702907
rect 362416 702843 362432 702907
rect 362496 702843 362512 702907
rect 362576 702843 362592 702907
rect 362656 702843 362672 702907
rect 362736 702843 362752 702907
rect 362816 702843 362822 702907
rect 362266 702827 362822 702843
rect 362266 702763 362272 702827
rect 362336 702763 362352 702827
rect 362416 702763 362432 702827
rect 362496 702763 362512 702827
rect 362576 702763 362592 702827
rect 362656 702763 362672 702827
rect 362736 702763 362752 702827
rect 362816 702763 362822 702827
rect 362266 702747 362822 702763
rect 362266 702683 362272 702747
rect 362336 702683 362352 702747
rect 362416 702683 362432 702747
rect 362496 702683 362512 702747
rect 362576 702683 362592 702747
rect 362656 702683 362672 702747
rect 362736 702683 362752 702747
rect 362816 702683 362822 702747
rect 362266 702667 362822 702683
rect 325026 702608 325582 702609
rect 253026 702568 253582 702569
rect 253026 702504 253032 702568
rect 253096 702504 253112 702568
rect 253176 702504 253192 702568
rect 253256 702504 253272 702568
rect 253336 702504 253352 702568
rect 253416 702504 253432 702568
rect 253496 702504 253512 702568
rect 253576 702504 253582 702568
rect 253026 702488 253582 702504
rect 253026 702424 253032 702488
rect 253096 702424 253112 702488
rect 253176 702424 253192 702488
rect 253256 702424 253272 702488
rect 253336 702424 253352 702488
rect 253416 702424 253432 702488
rect 253496 702424 253512 702488
rect 253576 702424 253582 702488
rect 253026 702408 253582 702424
rect 253026 702344 253032 702408
rect 253096 702344 253112 702408
rect 253176 702344 253192 702408
rect 253256 702344 253272 702408
rect 253336 702344 253352 702408
rect 253416 702344 253432 702408
rect 253496 702344 253512 702408
rect 253576 702344 253582 702408
rect 253026 702328 253582 702344
rect 253026 702264 253032 702328
rect 253096 702264 253112 702328
rect 253176 702264 253192 702328
rect 253256 702264 253272 702328
rect 253336 702264 253352 702328
rect 253416 702264 253432 702328
rect 253496 702264 253512 702328
rect 253576 702264 253582 702328
rect 325026 702544 325032 702608
rect 325096 702544 325112 702608
rect 325176 702544 325192 702608
rect 325256 702544 325272 702608
rect 325336 702544 325352 702608
rect 325416 702544 325432 702608
rect 325496 702544 325512 702608
rect 325576 702544 325582 702608
rect 362266 702603 362272 702667
rect 362336 702603 362352 702667
rect 362416 702603 362432 702667
rect 362496 702603 362512 702667
rect 362576 702603 362592 702667
rect 362656 702603 362672 702667
rect 362736 702603 362752 702667
rect 362816 702603 362822 702667
rect 362266 702602 362822 702603
rect 434266 702770 434822 702771
rect 434266 702706 434272 702770
rect 434336 702706 434352 702770
rect 434416 702706 434432 702770
rect 434496 702706 434512 702770
rect 434576 702706 434592 702770
rect 434656 702706 434672 702770
rect 434736 702706 434752 702770
rect 434816 702706 434822 702770
rect 434266 702690 434822 702706
rect 434266 702626 434272 702690
rect 434336 702626 434352 702690
rect 434416 702626 434432 702690
rect 434496 702626 434512 702690
rect 434576 702626 434592 702690
rect 434656 702626 434672 702690
rect 434736 702626 434752 702690
rect 434816 702626 434822 702690
rect 434266 702610 434822 702626
rect 325026 702528 325582 702544
rect 325026 702464 325032 702528
rect 325096 702464 325112 702528
rect 325176 702464 325192 702528
rect 325256 702464 325272 702528
rect 325336 702464 325352 702528
rect 325416 702464 325432 702528
rect 325496 702464 325512 702528
rect 325576 702464 325582 702528
rect 434266 702546 434272 702610
rect 434336 702546 434352 702610
rect 434416 702546 434432 702610
rect 434496 702546 434512 702610
rect 434576 702546 434592 702610
rect 434656 702546 434672 702610
rect 434736 702546 434752 702610
rect 434816 702546 434822 702610
rect 434266 702530 434822 702546
rect 434266 702466 434272 702530
rect 434336 702466 434352 702530
rect 434416 702466 434432 702530
rect 434496 702466 434512 702530
rect 434576 702466 434592 702530
rect 434656 702466 434672 702530
rect 434736 702466 434752 702530
rect 434816 702466 434822 702530
rect 434266 702465 434822 702466
rect 506266 702524 506822 702525
rect 325026 702448 325582 702464
rect 325026 702384 325032 702448
rect 325096 702384 325112 702448
rect 325176 702384 325192 702448
rect 325256 702384 325272 702448
rect 325336 702384 325352 702448
rect 325416 702384 325432 702448
rect 325496 702384 325512 702448
rect 325576 702384 325582 702448
rect 325026 702368 325582 702384
rect 325026 702304 325032 702368
rect 325096 702304 325112 702368
rect 325176 702304 325192 702368
rect 325256 702304 325272 702368
rect 325336 702304 325352 702368
rect 325416 702304 325432 702368
rect 325496 702304 325512 702368
rect 325576 702304 325582 702368
rect 325026 702303 325582 702304
rect 506266 702460 506272 702524
rect 506336 702460 506352 702524
rect 506416 702460 506432 702524
rect 506496 702460 506512 702524
rect 506576 702460 506592 702524
rect 506656 702460 506672 702524
rect 506736 702460 506752 702524
rect 506816 702460 506822 702524
rect 506266 702444 506822 702460
rect 506266 702380 506272 702444
rect 506336 702380 506352 702444
rect 506416 702380 506432 702444
rect 506496 702380 506512 702444
rect 506576 702380 506592 702444
rect 506656 702380 506672 702444
rect 506736 702380 506752 702444
rect 506816 702380 506822 702444
rect 506266 702364 506822 702380
rect 253026 702263 253582 702264
rect 506266 702300 506272 702364
rect 506336 702300 506352 702364
rect 506416 702300 506432 702364
rect 506496 702300 506512 702364
rect 506576 702300 506592 702364
rect 506656 702300 506672 702364
rect 506736 702300 506752 702364
rect 506816 702300 506822 702364
rect 506266 702284 506822 702300
rect 506266 702220 506272 702284
rect 506336 702220 506352 702284
rect 506416 702220 506432 702284
rect 506496 702220 506512 702284
rect 506576 702220 506592 702284
rect 506656 702220 506672 702284
rect 506736 702220 506752 702284
rect 506816 702220 506822 702284
rect 506266 702219 506822 702220
rect 361026 702139 361582 702140
rect 361026 702075 361032 702139
rect 361096 702075 361112 702139
rect 361176 702075 361192 702139
rect 361256 702075 361272 702139
rect 361336 702075 361352 702139
rect 361416 702075 361432 702139
rect 361496 702075 361512 702139
rect 361576 702075 361582 702139
rect 361026 702059 361582 702075
rect 361026 701995 361032 702059
rect 361096 701995 361112 702059
rect 361176 701995 361192 702059
rect 361256 701995 361272 702059
rect 361336 701995 361352 702059
rect 361416 701995 361432 702059
rect 361496 701995 361512 702059
rect 361576 701995 361582 702059
rect 361026 701979 361582 701995
rect 361026 701915 361032 701979
rect 361096 701915 361112 701979
rect 361176 701915 361192 701979
rect 361256 701915 361272 701979
rect 361336 701915 361352 701979
rect 361416 701915 361432 701979
rect 361496 701915 361512 701979
rect 361576 701915 361582 701979
rect 361026 701899 361582 701915
rect 361026 701835 361032 701899
rect 361096 701835 361112 701899
rect 361176 701835 361192 701899
rect 361256 701835 361272 701899
rect 361336 701835 361352 701899
rect 361416 701835 361432 701899
rect 361496 701835 361512 701899
rect 361576 701835 361582 701899
rect 361026 701834 361582 701835
rect 433026 702002 433582 702003
rect 433026 701938 433032 702002
rect 433096 701938 433112 702002
rect 433176 701938 433192 702002
rect 433256 701938 433272 702002
rect 433336 701938 433352 702002
rect 433416 701938 433432 702002
rect 433496 701938 433512 702002
rect 433576 701938 433582 702002
rect 433026 701922 433582 701938
rect 433026 701858 433032 701922
rect 433096 701858 433112 701922
rect 433176 701858 433192 701922
rect 433256 701858 433272 701922
rect 433336 701858 433352 701922
rect 433416 701858 433432 701922
rect 433496 701858 433512 701922
rect 433576 701858 433582 701922
rect 433026 701842 433582 701858
rect 433026 701778 433032 701842
rect 433096 701778 433112 701842
rect 433176 701778 433192 701842
rect 433256 701778 433272 701842
rect 433336 701778 433352 701842
rect 433416 701778 433432 701842
rect 433496 701778 433512 701842
rect 433576 701778 433582 701842
rect 433026 701762 433582 701778
rect 433026 701698 433032 701762
rect 433096 701698 433112 701762
rect 433176 701698 433192 701762
rect 433256 701698 433272 701762
rect 433336 701698 433352 701762
rect 433416 701698 433432 701762
rect 433496 701698 433512 701762
rect 433576 701698 433582 701762
rect 433026 701697 433582 701698
rect 505026 701756 505582 701757
rect 505026 701692 505032 701756
rect 505096 701692 505112 701756
rect 505176 701692 505192 701756
rect 505256 701692 505272 701756
rect 505336 701692 505352 701756
rect 505416 701692 505432 701756
rect 505496 701692 505512 701756
rect 505576 701692 505582 701756
rect 505026 701676 505582 701692
rect 505026 701612 505032 701676
rect 505096 701612 505112 701676
rect 505176 701612 505192 701676
rect 505256 701612 505272 701676
rect 505336 701612 505352 701676
rect 505416 701612 505432 701676
rect 505496 701612 505512 701676
rect 505576 701612 505582 701676
rect 505026 701596 505582 701612
rect 505026 701532 505032 701596
rect 505096 701532 505112 701596
rect 505176 701532 505192 701596
rect 505256 701532 505272 701596
rect 505336 701532 505352 701596
rect 505416 701532 505432 701596
rect 505496 701532 505512 701596
rect 505576 701532 505582 701596
rect 505026 701516 505582 701532
rect 505026 701452 505032 701516
rect 505096 701452 505112 701516
rect 505176 701452 505192 701516
rect 505256 701452 505272 701516
rect 505336 701452 505352 701516
rect 505416 701452 505432 701516
rect 505496 701452 505512 701516
rect 505576 701452 505582 701516
rect 505026 701451 505582 701452
rect 478505 700772 478571 700775
rect 547965 700772 548031 700775
rect 478505 700770 548031 700772
rect 478505 700714 478510 700770
rect 478566 700714 547970 700770
rect 548026 700714 548031 700770
rect 478505 700712 548031 700714
rect 478505 700709 478571 700712
rect 547965 700709 548031 700712
rect 413645 700636 413711 700639
rect 547873 700636 547939 700639
rect 413645 700634 547939 700636
rect 413645 700578 413650 700634
rect 413706 700578 547878 700634
rect 547934 700578 547939 700634
rect 413645 700576 547939 700578
rect 413645 700573 413711 700576
rect 547873 700573 547939 700576
rect 348785 700500 348851 700503
rect 547413 700500 547479 700503
rect 348785 700498 547479 700500
rect 348785 700442 348790 700498
rect 348846 700442 547418 700498
rect 547474 700442 547479 700498
rect 348785 700440 547479 700442
rect 348785 700437 348851 700440
rect 547413 700437 547479 700440
rect 283833 700364 283899 700367
rect 547321 700364 547387 700367
rect 283833 700362 547387 700364
rect 283833 700306 283838 700362
rect 283894 700306 547326 700362
rect 547382 700306 547387 700362
rect 283833 700304 547387 700306
rect 283833 700301 283899 700304
rect 547321 700301 547387 700304
rect 543457 699820 543523 699823
rect 548057 699820 548123 699823
rect 543457 699818 548123 699820
rect 543457 699762 543462 699818
rect 543518 699762 548062 699818
rect 548118 699762 548123 699818
rect 543457 699760 548123 699762
rect 543457 699757 543523 699760
rect 548057 699757 548123 699760
rect 577026 697910 577582 697911
rect 577026 697846 577032 697910
rect 577096 697846 577112 697910
rect 577176 697846 577192 697910
rect 577256 697846 577272 697910
rect 577336 697846 577352 697910
rect 577416 697846 577432 697910
rect 577496 697846 577512 697910
rect 577576 697846 577582 697910
rect 577026 697830 577582 697846
rect 577026 697766 577032 697830
rect 577096 697766 577112 697830
rect 577176 697766 577192 697830
rect 577256 697766 577272 697830
rect 577336 697766 577352 697830
rect 577416 697766 577432 697830
rect 577496 697766 577512 697830
rect 577576 697766 577582 697830
rect 577026 697750 577582 697766
rect 577026 697686 577032 697750
rect 577096 697686 577112 697750
rect 577176 697686 577192 697750
rect 577256 697686 577272 697750
rect 577336 697686 577352 697750
rect 577416 697686 577432 697750
rect 577496 697686 577512 697750
rect 577576 697686 577582 697750
rect 577026 697670 577582 697686
rect 577026 697606 577032 697670
rect 577096 697606 577112 697670
rect 577176 697606 577192 697670
rect 577256 697606 577272 697670
rect 577336 697606 577352 697670
rect 577416 697606 577432 697670
rect 577496 697606 577512 697670
rect 577576 697606 577582 697670
rect 577026 697605 577582 697606
rect -960 697222 480 697462
rect 576600 697238 576666 697240
rect 580901 697238 580967 697239
rect 576600 697236 581237 697238
rect 583520 697236 584960 697326
rect 576600 697235 584960 697236
rect 576600 697179 576605 697235
rect 576661 697234 584960 697235
rect 576661 697179 580906 697234
rect 576600 697178 580906 697179
rect 580962 697178 584960 697234
rect 576600 697176 584960 697178
rect 576600 697174 576666 697176
rect 580901 697173 580967 697176
rect 578266 697115 578822 697116
rect 578266 697051 578272 697115
rect 578336 697051 578352 697115
rect 578416 697051 578432 697115
rect 578496 697051 578512 697115
rect 578576 697051 578592 697115
rect 578656 697051 578672 697115
rect 578736 697051 578752 697115
rect 578816 697051 578822 697115
rect 583520 697086 584960 697176
rect 578266 697035 578822 697051
rect 578266 696971 578272 697035
rect 578336 696971 578352 697035
rect 578416 696971 578432 697035
rect 578496 696971 578512 697035
rect 578576 696971 578592 697035
rect 578656 696971 578672 697035
rect 578736 696971 578752 697035
rect 578816 696971 578822 697035
rect 578266 696955 578822 696971
rect 578266 696891 578272 696955
rect 578336 696891 578352 696955
rect 578416 696891 578432 696955
rect 578496 696891 578512 696955
rect 578576 696891 578592 696955
rect 578656 696891 578672 696955
rect 578736 696891 578752 696955
rect 578816 696891 578822 696955
rect 578266 696875 578822 696891
rect 578266 696811 578272 696875
rect 578336 696811 578352 696875
rect 578416 696811 578432 696875
rect 578496 696811 578512 696875
rect 578576 696811 578592 696875
rect 578656 696811 578672 696875
rect 578736 696811 578752 696875
rect 578816 696811 578822 696875
rect 578266 696810 578822 696811
rect -960 684166 480 684406
rect 583520 683758 584960 683998
rect -960 671110 480 671350
rect 580257 670716 580323 670719
rect 583520 670716 584960 670806
rect 580257 670714 584960 670716
rect 580257 670658 580262 670714
rect 580318 670658 584960 670714
rect 580257 670656 584960 670658
rect 580257 670653 580323 670656
rect 583520 670566 584960 670656
rect -960 658054 480 658294
rect 583520 657238 584960 657478
rect -960 644998 480 645238
rect 577026 644734 577582 644735
rect 577026 644670 577032 644734
rect 577096 644670 577112 644734
rect 577176 644670 577192 644734
rect 577256 644670 577272 644734
rect 577336 644670 577352 644734
rect 577416 644670 577432 644734
rect 577496 644670 577512 644734
rect 577576 644670 577582 644734
rect 577026 644654 577582 644670
rect 577026 644590 577032 644654
rect 577096 644590 577112 644654
rect 577176 644590 577192 644654
rect 577256 644590 577272 644654
rect 577336 644590 577352 644654
rect 577416 644590 577432 644654
rect 577496 644590 577512 644654
rect 577576 644590 577582 644654
rect 577026 644574 577582 644590
rect 577026 644510 577032 644574
rect 577096 644510 577112 644574
rect 577176 644510 577192 644574
rect 577256 644510 577272 644574
rect 577336 644510 577352 644574
rect 577416 644510 577432 644574
rect 577496 644510 577512 644574
rect 577576 644510 577582 644574
rect 577026 644494 577582 644510
rect 577026 644430 577032 644494
rect 577096 644430 577112 644494
rect 577176 644430 577192 644494
rect 577256 644430 577272 644494
rect 577336 644430 577352 644494
rect 577416 644430 577432 644494
rect 577496 644430 577512 644494
rect 577576 644430 577582 644494
rect 577026 644429 577582 644430
rect 576600 644062 576666 644064
rect 580901 644062 580967 644063
rect 576600 644060 581164 644062
rect 583520 644060 584960 644150
rect 576600 644059 584960 644060
rect 576600 644003 576605 644059
rect 576661 644058 584960 644059
rect 576661 644003 580906 644058
rect 576600 644002 580906 644003
rect 580962 644002 584960 644058
rect 576600 644000 584960 644002
rect 576600 643998 576666 644000
rect 580901 643997 580967 644000
rect 578266 643939 578822 643940
rect 578266 643875 578272 643939
rect 578336 643875 578352 643939
rect 578416 643875 578432 643939
rect 578496 643875 578512 643939
rect 578576 643875 578592 643939
rect 578656 643875 578672 643939
rect 578736 643875 578752 643939
rect 578816 643875 578822 643939
rect 583520 643910 584960 644000
rect 578266 643859 578822 643875
rect 578266 643795 578272 643859
rect 578336 643795 578352 643859
rect 578416 643795 578432 643859
rect 578496 643795 578512 643859
rect 578576 643795 578592 643859
rect 578656 643795 578672 643859
rect 578736 643795 578752 643859
rect 578816 643795 578822 643859
rect 578266 643779 578822 643795
rect 578266 643715 578272 643779
rect 578336 643715 578352 643779
rect 578416 643715 578432 643779
rect 578496 643715 578512 643779
rect 578576 643715 578592 643779
rect 578656 643715 578672 643779
rect 578736 643715 578752 643779
rect 578816 643715 578822 643779
rect 578266 643699 578822 643715
rect 578266 643635 578272 643699
rect 578336 643635 578352 643699
rect 578416 643635 578432 643699
rect 578496 643635 578512 643699
rect 578576 643635 578592 643699
rect 578656 643635 578672 643699
rect 578736 643635 578752 643699
rect 578816 643635 578822 643699
rect 578266 643634 578822 643635
rect -960 631942 480 632182
rect 583520 630718 584960 630958
rect -960 619022 480 619262
rect 580441 617540 580507 617543
rect 583520 617540 584960 617630
rect 580441 617538 584960 617540
rect 580441 617482 580446 617538
rect 580502 617482 584960 617538
rect 580441 617480 584960 617482
rect 580441 617477 580507 617480
rect 583520 617390 584960 617480
rect -960 605966 480 606206
rect 583520 604062 584960 604302
rect -960 592910 480 593150
rect 577026 591694 577582 591695
rect 577026 591630 577032 591694
rect 577096 591630 577112 591694
rect 577176 591630 577192 591694
rect 577256 591630 577272 591694
rect 577336 591630 577352 591694
rect 577416 591630 577432 591694
rect 577496 591630 577512 591694
rect 577576 591630 577582 591694
rect 577026 591614 577582 591630
rect 577026 591550 577032 591614
rect 577096 591550 577112 591614
rect 577176 591550 577192 591614
rect 577256 591550 577272 591614
rect 577336 591550 577352 591614
rect 577416 591550 577432 591614
rect 577496 591550 577512 591614
rect 577576 591550 577582 591614
rect 577026 591534 577582 591550
rect 577026 591470 577032 591534
rect 577096 591470 577112 591534
rect 577176 591470 577192 591534
rect 577256 591470 577272 591534
rect 577336 591470 577352 591534
rect 577416 591470 577432 591534
rect 577496 591470 577512 591534
rect 577576 591470 577582 591534
rect 577026 591454 577582 591470
rect 577026 591390 577032 591454
rect 577096 591390 577112 591454
rect 577176 591390 577192 591454
rect 577256 591390 577272 591454
rect 577336 591390 577352 591454
rect 577416 591390 577432 591454
rect 577496 591390 577512 591454
rect 577576 591390 577582 591454
rect 577026 591389 577582 591390
rect 576600 591022 576666 591024
rect 580901 591022 580967 591023
rect 576600 591020 581271 591022
rect 583520 591020 584960 591110
rect 576600 591019 584960 591020
rect 576600 590963 576605 591019
rect 576661 591018 584960 591019
rect 576661 590963 580906 591018
rect 576600 590962 580906 590963
rect 580962 590962 584960 591018
rect 576600 590960 584960 590962
rect 576600 590958 576666 590960
rect 580901 590957 580967 590960
rect 578266 590899 578822 590900
rect 578266 590835 578272 590899
rect 578336 590835 578352 590899
rect 578416 590835 578432 590899
rect 578496 590835 578512 590899
rect 578576 590835 578592 590899
rect 578656 590835 578672 590899
rect 578736 590835 578752 590899
rect 578816 590835 578822 590899
rect 583520 590870 584960 590960
rect 578266 590819 578822 590835
rect 578266 590755 578272 590819
rect 578336 590755 578352 590819
rect 578416 590755 578432 590819
rect 578496 590755 578512 590819
rect 578576 590755 578592 590819
rect 578656 590755 578672 590819
rect 578736 590755 578752 590819
rect 578816 590755 578822 590819
rect 578266 590739 578822 590755
rect 578266 590675 578272 590739
rect 578336 590675 578352 590739
rect 578416 590675 578432 590739
rect 578496 590675 578512 590739
rect 578576 590675 578592 590739
rect 578656 590675 578672 590739
rect 578736 590675 578752 590739
rect 578816 590675 578822 590739
rect 578266 590659 578822 590675
rect 578266 590595 578272 590659
rect 578336 590595 578352 590659
rect 578416 590595 578432 590659
rect 578496 590595 578512 590659
rect 578576 590595 578592 590659
rect 578656 590595 578672 590659
rect 578736 590595 578752 590659
rect 578816 590595 578822 590659
rect 578266 590594 578822 590595
rect -960 579854 480 580094
rect 583520 577542 584960 577782
rect -960 566798 480 567038
rect 580625 564364 580691 564367
rect 583520 564364 584960 564454
rect 580625 564362 584960 564364
rect 580625 564306 580630 564362
rect 580686 564306 584960 564362
rect 580625 564304 584960 564306
rect 580625 564301 580691 564304
rect 583520 564214 584960 564304
rect 505026 554602 505582 554603
rect 505026 554538 505032 554602
rect 505096 554538 505112 554602
rect 505176 554538 505192 554602
rect 505256 554538 505272 554602
rect 505336 554538 505352 554602
rect 505416 554538 505432 554602
rect 505496 554538 505512 554602
rect 505576 554538 505582 554602
rect 505026 554522 505582 554538
rect 505026 554458 505032 554522
rect 505096 554458 505112 554522
rect 505176 554458 505192 554522
rect 505256 554458 505272 554522
rect 505336 554458 505352 554522
rect 505416 554458 505432 554522
rect 505496 554458 505512 554522
rect 505576 554458 505582 554522
rect 505026 554442 505582 554458
rect 505026 554378 505032 554442
rect 505096 554378 505112 554442
rect 505176 554378 505192 554442
rect 505256 554378 505272 554442
rect 505336 554378 505352 554442
rect 505416 554378 505432 554442
rect 505496 554378 505512 554442
rect 505576 554378 505582 554442
rect 505026 554362 505582 554378
rect 505026 554298 505032 554362
rect 505096 554298 505112 554362
rect 505176 554298 505192 554362
rect 505256 554298 505272 554362
rect 505336 554298 505352 554362
rect 505416 554298 505432 554362
rect 505496 554298 505512 554362
rect 505576 554298 505582 554362
rect 505026 554297 505582 554298
rect -960 553742 480 553982
rect 506266 553807 506822 553808
rect 506266 553743 506272 553807
rect 506336 553743 506352 553807
rect 506416 553743 506432 553807
rect 506496 553743 506512 553807
rect 506576 553743 506592 553807
rect 506656 553743 506672 553807
rect 506736 553743 506752 553807
rect 506816 553743 506822 553807
rect 506266 553727 506822 553743
rect 506266 553663 506272 553727
rect 506336 553663 506352 553727
rect 506416 553663 506432 553727
rect 506496 553663 506512 553727
rect 506576 553663 506592 553727
rect 506656 553663 506672 553727
rect 506736 553663 506752 553727
rect 506816 553663 506822 553727
rect 506266 553647 506822 553663
rect 506266 553583 506272 553647
rect 506336 553583 506352 553647
rect 506416 553583 506432 553647
rect 506496 553583 506512 553647
rect 506576 553583 506592 553647
rect 506656 553583 506672 553647
rect 506736 553583 506752 553647
rect 506816 553583 506822 553647
rect 506266 553567 506822 553583
rect 506266 553503 506272 553567
rect 506336 553503 506352 553567
rect 506416 553503 506432 553567
rect 506496 553503 506512 553567
rect 506576 553503 506592 553567
rect 506656 553503 506672 553567
rect 506736 553503 506752 553567
rect 506816 553503 506822 553567
rect 506266 553502 506822 553503
rect 583520 551022 584960 551262
rect -960 540686 480 540926
rect 577026 538518 577582 538519
rect 577026 538454 577032 538518
rect 577096 538454 577112 538518
rect 577176 538454 577192 538518
rect 577256 538454 577272 538518
rect 577336 538454 577352 538518
rect 577416 538454 577432 538518
rect 577496 538454 577512 538518
rect 577576 538454 577582 538518
rect 577026 538438 577582 538454
rect 577026 538374 577032 538438
rect 577096 538374 577112 538438
rect 577176 538374 577192 538438
rect 577256 538374 577272 538438
rect 577336 538374 577352 538438
rect 577416 538374 577432 538438
rect 577496 538374 577512 538438
rect 577576 538374 577582 538438
rect 577026 538358 577582 538374
rect 577026 538294 577032 538358
rect 577096 538294 577112 538358
rect 577176 538294 577192 538358
rect 577256 538294 577272 538358
rect 577336 538294 577352 538358
rect 577416 538294 577432 538358
rect 577496 538294 577512 538358
rect 577576 538294 577582 538358
rect 577026 538278 577582 538294
rect 577026 538214 577032 538278
rect 577096 538214 577112 538278
rect 577176 538214 577192 538278
rect 577256 538214 577272 538278
rect 577336 538214 577352 538278
rect 577416 538214 577432 538278
rect 577496 538214 577512 538278
rect 577576 538214 577582 538278
rect 577026 538213 577582 538214
rect 576600 537846 576666 537848
rect 580901 537846 580967 537847
rect 576600 537844 581074 537846
rect 583520 537844 584960 537934
rect 576600 537843 584960 537844
rect 576600 537787 576605 537843
rect 576661 537842 584960 537843
rect 576661 537787 580906 537842
rect 576600 537786 580906 537787
rect 580962 537786 584960 537842
rect 576600 537784 584960 537786
rect 576600 537782 576666 537784
rect 580901 537781 580967 537784
rect 578266 537723 578822 537724
rect 578266 537659 578272 537723
rect 578336 537659 578352 537723
rect 578416 537659 578432 537723
rect 578496 537659 578512 537723
rect 578576 537659 578592 537723
rect 578656 537659 578672 537723
rect 578736 537659 578752 537723
rect 578816 537659 578822 537723
rect 583520 537694 584960 537784
rect 578266 537643 578822 537659
rect 578266 537579 578272 537643
rect 578336 537579 578352 537643
rect 578416 537579 578432 537643
rect 578496 537579 578512 537643
rect 578576 537579 578592 537643
rect 578656 537579 578672 537643
rect 578736 537579 578752 537643
rect 578816 537579 578822 537643
rect 578266 537563 578822 537579
rect 578266 537499 578272 537563
rect 578336 537499 578352 537563
rect 578416 537499 578432 537563
rect 578496 537499 578512 537563
rect 578576 537499 578592 537563
rect 578656 537499 578672 537563
rect 578736 537499 578752 537563
rect 578816 537499 578822 537563
rect 578266 537483 578822 537499
rect 578266 537419 578272 537483
rect 578336 537419 578352 537483
rect 578416 537419 578432 537483
rect 578496 537419 578512 537483
rect 578576 537419 578592 537483
rect 578656 537419 578672 537483
rect 578736 537419 578752 537483
rect 578816 537419 578822 537483
rect 578266 537418 578822 537419
rect -960 527766 480 528006
rect 583520 524366 584960 524606
rect -960 514710 480 514950
rect 580809 511324 580875 511327
rect 583520 511324 584960 511414
rect 580809 511322 584960 511324
rect 580809 511266 580814 511322
rect 580870 511266 584960 511322
rect 580809 511264 584960 511266
rect 580809 511261 580875 511264
rect 583520 511174 584960 511264
rect -960 501654 480 501894
rect 583520 497846 584960 498086
rect -960 488598 480 488838
rect 577026 485342 577582 485343
rect 577026 485278 577032 485342
rect 577096 485278 577112 485342
rect 577176 485278 577192 485342
rect 577256 485278 577272 485342
rect 577336 485278 577352 485342
rect 577416 485278 577432 485342
rect 577496 485278 577512 485342
rect 577576 485278 577582 485342
rect 577026 485262 577582 485278
rect 577026 485198 577032 485262
rect 577096 485198 577112 485262
rect 577176 485198 577192 485262
rect 577256 485198 577272 485262
rect 577336 485198 577352 485262
rect 577416 485198 577432 485262
rect 577496 485198 577512 485262
rect 577576 485198 577582 485262
rect 577026 485182 577582 485198
rect 577026 485118 577032 485182
rect 577096 485118 577112 485182
rect 577176 485118 577192 485182
rect 577256 485118 577272 485182
rect 577336 485118 577352 485182
rect 577416 485118 577432 485182
rect 577496 485118 577512 485182
rect 577576 485118 577582 485182
rect 577026 485102 577582 485118
rect 577026 485038 577032 485102
rect 577096 485038 577112 485102
rect 577176 485038 577192 485102
rect 577256 485038 577272 485102
rect 577336 485038 577352 485102
rect 577416 485038 577432 485102
rect 577496 485038 577512 485102
rect 577576 485038 577582 485102
rect 577026 485037 577582 485038
rect 576600 484670 576666 484672
rect 580901 484670 580967 484671
rect 576600 484668 581277 484670
rect 583520 484668 584960 484758
rect 576600 484667 584960 484668
rect 576600 484611 576605 484667
rect 576661 484666 584960 484667
rect 576661 484611 580906 484666
rect 576600 484610 580906 484611
rect 580962 484610 584960 484666
rect 576600 484608 584960 484610
rect 576600 484606 576666 484608
rect 580901 484605 580967 484608
rect 578266 484547 578822 484548
rect 578266 484483 578272 484547
rect 578336 484483 578352 484547
rect 578416 484483 578432 484547
rect 578496 484483 578512 484547
rect 578576 484483 578592 484547
rect 578656 484483 578672 484547
rect 578736 484483 578752 484547
rect 578816 484483 578822 484547
rect 583520 484518 584960 484608
rect 578266 484467 578822 484483
rect 578266 484403 578272 484467
rect 578336 484403 578352 484467
rect 578416 484403 578432 484467
rect 578496 484403 578512 484467
rect 578576 484403 578592 484467
rect 578656 484403 578672 484467
rect 578736 484403 578752 484467
rect 578816 484403 578822 484467
rect 578266 484387 578822 484403
rect 578266 484323 578272 484387
rect 578336 484323 578352 484387
rect 578416 484323 578432 484387
rect 578496 484323 578512 484387
rect 578576 484323 578592 484387
rect 578656 484323 578672 484387
rect 578736 484323 578752 484387
rect 578816 484323 578822 484387
rect 578266 484307 578822 484323
rect 578266 484243 578272 484307
rect 578336 484243 578352 484307
rect 578416 484243 578432 484307
rect 578496 484243 578512 484307
rect 578576 484243 578592 484307
rect 578656 484243 578672 484307
rect 578736 484243 578752 484307
rect 578816 484243 578822 484307
rect 578266 484242 578822 484243
rect -960 475542 480 475782
rect 583520 471326 584960 471566
rect -960 462486 480 462726
rect 580165 458148 580231 458151
rect 583520 458148 584960 458238
rect 580165 458146 584960 458148
rect 580165 458090 580170 458146
rect 580226 458090 584960 458146
rect 580165 458088 584960 458090
rect 580165 458085 580231 458088
rect 583520 457998 584960 458088
rect 470266 451485 470822 451486
rect 470266 451421 470272 451485
rect 470336 451421 470352 451485
rect 470416 451421 470432 451485
rect 470496 451421 470512 451485
rect 470576 451421 470592 451485
rect 470656 451421 470672 451485
rect 470736 451421 470752 451485
rect 470816 451421 470822 451485
rect 470266 451405 470822 451421
rect 470266 451341 470272 451405
rect 470336 451341 470352 451405
rect 470416 451341 470432 451405
rect 470496 451341 470512 451405
rect 470576 451341 470592 451405
rect 470656 451341 470672 451405
rect 470736 451341 470752 451405
rect 470816 451341 470822 451405
rect 470266 451325 470822 451341
rect 470266 451261 470272 451325
rect 470336 451261 470352 451325
rect 470416 451261 470432 451325
rect 470496 451261 470512 451325
rect 470576 451261 470592 451325
rect 470656 451261 470672 451325
rect 470736 451261 470752 451325
rect 470816 451261 470822 451325
rect 470266 451245 470822 451261
rect 470266 451181 470272 451245
rect 470336 451181 470352 451245
rect 470416 451181 470432 451245
rect 470496 451181 470512 451245
rect 470576 451181 470592 451245
rect 470656 451181 470672 451245
rect 470736 451181 470752 451245
rect 470816 451181 470822 451245
rect 470266 451180 470822 451181
rect 469026 450399 469582 450400
rect 469026 450335 469032 450399
rect 469096 450335 469112 450399
rect 469176 450335 469192 450399
rect 469256 450335 469272 450399
rect 469336 450335 469352 450399
rect 469416 450335 469432 450399
rect 469496 450335 469512 450399
rect 469576 450335 469582 450399
rect 469026 450319 469582 450335
rect 469026 450255 469032 450319
rect 469096 450255 469112 450319
rect 469176 450255 469192 450319
rect 469256 450255 469272 450319
rect 469336 450255 469352 450319
rect 469416 450255 469432 450319
rect 469496 450255 469512 450319
rect 469576 450255 469582 450319
rect 469026 450239 469582 450255
rect 469026 450175 469032 450239
rect 469096 450175 469112 450239
rect 469176 450175 469192 450239
rect 469256 450175 469272 450239
rect 469336 450175 469352 450239
rect 469416 450175 469432 450239
rect 469496 450175 469512 450239
rect 469576 450175 469582 450239
rect 477838 450260 477904 450263
rect 481155 450262 481221 450263
rect 487788 450262 487854 450263
rect 478454 450260 478460 450262
rect 477838 450258 478460 450260
rect 477838 450202 477843 450258
rect 477899 450202 478460 450258
rect 477838 450200 478460 450202
rect 477838 450197 477904 450200
rect 478454 450198 478460 450200
rect 478524 450198 478530 450262
rect 481155 450258 481220 450262
rect 481155 450202 481160 450258
rect 481216 450202 481220 450258
rect 481155 450198 481220 450202
rect 481284 450260 481290 450262
rect 481284 450200 481312 450260
rect 487788 450258 487844 450262
rect 487908 450260 487914 450262
rect 487788 450202 487793 450258
rect 481284 450198 481290 450200
rect 487788 450198 487844 450202
rect 487908 450200 487945 450260
rect 487908 450198 487914 450200
rect 481155 450197 481221 450198
rect 487788 450197 487854 450198
rect 469026 450159 469582 450175
rect 469026 450095 469032 450159
rect 469096 450095 469112 450159
rect 469176 450095 469192 450159
rect 469256 450095 469272 450159
rect 469336 450095 469352 450159
rect 469416 450095 469432 450159
rect 469496 450095 469512 450159
rect 469576 450095 469582 450159
rect 469026 450094 469582 450095
rect -960 449430 480 449670
rect 473670 449654 473676 449718
rect 473740 449716 473746 449718
rect 474089 449716 474155 449719
rect 473740 449714 474155 449716
rect 473740 449658 474094 449714
rect 474150 449658 474155 449714
rect 473740 449656 474155 449658
rect 473740 449654 473746 449656
rect 474089 449653 474155 449656
rect 470266 449314 470822 449315
rect 470266 449250 470272 449314
rect 470336 449250 470352 449314
rect 470416 449250 470432 449314
rect 470496 449250 470512 449314
rect 470576 449250 470592 449314
rect 470656 449250 470672 449314
rect 470736 449250 470752 449314
rect 470816 449250 470822 449314
rect 470266 449234 470822 449250
rect 470266 449170 470272 449234
rect 470336 449170 470352 449234
rect 470416 449170 470432 449234
rect 470496 449170 470512 449234
rect 470576 449170 470592 449234
rect 470656 449170 470672 449234
rect 470736 449170 470752 449234
rect 470816 449170 470822 449234
rect 470266 449154 470822 449170
rect 470266 449090 470272 449154
rect 470336 449090 470352 449154
rect 470416 449090 470432 449154
rect 470496 449090 470512 449154
rect 470576 449090 470592 449154
rect 470656 449090 470672 449154
rect 470736 449090 470752 449154
rect 470816 449090 470822 449154
rect 470266 449074 470822 449090
rect 470266 449010 470272 449074
rect 470336 449010 470352 449074
rect 470416 449010 470432 449074
rect 470496 449010 470512 449074
rect 470576 449010 470592 449074
rect 470656 449010 470672 449074
rect 470736 449010 470752 449074
rect 470816 449010 470822 449074
rect 470266 449009 470822 449010
rect 546677 448084 546743 448087
rect 580257 448084 580323 448087
rect 546677 448082 580323 448084
rect 546677 448026 546682 448082
rect 546738 448026 580262 448082
rect 580318 448026 580323 448082
rect 546677 448024 580323 448026
rect 546677 448021 546743 448024
rect 580257 448021 580323 448024
rect 544193 447948 544259 447951
rect 580441 447948 580507 447951
rect 544193 447946 580507 447948
rect 544193 447890 544198 447946
rect 544254 447890 580446 447946
rect 580502 447890 580507 447946
rect 544193 447888 580507 447890
rect 544193 447885 544259 447888
rect 580441 447885 580507 447888
rect 539225 447812 539291 447815
rect 580809 447812 580875 447815
rect 539225 447810 580875 447812
rect 539225 447754 539230 447810
rect 539286 447754 580814 447810
rect 580870 447754 580875 447810
rect 539225 447752 580875 447754
rect 539225 447749 539291 447752
rect 580809 447749 580875 447752
rect 541709 447268 541775 447271
rect 580625 447268 580691 447271
rect 541709 447266 580691 447268
rect 541709 447210 541714 447266
rect 541770 447210 580630 447266
rect 580686 447210 580691 447266
rect 541709 447208 580691 447210
rect 541709 447205 541775 447208
rect 580625 447205 580691 447208
rect 544193 445772 544259 445775
rect 544326 445772 544332 445774
rect 544193 445770 544332 445772
rect 544193 445714 544198 445770
rect 544254 445714 544332 445770
rect 544193 445712 544332 445714
rect 544193 445709 544259 445712
rect 544326 445710 544332 445712
rect 544396 445710 544402 445774
rect 541566 445302 541572 445366
rect 541636 445364 541642 445366
rect 541709 445364 541775 445367
rect 541636 445362 541775 445364
rect 541636 445306 541714 445362
rect 541770 445306 541775 445362
rect 541636 445304 541775 445306
rect 541636 445302 541642 445304
rect 541709 445301 541775 445304
rect 535453 444820 535519 444823
rect 535453 444818 538108 444820
rect 535453 444762 535458 444818
rect 535514 444762 538108 444818
rect 535453 444760 538108 444762
rect 535453 444757 535519 444760
rect 583520 444670 584960 444910
rect 535453 443460 535519 443463
rect 535453 443458 538108 443460
rect 535453 443402 535458 443458
rect 535514 443402 538108 443458
rect 535453 443400 538108 443402
rect 535453 443397 535519 443400
rect 535453 442100 535519 442103
rect 535453 442098 538108 442100
rect 535453 442042 535458 442098
rect 535514 442042 538108 442098
rect 535453 442040 538108 442042
rect 535453 442037 535519 442040
rect 535453 440740 535519 440743
rect 535453 440738 538108 440740
rect 535453 440682 535458 440738
rect 535514 440682 538108 440738
rect 535453 440680 538108 440682
rect 535453 440677 535519 440680
rect 535453 439380 535519 439383
rect 535453 439378 538108 439380
rect 535453 439322 535458 439378
rect 535514 439322 538108 439378
rect 535453 439320 538108 439322
rect 535453 439317 535519 439320
rect 535453 438020 535519 438023
rect 535453 438018 538108 438020
rect 535453 437962 535458 438018
rect 535514 437962 538108 438018
rect 535453 437960 538108 437962
rect 535453 437957 535519 437960
rect -960 436510 480 436750
rect 535453 436660 535519 436663
rect 535453 436658 538108 436660
rect 535453 436602 535458 436658
rect 535514 436602 538108 436658
rect 535453 436600 538108 436602
rect 535453 436597 535519 436600
rect 548057 435436 548123 435439
rect 547830 435434 548123 435436
rect 547830 435378 548062 435434
rect 548118 435378 548123 435434
rect 547830 435376 548123 435378
rect 535453 435300 535519 435303
rect 535453 435298 538108 435300
rect 535453 435242 535458 435298
rect 535514 435242 538108 435298
rect 535453 435240 538108 435242
rect 535453 435237 535519 435240
rect 547830 434726 547890 435376
rect 548057 435373 548123 435376
rect 535453 433940 535519 433943
rect 535453 433938 538108 433940
rect 535453 433882 535458 433938
rect 535514 433882 538108 433938
rect 535453 433880 538108 433882
rect 535453 433877 535519 433880
rect 470266 433086 470822 433087
rect 470266 433022 470272 433086
rect 470336 433022 470352 433086
rect 470416 433022 470432 433086
rect 470496 433022 470512 433086
rect 470576 433022 470592 433086
rect 470656 433022 470672 433086
rect 470736 433022 470752 433086
rect 470816 433022 470822 433086
rect 470266 433006 470822 433022
rect 470266 432942 470272 433006
rect 470336 432942 470352 433006
rect 470416 432942 470432 433006
rect 470496 432942 470512 433006
rect 470576 432942 470592 433006
rect 470656 432942 470672 433006
rect 470736 432942 470752 433006
rect 470816 432942 470822 433006
rect 470266 432926 470822 432942
rect 470266 432862 470272 432926
rect 470336 432862 470352 432926
rect 470416 432862 470432 432926
rect 470496 432862 470512 432926
rect 470576 432862 470592 432926
rect 470656 432862 470672 432926
rect 470736 432862 470752 432926
rect 470816 432862 470822 432926
rect 470266 432846 470822 432862
rect 483657 432854 483723 432855
rect 483606 432852 483612 432854
rect 470266 432782 470272 432846
rect 470336 432782 470352 432846
rect 470416 432782 470432 432846
rect 470496 432782 470512 432846
rect 470576 432782 470592 432846
rect 470656 432782 470672 432846
rect 470736 432782 470752 432846
rect 470816 432782 470822 432846
rect 483566 432792 483612 432852
rect 483676 432850 483723 432854
rect 483718 432794 483723 432850
rect 483606 432790 483612 432792
rect 483676 432790 483723 432794
rect 483657 432789 483723 432790
rect 470266 432781 470822 432782
rect 535453 432580 535519 432583
rect 535453 432578 538108 432580
rect 535453 432522 535458 432578
rect 535514 432522 538108 432578
rect 535453 432520 538108 432522
rect 535453 432517 535519 432520
rect 483565 432310 483631 432311
rect 483565 432308 483612 432310
rect 483520 432306 483612 432308
rect 483520 432250 483570 432306
rect 483520 432248 483612 432250
rect 483565 432246 483612 432248
rect 483676 432246 483682 432310
rect 577026 432302 577582 432303
rect 483565 432245 483631 432246
rect 577026 432238 577032 432302
rect 577096 432238 577112 432302
rect 577176 432238 577192 432302
rect 577256 432238 577272 432302
rect 577336 432238 577352 432302
rect 577416 432238 577432 432302
rect 577496 432238 577512 432302
rect 577576 432238 577582 432302
rect 577026 432222 577582 432238
rect 481265 432174 481331 432175
rect 481214 432110 481220 432174
rect 481284 432172 481331 432174
rect 481284 432170 481376 432172
rect 481326 432114 481376 432170
rect 481284 432112 481376 432114
rect 577026 432158 577032 432222
rect 577096 432158 577112 432222
rect 577176 432158 577192 432222
rect 577256 432158 577272 432222
rect 577336 432158 577352 432222
rect 577416 432158 577432 432222
rect 577496 432158 577512 432222
rect 577576 432158 577582 432222
rect 577026 432142 577582 432158
rect 481284 432110 481331 432112
rect 481265 432109 481331 432110
rect 577026 432078 577032 432142
rect 577096 432078 577112 432142
rect 577176 432078 577192 432142
rect 577256 432078 577272 432142
rect 577336 432078 577352 432142
rect 577416 432078 577432 432142
rect 577496 432078 577512 432142
rect 577576 432078 577582 432142
rect 577026 432062 577582 432078
rect 469026 431999 469582 432000
rect 469026 431935 469032 431999
rect 469096 431935 469112 431999
rect 469176 431935 469192 431999
rect 469256 431935 469272 431999
rect 469336 431935 469352 431999
rect 469416 431935 469432 431999
rect 469496 431935 469512 431999
rect 469576 431935 469582 431999
rect 577026 431998 577032 432062
rect 577096 431998 577112 432062
rect 577176 431998 577192 432062
rect 577256 431998 577272 432062
rect 577336 431998 577352 432062
rect 577416 431998 577432 432062
rect 577496 431998 577512 432062
rect 577576 431998 577582 432062
rect 577026 431997 577582 431998
rect 469026 431919 469582 431935
rect 469026 431855 469032 431919
rect 469096 431855 469112 431919
rect 469176 431855 469192 431919
rect 469256 431855 469272 431919
rect 469336 431855 469352 431919
rect 469416 431855 469432 431919
rect 469496 431855 469512 431919
rect 469576 431855 469582 431919
rect 469026 431839 469582 431855
rect 469026 431775 469032 431839
rect 469096 431775 469112 431839
rect 469176 431775 469192 431839
rect 469256 431775 469272 431839
rect 469336 431775 469352 431839
rect 469416 431775 469432 431839
rect 469496 431775 469512 431839
rect 469576 431775 469582 431839
rect 473670 431838 473676 431902
rect 473740 431900 473746 431902
rect 474273 431900 474339 431903
rect 473740 431898 474339 431900
rect 473740 431842 474278 431898
rect 474334 431842 474339 431898
rect 473740 431840 474339 431842
rect 473740 431838 473746 431840
rect 474273 431837 474339 431840
rect 469026 431759 469582 431775
rect 469026 431695 469032 431759
rect 469096 431695 469112 431759
rect 469176 431695 469192 431759
rect 469256 431695 469272 431759
rect 469336 431695 469352 431759
rect 469416 431695 469432 431759
rect 469496 431695 469512 431759
rect 469576 431695 469582 431759
rect 469026 431694 469582 431695
rect 478097 431628 478163 431631
rect 488428 431630 488494 431631
rect 478454 431628 478460 431630
rect 478097 431626 478460 431628
rect 478097 431570 478102 431626
rect 478158 431570 478460 431626
rect 478097 431568 478460 431570
rect 478097 431565 478163 431568
rect 478454 431566 478460 431568
rect 478524 431566 478530 431630
rect 488390 431566 488396 431630
rect 488460 431628 488494 431630
rect 576600 431630 576666 431632
rect 580901 431630 580967 431631
rect 576600 431628 581169 431630
rect 583520 431628 584960 431718
rect 488460 431626 488552 431628
rect 488489 431570 488552 431626
rect 488460 431568 488552 431570
rect 576600 431627 584960 431628
rect 576600 431571 576605 431627
rect 576661 431626 584960 431627
rect 576661 431571 580906 431626
rect 576600 431570 580906 431571
rect 580962 431570 584960 431626
rect 576600 431568 584960 431570
rect 488460 431566 488494 431568
rect 576600 431566 576666 431568
rect 488428 431565 488494 431566
rect 580901 431565 580967 431568
rect 578266 431507 578822 431508
rect 578266 431443 578272 431507
rect 578336 431443 578352 431507
rect 578416 431443 578432 431507
rect 578496 431443 578512 431507
rect 578576 431443 578592 431507
rect 578656 431443 578672 431507
rect 578736 431443 578752 431507
rect 578816 431443 578822 431507
rect 583520 431478 584960 431568
rect 578266 431427 578822 431443
rect 578266 431363 578272 431427
rect 578336 431363 578352 431427
rect 578416 431363 578432 431427
rect 578496 431363 578512 431427
rect 578576 431363 578592 431427
rect 578656 431363 578672 431427
rect 578736 431363 578752 431427
rect 578816 431363 578822 431427
rect 578266 431347 578822 431363
rect 578266 431283 578272 431347
rect 578336 431283 578352 431347
rect 578416 431283 578432 431347
rect 578496 431283 578512 431347
rect 578576 431283 578592 431347
rect 578656 431283 578672 431347
rect 578736 431283 578752 431347
rect 578816 431283 578822 431347
rect 578266 431267 578822 431283
rect 536097 431220 536163 431223
rect 536097 431218 538108 431220
rect 536097 431162 536102 431218
rect 536158 431190 538108 431218
rect 578266 431203 578272 431267
rect 578336 431203 578352 431267
rect 578416 431203 578432 431267
rect 578496 431203 578512 431267
rect 578576 431203 578592 431267
rect 578656 431203 578672 431267
rect 578736 431203 578752 431267
rect 578816 431203 578822 431267
rect 578266 431202 578822 431203
rect 536158 431162 538138 431190
rect 536097 431160 538138 431162
rect 536097 431157 536163 431160
rect 470266 430914 470822 430915
rect 470266 430850 470272 430914
rect 470336 430850 470352 430914
rect 470416 430850 470432 430914
rect 470496 430850 470512 430914
rect 470576 430850 470592 430914
rect 470656 430850 470672 430914
rect 470736 430850 470752 430914
rect 470816 430850 470822 430914
rect 470266 430834 470822 430850
rect 470266 430770 470272 430834
rect 470336 430770 470352 430834
rect 470416 430770 470432 430834
rect 470496 430770 470512 430834
rect 470576 430770 470592 430834
rect 470656 430770 470672 430834
rect 470736 430770 470752 430834
rect 470816 430770 470822 430834
rect 470266 430754 470822 430770
rect 470266 430690 470272 430754
rect 470336 430690 470352 430754
rect 470416 430690 470432 430754
rect 470496 430690 470512 430754
rect 470576 430690 470592 430754
rect 470656 430690 470672 430754
rect 470736 430690 470752 430754
rect 470816 430690 470822 430754
rect 470266 430674 470822 430690
rect 470266 430610 470272 430674
rect 470336 430610 470352 430674
rect 470416 430610 470432 430674
rect 470496 430610 470512 430674
rect 470576 430610 470592 430674
rect 470656 430610 470672 430674
rect 470736 430610 470752 430674
rect 470816 430610 470822 430674
rect 470266 430609 470822 430610
rect 478965 427956 479031 427959
rect 480110 427956 480116 427958
rect 478965 427954 480116 427956
rect 478965 427898 478970 427954
rect 479026 427898 480116 427954
rect 478965 427896 480116 427898
rect 478965 427893 479031 427896
rect 480110 427894 480116 427896
rect 480180 427894 480186 427958
rect 485773 427956 485839 427959
rect 486550 427956 486556 427958
rect 485773 427954 486556 427956
rect 485773 427898 485778 427954
rect 485834 427898 486556 427954
rect 485773 427896 486556 427898
rect 485773 427893 485839 427896
rect 486550 427894 486556 427896
rect 486620 427894 486626 427958
rect 536741 424420 536807 424423
rect 538078 424420 538138 431160
rect 536741 424418 538138 424420
rect 536741 424362 536746 424418
rect 536802 424390 538138 424418
rect 536802 424362 538108 424390
rect 536741 424360 538108 424362
rect 536741 424357 536807 424360
rect -960 423454 480 423694
rect 583520 418150 584960 418390
rect 488390 413886 488396 413950
rect 488460 413948 488466 413950
rect 488533 413948 488599 413951
rect 488460 413946 488599 413948
rect 488460 413890 488538 413946
rect 488594 413890 488599 413946
rect 488460 413888 488599 413890
rect 488460 413886 488466 413888
rect 488533 413885 488599 413888
rect 470266 412086 470822 412087
rect 470266 412022 470272 412086
rect 470336 412022 470352 412086
rect 470416 412022 470432 412086
rect 470496 412022 470512 412086
rect 470576 412022 470592 412086
rect 470656 412022 470672 412086
rect 470736 412022 470752 412086
rect 470816 412022 470822 412086
rect 470266 412006 470822 412022
rect 470266 411942 470272 412006
rect 470336 411942 470352 412006
rect 470416 411942 470432 412006
rect 470496 411942 470512 412006
rect 470576 411942 470592 412006
rect 470656 411942 470672 412006
rect 470736 411942 470752 412006
rect 470816 411942 470822 412006
rect 470266 411926 470822 411942
rect 470266 411862 470272 411926
rect 470336 411862 470352 411926
rect 470416 411862 470432 411926
rect 470496 411862 470512 411926
rect 470576 411862 470592 411926
rect 470656 411862 470672 411926
rect 470736 411862 470752 411926
rect 470816 411862 470822 411926
rect 470266 411846 470822 411862
rect 470266 411782 470272 411846
rect 470336 411782 470352 411846
rect 470416 411782 470432 411846
rect 470496 411782 470512 411846
rect 470576 411782 470592 411846
rect 470656 411782 470672 411846
rect 470736 411782 470752 411846
rect 470816 411782 470822 411846
rect 470266 411781 470822 411782
rect 469026 411000 469582 411001
rect 469026 410936 469032 411000
rect 469096 410936 469112 411000
rect 469176 410936 469192 411000
rect 469256 410936 469272 411000
rect 469336 410936 469352 411000
rect 469416 410936 469432 411000
rect 469496 410936 469512 411000
rect 469576 410936 469582 411000
rect 473721 410958 473787 410959
rect 469026 410920 469582 410936
rect 469026 410856 469032 410920
rect 469096 410856 469112 410920
rect 469176 410856 469192 410920
rect 469256 410856 469272 410920
rect 469336 410856 469352 410920
rect 469416 410856 469432 410920
rect 469496 410856 469512 410920
rect 469576 410856 469582 410920
rect 473670 410894 473676 410958
rect 473740 410956 473787 410958
rect 473740 410954 473832 410956
rect 473782 410898 473832 410954
rect 473740 410896 473832 410898
rect 473740 410894 473787 410896
rect 473721 410893 473787 410894
rect 469026 410840 469582 410856
rect 469026 410776 469032 410840
rect 469096 410776 469112 410840
rect 469176 410776 469192 410840
rect 469256 410776 469272 410840
rect 469336 410776 469352 410840
rect 469416 410776 469432 410840
rect 469496 410776 469512 410840
rect 469576 410776 469582 410840
rect 469026 410760 469582 410776
rect 469026 410696 469032 410760
rect 469096 410696 469112 410760
rect 469176 410696 469192 410760
rect 469256 410696 469272 410760
rect 469336 410696 469352 410760
rect 469416 410696 469432 410760
rect 469496 410696 469512 410760
rect 469576 410696 469582 410760
rect 469026 410695 469582 410696
rect -960 410398 480 410638
rect 484117 410414 484183 410415
rect 484117 410412 484164 410414
rect 484072 410410 484164 410412
rect 484072 410354 484122 410410
rect 484072 410352 484164 410354
rect 484117 410350 484164 410352
rect 484228 410350 484234 410414
rect 484117 410349 484183 410350
rect 478413 410142 478479 410143
rect 481357 410142 481423 410143
rect 478413 410140 478460 410142
rect 478368 410138 478460 410140
rect 478368 410082 478418 410138
rect 478368 410080 478460 410082
rect 478413 410078 478460 410080
rect 478524 410078 478530 410142
rect 481357 410140 481404 410142
rect 481312 410138 481404 410140
rect 481312 410082 481362 410138
rect 481312 410080 481404 410082
rect 481357 410078 481404 410080
rect 481468 410078 481474 410142
rect 478413 410077 478479 410078
rect 481357 410077 481423 410078
rect 487613 410004 487679 410007
rect 488533 410004 488599 410007
rect 489821 410004 489887 410007
rect 580165 410004 580231 410007
rect 487613 410002 580231 410004
rect 487613 409946 487618 410002
rect 487674 409946 488538 410002
rect 488594 409946 489826 410002
rect 489882 409946 580170 410002
rect 580226 409946 580231 410002
rect 487613 409944 580231 409946
rect 487613 409941 487679 409944
rect 488533 409941 488599 409944
rect 489821 409941 489887 409944
rect 580165 409941 580231 409944
rect 470266 409914 470822 409915
rect 470266 409850 470272 409914
rect 470336 409850 470352 409914
rect 470416 409850 470432 409914
rect 470496 409850 470512 409914
rect 470576 409850 470592 409914
rect 470656 409850 470672 409914
rect 470736 409850 470752 409914
rect 470816 409850 470822 409914
rect 470266 409834 470822 409850
rect 470266 409770 470272 409834
rect 470336 409770 470352 409834
rect 470416 409770 470432 409834
rect 470496 409770 470512 409834
rect 470576 409770 470592 409834
rect 470656 409770 470672 409834
rect 470736 409770 470752 409834
rect 470816 409770 470822 409834
rect 470266 409754 470822 409770
rect 470266 409690 470272 409754
rect 470336 409690 470352 409754
rect 470416 409690 470432 409754
rect 470496 409690 470512 409754
rect 470576 409690 470592 409754
rect 470656 409690 470672 409754
rect 470736 409690 470752 409754
rect 470816 409690 470822 409754
rect 470266 409674 470822 409690
rect 470266 409610 470272 409674
rect 470336 409610 470352 409674
rect 470416 409610 470432 409674
rect 470496 409610 470512 409674
rect 470576 409610 470592 409674
rect 470656 409610 470672 409674
rect 470736 409610 470752 409674
rect 470816 409610 470822 409674
rect 470266 409609 470822 409610
rect 535453 409324 535519 409327
rect 535453 409322 538138 409324
rect 535453 409266 535458 409322
rect 535514 409266 538138 409322
rect 535453 409264 538138 409266
rect 535453 409261 535519 409264
rect 538078 408818 538138 409264
rect 541566 409262 541572 409326
rect 541636 409324 541642 409326
rect 541709 409324 541775 409327
rect 544285 409326 544351 409327
rect 544285 409324 544332 409326
rect 541636 409322 541775 409324
rect 541636 409266 541714 409322
rect 541770 409266 541775 409322
rect 541636 409264 541775 409266
rect 544240 409322 544332 409324
rect 544240 409266 544290 409322
rect 544240 409264 544332 409266
rect 541636 409262 541642 409264
rect 541709 409261 541775 409264
rect 544285 409262 544332 409264
rect 544396 409262 544402 409326
rect 544285 409261 544351 409262
rect 480110 407494 480116 407558
rect 480180 407556 480186 407558
rect 480180 407496 538138 407556
rect 480180 407494 480186 407496
rect 538078 407458 538138 407496
rect 481817 407148 481883 407151
rect 482870 407148 482876 407150
rect 481817 407146 482876 407148
rect 481817 407090 481822 407146
rect 481878 407090 482876 407146
rect 481817 407088 482876 407090
rect 481817 407085 481883 407088
rect 482870 407086 482876 407088
rect 482940 407086 482946 407150
rect 485129 407148 485195 407151
rect 485630 407148 485636 407150
rect 485129 407146 485636 407148
rect 485129 407090 485134 407146
rect 485190 407090 485636 407146
rect 485129 407088 485636 407090
rect 485129 407085 485195 407088
rect 485630 407086 485636 407088
rect 485700 407086 485706 407150
rect 535453 406604 535519 406607
rect 535453 406602 538138 406604
rect 535453 406546 535458 406602
rect 535514 406546 538138 406602
rect 535453 406544 538138 406546
rect 535453 406541 535519 406544
rect 538078 406098 538138 406544
rect 580165 404972 580231 404975
rect 583520 404972 584960 405062
rect 580165 404970 584960 404972
rect 580165 404914 580170 404970
rect 580226 404914 584960 404970
rect 580165 404912 584960 404914
rect 580165 404909 580231 404912
rect 583520 404822 584960 404912
rect 535453 404564 535519 404567
rect 538078 404564 538138 404738
rect 535453 404562 538138 404564
rect 535453 404506 535458 404562
rect 535514 404506 538138 404562
rect 535453 404504 538138 404506
rect 535453 404501 535519 404504
rect 535453 403204 535519 403207
rect 538078 403204 538138 403378
rect 535453 403202 538138 403204
rect 535453 403146 535458 403202
rect 535514 403146 538138 403202
rect 535453 403144 538138 403146
rect 535453 403141 535519 403144
rect 536373 401708 536439 401711
rect 538078 401708 538138 402018
rect 536373 401706 538138 401708
rect 536373 401650 536378 401706
rect 536434 401650 538138 401706
rect 536373 401648 538138 401650
rect 536373 401645 536439 401648
rect 536281 400348 536347 400351
rect 538078 400348 538138 400658
rect 536281 400346 538138 400348
rect 536281 400290 536286 400346
rect 536342 400290 538138 400346
rect 536281 400288 538138 400290
rect 536281 400285 536347 400288
rect 535453 399124 535519 399127
rect 538078 399124 538138 399298
rect 535453 399122 538138 399124
rect 535453 399066 535458 399122
rect 535514 399066 538138 399122
rect 535453 399064 538138 399066
rect 535453 399061 535519 399064
rect 547830 398580 547890 398754
rect 547965 398580 548031 398583
rect 547830 398578 548031 398580
rect 547830 398522 547970 398578
rect 548026 398522 548031 398578
rect 547830 398520 548031 398522
rect 547965 398517 548031 398520
rect -960 397342 480 397582
rect 536097 397492 536163 397495
rect 538078 397492 538138 397938
rect 536097 397490 538138 397492
rect 536097 397434 536102 397490
rect 536158 397434 538138 397490
rect 536097 397432 538138 397434
rect 536097 397429 536163 397432
rect 535453 396404 535519 396407
rect 538078 396404 538138 396578
rect 535453 396402 538138 396404
rect 535453 396346 535458 396402
rect 535514 396346 538138 396402
rect 535453 396344 538138 396346
rect 535453 396341 535519 396344
rect 536741 395996 536807 395999
rect 536741 395994 538138 395996
rect 536741 395938 536746 395994
rect 536802 395938 538138 395994
rect 536741 395936 538138 395938
rect 536741 395933 536807 395936
rect 473670 391990 473676 392054
rect 473740 392052 473746 392054
rect 474958 392052 474964 392054
rect 473740 391992 474964 392052
rect 473740 391990 473746 391992
rect 474958 391990 474964 391992
rect 475028 391990 475034 392054
rect 489310 391990 489316 392054
rect 489380 392052 489386 392054
rect 489821 392052 489887 392055
rect 489380 392050 489887 392052
rect 489380 391994 489826 392050
rect 489882 391994 489887 392050
rect 489380 391992 489887 391994
rect 489380 391990 489386 391992
rect 489821 391989 489887 391992
rect 470266 391087 470822 391088
rect 470266 391023 470272 391087
rect 470336 391023 470352 391087
rect 470416 391023 470432 391087
rect 470496 391023 470512 391087
rect 470576 391023 470592 391087
rect 470656 391023 470672 391087
rect 470736 391023 470752 391087
rect 470816 391023 470822 391087
rect 470266 391007 470822 391023
rect 470266 390943 470272 391007
rect 470336 390943 470352 391007
rect 470416 390943 470432 391007
rect 470496 390943 470512 391007
rect 470576 390943 470592 391007
rect 470656 390943 470672 391007
rect 470736 390943 470752 391007
rect 470816 390943 470822 391007
rect 470266 390927 470822 390943
rect 470266 390863 470272 390927
rect 470336 390863 470352 390927
rect 470416 390863 470432 390927
rect 470496 390863 470512 390927
rect 470576 390863 470592 390927
rect 470656 390863 470672 390927
rect 470736 390863 470752 390927
rect 470816 390863 470822 390927
rect 470266 390847 470822 390863
rect 470266 390783 470272 390847
rect 470336 390783 470352 390847
rect 470416 390783 470432 390847
rect 470496 390783 470512 390847
rect 470576 390783 470592 390847
rect 470656 390783 470672 390847
rect 470736 390783 470752 390847
rect 470816 390783 470822 390847
rect 470266 390782 470822 390783
rect 484900 390299 484964 390305
rect 484900 390229 484964 390235
rect 469026 390004 469582 390005
rect 469026 389940 469032 390004
rect 469096 389940 469112 390004
rect 469176 389940 469192 390004
rect 469256 389940 469272 390004
rect 469336 389940 469352 390004
rect 469416 389940 469432 390004
rect 469496 389940 469512 390004
rect 469576 389940 469582 390004
rect 469026 389924 469582 389940
rect 469026 389860 469032 389924
rect 469096 389860 469112 389924
rect 469176 389860 469192 389924
rect 469256 389860 469272 389924
rect 469336 389860 469352 389924
rect 469416 389860 469432 389924
rect 469496 389860 469512 389924
rect 469576 389860 469582 389924
rect 469026 389844 469582 389860
rect 469026 389780 469032 389844
rect 469096 389780 469112 389844
rect 469176 389780 469192 389844
rect 469256 389780 469272 389844
rect 469336 389780 469352 389844
rect 469416 389780 469432 389844
rect 469496 389780 469512 389844
rect 469576 389780 469582 389844
rect 469026 389764 469582 389780
rect 469026 389700 469032 389764
rect 469096 389700 469112 389764
rect 469176 389700 469192 389764
rect 469256 389700 469272 389764
rect 469336 389700 469352 389764
rect 469416 389700 469432 389764
rect 469496 389700 469512 389764
rect 469576 389700 469582 389764
rect 469026 389699 469582 389700
rect 481766 389406 481772 389470
rect 481836 389468 481842 389470
rect 482093 389468 482159 389471
rect 489361 389470 489427 389471
rect 481836 389466 482159 389468
rect 481836 389410 482098 389466
rect 482154 389410 482159 389466
rect 481836 389408 482159 389410
rect 481836 389406 481842 389408
rect 482093 389405 482159 389408
rect 489310 389406 489316 389470
rect 489380 389468 489427 389470
rect 489380 389466 489472 389468
rect 489422 389410 489472 389466
rect 489380 389408 489472 389410
rect 489380 389406 489427 389408
rect 489361 389405 489427 389406
rect 474917 389334 474983 389335
rect 478629 389334 478695 389335
rect 474917 389332 474964 389334
rect 474872 389330 474964 389332
rect 474872 389274 474922 389330
rect 474872 389272 474964 389274
rect 474917 389270 474964 389272
rect 475028 389270 475034 389334
rect 478629 389332 478644 389334
rect 478552 389330 478644 389332
rect 478552 389274 478634 389330
rect 478552 389272 478644 389274
rect 478629 389270 478644 389272
rect 478708 389270 478714 389334
rect 474917 389269 474983 389270
rect 478629 389269 478695 389270
rect 470266 388914 470822 388915
rect 470266 388850 470272 388914
rect 470336 388850 470352 388914
rect 470416 388850 470432 388914
rect 470496 388850 470512 388914
rect 470576 388850 470592 388914
rect 470656 388850 470672 388914
rect 470736 388850 470752 388914
rect 470816 388850 470822 388914
rect 470266 388834 470822 388850
rect 470266 388770 470272 388834
rect 470336 388770 470352 388834
rect 470416 388770 470432 388834
rect 470496 388770 470512 388834
rect 470576 388770 470592 388834
rect 470656 388770 470672 388834
rect 470736 388770 470752 388834
rect 470816 388770 470822 388834
rect 470266 388754 470822 388770
rect 470266 388690 470272 388754
rect 470336 388690 470352 388754
rect 470416 388690 470432 388754
rect 470496 388690 470512 388754
rect 470576 388690 470592 388754
rect 470656 388690 470672 388754
rect 470736 388690 470752 388754
rect 470816 388690 470822 388754
rect 470266 388674 470822 388690
rect 470266 388610 470272 388674
rect 470336 388610 470352 388674
rect 470416 388610 470432 388674
rect 470496 388610 470512 388674
rect 470576 388610 470592 388674
rect 470656 388610 470672 388674
rect 470736 388610 470752 388674
rect 470816 388610 470822 388674
rect 470266 388609 470822 388610
rect 536741 388380 536807 388383
rect 538078 388380 538138 395936
rect 583520 391630 584960 391870
rect 536741 388378 538138 388380
rect 536741 388322 536746 388378
rect 536802 388322 538138 388378
rect 536741 388320 538138 388322
rect 536741 388317 536807 388320
rect 486734 386414 486740 386478
rect 486804 386476 486810 386478
rect 486877 386476 486943 386479
rect 486804 386474 486943 386476
rect 486804 386418 486882 386474
rect 486938 386418 486943 386474
rect 486804 386416 486943 386418
rect 486804 386414 486810 386416
rect 486877 386413 486943 386416
rect -960 384286 480 384526
rect 577026 379126 577582 379127
rect 577026 379062 577032 379126
rect 577096 379062 577112 379126
rect 577176 379062 577192 379126
rect 577256 379062 577272 379126
rect 577336 379062 577352 379126
rect 577416 379062 577432 379126
rect 577496 379062 577512 379126
rect 577576 379062 577582 379126
rect 577026 379046 577582 379062
rect 577026 378982 577032 379046
rect 577096 378982 577112 379046
rect 577176 378982 577192 379046
rect 577256 378982 577272 379046
rect 577336 378982 577352 379046
rect 577416 378982 577432 379046
rect 577496 378982 577512 379046
rect 577576 378982 577582 379046
rect 577026 378966 577582 378982
rect 577026 378902 577032 378966
rect 577096 378902 577112 378966
rect 577176 378902 577192 378966
rect 577256 378902 577272 378966
rect 577336 378902 577352 378966
rect 577416 378902 577432 378966
rect 577496 378902 577512 378966
rect 577576 378902 577582 378966
rect 577026 378886 577582 378902
rect 577026 378822 577032 378886
rect 577096 378822 577112 378886
rect 577176 378822 577192 378886
rect 577256 378822 577272 378886
rect 577336 378822 577352 378886
rect 577416 378822 577432 378886
rect 577496 378822 577512 378886
rect 577576 378822 577582 378886
rect 577026 378821 577582 378822
rect 576600 378454 576666 378456
rect 580901 378454 580967 378455
rect 576600 378452 581533 378454
rect 583520 378452 584960 378542
rect 576600 378451 584960 378452
rect 576600 378395 576605 378451
rect 576661 378450 584960 378451
rect 576661 378395 580906 378450
rect 576600 378394 580906 378395
rect 580962 378394 584960 378450
rect 576600 378392 584960 378394
rect 576600 378390 576666 378392
rect 580901 378389 580967 378392
rect 578266 378331 578822 378332
rect 578266 378267 578272 378331
rect 578336 378267 578352 378331
rect 578416 378267 578432 378331
rect 578496 378267 578512 378331
rect 578576 378267 578592 378331
rect 578656 378267 578672 378331
rect 578736 378267 578752 378331
rect 578816 378267 578822 378331
rect 583520 378302 584960 378392
rect 578266 378251 578822 378267
rect 578266 378187 578272 378251
rect 578336 378187 578352 378251
rect 578416 378187 578432 378251
rect 578496 378187 578512 378251
rect 578576 378187 578592 378251
rect 578656 378187 578672 378251
rect 578736 378187 578752 378251
rect 578816 378187 578822 378251
rect 578266 378171 578822 378187
rect 578266 378107 578272 378171
rect 578336 378107 578352 378171
rect 578416 378107 578432 378171
rect 578496 378107 578512 378171
rect 578576 378107 578592 378171
rect 578656 378107 578672 378171
rect 578736 378107 578752 378171
rect 578816 378107 578822 378171
rect 578266 378091 578822 378107
rect 578266 378027 578272 378091
rect 578336 378027 578352 378091
rect 578416 378027 578432 378091
rect 578496 378027 578512 378091
rect 578576 378027 578592 378091
rect 578656 378027 578672 378091
rect 578736 378027 578752 378091
rect 578816 378027 578822 378091
rect 578266 378026 578822 378027
rect 541566 373086 541572 373150
rect 541636 373148 541642 373150
rect 541709 373148 541775 373151
rect 541636 373146 541775 373148
rect 541636 373090 541714 373146
rect 541770 373090 541775 373146
rect 541636 373088 541775 373090
rect 541636 373086 541642 373088
rect 541709 373085 541775 373088
rect 544193 373148 544259 373151
rect 544326 373148 544332 373150
rect 544193 373146 544332 373148
rect 544193 373090 544198 373146
rect 544254 373090 544332 373146
rect 544193 373088 544332 373090
rect 544193 373085 544259 373088
rect 544326 373086 544332 373088
rect 544396 373086 544402 373150
rect 535453 372876 535519 372879
rect 535453 372874 538108 372876
rect 535453 372818 535458 372874
rect 535514 372818 538108 372874
rect 535453 372816 538108 372818
rect 535453 372813 535519 372816
rect 535453 371516 535519 371519
rect 535453 371514 538108 371516
rect -960 371230 480 371470
rect 535453 371458 535458 371514
rect 535514 371458 538108 371514
rect 535453 371456 538108 371458
rect 535453 371453 535519 371456
rect 482870 370094 482876 370158
rect 482940 370156 482946 370158
rect 482940 370096 538108 370156
rect 482940 370094 482946 370096
rect 535453 368796 535519 368799
rect 535453 368794 538108 368796
rect 535453 368738 535458 368794
rect 535514 368738 538108 368794
rect 535453 368736 538108 368738
rect 535453 368733 535519 368736
rect 535453 367436 535519 367439
rect 535453 367434 538108 367436
rect 535453 367378 535458 367434
rect 535514 367378 538108 367434
rect 535453 367376 538108 367378
rect 535453 367373 535519 367376
rect 535453 366076 535519 366079
rect 535453 366074 538108 366076
rect 535453 366018 535458 366074
rect 535514 366018 538108 366074
rect 535453 366016 538108 366018
rect 535453 366013 535519 366016
rect 583520 364974 584960 365214
rect 536557 364716 536623 364719
rect 536557 364714 538108 364716
rect 536557 364658 536562 364714
rect 536618 364658 538108 364714
rect 536557 364656 538108 364658
rect 536557 364653 536623 364656
rect 536465 363356 536531 363359
rect 536465 363354 538108 363356
rect 536465 363298 536470 363354
rect 536526 363298 538108 363354
rect 536465 363296 538108 363298
rect 536465 363293 536531 363296
rect 547873 362948 547939 362951
rect 547830 362946 547939 362948
rect 547830 362890 547878 362946
rect 547934 362890 547939 362946
rect 547830 362885 547939 362890
rect 547830 362782 547890 362885
rect 535453 361996 535519 361999
rect 535453 361994 538108 361996
rect 535453 361938 535458 361994
rect 535514 361938 538108 361994
rect 535453 361936 538108 361938
rect 535453 361933 535519 361936
rect 536189 360636 536255 360639
rect 536189 360634 538108 360636
rect 536189 360578 536194 360634
rect 536250 360578 538108 360634
rect 536189 360576 538108 360578
rect 536189 360573 536255 360576
rect 536741 359276 536807 359279
rect 536741 359274 538108 359276
rect 536741 359218 536746 359274
rect 536802 359246 538108 359274
rect 536802 359218 538138 359246
rect 536741 359216 538138 359218
rect 536741 359213 536807 359216
rect -960 358310 480 358550
rect 470266 358487 470822 358488
rect 470266 358423 470272 358487
rect 470336 358423 470352 358487
rect 470416 358423 470432 358487
rect 470496 358423 470512 358487
rect 470576 358423 470592 358487
rect 470656 358423 470672 358487
rect 470736 358423 470752 358487
rect 470816 358423 470822 358487
rect 470266 358407 470822 358423
rect 470266 358343 470272 358407
rect 470336 358343 470352 358407
rect 470416 358343 470432 358407
rect 470496 358343 470512 358407
rect 470576 358343 470592 358407
rect 470656 358343 470672 358407
rect 470736 358343 470752 358407
rect 470816 358343 470822 358407
rect 470266 358327 470822 358343
rect 470266 358263 470272 358327
rect 470336 358263 470352 358327
rect 470416 358263 470432 358327
rect 470496 358263 470512 358327
rect 470576 358263 470592 358327
rect 470656 358263 470672 358327
rect 470736 358263 470752 358327
rect 470816 358263 470822 358327
rect 470266 358247 470822 358263
rect 470266 358183 470272 358247
rect 470336 358183 470352 358247
rect 470416 358183 470432 358247
rect 470496 358183 470512 358247
rect 470576 358183 470592 358247
rect 470656 358183 470672 358247
rect 470736 358183 470752 358247
rect 470816 358183 470822 358247
rect 470266 358182 470822 358183
rect 478638 357990 478644 358054
rect 478708 358052 478714 358054
rect 478873 358052 478939 358055
rect 481817 358054 481883 358055
rect 484945 358054 485011 358055
rect 488441 358054 488507 358055
rect 478708 358050 478939 358052
rect 478708 357994 478878 358050
rect 478934 357994 478939 358050
rect 478708 357992 478939 357994
rect 478708 357990 478714 357992
rect 478873 357989 478939 357992
rect 481766 357990 481772 358054
rect 481836 358052 481883 358054
rect 481836 358050 481928 358052
rect 481878 357994 481928 358050
rect 481836 357992 481928 357994
rect 481836 357990 481883 357992
rect 484894 357990 484900 358054
rect 484964 358052 485011 358054
rect 488390 358052 488396 358054
rect 484964 358050 485056 358052
rect 485006 357994 485056 358050
rect 484964 357992 485056 357994
rect 488314 357992 488396 358052
rect 488460 358052 488507 358054
rect 489310 358052 489316 358054
rect 488460 358050 489316 358052
rect 488502 357994 489316 358050
rect 484964 357990 485011 357992
rect 488390 357990 488396 357992
rect 488460 357992 489316 357994
rect 488460 357990 488507 357992
rect 489310 357990 489316 357992
rect 489380 357990 489386 358054
rect 481817 357989 481883 357990
rect 484945 357989 485011 357990
rect 488441 357989 488507 357990
rect 475009 357510 475075 357511
rect 474958 357446 474964 357510
rect 475028 357508 475075 357510
rect 475028 357506 475120 357508
rect 475070 357450 475120 357506
rect 475028 357448 475120 357450
rect 475028 357446 475075 357448
rect 475009 357445 475075 357446
rect 469026 357401 469582 357402
rect 469026 357337 469032 357401
rect 469096 357337 469112 357401
rect 469176 357337 469192 357401
rect 469256 357337 469272 357401
rect 469336 357337 469352 357401
rect 469416 357337 469432 357401
rect 469496 357337 469512 357401
rect 469576 357337 469582 357401
rect 469026 357321 469582 357337
rect 469026 357257 469032 357321
rect 469096 357257 469112 357321
rect 469176 357257 469192 357321
rect 469256 357257 469272 357321
rect 469336 357257 469352 357321
rect 469416 357257 469432 357321
rect 469496 357257 469512 357321
rect 469576 357257 469582 357321
rect 469026 357241 469582 357257
rect 469026 357177 469032 357241
rect 469096 357177 469112 357241
rect 469176 357177 469192 357241
rect 469256 357177 469272 357241
rect 469336 357177 469352 357241
rect 469416 357177 469432 357241
rect 469496 357177 469512 357241
rect 469576 357177 469582 357241
rect 469026 357161 469582 357177
rect 469026 357097 469032 357161
rect 469096 357097 469112 357161
rect 469176 357097 469192 357161
rect 469256 357097 469272 357161
rect 469336 357097 469352 357161
rect 469416 357097 469432 357161
rect 469496 357097 469512 357161
rect 469576 357097 469582 357161
rect 469026 357096 469582 357097
rect 470266 356314 470822 356315
rect 470266 356250 470272 356314
rect 470336 356250 470352 356314
rect 470416 356250 470432 356314
rect 470496 356250 470512 356314
rect 470576 356250 470592 356314
rect 470656 356250 470672 356314
rect 470736 356250 470752 356314
rect 470816 356250 470822 356314
rect 470266 356234 470822 356250
rect 470266 356170 470272 356234
rect 470336 356170 470352 356234
rect 470416 356170 470432 356234
rect 470496 356170 470512 356234
rect 470576 356170 470592 356234
rect 470656 356170 470672 356234
rect 470736 356170 470752 356234
rect 470816 356170 470822 356234
rect 470266 356154 470822 356170
rect 470266 356090 470272 356154
rect 470336 356090 470352 356154
rect 470416 356090 470432 356154
rect 470496 356090 470512 356154
rect 470576 356090 470592 356154
rect 470656 356090 470672 356154
rect 470736 356090 470752 356154
rect 470816 356090 470822 356154
rect 470266 356074 470822 356090
rect 470266 356010 470272 356074
rect 470336 356010 470352 356074
rect 470416 356010 470432 356074
rect 470496 356010 470512 356074
rect 470576 356010 470592 356074
rect 470656 356010 470672 356074
rect 470736 356010 470752 356074
rect 470816 356010 470822 356074
rect 470266 356009 470822 356010
rect 536741 352476 536807 352479
rect 538078 352476 538138 359216
rect 536741 352474 538138 352476
rect 536741 352418 536746 352474
rect 536802 352446 538138 352474
rect 536802 352418 538108 352446
rect 536741 352416 538108 352418
rect 536741 352413 536807 352416
rect 484577 351932 484643 351935
rect 485446 351932 485452 351934
rect 484577 351930 485452 351932
rect 484577 351874 484582 351930
rect 484638 351874 485452 351930
rect 484577 351872 485452 351874
rect 484577 351869 484643 351872
rect 485446 351870 485452 351872
rect 485516 351932 485522 351934
rect 583520 351932 584960 352022
rect 485516 351872 584960 351932
rect 485516 351870 485522 351872
rect 583520 351782 584960 351872
rect -960 345254 480 345494
rect 473670 343710 473676 343774
rect 473740 343772 473746 343774
rect 474958 343772 474964 343774
rect 473740 343712 474964 343772
rect 473740 343710 473746 343712
rect 474958 343710 474964 343712
rect 475028 343710 475034 343774
rect 470266 342486 470822 342487
rect 470266 342422 470272 342486
rect 470336 342422 470352 342486
rect 470416 342422 470432 342486
rect 470496 342422 470512 342486
rect 470576 342422 470592 342486
rect 470656 342422 470672 342486
rect 470736 342422 470752 342486
rect 470816 342422 470822 342486
rect 470266 342406 470822 342422
rect 470266 342342 470272 342406
rect 470336 342342 470352 342406
rect 470416 342342 470432 342406
rect 470496 342342 470512 342406
rect 470576 342342 470592 342406
rect 470656 342342 470672 342406
rect 470736 342342 470752 342406
rect 470816 342342 470822 342406
rect 470266 342326 470822 342342
rect 470266 342262 470272 342326
rect 470336 342262 470352 342326
rect 470416 342262 470432 342326
rect 470496 342262 470512 342326
rect 470576 342262 470592 342326
rect 470656 342262 470672 342326
rect 470736 342262 470752 342326
rect 470816 342262 470822 342326
rect 484577 342276 484643 342279
rect 470266 342246 470822 342262
rect 470266 342182 470272 342246
rect 470336 342182 470352 342246
rect 470416 342182 470432 342246
rect 470496 342182 470512 342246
rect 470576 342182 470592 342246
rect 470656 342182 470672 342246
rect 470736 342182 470752 342246
rect 470816 342182 470822 342246
rect 470266 342181 470822 342182
rect 484534 342274 484643 342276
rect 484534 342218 484582 342274
rect 484638 342218 484643 342274
rect 484534 342213 484643 342218
rect 484393 341732 484459 341735
rect 484534 341732 484594 342213
rect 484393 341730 484594 341732
rect 484393 341674 484398 341730
rect 484454 341674 484594 341730
rect 484393 341672 484594 341674
rect 484393 341669 484459 341672
rect 469026 341399 469582 341400
rect 469026 341335 469032 341399
rect 469096 341335 469112 341399
rect 469176 341335 469192 341399
rect 469256 341335 469272 341399
rect 469336 341335 469352 341399
rect 469416 341335 469432 341399
rect 469496 341335 469512 341399
rect 469576 341335 469582 341399
rect 469026 341319 469582 341335
rect 469026 341255 469032 341319
rect 469096 341255 469112 341319
rect 469176 341255 469192 341319
rect 469256 341255 469272 341319
rect 469336 341255 469352 341319
rect 469416 341255 469432 341319
rect 469496 341255 469512 341319
rect 469576 341255 469582 341319
rect 469026 341239 469582 341255
rect 469026 341175 469032 341239
rect 469096 341175 469112 341239
rect 469176 341175 469192 341239
rect 469256 341175 469272 341239
rect 469336 341175 469352 341239
rect 469416 341175 469432 341239
rect 469496 341175 469512 341239
rect 469576 341175 469582 341239
rect 469026 341159 469582 341175
rect 469026 341095 469032 341159
rect 469096 341095 469112 341159
rect 469176 341095 469192 341159
rect 469256 341095 469272 341159
rect 469336 341095 469352 341159
rect 469416 341095 469432 341159
rect 469496 341095 469512 341159
rect 469576 341095 469582 341159
rect 469026 341094 469582 341095
rect 477910 341052 477976 341055
rect 478454 341052 478460 341054
rect 477910 341050 478460 341052
rect 477910 340994 477915 341050
rect 477971 340994 478460 341050
rect 477910 340992 478460 340994
rect 477910 340989 477976 340992
rect 478454 340990 478460 340992
rect 478524 340990 478530 341054
rect 481227 341052 481293 341055
rect 481398 341052 481404 341054
rect 481227 341050 481404 341052
rect 481227 340994 481232 341050
rect 481288 340994 481404 341050
rect 481227 340992 481404 340994
rect 481227 340989 481293 340992
rect 481398 340990 481404 340992
rect 481468 340990 481474 341054
rect 487889 341052 487955 341055
rect 488022 341052 488028 341054
rect 487889 341050 488028 341052
rect 487889 340994 487894 341050
rect 487950 340994 488028 341050
rect 487889 340992 488028 340994
rect 487889 340989 487955 340992
rect 488022 340990 488028 340992
rect 488092 340990 488098 341054
rect 473670 340446 473676 340510
rect 473740 340508 473746 340510
rect 474549 340508 474615 340511
rect 473740 340506 474615 340508
rect 473740 340450 474554 340506
rect 474610 340450 474615 340506
rect 473740 340448 474615 340450
rect 473740 340446 473746 340448
rect 474549 340445 474615 340448
rect 470266 340314 470822 340315
rect 470266 340250 470272 340314
rect 470336 340250 470352 340314
rect 470416 340250 470432 340314
rect 470496 340250 470512 340314
rect 470576 340250 470592 340314
rect 470656 340250 470672 340314
rect 470736 340250 470752 340314
rect 470816 340250 470822 340314
rect 470266 340234 470822 340250
rect 470266 340170 470272 340234
rect 470336 340170 470352 340234
rect 470416 340170 470432 340234
rect 470496 340170 470512 340234
rect 470576 340170 470592 340234
rect 470656 340170 470672 340234
rect 470736 340170 470752 340234
rect 470816 340170 470822 340234
rect 470266 340154 470822 340170
rect 470266 340090 470272 340154
rect 470336 340090 470352 340154
rect 470416 340090 470432 340154
rect 470496 340090 470512 340154
rect 470576 340090 470592 340154
rect 470656 340090 470672 340154
rect 470736 340090 470752 340154
rect 470816 340090 470822 340154
rect 470266 340074 470822 340090
rect 470266 340010 470272 340074
rect 470336 340010 470352 340074
rect 470416 340010 470432 340074
rect 470496 340010 470512 340074
rect 470576 340010 470592 340074
rect 470656 340010 470672 340074
rect 470736 340010 470752 340074
rect 470816 340010 470822 340074
rect 470266 340009 470822 340010
rect 541566 339494 541572 339558
rect 541636 339556 541642 339558
rect 541709 339556 541775 339559
rect 541636 339554 541775 339556
rect 541636 339498 541714 339554
rect 541770 339498 541775 339554
rect 541636 339496 541775 339498
rect 541636 339494 541642 339496
rect 541709 339493 541775 339496
rect 544193 339556 544259 339559
rect 544326 339556 544332 339558
rect 544193 339554 544332 339556
rect 544193 339498 544198 339554
rect 544254 339498 544332 339554
rect 544193 339496 544332 339498
rect 544193 339493 544259 339496
rect 544326 339494 544332 339496
rect 544396 339494 544402 339558
rect 583520 338454 584960 338694
rect 535453 336836 535519 336839
rect 535453 336834 538108 336836
rect 535453 336778 535458 336834
rect 535514 336778 538108 336834
rect 535453 336776 538108 336778
rect 535453 336773 535519 336776
rect 486550 335414 486556 335478
rect 486620 335476 486626 335478
rect 486620 335416 538108 335476
rect 486620 335414 486626 335416
rect 485630 334054 485636 334118
rect 485700 334116 485706 334118
rect 485700 334056 538108 334116
rect 485700 334054 485706 334056
rect 486734 332694 486740 332758
rect 486804 332756 486810 332758
rect 486804 332696 538108 332756
rect 486804 332694 486810 332696
rect -960 332198 480 332438
rect 535453 331396 535519 331399
rect 535453 331394 538108 331396
rect 535453 331338 535458 331394
rect 535514 331338 538108 331394
rect 535453 331336 538108 331338
rect 535453 331333 535519 331336
rect 535453 330036 535519 330039
rect 535453 330034 538108 330036
rect 535453 329978 535458 330034
rect 535514 329978 538108 330034
rect 535453 329976 538108 329978
rect 535453 329973 535519 329976
rect 536005 328676 536071 328679
rect 536005 328674 538108 328676
rect 536005 328618 536010 328674
rect 536066 328618 538108 328674
rect 536005 328616 538108 328618
rect 536005 328613 536071 328616
rect 536649 327316 536715 327319
rect 536649 327314 538108 327316
rect 536649 327258 536654 327314
rect 536710 327258 538108 327314
rect 536649 327256 538108 327258
rect 536649 327253 536715 327256
rect 547413 327044 547479 327047
rect 547413 327042 547522 327044
rect 547413 326986 547418 327042
rect 547474 326986 547522 327042
rect 547413 326981 547522 326986
rect 547462 326742 547522 326981
rect 535453 325956 535519 325959
rect 535453 325954 538108 325956
rect 535453 325898 535458 325954
rect 535514 325898 538108 325954
rect 535453 325896 538108 325898
rect 577026 325950 577582 325951
rect 535453 325893 535519 325896
rect 577026 325886 577032 325950
rect 577096 325886 577112 325950
rect 577176 325886 577192 325950
rect 577256 325886 577272 325950
rect 577336 325886 577352 325950
rect 577416 325886 577432 325950
rect 577496 325886 577512 325950
rect 577576 325886 577582 325950
rect 577026 325870 577582 325886
rect 577026 325806 577032 325870
rect 577096 325806 577112 325870
rect 577176 325806 577192 325870
rect 577256 325806 577272 325870
rect 577336 325806 577352 325870
rect 577416 325806 577432 325870
rect 577496 325806 577512 325870
rect 577576 325806 577582 325870
rect 577026 325790 577582 325806
rect 577026 325726 577032 325790
rect 577096 325726 577112 325790
rect 577176 325726 577192 325790
rect 577256 325726 577272 325790
rect 577336 325726 577352 325790
rect 577416 325726 577432 325790
rect 577496 325726 577512 325790
rect 577576 325726 577582 325790
rect 577026 325710 577582 325726
rect 577026 325646 577032 325710
rect 577096 325646 577112 325710
rect 577176 325646 577192 325710
rect 577256 325646 577272 325710
rect 577336 325646 577352 325710
rect 577416 325646 577432 325710
rect 577496 325646 577512 325710
rect 577576 325646 577582 325710
rect 577026 325645 577582 325646
rect 576600 325278 576666 325280
rect 580901 325278 580967 325279
rect 576600 325276 581156 325278
rect 583520 325276 584960 325366
rect 576600 325275 584960 325276
rect 576600 325219 576605 325275
rect 576661 325274 584960 325275
rect 576661 325219 580906 325274
rect 576600 325218 580906 325219
rect 580962 325218 584960 325274
rect 576600 325216 584960 325218
rect 576600 325214 576666 325216
rect 580901 325213 580967 325216
rect 578266 325155 578822 325156
rect 578266 325091 578272 325155
rect 578336 325091 578352 325155
rect 578416 325091 578432 325155
rect 578496 325091 578512 325155
rect 578576 325091 578592 325155
rect 578656 325091 578672 325155
rect 578736 325091 578752 325155
rect 578816 325091 578822 325155
rect 583520 325126 584960 325216
rect 578266 325075 578822 325091
rect 578266 325011 578272 325075
rect 578336 325011 578352 325075
rect 578416 325011 578432 325075
rect 578496 325011 578512 325075
rect 578576 325011 578592 325075
rect 578656 325011 578672 325075
rect 578736 325011 578752 325075
rect 578816 325011 578822 325075
rect 578266 324995 578822 325011
rect 578266 324931 578272 324995
rect 578336 324931 578352 324995
rect 578416 324931 578432 324995
rect 578496 324931 578512 324995
rect 578576 324931 578592 324995
rect 578656 324931 578672 324995
rect 578736 324931 578752 324995
rect 578816 324931 578822 324995
rect 578266 324915 578822 324931
rect 578266 324851 578272 324915
rect 578336 324851 578352 324915
rect 578416 324851 578432 324915
rect 578496 324851 578512 324915
rect 578576 324851 578592 324915
rect 578656 324851 578672 324915
rect 578736 324851 578752 324915
rect 578816 324851 578822 324915
rect 578266 324850 578822 324851
rect 536373 324596 536439 324599
rect 536373 324594 538108 324596
rect 536373 324538 536378 324594
rect 536434 324538 538108 324594
rect 536373 324536 538108 324538
rect 536373 324533 536439 324536
rect 536741 323236 536807 323239
rect 536741 323234 538108 323236
rect 536741 323178 536746 323234
rect 536802 323206 538108 323234
rect 536802 323178 538138 323206
rect 536741 323176 538138 323178
rect 536741 323173 536807 323176
rect 470266 322486 470822 322487
rect 470266 322422 470272 322486
rect 470336 322422 470352 322486
rect 470416 322422 470432 322486
rect 470496 322422 470512 322486
rect 470576 322422 470592 322486
rect 470656 322422 470672 322486
rect 470736 322422 470752 322486
rect 470816 322422 470822 322486
rect 470266 322406 470822 322422
rect 470266 322342 470272 322406
rect 470336 322342 470352 322406
rect 470416 322342 470432 322406
rect 470496 322342 470512 322406
rect 470576 322342 470592 322406
rect 470656 322342 470672 322406
rect 470736 322342 470752 322406
rect 470816 322342 470822 322406
rect 470266 322326 470822 322342
rect 470266 322262 470272 322326
rect 470336 322262 470352 322326
rect 470416 322262 470432 322326
rect 470496 322262 470512 322326
rect 470576 322262 470592 322326
rect 470656 322262 470672 322326
rect 470736 322262 470752 322326
rect 470816 322262 470822 322326
rect 470266 322246 470822 322262
rect 470266 322182 470272 322246
rect 470336 322182 470352 322246
rect 470416 322182 470432 322246
rect 470496 322182 470512 322246
rect 470576 322182 470592 322246
rect 470656 322182 470672 322246
rect 470736 322182 470752 322246
rect 470816 322182 470822 322246
rect 470266 322181 470822 322182
rect 483606 322086 483612 322150
rect 483676 322148 483682 322150
rect 484301 322148 484367 322151
rect 483676 322146 484367 322148
rect 483676 322090 484306 322146
rect 484362 322090 484367 322146
rect 483676 322088 484367 322090
rect 483676 322086 483682 322088
rect 484301 322085 484367 322088
rect 483473 321604 483539 321607
rect 483606 321604 483612 321606
rect 483473 321602 483612 321604
rect 483473 321546 483478 321602
rect 483534 321546 483612 321602
rect 483473 321544 483612 321546
rect 483473 321541 483539 321544
rect 483606 321542 483612 321544
rect 483676 321542 483682 321606
rect 469026 321399 469582 321400
rect 469026 321335 469032 321399
rect 469096 321335 469112 321399
rect 469176 321335 469192 321399
rect 469256 321335 469272 321399
rect 469336 321335 469352 321399
rect 469416 321335 469432 321399
rect 469496 321335 469512 321399
rect 469576 321335 469582 321399
rect 469026 321319 469582 321335
rect 469026 321255 469032 321319
rect 469096 321255 469112 321319
rect 469176 321255 469192 321319
rect 469256 321255 469272 321319
rect 469336 321255 469352 321319
rect 469416 321255 469432 321319
rect 469496 321255 469512 321319
rect 469576 321255 469582 321319
rect 473670 321270 473676 321334
rect 473740 321332 473746 321334
rect 474273 321332 474339 321335
rect 473740 321330 474339 321332
rect 473740 321274 474278 321330
rect 474334 321274 474339 321330
rect 473740 321272 474339 321274
rect 473740 321270 473746 321272
rect 474273 321269 474339 321272
rect 469026 321239 469582 321255
rect 469026 321175 469032 321239
rect 469096 321175 469112 321239
rect 469176 321175 469192 321239
rect 469256 321175 469272 321239
rect 469336 321175 469352 321239
rect 469416 321175 469432 321239
rect 469496 321175 469512 321239
rect 469576 321175 469582 321239
rect 469026 321159 469582 321175
rect 469026 321095 469032 321159
rect 469096 321095 469112 321159
rect 469176 321095 469192 321159
rect 469256 321095 469272 321159
rect 469336 321095 469352 321159
rect 469416 321095 469432 321159
rect 469496 321095 469512 321159
rect 469576 321095 469582 321159
rect 469026 321094 469582 321095
rect 481030 320998 481036 321062
rect 481100 321060 481106 321062
rect 481173 321060 481239 321063
rect 481100 321058 481239 321060
rect 481100 321002 481178 321058
rect 481234 321002 481239 321058
rect 481100 321000 481239 321002
rect 481100 320998 481106 321000
rect 481173 320997 481239 321000
rect 488022 320998 488028 321062
rect 488092 321060 488098 321062
rect 488165 321060 488231 321063
rect 488092 321058 488231 321060
rect 488092 321002 488170 321058
rect 488226 321002 488231 321058
rect 488092 321000 488231 321002
rect 488092 320998 488098 321000
rect 488165 320997 488231 321000
rect 478137 320924 478203 320927
rect 478638 320924 478644 320926
rect 478137 320922 478644 320924
rect 478137 320866 478142 320922
rect 478198 320866 478644 320922
rect 478137 320864 478644 320866
rect 478137 320861 478203 320864
rect 478638 320862 478644 320864
rect 478708 320862 478714 320926
rect 470266 320314 470822 320315
rect 470266 320250 470272 320314
rect 470336 320250 470352 320314
rect 470416 320250 470432 320314
rect 470496 320250 470512 320314
rect 470576 320250 470592 320314
rect 470656 320250 470672 320314
rect 470736 320250 470752 320314
rect 470816 320250 470822 320314
rect 470266 320234 470822 320250
rect 470266 320170 470272 320234
rect 470336 320170 470352 320234
rect 470416 320170 470432 320234
rect 470496 320170 470512 320234
rect 470576 320170 470592 320234
rect 470656 320170 470672 320234
rect 470736 320170 470752 320234
rect 470816 320170 470822 320234
rect 470266 320154 470822 320170
rect 470266 320090 470272 320154
rect 470336 320090 470352 320154
rect 470416 320090 470432 320154
rect 470496 320090 470512 320154
rect 470576 320090 470592 320154
rect 470656 320090 470672 320154
rect 470736 320090 470752 320154
rect 470816 320090 470822 320154
rect 470266 320074 470822 320090
rect 470266 320010 470272 320074
rect 470336 320010 470352 320074
rect 470416 320010 470432 320074
rect 470496 320010 470512 320074
rect 470576 320010 470592 320074
rect 470656 320010 470672 320074
rect 470736 320010 470752 320074
rect 470816 320010 470822 320074
rect 470266 320009 470822 320010
rect -960 319142 480 319382
rect 536741 316436 536807 316439
rect 538078 316436 538138 323176
rect 536741 316434 538138 316436
rect 536741 316378 536746 316434
rect 536802 316406 538138 316434
rect 536802 316378 538108 316406
rect 536741 316376 538108 316378
rect 536741 316373 536807 316376
rect 583520 311934 584960 312174
rect 470266 307086 470822 307087
rect 470266 307022 470272 307086
rect 470336 307022 470352 307086
rect 470416 307022 470432 307086
rect 470496 307022 470512 307086
rect 470576 307022 470592 307086
rect 470656 307022 470672 307086
rect 470736 307022 470752 307086
rect 470816 307022 470822 307086
rect 470266 307006 470822 307022
rect 470266 306942 470272 307006
rect 470336 306942 470352 307006
rect 470416 306942 470432 307006
rect 470496 306942 470512 307006
rect 470576 306942 470592 307006
rect 470656 306942 470672 307006
rect 470736 306942 470752 307006
rect 470816 306942 470822 307006
rect 470266 306926 470822 306942
rect 470266 306862 470272 306926
rect 470336 306862 470352 306926
rect 470416 306862 470432 306926
rect 470496 306862 470512 306926
rect 470576 306862 470592 306926
rect 470656 306862 470672 306926
rect 470736 306862 470752 306926
rect 470816 306862 470822 306926
rect 470266 306846 470822 306862
rect 470266 306782 470272 306846
rect 470336 306782 470352 306846
rect 470416 306782 470432 306846
rect 470496 306782 470512 306846
rect 470576 306782 470592 306846
rect 470656 306782 470672 306846
rect 470736 306782 470752 306846
rect 470816 306782 470822 306846
rect 470266 306781 470822 306782
rect 480897 306510 480963 306511
rect 480846 306446 480852 306510
rect 480916 306508 480963 306510
rect 480916 306506 481008 306508
rect 480958 306450 481008 306506
rect 480916 306448 481008 306450
rect 480916 306446 480963 306448
rect 480897 306445 480963 306446
rect -960 306086 480 306326
rect 487654 306310 487660 306374
rect 487724 306310 487730 306374
rect 487529 306236 487595 306239
rect 487662 306236 487722 306310
rect 487529 306234 487722 306236
rect 487529 306178 487534 306234
rect 487590 306178 487722 306234
rect 487529 306176 487722 306178
rect 487529 306173 487595 306176
rect 469026 306001 469582 306002
rect 469026 305937 469032 306001
rect 469096 305937 469112 306001
rect 469176 305937 469192 306001
rect 469256 305937 469272 306001
rect 469336 305937 469352 306001
rect 469416 305937 469432 306001
rect 469496 305937 469512 306001
rect 469576 305937 469582 306001
rect 473721 305966 473787 305967
rect 469026 305921 469582 305937
rect 469026 305857 469032 305921
rect 469096 305857 469112 305921
rect 469176 305857 469192 305921
rect 469256 305857 469272 305921
rect 469336 305857 469352 305921
rect 469416 305857 469432 305921
rect 469496 305857 469512 305921
rect 469576 305857 469582 305921
rect 473670 305902 473676 305966
rect 473740 305964 473787 305966
rect 473740 305962 473832 305964
rect 473782 305906 473832 305962
rect 473740 305904 473832 305906
rect 473740 305902 473787 305904
rect 473721 305901 473787 305902
rect 469026 305841 469582 305857
rect 469026 305777 469032 305841
rect 469096 305777 469112 305841
rect 469176 305777 469192 305841
rect 469256 305777 469272 305841
rect 469336 305777 469352 305841
rect 469416 305777 469432 305841
rect 469496 305777 469512 305841
rect 469576 305777 469582 305841
rect 469026 305761 469582 305777
rect 469026 305697 469032 305761
rect 469096 305697 469112 305761
rect 469176 305697 469192 305761
rect 469256 305697 469272 305761
rect 469336 305697 469352 305761
rect 469416 305697 469432 305761
rect 469496 305697 469512 305761
rect 469576 305697 469582 305761
rect 469026 305696 469582 305697
rect 477734 305692 477800 305695
rect 478822 305692 478828 305694
rect 477734 305690 478828 305692
rect 477734 305634 477739 305690
rect 477795 305634 478828 305690
rect 477734 305632 478828 305634
rect 477734 305629 477800 305632
rect 478822 305630 478828 305632
rect 478892 305630 478898 305694
rect 484117 305558 484183 305559
rect 484117 305556 484164 305558
rect 484072 305554 484164 305556
rect 484072 305498 484122 305554
rect 484072 305496 484164 305498
rect 484117 305494 484164 305496
rect 484228 305494 484234 305558
rect 484117 305493 484183 305494
rect 470266 304914 470822 304915
rect 470266 304850 470272 304914
rect 470336 304850 470352 304914
rect 470416 304850 470432 304914
rect 470496 304850 470512 304914
rect 470576 304850 470592 304914
rect 470656 304850 470672 304914
rect 470736 304850 470752 304914
rect 470816 304850 470822 304914
rect 470266 304834 470822 304850
rect 470266 304770 470272 304834
rect 470336 304770 470352 304834
rect 470416 304770 470432 304834
rect 470496 304770 470512 304834
rect 470576 304770 470592 304834
rect 470656 304770 470672 304834
rect 470736 304770 470752 304834
rect 470816 304770 470822 304834
rect 470266 304754 470822 304770
rect 470266 304690 470272 304754
rect 470336 304690 470352 304754
rect 470416 304690 470432 304754
rect 470496 304690 470512 304754
rect 470576 304690 470592 304754
rect 470656 304690 470672 304754
rect 470736 304690 470752 304754
rect 470816 304690 470822 304754
rect 470266 304674 470822 304690
rect 470266 304610 470272 304674
rect 470336 304610 470352 304674
rect 470416 304610 470432 304674
rect 470496 304610 470512 304674
rect 470576 304610 470592 304674
rect 470656 304610 470672 304674
rect 470736 304610 470752 304674
rect 470816 304610 470822 304674
rect 470266 304609 470822 304610
rect 541566 303726 541572 303790
rect 541636 303788 541642 303790
rect 541709 303788 541775 303791
rect 541636 303786 541775 303788
rect 541636 303730 541714 303786
rect 541770 303730 541775 303786
rect 541636 303728 541775 303730
rect 541636 303726 541642 303728
rect 541709 303725 541775 303728
rect 544193 303788 544259 303791
rect 544326 303788 544332 303790
rect 544193 303786 544332 303788
rect 544193 303730 544198 303786
rect 544254 303730 544332 303786
rect 544193 303728 544332 303730
rect 544193 303725 544259 303728
rect 544326 303726 544332 303728
rect 544396 303726 544402 303790
rect 480846 302230 480852 302294
rect 480916 302292 480922 302294
rect 482277 302292 482343 302295
rect 580165 302292 580231 302295
rect 480916 302290 580231 302292
rect 480916 302234 482282 302290
rect 482338 302234 580170 302290
rect 580226 302234 580231 302290
rect 480916 302232 580231 302234
rect 480916 302230 480922 302232
rect 482277 302229 482343 302232
rect 580165 302229 580231 302232
rect 535453 300796 535519 300799
rect 535453 300794 538108 300796
rect 535453 300738 535458 300794
rect 535514 300738 538108 300794
rect 535453 300736 538108 300738
rect 535453 300733 535519 300736
rect 535453 299436 535519 299439
rect 535453 299434 538108 299436
rect 535453 299378 535458 299434
rect 535514 299378 538108 299434
rect 535453 299376 538108 299378
rect 535453 299373 535519 299376
rect 580165 298756 580231 298759
rect 583520 298756 584960 298846
rect 580165 298754 584960 298756
rect 580165 298698 580170 298754
rect 580226 298698 584960 298754
rect 580165 298696 584960 298698
rect 580165 298693 580231 298696
rect 583520 298606 584960 298696
rect 535453 298076 535519 298079
rect 535453 298074 538108 298076
rect 535453 298018 535458 298074
rect 535514 298018 538108 298074
rect 535453 298016 538108 298018
rect 535453 298013 535519 298016
rect 535453 296716 535519 296719
rect 535453 296714 538108 296716
rect 535453 296658 535458 296714
rect 535514 296658 538108 296714
rect 535453 296656 538108 296658
rect 535453 296653 535519 296656
rect 535545 295356 535611 295359
rect 535545 295354 538108 295356
rect 535545 295298 535550 295354
rect 535606 295298 538108 295354
rect 535545 295296 538108 295298
rect 535545 295293 535611 295296
rect 535453 293996 535519 293999
rect 535453 293994 538108 293996
rect 535453 293938 535458 293994
rect 535514 293938 538108 293994
rect 535453 293936 538108 293938
rect 535453 293933 535519 293936
rect -960 293030 480 293270
rect 535545 292636 535611 292639
rect 535545 292634 538108 292636
rect 535545 292578 535550 292634
rect 535606 292578 538108 292634
rect 535545 292576 538108 292578
rect 535545 292573 535611 292576
rect 535453 291276 535519 291279
rect 535453 291274 538108 291276
rect 535453 291218 535458 291274
rect 535514 291218 538108 291274
rect 535453 291216 538108 291218
rect 535453 291213 535519 291216
rect 547321 291140 547387 291143
rect 547278 291138 547387 291140
rect 547278 291082 547326 291138
rect 547382 291082 547387 291138
rect 547278 291077 547387 291082
rect 547278 290702 547338 291077
rect 535453 289916 535519 289919
rect 535453 289914 538108 289916
rect 535453 289858 535458 289914
rect 535514 289858 538108 289914
rect 535453 289856 538108 289858
rect 535453 289853 535519 289856
rect 473670 289718 473676 289782
rect 473740 289780 473746 289782
rect 476062 289780 476068 289782
rect 473740 289720 476068 289780
rect 473740 289718 473746 289720
rect 476062 289718 476068 289720
rect 476132 289718 476138 289782
rect 535453 288556 535519 288559
rect 535453 288554 538108 288556
rect 535453 288498 535458 288554
rect 535514 288498 538108 288554
rect 535453 288496 538108 288498
rect 535453 288493 535519 288496
rect 482134 288358 482140 288422
rect 482204 288420 482210 288422
rect 482277 288420 482343 288423
rect 482204 288418 482343 288420
rect 482204 288362 482282 288418
rect 482338 288362 482343 288418
rect 482204 288360 482343 288362
rect 482204 288358 482210 288360
rect 482277 288357 482343 288360
rect 470266 287487 470822 287488
rect 470266 287423 470272 287487
rect 470336 287423 470352 287487
rect 470416 287423 470432 287487
rect 470496 287423 470512 287487
rect 470576 287423 470592 287487
rect 470656 287423 470672 287487
rect 470736 287423 470752 287487
rect 470816 287423 470822 287487
rect 470266 287407 470822 287423
rect 470266 287343 470272 287407
rect 470336 287343 470352 287407
rect 470416 287343 470432 287407
rect 470496 287343 470512 287407
rect 470576 287343 470592 287407
rect 470656 287343 470672 287407
rect 470736 287343 470752 287407
rect 470816 287343 470822 287407
rect 470266 287327 470822 287343
rect 470266 287263 470272 287327
rect 470336 287263 470352 287327
rect 470416 287263 470432 287327
rect 470496 287263 470512 287327
rect 470576 287263 470592 287327
rect 470656 287263 470672 287327
rect 470736 287263 470752 287327
rect 470816 287263 470822 287327
rect 470266 287247 470822 287263
rect 470266 287183 470272 287247
rect 470336 287183 470352 287247
rect 470416 287183 470432 287247
rect 470496 287183 470512 287247
rect 470576 287183 470592 287247
rect 470656 287183 470672 287247
rect 470736 287183 470752 287247
rect 470816 287183 470822 287247
rect 470266 287182 470822 287183
rect 536741 287196 536807 287199
rect 536741 287194 538108 287196
rect 536741 287138 536746 287194
rect 536802 287166 538108 287194
rect 536802 287138 538138 287166
rect 536741 287136 538138 287138
rect 536741 287133 536807 287136
rect 478628 286924 478694 286927
rect 478822 286924 478828 286926
rect 478628 286922 478828 286924
rect 478628 286866 478633 286922
rect 478689 286866 478828 286922
rect 478628 286864 478828 286866
rect 478628 286861 478694 286864
rect 478822 286862 478828 286864
rect 478892 286862 478898 286926
rect 488390 286726 488396 286790
rect 488460 286726 488466 286790
rect 474916 286652 474982 286655
rect 476062 286652 476068 286654
rect 474916 286650 476068 286652
rect 474916 286594 474921 286650
rect 474977 286594 476068 286650
rect 474916 286592 476068 286594
rect 474916 286589 474982 286592
rect 476062 286590 476068 286592
rect 476132 286590 476138 286654
rect 484158 286590 484164 286654
rect 484228 286652 484234 286654
rect 484761 286652 484827 286655
rect 484228 286650 484827 286652
rect 484228 286594 484766 286650
rect 484822 286594 484827 286650
rect 484228 286592 484827 286594
rect 488398 286652 488458 286726
rect 488533 286652 488599 286655
rect 488398 286650 488599 286652
rect 488398 286594 488538 286650
rect 488594 286594 488599 286650
rect 488398 286592 488599 286594
rect 484228 286590 484234 286592
rect 484761 286589 484827 286592
rect 488533 286589 488599 286592
rect 469026 286402 469582 286403
rect 469026 286338 469032 286402
rect 469096 286338 469112 286402
rect 469176 286338 469192 286402
rect 469256 286338 469272 286402
rect 469336 286338 469352 286402
rect 469416 286338 469432 286402
rect 469496 286338 469512 286402
rect 469576 286338 469582 286402
rect 469026 286322 469582 286338
rect 469026 286258 469032 286322
rect 469096 286258 469112 286322
rect 469176 286258 469192 286322
rect 469256 286258 469272 286322
rect 469336 286258 469352 286322
rect 469416 286258 469432 286322
rect 469496 286258 469512 286322
rect 469576 286258 469582 286322
rect 469026 286242 469582 286258
rect 469026 286178 469032 286242
rect 469096 286178 469112 286242
rect 469176 286178 469192 286242
rect 469256 286178 469272 286242
rect 469336 286178 469352 286242
rect 469416 286178 469432 286242
rect 469496 286178 469512 286242
rect 469576 286178 469582 286242
rect 469026 286162 469582 286178
rect 469026 286098 469032 286162
rect 469096 286098 469112 286162
rect 469176 286098 469192 286162
rect 469256 286098 469272 286162
rect 469336 286098 469352 286162
rect 469416 286098 469432 286162
rect 469496 286098 469512 286162
rect 469576 286098 469582 286162
rect 469026 286097 469582 286098
rect 482185 285702 482251 285703
rect 482134 285638 482140 285702
rect 482204 285700 482251 285702
rect 482204 285698 482296 285700
rect 482246 285642 482296 285698
rect 482204 285640 482296 285642
rect 482204 285638 482251 285640
rect 482185 285637 482251 285638
rect 470266 285314 470822 285315
rect 470266 285250 470272 285314
rect 470336 285250 470352 285314
rect 470416 285250 470432 285314
rect 470496 285250 470512 285314
rect 470576 285250 470592 285314
rect 470656 285250 470672 285314
rect 470736 285250 470752 285314
rect 470816 285250 470822 285314
rect 470266 285234 470822 285250
rect 470266 285170 470272 285234
rect 470336 285170 470352 285234
rect 470416 285170 470432 285234
rect 470496 285170 470512 285234
rect 470576 285170 470592 285234
rect 470656 285170 470672 285234
rect 470736 285170 470752 285234
rect 470816 285170 470822 285234
rect 470266 285154 470822 285170
rect 470266 285090 470272 285154
rect 470336 285090 470352 285154
rect 470416 285090 470432 285154
rect 470496 285090 470512 285154
rect 470576 285090 470592 285154
rect 470656 285090 470672 285154
rect 470736 285090 470752 285154
rect 470816 285090 470822 285154
rect 470266 285074 470822 285090
rect 470266 285010 470272 285074
rect 470336 285010 470352 285074
rect 470416 285010 470432 285074
rect 470496 285010 470512 285074
rect 470576 285010 470592 285074
rect 470656 285010 470672 285074
rect 470736 285010 470752 285074
rect 470816 285010 470822 285074
rect 470266 285009 470822 285010
rect 538078 280366 538138 287136
rect 583520 285278 584960 285518
rect -960 279974 480 280214
rect 482134 273262 482140 273326
rect 482204 273324 482210 273326
rect 482369 273324 482435 273327
rect 482204 273322 482435 273324
rect 482204 273266 482374 273322
rect 482430 273266 482435 273322
rect 482204 273264 482435 273266
rect 482204 273262 482210 273264
rect 482369 273261 482435 273264
rect 577026 272910 577582 272911
rect 577026 272846 577032 272910
rect 577096 272846 577112 272910
rect 577176 272846 577192 272910
rect 577256 272846 577272 272910
rect 577336 272846 577352 272910
rect 577416 272846 577432 272910
rect 577496 272846 577512 272910
rect 577576 272846 577582 272910
rect 577026 272830 577582 272846
rect 577026 272766 577032 272830
rect 577096 272766 577112 272830
rect 577176 272766 577192 272830
rect 577256 272766 577272 272830
rect 577336 272766 577352 272830
rect 577416 272766 577432 272830
rect 577496 272766 577512 272830
rect 577576 272766 577582 272830
rect 577026 272750 577582 272766
rect 577026 272686 577032 272750
rect 577096 272686 577112 272750
rect 577176 272686 577192 272750
rect 577256 272686 577272 272750
rect 577336 272686 577352 272750
rect 577416 272686 577432 272750
rect 577496 272686 577512 272750
rect 577576 272686 577582 272750
rect 577026 272670 577582 272686
rect 484158 272582 484164 272646
rect 484228 272644 484234 272646
rect 485497 272644 485563 272647
rect 484228 272642 485563 272644
rect 484228 272586 485502 272642
rect 485558 272586 485563 272642
rect 577026 272606 577032 272670
rect 577096 272606 577112 272670
rect 577176 272606 577192 272670
rect 577256 272606 577272 272670
rect 577336 272606 577352 272670
rect 577416 272606 577432 272670
rect 577496 272606 577512 272670
rect 577576 272606 577582 272670
rect 577026 272605 577582 272606
rect 484228 272584 485563 272586
rect 484228 272582 484234 272584
rect 485497 272581 485563 272584
rect 576600 272238 576666 272240
rect 580901 272238 580967 272239
rect 576600 272236 581040 272238
rect 583520 272236 584960 272326
rect 576600 272235 584960 272236
rect 576600 272179 576605 272235
rect 576661 272234 584960 272235
rect 576661 272179 580906 272234
rect 576600 272178 580906 272179
rect 580962 272178 584960 272234
rect 576600 272176 584960 272178
rect 576600 272174 576666 272176
rect 580901 272173 580967 272176
rect 578266 272115 578822 272116
rect 578266 272051 578272 272115
rect 578336 272051 578352 272115
rect 578416 272051 578432 272115
rect 578496 272051 578512 272115
rect 578576 272051 578592 272115
rect 578656 272051 578672 272115
rect 578736 272051 578752 272115
rect 578816 272051 578822 272115
rect 583520 272086 584960 272176
rect 578266 272035 578822 272051
rect 578266 271971 578272 272035
rect 578336 271971 578352 272035
rect 578416 271971 578432 272035
rect 578496 271971 578512 272035
rect 578576 271971 578592 272035
rect 578656 271971 578672 272035
rect 578736 271971 578752 272035
rect 578816 271971 578822 272035
rect 578266 271955 578822 271971
rect 578266 271891 578272 271955
rect 578336 271891 578352 271955
rect 578416 271891 578432 271955
rect 578496 271891 578512 271955
rect 578576 271891 578592 271955
rect 578656 271891 578672 271955
rect 578736 271891 578752 271955
rect 578816 271891 578822 271955
rect 578266 271875 578822 271891
rect 578266 271811 578272 271875
rect 578336 271811 578352 271875
rect 578416 271811 578432 271875
rect 578496 271811 578512 271875
rect 578576 271811 578592 271875
rect 578656 271811 578672 271875
rect 578736 271811 578752 271875
rect 578816 271811 578822 271875
rect 578266 271810 578822 271811
rect 470266 267487 470822 267488
rect 470266 267423 470272 267487
rect 470336 267423 470352 267487
rect 470416 267423 470432 267487
rect 470496 267423 470512 267487
rect 470576 267423 470592 267487
rect 470656 267423 470672 267487
rect 470736 267423 470752 267487
rect 470816 267423 470822 267487
rect 470266 267407 470822 267423
rect 470266 267343 470272 267407
rect 470336 267343 470352 267407
rect 470416 267343 470432 267407
rect 470496 267343 470512 267407
rect 470576 267343 470592 267407
rect 470656 267343 470672 267407
rect 470736 267343 470752 267407
rect 470816 267343 470822 267407
rect 470266 267327 470822 267343
rect 482369 267340 482435 267343
rect 485497 267340 485563 267343
rect -960 267054 480 267294
rect 470266 267263 470272 267327
rect 470336 267263 470352 267327
rect 470416 267263 470432 267327
rect 470496 267263 470512 267327
rect 470576 267263 470592 267327
rect 470656 267263 470672 267327
rect 470736 267263 470752 267327
rect 470816 267263 470822 267327
rect 470266 267247 470822 267263
rect 470266 267183 470272 267247
rect 470336 267183 470352 267247
rect 470416 267183 470432 267247
rect 470496 267183 470512 267247
rect 470576 267183 470592 267247
rect 470656 267183 470672 267247
rect 470736 267183 470752 267247
rect 470816 267183 470822 267247
rect 470266 267182 470822 267183
rect 482326 267338 482435 267340
rect 482326 267282 482374 267338
rect 482430 267282 482435 267338
rect 482326 267277 482435 267282
rect 485454 267338 485563 267340
rect 485454 267282 485502 267338
rect 485558 267282 485563 267338
rect 485454 267277 485563 267282
rect 482326 267071 482386 267277
rect 485454 267071 485514 267277
rect 482326 267066 482435 267071
rect 482326 267010 482374 267066
rect 482430 267010 482435 267066
rect 482326 267008 482435 267010
rect 482369 267005 482435 267008
rect 485405 267066 485514 267071
rect 488441 267070 488507 267071
rect 488390 267068 488396 267070
rect 485405 267010 485410 267066
rect 485466 267010 485514 267066
rect 485405 267008 485514 267010
rect 488350 267008 488396 267068
rect 488460 267066 488507 267070
rect 488502 267010 488507 267066
rect 485405 267005 485471 267008
rect 488390 267006 488396 267008
rect 488460 267006 488507 267010
rect 488441 267005 488507 267006
rect 469026 266401 469582 266402
rect 469026 266337 469032 266401
rect 469096 266337 469112 266401
rect 469176 266337 469192 266401
rect 469256 266337 469272 266401
rect 469336 266337 469352 266401
rect 469416 266337 469432 266401
rect 469496 266337 469512 266401
rect 469576 266337 469582 266401
rect 469026 266321 469582 266337
rect 469026 266257 469032 266321
rect 469096 266257 469112 266321
rect 469176 266257 469192 266321
rect 469256 266257 469272 266321
rect 469336 266257 469352 266321
rect 469416 266257 469432 266321
rect 469496 266257 469512 266321
rect 469576 266257 469582 266321
rect 469026 266241 469582 266257
rect 469026 266177 469032 266241
rect 469096 266177 469112 266241
rect 469176 266177 469192 266241
rect 469256 266177 469272 266241
rect 469336 266177 469352 266241
rect 469416 266177 469432 266241
rect 469496 266177 469512 266241
rect 469576 266177 469582 266241
rect 469026 266161 469582 266177
rect 469026 266097 469032 266161
rect 469096 266097 469112 266161
rect 469176 266097 469192 266161
rect 469256 266097 469272 266161
rect 469336 266097 469352 266161
rect 469416 266097 469432 266161
rect 469496 266097 469512 266161
rect 469576 266097 469582 266161
rect 469026 266096 469582 266097
rect 479057 265982 479123 265983
rect 479006 265980 479012 265982
rect 478966 265920 479012 265980
rect 479076 265978 479123 265982
rect 479118 265922 479123 265978
rect 479006 265918 479012 265920
rect 479076 265918 479123 265922
rect 479057 265917 479123 265918
rect 470266 265314 470822 265315
rect 470266 265250 470272 265314
rect 470336 265250 470352 265314
rect 470416 265250 470432 265314
rect 470496 265250 470512 265314
rect 470576 265250 470592 265314
rect 470656 265250 470672 265314
rect 470736 265250 470752 265314
rect 470816 265250 470822 265314
rect 470266 265234 470822 265250
rect 470266 265170 470272 265234
rect 470336 265170 470352 265234
rect 470416 265170 470432 265234
rect 470496 265170 470512 265234
rect 470576 265170 470592 265234
rect 470656 265170 470672 265234
rect 470736 265170 470752 265234
rect 470816 265170 470822 265234
rect 470266 265154 470822 265170
rect 470266 265090 470272 265154
rect 470336 265090 470352 265154
rect 470416 265090 470432 265154
rect 470496 265090 470512 265154
rect 470576 265090 470592 265154
rect 470656 265090 470672 265154
rect 470736 265090 470752 265154
rect 470816 265090 470822 265154
rect 470266 265074 470822 265090
rect 470266 265010 470272 265074
rect 470336 265010 470352 265074
rect 470416 265010 470432 265074
rect 470496 265010 470512 265074
rect 470576 265010 470592 265074
rect 470656 265010 470672 265074
rect 470736 265010 470752 265074
rect 470816 265010 470822 265074
rect 476481 265030 476547 265031
rect 476430 265028 476436 265030
rect 470266 265009 470822 265010
rect 476354 264968 476436 265028
rect 476500 265028 476547 265030
rect 477350 265028 477356 265030
rect 476500 265026 477356 265028
rect 476542 264970 477356 265026
rect 476430 264966 476436 264968
rect 476500 264968 477356 264970
rect 476500 264966 476547 264968
rect 477350 264966 477356 264968
rect 477420 264966 477426 265030
rect 479517 265028 479583 265031
rect 480110 265028 480116 265030
rect 479517 265026 480116 265028
rect 479517 264970 479522 265026
rect 479578 264970 480116 265026
rect 479517 264968 480116 264970
rect 476481 264965 476547 264966
rect 479517 264965 479583 264968
rect 480110 264966 480116 264968
rect 480180 264966 480186 265030
rect 583520 258758 584960 258998
rect -960 253998 480 254238
rect 480110 245518 480116 245582
rect 480180 245580 480186 245582
rect 583520 245580 584960 245670
rect 480180 245520 584960 245580
rect 480180 245518 480186 245520
rect 583520 245430 584960 245520
rect -960 240942 480 241182
rect 577026 233063 577582 233064
rect 577026 232999 577032 233063
rect 577096 232999 577112 233063
rect 577176 232999 577192 233063
rect 577256 232999 577272 233063
rect 577336 232999 577352 233063
rect 577416 232999 577432 233063
rect 577496 232999 577512 233063
rect 577576 232999 577582 233063
rect 577026 232983 577582 232999
rect 577026 232919 577032 232983
rect 577096 232919 577112 232983
rect 577176 232919 577192 232983
rect 577256 232919 577272 232983
rect 577336 232919 577352 232983
rect 577416 232919 577432 232983
rect 577496 232919 577512 232983
rect 577576 232919 577582 232983
rect 577026 232903 577582 232919
rect 577026 232839 577032 232903
rect 577096 232839 577112 232903
rect 577176 232839 577192 232903
rect 577256 232839 577272 232903
rect 577336 232839 577352 232903
rect 577416 232839 577432 232903
rect 577496 232839 577512 232903
rect 577576 232839 577582 232903
rect 577026 232823 577582 232839
rect 577026 232759 577032 232823
rect 577096 232759 577112 232823
rect 577176 232759 577192 232823
rect 577256 232759 577272 232823
rect 577336 232759 577352 232823
rect 577416 232759 577432 232823
rect 577496 232759 577512 232823
rect 577576 232759 577582 232823
rect 577026 232758 577582 232759
rect 576600 232391 576666 232393
rect 576600 232388 582156 232391
rect 583520 232388 584960 232478
rect 576600 232332 576605 232388
rect 576661 232386 584960 232388
rect 576661 232332 580906 232386
rect 576600 232330 580906 232332
rect 580962 232330 584960 232386
rect 576600 232329 584960 232330
rect 576600 232327 576666 232329
rect 580901 232328 584960 232329
rect 580901 232325 580967 232328
rect 578266 232268 578822 232269
rect 578266 232204 578272 232268
rect 578336 232204 578352 232268
rect 578416 232204 578432 232268
rect 578496 232204 578512 232268
rect 578576 232204 578592 232268
rect 578656 232204 578672 232268
rect 578736 232204 578752 232268
rect 578816 232204 578822 232268
rect 583520 232238 584960 232328
rect 578266 232188 578822 232204
rect 578266 232124 578272 232188
rect 578336 232124 578352 232188
rect 578416 232124 578432 232188
rect 578496 232124 578512 232188
rect 578576 232124 578592 232188
rect 578656 232124 578672 232188
rect 578736 232124 578752 232188
rect 578816 232124 578822 232188
rect 578266 232108 578822 232124
rect 578266 232044 578272 232108
rect 578336 232044 578352 232108
rect 578416 232044 578432 232108
rect 578496 232044 578512 232108
rect 578576 232044 578592 232108
rect 578656 232044 578672 232108
rect 578736 232044 578752 232108
rect 578816 232044 578822 232108
rect 578266 232028 578822 232044
rect 578266 231964 578272 232028
rect 578336 231964 578352 232028
rect 578416 231964 578432 232028
rect 578496 231964 578512 232028
rect 578576 231964 578592 232028
rect 578656 231964 578672 232028
rect 578736 231964 578752 232028
rect 578816 231964 578822 232028
rect 578266 231963 578822 231964
rect -960 227886 480 228126
rect 583520 218910 584960 219150
rect -960 214830 480 215070
rect 477350 205670 477356 205734
rect 477420 205732 477426 205734
rect 583520 205732 584960 205822
rect 477420 205672 584960 205732
rect 477420 205670 477426 205672
rect 583520 205582 584960 205672
rect -960 201774 480 202014
rect 583520 192390 584960 192630
rect -960 188718 480 188958
rect 583520 179062 584960 179302
rect -960 175798 480 176038
rect 583520 165734 584960 165974
rect -960 162742 480 162982
rect 583520 152542 584960 152782
rect -960 149686 480 149926
rect 583520 139214 584960 139454
rect -960 136630 480 136870
rect 583520 125886 584960 126126
rect -960 123574 480 123814
rect 583520 112694 584960 112934
rect -960 110518 480 110758
rect 583520 99366 584960 99606
rect -960 97462 480 97702
rect 583520 86038 584960 86278
rect -960 84542 480 84782
rect 583520 72846 584960 73086
rect -960 71486 480 71726
rect 583520 59518 584960 59758
rect -960 58430 480 58670
rect 583520 46190 584960 46430
rect -960 45374 480 45614
rect 583520 32998 584960 33238
rect -960 32318 480 32558
rect 583520 19670 584960 19910
rect -960 19262 480 19502
rect -960 6342 480 6582
rect 583520 6478 584960 6718
<< via3 >>
rect 254272 703332 254336 703336
rect 254272 703276 254276 703332
rect 254276 703276 254332 703332
rect 254332 703276 254336 703332
rect 254272 703272 254336 703276
rect 254352 703332 254416 703336
rect 254352 703276 254356 703332
rect 254356 703276 254412 703332
rect 254412 703276 254416 703332
rect 254352 703272 254416 703276
rect 254432 703332 254496 703336
rect 254432 703276 254436 703332
rect 254436 703276 254492 703332
rect 254492 703276 254496 703332
rect 254432 703272 254496 703276
rect 254512 703332 254576 703336
rect 254512 703276 254516 703332
rect 254516 703276 254572 703332
rect 254572 703276 254576 703332
rect 254512 703272 254576 703276
rect 254592 703332 254656 703336
rect 254592 703276 254596 703332
rect 254596 703276 254652 703332
rect 254652 703276 254656 703332
rect 254592 703272 254656 703276
rect 254672 703332 254736 703336
rect 254672 703276 254676 703332
rect 254676 703276 254732 703332
rect 254732 703276 254736 703332
rect 254672 703272 254736 703276
rect 254752 703332 254816 703336
rect 254752 703276 254756 703332
rect 254756 703276 254812 703332
rect 254812 703276 254816 703332
rect 254752 703272 254816 703276
rect 254272 703252 254336 703256
rect 254272 703196 254276 703252
rect 254276 703196 254332 703252
rect 254332 703196 254336 703252
rect 254272 703192 254336 703196
rect 254352 703252 254416 703256
rect 254352 703196 254356 703252
rect 254356 703196 254412 703252
rect 254412 703196 254416 703252
rect 254352 703192 254416 703196
rect 254432 703252 254496 703256
rect 254432 703196 254436 703252
rect 254436 703196 254492 703252
rect 254492 703196 254496 703252
rect 254432 703192 254496 703196
rect 254512 703252 254576 703256
rect 254512 703196 254516 703252
rect 254516 703196 254572 703252
rect 254572 703196 254576 703252
rect 254512 703192 254576 703196
rect 254592 703252 254656 703256
rect 254592 703196 254596 703252
rect 254596 703196 254652 703252
rect 254652 703196 254656 703252
rect 254592 703192 254656 703196
rect 254672 703252 254736 703256
rect 254672 703196 254676 703252
rect 254676 703196 254732 703252
rect 254732 703196 254736 703252
rect 254672 703192 254736 703196
rect 254752 703252 254816 703256
rect 254752 703196 254756 703252
rect 254756 703196 254812 703252
rect 254812 703196 254816 703252
rect 254752 703192 254816 703196
rect 254272 703172 254336 703176
rect 254272 703116 254276 703172
rect 254276 703116 254332 703172
rect 254332 703116 254336 703172
rect 254272 703112 254336 703116
rect 254352 703172 254416 703176
rect 254352 703116 254356 703172
rect 254356 703116 254412 703172
rect 254412 703116 254416 703172
rect 254352 703112 254416 703116
rect 254432 703172 254496 703176
rect 254432 703116 254436 703172
rect 254436 703116 254492 703172
rect 254492 703116 254496 703172
rect 254432 703112 254496 703116
rect 254512 703172 254576 703176
rect 254512 703116 254516 703172
rect 254516 703116 254572 703172
rect 254572 703116 254576 703172
rect 254512 703112 254576 703116
rect 254592 703172 254656 703176
rect 254592 703116 254596 703172
rect 254596 703116 254652 703172
rect 254652 703116 254656 703172
rect 254592 703112 254656 703116
rect 254672 703172 254736 703176
rect 254672 703116 254676 703172
rect 254676 703116 254732 703172
rect 254732 703116 254736 703172
rect 254672 703112 254736 703116
rect 254752 703172 254816 703176
rect 254752 703116 254756 703172
rect 254756 703116 254812 703172
rect 254812 703116 254816 703172
rect 254752 703112 254816 703116
rect 254272 703092 254336 703096
rect 254272 703036 254276 703092
rect 254276 703036 254332 703092
rect 254332 703036 254336 703092
rect 254272 703032 254336 703036
rect 254352 703092 254416 703096
rect 254352 703036 254356 703092
rect 254356 703036 254412 703092
rect 254412 703036 254416 703092
rect 254352 703032 254416 703036
rect 254432 703092 254496 703096
rect 254432 703036 254436 703092
rect 254436 703036 254492 703092
rect 254492 703036 254496 703092
rect 254432 703032 254496 703036
rect 254512 703092 254576 703096
rect 254512 703036 254516 703092
rect 254516 703036 254572 703092
rect 254572 703036 254576 703092
rect 254512 703032 254576 703036
rect 254592 703092 254656 703096
rect 254592 703036 254596 703092
rect 254596 703036 254652 703092
rect 254652 703036 254656 703092
rect 254592 703032 254656 703036
rect 254672 703092 254736 703096
rect 254672 703036 254676 703092
rect 254676 703036 254732 703092
rect 254732 703036 254736 703092
rect 254672 703032 254736 703036
rect 254752 703092 254816 703096
rect 254752 703036 254756 703092
rect 254756 703036 254812 703092
rect 254812 703036 254816 703092
rect 254752 703032 254816 703036
rect 326272 703372 326336 703376
rect 326272 703316 326276 703372
rect 326276 703316 326332 703372
rect 326332 703316 326336 703372
rect 326272 703312 326336 703316
rect 326352 703372 326416 703376
rect 326352 703316 326356 703372
rect 326356 703316 326412 703372
rect 326412 703316 326416 703372
rect 326352 703312 326416 703316
rect 326432 703372 326496 703376
rect 326432 703316 326436 703372
rect 326436 703316 326492 703372
rect 326492 703316 326496 703372
rect 326432 703312 326496 703316
rect 326512 703372 326576 703376
rect 326512 703316 326516 703372
rect 326516 703316 326572 703372
rect 326572 703316 326576 703372
rect 326512 703312 326576 703316
rect 326592 703372 326656 703376
rect 326592 703316 326596 703372
rect 326596 703316 326652 703372
rect 326652 703316 326656 703372
rect 326592 703312 326656 703316
rect 326672 703372 326736 703376
rect 326672 703316 326676 703372
rect 326676 703316 326732 703372
rect 326732 703316 326736 703372
rect 326672 703312 326736 703316
rect 326752 703372 326816 703376
rect 326752 703316 326756 703372
rect 326756 703316 326812 703372
rect 326812 703316 326816 703372
rect 326752 703312 326816 703316
rect 326272 703292 326336 703296
rect 326272 703236 326276 703292
rect 326276 703236 326332 703292
rect 326332 703236 326336 703292
rect 326272 703232 326336 703236
rect 326352 703292 326416 703296
rect 326352 703236 326356 703292
rect 326356 703236 326412 703292
rect 326412 703236 326416 703292
rect 326352 703232 326416 703236
rect 326432 703292 326496 703296
rect 326432 703236 326436 703292
rect 326436 703236 326492 703292
rect 326492 703236 326496 703292
rect 326432 703232 326496 703236
rect 326512 703292 326576 703296
rect 326512 703236 326516 703292
rect 326516 703236 326572 703292
rect 326572 703236 326576 703292
rect 326512 703232 326576 703236
rect 326592 703292 326656 703296
rect 326592 703236 326596 703292
rect 326596 703236 326652 703292
rect 326652 703236 326656 703292
rect 326592 703232 326656 703236
rect 326672 703292 326736 703296
rect 326672 703236 326676 703292
rect 326676 703236 326732 703292
rect 326732 703236 326736 703292
rect 326672 703232 326736 703236
rect 326752 703292 326816 703296
rect 326752 703236 326756 703292
rect 326756 703236 326812 703292
rect 326812 703236 326816 703292
rect 326752 703232 326816 703236
rect 326272 703212 326336 703216
rect 326272 703156 326276 703212
rect 326276 703156 326332 703212
rect 326332 703156 326336 703212
rect 326272 703152 326336 703156
rect 326352 703212 326416 703216
rect 326352 703156 326356 703212
rect 326356 703156 326412 703212
rect 326412 703156 326416 703212
rect 326352 703152 326416 703156
rect 326432 703212 326496 703216
rect 326432 703156 326436 703212
rect 326436 703156 326492 703212
rect 326492 703156 326496 703212
rect 326432 703152 326496 703156
rect 326512 703212 326576 703216
rect 326512 703156 326516 703212
rect 326516 703156 326572 703212
rect 326572 703156 326576 703212
rect 326512 703152 326576 703156
rect 326592 703212 326656 703216
rect 326592 703156 326596 703212
rect 326596 703156 326652 703212
rect 326652 703156 326656 703212
rect 326592 703152 326656 703156
rect 326672 703212 326736 703216
rect 326672 703156 326676 703212
rect 326676 703156 326732 703212
rect 326732 703156 326736 703212
rect 326672 703152 326736 703156
rect 326752 703212 326816 703216
rect 326752 703156 326756 703212
rect 326756 703156 326812 703212
rect 326812 703156 326816 703212
rect 326752 703152 326816 703156
rect 326272 703132 326336 703136
rect 326272 703076 326276 703132
rect 326276 703076 326332 703132
rect 326332 703076 326336 703132
rect 326272 703072 326336 703076
rect 326352 703132 326416 703136
rect 326352 703076 326356 703132
rect 326356 703076 326412 703132
rect 326412 703076 326416 703132
rect 326352 703072 326416 703076
rect 326432 703132 326496 703136
rect 326432 703076 326436 703132
rect 326436 703076 326492 703132
rect 326492 703076 326496 703132
rect 326432 703072 326496 703076
rect 326512 703132 326576 703136
rect 326512 703076 326516 703132
rect 326516 703076 326572 703132
rect 326572 703076 326576 703132
rect 326512 703072 326576 703076
rect 326592 703132 326656 703136
rect 326592 703076 326596 703132
rect 326596 703076 326652 703132
rect 326652 703076 326656 703132
rect 326592 703072 326656 703076
rect 326672 703132 326736 703136
rect 326672 703076 326676 703132
rect 326676 703076 326732 703132
rect 326732 703076 326736 703132
rect 326672 703072 326736 703076
rect 326752 703132 326816 703136
rect 326752 703076 326756 703132
rect 326756 703076 326812 703132
rect 326812 703076 326816 703132
rect 326752 703072 326816 703076
rect 362272 702903 362336 702907
rect 362272 702847 362276 702903
rect 362276 702847 362332 702903
rect 362332 702847 362336 702903
rect 362272 702843 362336 702847
rect 362352 702903 362416 702907
rect 362352 702847 362356 702903
rect 362356 702847 362412 702903
rect 362412 702847 362416 702903
rect 362352 702843 362416 702847
rect 362432 702903 362496 702907
rect 362432 702847 362436 702903
rect 362436 702847 362492 702903
rect 362492 702847 362496 702903
rect 362432 702843 362496 702847
rect 362512 702903 362576 702907
rect 362512 702847 362516 702903
rect 362516 702847 362572 702903
rect 362572 702847 362576 702903
rect 362512 702843 362576 702847
rect 362592 702903 362656 702907
rect 362592 702847 362596 702903
rect 362596 702847 362652 702903
rect 362652 702847 362656 702903
rect 362592 702843 362656 702847
rect 362672 702903 362736 702907
rect 362672 702847 362676 702903
rect 362676 702847 362732 702903
rect 362732 702847 362736 702903
rect 362672 702843 362736 702847
rect 362752 702903 362816 702907
rect 362752 702847 362756 702903
rect 362756 702847 362812 702903
rect 362812 702847 362816 702903
rect 362752 702843 362816 702847
rect 362272 702823 362336 702827
rect 362272 702767 362276 702823
rect 362276 702767 362332 702823
rect 362332 702767 362336 702823
rect 362272 702763 362336 702767
rect 362352 702823 362416 702827
rect 362352 702767 362356 702823
rect 362356 702767 362412 702823
rect 362412 702767 362416 702823
rect 362352 702763 362416 702767
rect 362432 702823 362496 702827
rect 362432 702767 362436 702823
rect 362436 702767 362492 702823
rect 362492 702767 362496 702823
rect 362432 702763 362496 702767
rect 362512 702823 362576 702827
rect 362512 702767 362516 702823
rect 362516 702767 362572 702823
rect 362572 702767 362576 702823
rect 362512 702763 362576 702767
rect 362592 702823 362656 702827
rect 362592 702767 362596 702823
rect 362596 702767 362652 702823
rect 362652 702767 362656 702823
rect 362592 702763 362656 702767
rect 362672 702823 362736 702827
rect 362672 702767 362676 702823
rect 362676 702767 362732 702823
rect 362732 702767 362736 702823
rect 362672 702763 362736 702767
rect 362752 702823 362816 702827
rect 362752 702767 362756 702823
rect 362756 702767 362812 702823
rect 362812 702767 362816 702823
rect 362752 702763 362816 702767
rect 362272 702743 362336 702747
rect 362272 702687 362276 702743
rect 362276 702687 362332 702743
rect 362332 702687 362336 702743
rect 362272 702683 362336 702687
rect 362352 702743 362416 702747
rect 362352 702687 362356 702743
rect 362356 702687 362412 702743
rect 362412 702687 362416 702743
rect 362352 702683 362416 702687
rect 362432 702743 362496 702747
rect 362432 702687 362436 702743
rect 362436 702687 362492 702743
rect 362492 702687 362496 702743
rect 362432 702683 362496 702687
rect 362512 702743 362576 702747
rect 362512 702687 362516 702743
rect 362516 702687 362572 702743
rect 362572 702687 362576 702743
rect 362512 702683 362576 702687
rect 362592 702743 362656 702747
rect 362592 702687 362596 702743
rect 362596 702687 362652 702743
rect 362652 702687 362656 702743
rect 362592 702683 362656 702687
rect 362672 702743 362736 702747
rect 362672 702687 362676 702743
rect 362676 702687 362732 702743
rect 362732 702687 362736 702743
rect 362672 702683 362736 702687
rect 362752 702743 362816 702747
rect 362752 702687 362756 702743
rect 362756 702687 362812 702743
rect 362812 702687 362816 702743
rect 362752 702683 362816 702687
rect 253032 702564 253096 702568
rect 253032 702508 253036 702564
rect 253036 702508 253092 702564
rect 253092 702508 253096 702564
rect 253032 702504 253096 702508
rect 253112 702564 253176 702568
rect 253112 702508 253116 702564
rect 253116 702508 253172 702564
rect 253172 702508 253176 702564
rect 253112 702504 253176 702508
rect 253192 702564 253256 702568
rect 253192 702508 253196 702564
rect 253196 702508 253252 702564
rect 253252 702508 253256 702564
rect 253192 702504 253256 702508
rect 253272 702564 253336 702568
rect 253272 702508 253276 702564
rect 253276 702508 253332 702564
rect 253332 702508 253336 702564
rect 253272 702504 253336 702508
rect 253352 702564 253416 702568
rect 253352 702508 253356 702564
rect 253356 702508 253412 702564
rect 253412 702508 253416 702564
rect 253352 702504 253416 702508
rect 253432 702564 253496 702568
rect 253432 702508 253436 702564
rect 253436 702508 253492 702564
rect 253492 702508 253496 702564
rect 253432 702504 253496 702508
rect 253512 702564 253576 702568
rect 253512 702508 253516 702564
rect 253516 702508 253572 702564
rect 253572 702508 253576 702564
rect 253512 702504 253576 702508
rect 253032 702484 253096 702488
rect 253032 702428 253036 702484
rect 253036 702428 253092 702484
rect 253092 702428 253096 702484
rect 253032 702424 253096 702428
rect 253112 702484 253176 702488
rect 253112 702428 253116 702484
rect 253116 702428 253172 702484
rect 253172 702428 253176 702484
rect 253112 702424 253176 702428
rect 253192 702484 253256 702488
rect 253192 702428 253196 702484
rect 253196 702428 253252 702484
rect 253252 702428 253256 702484
rect 253192 702424 253256 702428
rect 253272 702484 253336 702488
rect 253272 702428 253276 702484
rect 253276 702428 253332 702484
rect 253332 702428 253336 702484
rect 253272 702424 253336 702428
rect 253352 702484 253416 702488
rect 253352 702428 253356 702484
rect 253356 702428 253412 702484
rect 253412 702428 253416 702484
rect 253352 702424 253416 702428
rect 253432 702484 253496 702488
rect 253432 702428 253436 702484
rect 253436 702428 253492 702484
rect 253492 702428 253496 702484
rect 253432 702424 253496 702428
rect 253512 702484 253576 702488
rect 253512 702428 253516 702484
rect 253516 702428 253572 702484
rect 253572 702428 253576 702484
rect 253512 702424 253576 702428
rect 253032 702404 253096 702408
rect 253032 702348 253036 702404
rect 253036 702348 253092 702404
rect 253092 702348 253096 702404
rect 253032 702344 253096 702348
rect 253112 702404 253176 702408
rect 253112 702348 253116 702404
rect 253116 702348 253172 702404
rect 253172 702348 253176 702404
rect 253112 702344 253176 702348
rect 253192 702404 253256 702408
rect 253192 702348 253196 702404
rect 253196 702348 253252 702404
rect 253252 702348 253256 702404
rect 253192 702344 253256 702348
rect 253272 702404 253336 702408
rect 253272 702348 253276 702404
rect 253276 702348 253332 702404
rect 253332 702348 253336 702404
rect 253272 702344 253336 702348
rect 253352 702404 253416 702408
rect 253352 702348 253356 702404
rect 253356 702348 253412 702404
rect 253412 702348 253416 702404
rect 253352 702344 253416 702348
rect 253432 702404 253496 702408
rect 253432 702348 253436 702404
rect 253436 702348 253492 702404
rect 253492 702348 253496 702404
rect 253432 702344 253496 702348
rect 253512 702404 253576 702408
rect 253512 702348 253516 702404
rect 253516 702348 253572 702404
rect 253572 702348 253576 702404
rect 253512 702344 253576 702348
rect 253032 702324 253096 702328
rect 253032 702268 253036 702324
rect 253036 702268 253092 702324
rect 253092 702268 253096 702324
rect 253032 702264 253096 702268
rect 253112 702324 253176 702328
rect 253112 702268 253116 702324
rect 253116 702268 253172 702324
rect 253172 702268 253176 702324
rect 253112 702264 253176 702268
rect 253192 702324 253256 702328
rect 253192 702268 253196 702324
rect 253196 702268 253252 702324
rect 253252 702268 253256 702324
rect 253192 702264 253256 702268
rect 253272 702324 253336 702328
rect 253272 702268 253276 702324
rect 253276 702268 253332 702324
rect 253332 702268 253336 702324
rect 253272 702264 253336 702268
rect 253352 702324 253416 702328
rect 253352 702268 253356 702324
rect 253356 702268 253412 702324
rect 253412 702268 253416 702324
rect 253352 702264 253416 702268
rect 253432 702324 253496 702328
rect 253432 702268 253436 702324
rect 253436 702268 253492 702324
rect 253492 702268 253496 702324
rect 253432 702264 253496 702268
rect 253512 702324 253576 702328
rect 253512 702268 253516 702324
rect 253516 702268 253572 702324
rect 253572 702268 253576 702324
rect 253512 702264 253576 702268
rect 325032 702604 325096 702608
rect 325032 702548 325036 702604
rect 325036 702548 325092 702604
rect 325092 702548 325096 702604
rect 325032 702544 325096 702548
rect 325112 702604 325176 702608
rect 325112 702548 325116 702604
rect 325116 702548 325172 702604
rect 325172 702548 325176 702604
rect 325112 702544 325176 702548
rect 325192 702604 325256 702608
rect 325192 702548 325196 702604
rect 325196 702548 325252 702604
rect 325252 702548 325256 702604
rect 325192 702544 325256 702548
rect 325272 702604 325336 702608
rect 325272 702548 325276 702604
rect 325276 702548 325332 702604
rect 325332 702548 325336 702604
rect 325272 702544 325336 702548
rect 325352 702604 325416 702608
rect 325352 702548 325356 702604
rect 325356 702548 325412 702604
rect 325412 702548 325416 702604
rect 325352 702544 325416 702548
rect 325432 702604 325496 702608
rect 325432 702548 325436 702604
rect 325436 702548 325492 702604
rect 325492 702548 325496 702604
rect 325432 702544 325496 702548
rect 325512 702604 325576 702608
rect 325512 702548 325516 702604
rect 325516 702548 325572 702604
rect 325572 702548 325576 702604
rect 325512 702544 325576 702548
rect 362272 702663 362336 702667
rect 362272 702607 362276 702663
rect 362276 702607 362332 702663
rect 362332 702607 362336 702663
rect 362272 702603 362336 702607
rect 362352 702663 362416 702667
rect 362352 702607 362356 702663
rect 362356 702607 362412 702663
rect 362412 702607 362416 702663
rect 362352 702603 362416 702607
rect 362432 702663 362496 702667
rect 362432 702607 362436 702663
rect 362436 702607 362492 702663
rect 362492 702607 362496 702663
rect 362432 702603 362496 702607
rect 362512 702663 362576 702667
rect 362512 702607 362516 702663
rect 362516 702607 362572 702663
rect 362572 702607 362576 702663
rect 362512 702603 362576 702607
rect 362592 702663 362656 702667
rect 362592 702607 362596 702663
rect 362596 702607 362652 702663
rect 362652 702607 362656 702663
rect 362592 702603 362656 702607
rect 362672 702663 362736 702667
rect 362672 702607 362676 702663
rect 362676 702607 362732 702663
rect 362732 702607 362736 702663
rect 362672 702603 362736 702607
rect 362752 702663 362816 702667
rect 362752 702607 362756 702663
rect 362756 702607 362812 702663
rect 362812 702607 362816 702663
rect 362752 702603 362816 702607
rect 434272 702766 434336 702770
rect 434272 702710 434276 702766
rect 434276 702710 434332 702766
rect 434332 702710 434336 702766
rect 434272 702706 434336 702710
rect 434352 702766 434416 702770
rect 434352 702710 434356 702766
rect 434356 702710 434412 702766
rect 434412 702710 434416 702766
rect 434352 702706 434416 702710
rect 434432 702766 434496 702770
rect 434432 702710 434436 702766
rect 434436 702710 434492 702766
rect 434492 702710 434496 702766
rect 434432 702706 434496 702710
rect 434512 702766 434576 702770
rect 434512 702710 434516 702766
rect 434516 702710 434572 702766
rect 434572 702710 434576 702766
rect 434512 702706 434576 702710
rect 434592 702766 434656 702770
rect 434592 702710 434596 702766
rect 434596 702710 434652 702766
rect 434652 702710 434656 702766
rect 434592 702706 434656 702710
rect 434672 702766 434736 702770
rect 434672 702710 434676 702766
rect 434676 702710 434732 702766
rect 434732 702710 434736 702766
rect 434672 702706 434736 702710
rect 434752 702766 434816 702770
rect 434752 702710 434756 702766
rect 434756 702710 434812 702766
rect 434812 702710 434816 702766
rect 434752 702706 434816 702710
rect 434272 702686 434336 702690
rect 434272 702630 434276 702686
rect 434276 702630 434332 702686
rect 434332 702630 434336 702686
rect 434272 702626 434336 702630
rect 434352 702686 434416 702690
rect 434352 702630 434356 702686
rect 434356 702630 434412 702686
rect 434412 702630 434416 702686
rect 434352 702626 434416 702630
rect 434432 702686 434496 702690
rect 434432 702630 434436 702686
rect 434436 702630 434492 702686
rect 434492 702630 434496 702686
rect 434432 702626 434496 702630
rect 434512 702686 434576 702690
rect 434512 702630 434516 702686
rect 434516 702630 434572 702686
rect 434572 702630 434576 702686
rect 434512 702626 434576 702630
rect 434592 702686 434656 702690
rect 434592 702630 434596 702686
rect 434596 702630 434652 702686
rect 434652 702630 434656 702686
rect 434592 702626 434656 702630
rect 434672 702686 434736 702690
rect 434672 702630 434676 702686
rect 434676 702630 434732 702686
rect 434732 702630 434736 702686
rect 434672 702626 434736 702630
rect 434752 702686 434816 702690
rect 434752 702630 434756 702686
rect 434756 702630 434812 702686
rect 434812 702630 434816 702686
rect 434752 702626 434816 702630
rect 325032 702524 325096 702528
rect 325032 702468 325036 702524
rect 325036 702468 325092 702524
rect 325092 702468 325096 702524
rect 325032 702464 325096 702468
rect 325112 702524 325176 702528
rect 325112 702468 325116 702524
rect 325116 702468 325172 702524
rect 325172 702468 325176 702524
rect 325112 702464 325176 702468
rect 325192 702524 325256 702528
rect 325192 702468 325196 702524
rect 325196 702468 325252 702524
rect 325252 702468 325256 702524
rect 325192 702464 325256 702468
rect 325272 702524 325336 702528
rect 325272 702468 325276 702524
rect 325276 702468 325332 702524
rect 325332 702468 325336 702524
rect 325272 702464 325336 702468
rect 325352 702524 325416 702528
rect 325352 702468 325356 702524
rect 325356 702468 325412 702524
rect 325412 702468 325416 702524
rect 325352 702464 325416 702468
rect 325432 702524 325496 702528
rect 325432 702468 325436 702524
rect 325436 702468 325492 702524
rect 325492 702468 325496 702524
rect 325432 702464 325496 702468
rect 325512 702524 325576 702528
rect 325512 702468 325516 702524
rect 325516 702468 325572 702524
rect 325572 702468 325576 702524
rect 325512 702464 325576 702468
rect 434272 702606 434336 702610
rect 434272 702550 434276 702606
rect 434276 702550 434332 702606
rect 434332 702550 434336 702606
rect 434272 702546 434336 702550
rect 434352 702606 434416 702610
rect 434352 702550 434356 702606
rect 434356 702550 434412 702606
rect 434412 702550 434416 702606
rect 434352 702546 434416 702550
rect 434432 702606 434496 702610
rect 434432 702550 434436 702606
rect 434436 702550 434492 702606
rect 434492 702550 434496 702606
rect 434432 702546 434496 702550
rect 434512 702606 434576 702610
rect 434512 702550 434516 702606
rect 434516 702550 434572 702606
rect 434572 702550 434576 702606
rect 434512 702546 434576 702550
rect 434592 702606 434656 702610
rect 434592 702550 434596 702606
rect 434596 702550 434652 702606
rect 434652 702550 434656 702606
rect 434592 702546 434656 702550
rect 434672 702606 434736 702610
rect 434672 702550 434676 702606
rect 434676 702550 434732 702606
rect 434732 702550 434736 702606
rect 434672 702546 434736 702550
rect 434752 702606 434816 702610
rect 434752 702550 434756 702606
rect 434756 702550 434812 702606
rect 434812 702550 434816 702606
rect 434752 702546 434816 702550
rect 434272 702526 434336 702530
rect 434272 702470 434276 702526
rect 434276 702470 434332 702526
rect 434332 702470 434336 702526
rect 434272 702466 434336 702470
rect 434352 702526 434416 702530
rect 434352 702470 434356 702526
rect 434356 702470 434412 702526
rect 434412 702470 434416 702526
rect 434352 702466 434416 702470
rect 434432 702526 434496 702530
rect 434432 702470 434436 702526
rect 434436 702470 434492 702526
rect 434492 702470 434496 702526
rect 434432 702466 434496 702470
rect 434512 702526 434576 702530
rect 434512 702470 434516 702526
rect 434516 702470 434572 702526
rect 434572 702470 434576 702526
rect 434512 702466 434576 702470
rect 434592 702526 434656 702530
rect 434592 702470 434596 702526
rect 434596 702470 434652 702526
rect 434652 702470 434656 702526
rect 434592 702466 434656 702470
rect 434672 702526 434736 702530
rect 434672 702470 434676 702526
rect 434676 702470 434732 702526
rect 434732 702470 434736 702526
rect 434672 702466 434736 702470
rect 434752 702526 434816 702530
rect 434752 702470 434756 702526
rect 434756 702470 434812 702526
rect 434812 702470 434816 702526
rect 434752 702466 434816 702470
rect 325032 702444 325096 702448
rect 325032 702388 325036 702444
rect 325036 702388 325092 702444
rect 325092 702388 325096 702444
rect 325032 702384 325096 702388
rect 325112 702444 325176 702448
rect 325112 702388 325116 702444
rect 325116 702388 325172 702444
rect 325172 702388 325176 702444
rect 325112 702384 325176 702388
rect 325192 702444 325256 702448
rect 325192 702388 325196 702444
rect 325196 702388 325252 702444
rect 325252 702388 325256 702444
rect 325192 702384 325256 702388
rect 325272 702444 325336 702448
rect 325272 702388 325276 702444
rect 325276 702388 325332 702444
rect 325332 702388 325336 702444
rect 325272 702384 325336 702388
rect 325352 702444 325416 702448
rect 325352 702388 325356 702444
rect 325356 702388 325412 702444
rect 325412 702388 325416 702444
rect 325352 702384 325416 702388
rect 325432 702444 325496 702448
rect 325432 702388 325436 702444
rect 325436 702388 325492 702444
rect 325492 702388 325496 702444
rect 325432 702384 325496 702388
rect 325512 702444 325576 702448
rect 325512 702388 325516 702444
rect 325516 702388 325572 702444
rect 325572 702388 325576 702444
rect 325512 702384 325576 702388
rect 325032 702364 325096 702368
rect 325032 702308 325036 702364
rect 325036 702308 325092 702364
rect 325092 702308 325096 702364
rect 325032 702304 325096 702308
rect 325112 702364 325176 702368
rect 325112 702308 325116 702364
rect 325116 702308 325172 702364
rect 325172 702308 325176 702364
rect 325112 702304 325176 702308
rect 325192 702364 325256 702368
rect 325192 702308 325196 702364
rect 325196 702308 325252 702364
rect 325252 702308 325256 702364
rect 325192 702304 325256 702308
rect 325272 702364 325336 702368
rect 325272 702308 325276 702364
rect 325276 702308 325332 702364
rect 325332 702308 325336 702364
rect 325272 702304 325336 702308
rect 325352 702364 325416 702368
rect 325352 702308 325356 702364
rect 325356 702308 325412 702364
rect 325412 702308 325416 702364
rect 325352 702304 325416 702308
rect 325432 702364 325496 702368
rect 325432 702308 325436 702364
rect 325436 702308 325492 702364
rect 325492 702308 325496 702364
rect 325432 702304 325496 702308
rect 325512 702364 325576 702368
rect 325512 702308 325516 702364
rect 325516 702308 325572 702364
rect 325572 702308 325576 702364
rect 325512 702304 325576 702308
rect 506272 702520 506336 702524
rect 506272 702464 506276 702520
rect 506276 702464 506332 702520
rect 506332 702464 506336 702520
rect 506272 702460 506336 702464
rect 506352 702520 506416 702524
rect 506352 702464 506356 702520
rect 506356 702464 506412 702520
rect 506412 702464 506416 702520
rect 506352 702460 506416 702464
rect 506432 702520 506496 702524
rect 506432 702464 506436 702520
rect 506436 702464 506492 702520
rect 506492 702464 506496 702520
rect 506432 702460 506496 702464
rect 506512 702520 506576 702524
rect 506512 702464 506516 702520
rect 506516 702464 506572 702520
rect 506572 702464 506576 702520
rect 506512 702460 506576 702464
rect 506592 702520 506656 702524
rect 506592 702464 506596 702520
rect 506596 702464 506652 702520
rect 506652 702464 506656 702520
rect 506592 702460 506656 702464
rect 506672 702520 506736 702524
rect 506672 702464 506676 702520
rect 506676 702464 506732 702520
rect 506732 702464 506736 702520
rect 506672 702460 506736 702464
rect 506752 702520 506816 702524
rect 506752 702464 506756 702520
rect 506756 702464 506812 702520
rect 506812 702464 506816 702520
rect 506752 702460 506816 702464
rect 506272 702440 506336 702444
rect 506272 702384 506276 702440
rect 506276 702384 506332 702440
rect 506332 702384 506336 702440
rect 506272 702380 506336 702384
rect 506352 702440 506416 702444
rect 506352 702384 506356 702440
rect 506356 702384 506412 702440
rect 506412 702384 506416 702440
rect 506352 702380 506416 702384
rect 506432 702440 506496 702444
rect 506432 702384 506436 702440
rect 506436 702384 506492 702440
rect 506492 702384 506496 702440
rect 506432 702380 506496 702384
rect 506512 702440 506576 702444
rect 506512 702384 506516 702440
rect 506516 702384 506572 702440
rect 506572 702384 506576 702440
rect 506512 702380 506576 702384
rect 506592 702440 506656 702444
rect 506592 702384 506596 702440
rect 506596 702384 506652 702440
rect 506652 702384 506656 702440
rect 506592 702380 506656 702384
rect 506672 702440 506736 702444
rect 506672 702384 506676 702440
rect 506676 702384 506732 702440
rect 506732 702384 506736 702440
rect 506672 702380 506736 702384
rect 506752 702440 506816 702444
rect 506752 702384 506756 702440
rect 506756 702384 506812 702440
rect 506812 702384 506816 702440
rect 506752 702380 506816 702384
rect 506272 702360 506336 702364
rect 506272 702304 506276 702360
rect 506276 702304 506332 702360
rect 506332 702304 506336 702360
rect 506272 702300 506336 702304
rect 506352 702360 506416 702364
rect 506352 702304 506356 702360
rect 506356 702304 506412 702360
rect 506412 702304 506416 702360
rect 506352 702300 506416 702304
rect 506432 702360 506496 702364
rect 506432 702304 506436 702360
rect 506436 702304 506492 702360
rect 506492 702304 506496 702360
rect 506432 702300 506496 702304
rect 506512 702360 506576 702364
rect 506512 702304 506516 702360
rect 506516 702304 506572 702360
rect 506572 702304 506576 702360
rect 506512 702300 506576 702304
rect 506592 702360 506656 702364
rect 506592 702304 506596 702360
rect 506596 702304 506652 702360
rect 506652 702304 506656 702360
rect 506592 702300 506656 702304
rect 506672 702360 506736 702364
rect 506672 702304 506676 702360
rect 506676 702304 506732 702360
rect 506732 702304 506736 702360
rect 506672 702300 506736 702304
rect 506752 702360 506816 702364
rect 506752 702304 506756 702360
rect 506756 702304 506812 702360
rect 506812 702304 506816 702360
rect 506752 702300 506816 702304
rect 506272 702280 506336 702284
rect 506272 702224 506276 702280
rect 506276 702224 506332 702280
rect 506332 702224 506336 702280
rect 506272 702220 506336 702224
rect 506352 702280 506416 702284
rect 506352 702224 506356 702280
rect 506356 702224 506412 702280
rect 506412 702224 506416 702280
rect 506352 702220 506416 702224
rect 506432 702280 506496 702284
rect 506432 702224 506436 702280
rect 506436 702224 506492 702280
rect 506492 702224 506496 702280
rect 506432 702220 506496 702224
rect 506512 702280 506576 702284
rect 506512 702224 506516 702280
rect 506516 702224 506572 702280
rect 506572 702224 506576 702280
rect 506512 702220 506576 702224
rect 506592 702280 506656 702284
rect 506592 702224 506596 702280
rect 506596 702224 506652 702280
rect 506652 702224 506656 702280
rect 506592 702220 506656 702224
rect 506672 702280 506736 702284
rect 506672 702224 506676 702280
rect 506676 702224 506732 702280
rect 506732 702224 506736 702280
rect 506672 702220 506736 702224
rect 506752 702280 506816 702284
rect 506752 702224 506756 702280
rect 506756 702224 506812 702280
rect 506812 702224 506816 702280
rect 506752 702220 506816 702224
rect 361032 702135 361096 702139
rect 361032 702079 361036 702135
rect 361036 702079 361092 702135
rect 361092 702079 361096 702135
rect 361032 702075 361096 702079
rect 361112 702135 361176 702139
rect 361112 702079 361116 702135
rect 361116 702079 361172 702135
rect 361172 702079 361176 702135
rect 361112 702075 361176 702079
rect 361192 702135 361256 702139
rect 361192 702079 361196 702135
rect 361196 702079 361252 702135
rect 361252 702079 361256 702135
rect 361192 702075 361256 702079
rect 361272 702135 361336 702139
rect 361272 702079 361276 702135
rect 361276 702079 361332 702135
rect 361332 702079 361336 702135
rect 361272 702075 361336 702079
rect 361352 702135 361416 702139
rect 361352 702079 361356 702135
rect 361356 702079 361412 702135
rect 361412 702079 361416 702135
rect 361352 702075 361416 702079
rect 361432 702135 361496 702139
rect 361432 702079 361436 702135
rect 361436 702079 361492 702135
rect 361492 702079 361496 702135
rect 361432 702075 361496 702079
rect 361512 702135 361576 702139
rect 361512 702079 361516 702135
rect 361516 702079 361572 702135
rect 361572 702079 361576 702135
rect 361512 702075 361576 702079
rect 361032 702055 361096 702059
rect 361032 701999 361036 702055
rect 361036 701999 361092 702055
rect 361092 701999 361096 702055
rect 361032 701995 361096 701999
rect 361112 702055 361176 702059
rect 361112 701999 361116 702055
rect 361116 701999 361172 702055
rect 361172 701999 361176 702055
rect 361112 701995 361176 701999
rect 361192 702055 361256 702059
rect 361192 701999 361196 702055
rect 361196 701999 361252 702055
rect 361252 701999 361256 702055
rect 361192 701995 361256 701999
rect 361272 702055 361336 702059
rect 361272 701999 361276 702055
rect 361276 701999 361332 702055
rect 361332 701999 361336 702055
rect 361272 701995 361336 701999
rect 361352 702055 361416 702059
rect 361352 701999 361356 702055
rect 361356 701999 361412 702055
rect 361412 701999 361416 702055
rect 361352 701995 361416 701999
rect 361432 702055 361496 702059
rect 361432 701999 361436 702055
rect 361436 701999 361492 702055
rect 361492 701999 361496 702055
rect 361432 701995 361496 701999
rect 361512 702055 361576 702059
rect 361512 701999 361516 702055
rect 361516 701999 361572 702055
rect 361572 701999 361576 702055
rect 361512 701995 361576 701999
rect 361032 701975 361096 701979
rect 361032 701919 361036 701975
rect 361036 701919 361092 701975
rect 361092 701919 361096 701975
rect 361032 701915 361096 701919
rect 361112 701975 361176 701979
rect 361112 701919 361116 701975
rect 361116 701919 361172 701975
rect 361172 701919 361176 701975
rect 361112 701915 361176 701919
rect 361192 701975 361256 701979
rect 361192 701919 361196 701975
rect 361196 701919 361252 701975
rect 361252 701919 361256 701975
rect 361192 701915 361256 701919
rect 361272 701975 361336 701979
rect 361272 701919 361276 701975
rect 361276 701919 361332 701975
rect 361332 701919 361336 701975
rect 361272 701915 361336 701919
rect 361352 701975 361416 701979
rect 361352 701919 361356 701975
rect 361356 701919 361412 701975
rect 361412 701919 361416 701975
rect 361352 701915 361416 701919
rect 361432 701975 361496 701979
rect 361432 701919 361436 701975
rect 361436 701919 361492 701975
rect 361492 701919 361496 701975
rect 361432 701915 361496 701919
rect 361512 701975 361576 701979
rect 361512 701919 361516 701975
rect 361516 701919 361572 701975
rect 361572 701919 361576 701975
rect 361512 701915 361576 701919
rect 361032 701895 361096 701899
rect 361032 701839 361036 701895
rect 361036 701839 361092 701895
rect 361092 701839 361096 701895
rect 361032 701835 361096 701839
rect 361112 701895 361176 701899
rect 361112 701839 361116 701895
rect 361116 701839 361172 701895
rect 361172 701839 361176 701895
rect 361112 701835 361176 701839
rect 361192 701895 361256 701899
rect 361192 701839 361196 701895
rect 361196 701839 361252 701895
rect 361252 701839 361256 701895
rect 361192 701835 361256 701839
rect 361272 701895 361336 701899
rect 361272 701839 361276 701895
rect 361276 701839 361332 701895
rect 361332 701839 361336 701895
rect 361272 701835 361336 701839
rect 361352 701895 361416 701899
rect 361352 701839 361356 701895
rect 361356 701839 361412 701895
rect 361412 701839 361416 701895
rect 361352 701835 361416 701839
rect 361432 701895 361496 701899
rect 361432 701839 361436 701895
rect 361436 701839 361492 701895
rect 361492 701839 361496 701895
rect 361432 701835 361496 701839
rect 361512 701895 361576 701899
rect 361512 701839 361516 701895
rect 361516 701839 361572 701895
rect 361572 701839 361576 701895
rect 361512 701835 361576 701839
rect 433032 701998 433096 702002
rect 433032 701942 433036 701998
rect 433036 701942 433092 701998
rect 433092 701942 433096 701998
rect 433032 701938 433096 701942
rect 433112 701998 433176 702002
rect 433112 701942 433116 701998
rect 433116 701942 433172 701998
rect 433172 701942 433176 701998
rect 433112 701938 433176 701942
rect 433192 701998 433256 702002
rect 433192 701942 433196 701998
rect 433196 701942 433252 701998
rect 433252 701942 433256 701998
rect 433192 701938 433256 701942
rect 433272 701998 433336 702002
rect 433272 701942 433276 701998
rect 433276 701942 433332 701998
rect 433332 701942 433336 701998
rect 433272 701938 433336 701942
rect 433352 701998 433416 702002
rect 433352 701942 433356 701998
rect 433356 701942 433412 701998
rect 433412 701942 433416 701998
rect 433352 701938 433416 701942
rect 433432 701998 433496 702002
rect 433432 701942 433436 701998
rect 433436 701942 433492 701998
rect 433492 701942 433496 701998
rect 433432 701938 433496 701942
rect 433512 701998 433576 702002
rect 433512 701942 433516 701998
rect 433516 701942 433572 701998
rect 433572 701942 433576 701998
rect 433512 701938 433576 701942
rect 433032 701918 433096 701922
rect 433032 701862 433036 701918
rect 433036 701862 433092 701918
rect 433092 701862 433096 701918
rect 433032 701858 433096 701862
rect 433112 701918 433176 701922
rect 433112 701862 433116 701918
rect 433116 701862 433172 701918
rect 433172 701862 433176 701918
rect 433112 701858 433176 701862
rect 433192 701918 433256 701922
rect 433192 701862 433196 701918
rect 433196 701862 433252 701918
rect 433252 701862 433256 701918
rect 433192 701858 433256 701862
rect 433272 701918 433336 701922
rect 433272 701862 433276 701918
rect 433276 701862 433332 701918
rect 433332 701862 433336 701918
rect 433272 701858 433336 701862
rect 433352 701918 433416 701922
rect 433352 701862 433356 701918
rect 433356 701862 433412 701918
rect 433412 701862 433416 701918
rect 433352 701858 433416 701862
rect 433432 701918 433496 701922
rect 433432 701862 433436 701918
rect 433436 701862 433492 701918
rect 433492 701862 433496 701918
rect 433432 701858 433496 701862
rect 433512 701918 433576 701922
rect 433512 701862 433516 701918
rect 433516 701862 433572 701918
rect 433572 701862 433576 701918
rect 433512 701858 433576 701862
rect 433032 701838 433096 701842
rect 433032 701782 433036 701838
rect 433036 701782 433092 701838
rect 433092 701782 433096 701838
rect 433032 701778 433096 701782
rect 433112 701838 433176 701842
rect 433112 701782 433116 701838
rect 433116 701782 433172 701838
rect 433172 701782 433176 701838
rect 433112 701778 433176 701782
rect 433192 701838 433256 701842
rect 433192 701782 433196 701838
rect 433196 701782 433252 701838
rect 433252 701782 433256 701838
rect 433192 701778 433256 701782
rect 433272 701838 433336 701842
rect 433272 701782 433276 701838
rect 433276 701782 433332 701838
rect 433332 701782 433336 701838
rect 433272 701778 433336 701782
rect 433352 701838 433416 701842
rect 433352 701782 433356 701838
rect 433356 701782 433412 701838
rect 433412 701782 433416 701838
rect 433352 701778 433416 701782
rect 433432 701838 433496 701842
rect 433432 701782 433436 701838
rect 433436 701782 433492 701838
rect 433492 701782 433496 701838
rect 433432 701778 433496 701782
rect 433512 701838 433576 701842
rect 433512 701782 433516 701838
rect 433516 701782 433572 701838
rect 433572 701782 433576 701838
rect 433512 701778 433576 701782
rect 433032 701758 433096 701762
rect 433032 701702 433036 701758
rect 433036 701702 433092 701758
rect 433092 701702 433096 701758
rect 433032 701698 433096 701702
rect 433112 701758 433176 701762
rect 433112 701702 433116 701758
rect 433116 701702 433172 701758
rect 433172 701702 433176 701758
rect 433112 701698 433176 701702
rect 433192 701758 433256 701762
rect 433192 701702 433196 701758
rect 433196 701702 433252 701758
rect 433252 701702 433256 701758
rect 433192 701698 433256 701702
rect 433272 701758 433336 701762
rect 433272 701702 433276 701758
rect 433276 701702 433332 701758
rect 433332 701702 433336 701758
rect 433272 701698 433336 701702
rect 433352 701758 433416 701762
rect 433352 701702 433356 701758
rect 433356 701702 433412 701758
rect 433412 701702 433416 701758
rect 433352 701698 433416 701702
rect 433432 701758 433496 701762
rect 433432 701702 433436 701758
rect 433436 701702 433492 701758
rect 433492 701702 433496 701758
rect 433432 701698 433496 701702
rect 433512 701758 433576 701762
rect 433512 701702 433516 701758
rect 433516 701702 433572 701758
rect 433572 701702 433576 701758
rect 433512 701698 433576 701702
rect 505032 701752 505096 701756
rect 505032 701696 505036 701752
rect 505036 701696 505092 701752
rect 505092 701696 505096 701752
rect 505032 701692 505096 701696
rect 505112 701752 505176 701756
rect 505112 701696 505116 701752
rect 505116 701696 505172 701752
rect 505172 701696 505176 701752
rect 505112 701692 505176 701696
rect 505192 701752 505256 701756
rect 505192 701696 505196 701752
rect 505196 701696 505252 701752
rect 505252 701696 505256 701752
rect 505192 701692 505256 701696
rect 505272 701752 505336 701756
rect 505272 701696 505276 701752
rect 505276 701696 505332 701752
rect 505332 701696 505336 701752
rect 505272 701692 505336 701696
rect 505352 701752 505416 701756
rect 505352 701696 505356 701752
rect 505356 701696 505412 701752
rect 505412 701696 505416 701752
rect 505352 701692 505416 701696
rect 505432 701752 505496 701756
rect 505432 701696 505436 701752
rect 505436 701696 505492 701752
rect 505492 701696 505496 701752
rect 505432 701692 505496 701696
rect 505512 701752 505576 701756
rect 505512 701696 505516 701752
rect 505516 701696 505572 701752
rect 505572 701696 505576 701752
rect 505512 701692 505576 701696
rect 505032 701672 505096 701676
rect 505032 701616 505036 701672
rect 505036 701616 505092 701672
rect 505092 701616 505096 701672
rect 505032 701612 505096 701616
rect 505112 701672 505176 701676
rect 505112 701616 505116 701672
rect 505116 701616 505172 701672
rect 505172 701616 505176 701672
rect 505112 701612 505176 701616
rect 505192 701672 505256 701676
rect 505192 701616 505196 701672
rect 505196 701616 505252 701672
rect 505252 701616 505256 701672
rect 505192 701612 505256 701616
rect 505272 701672 505336 701676
rect 505272 701616 505276 701672
rect 505276 701616 505332 701672
rect 505332 701616 505336 701672
rect 505272 701612 505336 701616
rect 505352 701672 505416 701676
rect 505352 701616 505356 701672
rect 505356 701616 505412 701672
rect 505412 701616 505416 701672
rect 505352 701612 505416 701616
rect 505432 701672 505496 701676
rect 505432 701616 505436 701672
rect 505436 701616 505492 701672
rect 505492 701616 505496 701672
rect 505432 701612 505496 701616
rect 505512 701672 505576 701676
rect 505512 701616 505516 701672
rect 505516 701616 505572 701672
rect 505572 701616 505576 701672
rect 505512 701612 505576 701616
rect 505032 701592 505096 701596
rect 505032 701536 505036 701592
rect 505036 701536 505092 701592
rect 505092 701536 505096 701592
rect 505032 701532 505096 701536
rect 505112 701592 505176 701596
rect 505112 701536 505116 701592
rect 505116 701536 505172 701592
rect 505172 701536 505176 701592
rect 505112 701532 505176 701536
rect 505192 701592 505256 701596
rect 505192 701536 505196 701592
rect 505196 701536 505252 701592
rect 505252 701536 505256 701592
rect 505192 701532 505256 701536
rect 505272 701592 505336 701596
rect 505272 701536 505276 701592
rect 505276 701536 505332 701592
rect 505332 701536 505336 701592
rect 505272 701532 505336 701536
rect 505352 701592 505416 701596
rect 505352 701536 505356 701592
rect 505356 701536 505412 701592
rect 505412 701536 505416 701592
rect 505352 701532 505416 701536
rect 505432 701592 505496 701596
rect 505432 701536 505436 701592
rect 505436 701536 505492 701592
rect 505492 701536 505496 701592
rect 505432 701532 505496 701536
rect 505512 701592 505576 701596
rect 505512 701536 505516 701592
rect 505516 701536 505572 701592
rect 505572 701536 505576 701592
rect 505512 701532 505576 701536
rect 505032 701512 505096 701516
rect 505032 701456 505036 701512
rect 505036 701456 505092 701512
rect 505092 701456 505096 701512
rect 505032 701452 505096 701456
rect 505112 701512 505176 701516
rect 505112 701456 505116 701512
rect 505116 701456 505172 701512
rect 505172 701456 505176 701512
rect 505112 701452 505176 701456
rect 505192 701512 505256 701516
rect 505192 701456 505196 701512
rect 505196 701456 505252 701512
rect 505252 701456 505256 701512
rect 505192 701452 505256 701456
rect 505272 701512 505336 701516
rect 505272 701456 505276 701512
rect 505276 701456 505332 701512
rect 505332 701456 505336 701512
rect 505272 701452 505336 701456
rect 505352 701512 505416 701516
rect 505352 701456 505356 701512
rect 505356 701456 505412 701512
rect 505412 701456 505416 701512
rect 505352 701452 505416 701456
rect 505432 701512 505496 701516
rect 505432 701456 505436 701512
rect 505436 701456 505492 701512
rect 505492 701456 505496 701512
rect 505432 701452 505496 701456
rect 505512 701512 505576 701516
rect 505512 701456 505516 701512
rect 505516 701456 505572 701512
rect 505572 701456 505576 701512
rect 505512 701452 505576 701456
rect 577032 697906 577096 697910
rect 577032 697850 577036 697906
rect 577036 697850 577092 697906
rect 577092 697850 577096 697906
rect 577032 697846 577096 697850
rect 577112 697906 577176 697910
rect 577112 697850 577116 697906
rect 577116 697850 577172 697906
rect 577172 697850 577176 697906
rect 577112 697846 577176 697850
rect 577192 697906 577256 697910
rect 577192 697850 577196 697906
rect 577196 697850 577252 697906
rect 577252 697850 577256 697906
rect 577192 697846 577256 697850
rect 577272 697906 577336 697910
rect 577272 697850 577276 697906
rect 577276 697850 577332 697906
rect 577332 697850 577336 697906
rect 577272 697846 577336 697850
rect 577352 697906 577416 697910
rect 577352 697850 577356 697906
rect 577356 697850 577412 697906
rect 577412 697850 577416 697906
rect 577352 697846 577416 697850
rect 577432 697906 577496 697910
rect 577432 697850 577436 697906
rect 577436 697850 577492 697906
rect 577492 697850 577496 697906
rect 577432 697846 577496 697850
rect 577512 697906 577576 697910
rect 577512 697850 577516 697906
rect 577516 697850 577572 697906
rect 577572 697850 577576 697906
rect 577512 697846 577576 697850
rect 577032 697826 577096 697830
rect 577032 697770 577036 697826
rect 577036 697770 577092 697826
rect 577092 697770 577096 697826
rect 577032 697766 577096 697770
rect 577112 697826 577176 697830
rect 577112 697770 577116 697826
rect 577116 697770 577172 697826
rect 577172 697770 577176 697826
rect 577112 697766 577176 697770
rect 577192 697826 577256 697830
rect 577192 697770 577196 697826
rect 577196 697770 577252 697826
rect 577252 697770 577256 697826
rect 577192 697766 577256 697770
rect 577272 697826 577336 697830
rect 577272 697770 577276 697826
rect 577276 697770 577332 697826
rect 577332 697770 577336 697826
rect 577272 697766 577336 697770
rect 577352 697826 577416 697830
rect 577352 697770 577356 697826
rect 577356 697770 577412 697826
rect 577412 697770 577416 697826
rect 577352 697766 577416 697770
rect 577432 697826 577496 697830
rect 577432 697770 577436 697826
rect 577436 697770 577492 697826
rect 577492 697770 577496 697826
rect 577432 697766 577496 697770
rect 577512 697826 577576 697830
rect 577512 697770 577516 697826
rect 577516 697770 577572 697826
rect 577572 697770 577576 697826
rect 577512 697766 577576 697770
rect 577032 697746 577096 697750
rect 577032 697690 577036 697746
rect 577036 697690 577092 697746
rect 577092 697690 577096 697746
rect 577032 697686 577096 697690
rect 577112 697746 577176 697750
rect 577112 697690 577116 697746
rect 577116 697690 577172 697746
rect 577172 697690 577176 697746
rect 577112 697686 577176 697690
rect 577192 697746 577256 697750
rect 577192 697690 577196 697746
rect 577196 697690 577252 697746
rect 577252 697690 577256 697746
rect 577192 697686 577256 697690
rect 577272 697746 577336 697750
rect 577272 697690 577276 697746
rect 577276 697690 577332 697746
rect 577332 697690 577336 697746
rect 577272 697686 577336 697690
rect 577352 697746 577416 697750
rect 577352 697690 577356 697746
rect 577356 697690 577412 697746
rect 577412 697690 577416 697746
rect 577352 697686 577416 697690
rect 577432 697746 577496 697750
rect 577432 697690 577436 697746
rect 577436 697690 577492 697746
rect 577492 697690 577496 697746
rect 577432 697686 577496 697690
rect 577512 697746 577576 697750
rect 577512 697690 577516 697746
rect 577516 697690 577572 697746
rect 577572 697690 577576 697746
rect 577512 697686 577576 697690
rect 577032 697666 577096 697670
rect 577032 697610 577036 697666
rect 577036 697610 577092 697666
rect 577092 697610 577096 697666
rect 577032 697606 577096 697610
rect 577112 697666 577176 697670
rect 577112 697610 577116 697666
rect 577116 697610 577172 697666
rect 577172 697610 577176 697666
rect 577112 697606 577176 697610
rect 577192 697666 577256 697670
rect 577192 697610 577196 697666
rect 577196 697610 577252 697666
rect 577252 697610 577256 697666
rect 577192 697606 577256 697610
rect 577272 697666 577336 697670
rect 577272 697610 577276 697666
rect 577276 697610 577332 697666
rect 577332 697610 577336 697666
rect 577272 697606 577336 697610
rect 577352 697666 577416 697670
rect 577352 697610 577356 697666
rect 577356 697610 577412 697666
rect 577412 697610 577416 697666
rect 577352 697606 577416 697610
rect 577432 697666 577496 697670
rect 577432 697610 577436 697666
rect 577436 697610 577492 697666
rect 577492 697610 577496 697666
rect 577432 697606 577496 697610
rect 577512 697666 577576 697670
rect 577512 697610 577516 697666
rect 577516 697610 577572 697666
rect 577572 697610 577576 697666
rect 577512 697606 577576 697610
rect 578272 697111 578336 697115
rect 578272 697055 578276 697111
rect 578276 697055 578332 697111
rect 578332 697055 578336 697111
rect 578272 697051 578336 697055
rect 578352 697111 578416 697115
rect 578352 697055 578356 697111
rect 578356 697055 578412 697111
rect 578412 697055 578416 697111
rect 578352 697051 578416 697055
rect 578432 697111 578496 697115
rect 578432 697055 578436 697111
rect 578436 697055 578492 697111
rect 578492 697055 578496 697111
rect 578432 697051 578496 697055
rect 578512 697111 578576 697115
rect 578512 697055 578516 697111
rect 578516 697055 578572 697111
rect 578572 697055 578576 697111
rect 578512 697051 578576 697055
rect 578592 697111 578656 697115
rect 578592 697055 578596 697111
rect 578596 697055 578652 697111
rect 578652 697055 578656 697111
rect 578592 697051 578656 697055
rect 578672 697111 578736 697115
rect 578672 697055 578676 697111
rect 578676 697055 578732 697111
rect 578732 697055 578736 697111
rect 578672 697051 578736 697055
rect 578752 697111 578816 697115
rect 578752 697055 578756 697111
rect 578756 697055 578812 697111
rect 578812 697055 578816 697111
rect 578752 697051 578816 697055
rect 578272 697031 578336 697035
rect 578272 696975 578276 697031
rect 578276 696975 578332 697031
rect 578332 696975 578336 697031
rect 578272 696971 578336 696975
rect 578352 697031 578416 697035
rect 578352 696975 578356 697031
rect 578356 696975 578412 697031
rect 578412 696975 578416 697031
rect 578352 696971 578416 696975
rect 578432 697031 578496 697035
rect 578432 696975 578436 697031
rect 578436 696975 578492 697031
rect 578492 696975 578496 697031
rect 578432 696971 578496 696975
rect 578512 697031 578576 697035
rect 578512 696975 578516 697031
rect 578516 696975 578572 697031
rect 578572 696975 578576 697031
rect 578512 696971 578576 696975
rect 578592 697031 578656 697035
rect 578592 696975 578596 697031
rect 578596 696975 578652 697031
rect 578652 696975 578656 697031
rect 578592 696971 578656 696975
rect 578672 697031 578736 697035
rect 578672 696975 578676 697031
rect 578676 696975 578732 697031
rect 578732 696975 578736 697031
rect 578672 696971 578736 696975
rect 578752 697031 578816 697035
rect 578752 696975 578756 697031
rect 578756 696975 578812 697031
rect 578812 696975 578816 697031
rect 578752 696971 578816 696975
rect 578272 696951 578336 696955
rect 578272 696895 578276 696951
rect 578276 696895 578332 696951
rect 578332 696895 578336 696951
rect 578272 696891 578336 696895
rect 578352 696951 578416 696955
rect 578352 696895 578356 696951
rect 578356 696895 578412 696951
rect 578412 696895 578416 696951
rect 578352 696891 578416 696895
rect 578432 696951 578496 696955
rect 578432 696895 578436 696951
rect 578436 696895 578492 696951
rect 578492 696895 578496 696951
rect 578432 696891 578496 696895
rect 578512 696951 578576 696955
rect 578512 696895 578516 696951
rect 578516 696895 578572 696951
rect 578572 696895 578576 696951
rect 578512 696891 578576 696895
rect 578592 696951 578656 696955
rect 578592 696895 578596 696951
rect 578596 696895 578652 696951
rect 578652 696895 578656 696951
rect 578592 696891 578656 696895
rect 578672 696951 578736 696955
rect 578672 696895 578676 696951
rect 578676 696895 578732 696951
rect 578732 696895 578736 696951
rect 578672 696891 578736 696895
rect 578752 696951 578816 696955
rect 578752 696895 578756 696951
rect 578756 696895 578812 696951
rect 578812 696895 578816 696951
rect 578752 696891 578816 696895
rect 578272 696871 578336 696875
rect 578272 696815 578276 696871
rect 578276 696815 578332 696871
rect 578332 696815 578336 696871
rect 578272 696811 578336 696815
rect 578352 696871 578416 696875
rect 578352 696815 578356 696871
rect 578356 696815 578412 696871
rect 578412 696815 578416 696871
rect 578352 696811 578416 696815
rect 578432 696871 578496 696875
rect 578432 696815 578436 696871
rect 578436 696815 578492 696871
rect 578492 696815 578496 696871
rect 578432 696811 578496 696815
rect 578512 696871 578576 696875
rect 578512 696815 578516 696871
rect 578516 696815 578572 696871
rect 578572 696815 578576 696871
rect 578512 696811 578576 696815
rect 578592 696871 578656 696875
rect 578592 696815 578596 696871
rect 578596 696815 578652 696871
rect 578652 696815 578656 696871
rect 578592 696811 578656 696815
rect 578672 696871 578736 696875
rect 578672 696815 578676 696871
rect 578676 696815 578732 696871
rect 578732 696815 578736 696871
rect 578672 696811 578736 696815
rect 578752 696871 578816 696875
rect 578752 696815 578756 696871
rect 578756 696815 578812 696871
rect 578812 696815 578816 696871
rect 578752 696811 578816 696815
rect 577032 644730 577096 644734
rect 577032 644674 577036 644730
rect 577036 644674 577092 644730
rect 577092 644674 577096 644730
rect 577032 644670 577096 644674
rect 577112 644730 577176 644734
rect 577112 644674 577116 644730
rect 577116 644674 577172 644730
rect 577172 644674 577176 644730
rect 577112 644670 577176 644674
rect 577192 644730 577256 644734
rect 577192 644674 577196 644730
rect 577196 644674 577252 644730
rect 577252 644674 577256 644730
rect 577192 644670 577256 644674
rect 577272 644730 577336 644734
rect 577272 644674 577276 644730
rect 577276 644674 577332 644730
rect 577332 644674 577336 644730
rect 577272 644670 577336 644674
rect 577352 644730 577416 644734
rect 577352 644674 577356 644730
rect 577356 644674 577412 644730
rect 577412 644674 577416 644730
rect 577352 644670 577416 644674
rect 577432 644730 577496 644734
rect 577432 644674 577436 644730
rect 577436 644674 577492 644730
rect 577492 644674 577496 644730
rect 577432 644670 577496 644674
rect 577512 644730 577576 644734
rect 577512 644674 577516 644730
rect 577516 644674 577572 644730
rect 577572 644674 577576 644730
rect 577512 644670 577576 644674
rect 577032 644650 577096 644654
rect 577032 644594 577036 644650
rect 577036 644594 577092 644650
rect 577092 644594 577096 644650
rect 577032 644590 577096 644594
rect 577112 644650 577176 644654
rect 577112 644594 577116 644650
rect 577116 644594 577172 644650
rect 577172 644594 577176 644650
rect 577112 644590 577176 644594
rect 577192 644650 577256 644654
rect 577192 644594 577196 644650
rect 577196 644594 577252 644650
rect 577252 644594 577256 644650
rect 577192 644590 577256 644594
rect 577272 644650 577336 644654
rect 577272 644594 577276 644650
rect 577276 644594 577332 644650
rect 577332 644594 577336 644650
rect 577272 644590 577336 644594
rect 577352 644650 577416 644654
rect 577352 644594 577356 644650
rect 577356 644594 577412 644650
rect 577412 644594 577416 644650
rect 577352 644590 577416 644594
rect 577432 644650 577496 644654
rect 577432 644594 577436 644650
rect 577436 644594 577492 644650
rect 577492 644594 577496 644650
rect 577432 644590 577496 644594
rect 577512 644650 577576 644654
rect 577512 644594 577516 644650
rect 577516 644594 577572 644650
rect 577572 644594 577576 644650
rect 577512 644590 577576 644594
rect 577032 644570 577096 644574
rect 577032 644514 577036 644570
rect 577036 644514 577092 644570
rect 577092 644514 577096 644570
rect 577032 644510 577096 644514
rect 577112 644570 577176 644574
rect 577112 644514 577116 644570
rect 577116 644514 577172 644570
rect 577172 644514 577176 644570
rect 577112 644510 577176 644514
rect 577192 644570 577256 644574
rect 577192 644514 577196 644570
rect 577196 644514 577252 644570
rect 577252 644514 577256 644570
rect 577192 644510 577256 644514
rect 577272 644570 577336 644574
rect 577272 644514 577276 644570
rect 577276 644514 577332 644570
rect 577332 644514 577336 644570
rect 577272 644510 577336 644514
rect 577352 644570 577416 644574
rect 577352 644514 577356 644570
rect 577356 644514 577412 644570
rect 577412 644514 577416 644570
rect 577352 644510 577416 644514
rect 577432 644570 577496 644574
rect 577432 644514 577436 644570
rect 577436 644514 577492 644570
rect 577492 644514 577496 644570
rect 577432 644510 577496 644514
rect 577512 644570 577576 644574
rect 577512 644514 577516 644570
rect 577516 644514 577572 644570
rect 577572 644514 577576 644570
rect 577512 644510 577576 644514
rect 577032 644490 577096 644494
rect 577032 644434 577036 644490
rect 577036 644434 577092 644490
rect 577092 644434 577096 644490
rect 577032 644430 577096 644434
rect 577112 644490 577176 644494
rect 577112 644434 577116 644490
rect 577116 644434 577172 644490
rect 577172 644434 577176 644490
rect 577112 644430 577176 644434
rect 577192 644490 577256 644494
rect 577192 644434 577196 644490
rect 577196 644434 577252 644490
rect 577252 644434 577256 644490
rect 577192 644430 577256 644434
rect 577272 644490 577336 644494
rect 577272 644434 577276 644490
rect 577276 644434 577332 644490
rect 577332 644434 577336 644490
rect 577272 644430 577336 644434
rect 577352 644490 577416 644494
rect 577352 644434 577356 644490
rect 577356 644434 577412 644490
rect 577412 644434 577416 644490
rect 577352 644430 577416 644434
rect 577432 644490 577496 644494
rect 577432 644434 577436 644490
rect 577436 644434 577492 644490
rect 577492 644434 577496 644490
rect 577432 644430 577496 644434
rect 577512 644490 577576 644494
rect 577512 644434 577516 644490
rect 577516 644434 577572 644490
rect 577572 644434 577576 644490
rect 577512 644430 577576 644434
rect 578272 643935 578336 643939
rect 578272 643879 578276 643935
rect 578276 643879 578332 643935
rect 578332 643879 578336 643935
rect 578272 643875 578336 643879
rect 578352 643935 578416 643939
rect 578352 643879 578356 643935
rect 578356 643879 578412 643935
rect 578412 643879 578416 643935
rect 578352 643875 578416 643879
rect 578432 643935 578496 643939
rect 578432 643879 578436 643935
rect 578436 643879 578492 643935
rect 578492 643879 578496 643935
rect 578432 643875 578496 643879
rect 578512 643935 578576 643939
rect 578512 643879 578516 643935
rect 578516 643879 578572 643935
rect 578572 643879 578576 643935
rect 578512 643875 578576 643879
rect 578592 643935 578656 643939
rect 578592 643879 578596 643935
rect 578596 643879 578652 643935
rect 578652 643879 578656 643935
rect 578592 643875 578656 643879
rect 578672 643935 578736 643939
rect 578672 643879 578676 643935
rect 578676 643879 578732 643935
rect 578732 643879 578736 643935
rect 578672 643875 578736 643879
rect 578752 643935 578816 643939
rect 578752 643879 578756 643935
rect 578756 643879 578812 643935
rect 578812 643879 578816 643935
rect 578752 643875 578816 643879
rect 578272 643855 578336 643859
rect 578272 643799 578276 643855
rect 578276 643799 578332 643855
rect 578332 643799 578336 643855
rect 578272 643795 578336 643799
rect 578352 643855 578416 643859
rect 578352 643799 578356 643855
rect 578356 643799 578412 643855
rect 578412 643799 578416 643855
rect 578352 643795 578416 643799
rect 578432 643855 578496 643859
rect 578432 643799 578436 643855
rect 578436 643799 578492 643855
rect 578492 643799 578496 643855
rect 578432 643795 578496 643799
rect 578512 643855 578576 643859
rect 578512 643799 578516 643855
rect 578516 643799 578572 643855
rect 578572 643799 578576 643855
rect 578512 643795 578576 643799
rect 578592 643855 578656 643859
rect 578592 643799 578596 643855
rect 578596 643799 578652 643855
rect 578652 643799 578656 643855
rect 578592 643795 578656 643799
rect 578672 643855 578736 643859
rect 578672 643799 578676 643855
rect 578676 643799 578732 643855
rect 578732 643799 578736 643855
rect 578672 643795 578736 643799
rect 578752 643855 578816 643859
rect 578752 643799 578756 643855
rect 578756 643799 578812 643855
rect 578812 643799 578816 643855
rect 578752 643795 578816 643799
rect 578272 643775 578336 643779
rect 578272 643719 578276 643775
rect 578276 643719 578332 643775
rect 578332 643719 578336 643775
rect 578272 643715 578336 643719
rect 578352 643775 578416 643779
rect 578352 643719 578356 643775
rect 578356 643719 578412 643775
rect 578412 643719 578416 643775
rect 578352 643715 578416 643719
rect 578432 643775 578496 643779
rect 578432 643719 578436 643775
rect 578436 643719 578492 643775
rect 578492 643719 578496 643775
rect 578432 643715 578496 643719
rect 578512 643775 578576 643779
rect 578512 643719 578516 643775
rect 578516 643719 578572 643775
rect 578572 643719 578576 643775
rect 578512 643715 578576 643719
rect 578592 643775 578656 643779
rect 578592 643719 578596 643775
rect 578596 643719 578652 643775
rect 578652 643719 578656 643775
rect 578592 643715 578656 643719
rect 578672 643775 578736 643779
rect 578672 643719 578676 643775
rect 578676 643719 578732 643775
rect 578732 643719 578736 643775
rect 578672 643715 578736 643719
rect 578752 643775 578816 643779
rect 578752 643719 578756 643775
rect 578756 643719 578812 643775
rect 578812 643719 578816 643775
rect 578752 643715 578816 643719
rect 578272 643695 578336 643699
rect 578272 643639 578276 643695
rect 578276 643639 578332 643695
rect 578332 643639 578336 643695
rect 578272 643635 578336 643639
rect 578352 643695 578416 643699
rect 578352 643639 578356 643695
rect 578356 643639 578412 643695
rect 578412 643639 578416 643695
rect 578352 643635 578416 643639
rect 578432 643695 578496 643699
rect 578432 643639 578436 643695
rect 578436 643639 578492 643695
rect 578492 643639 578496 643695
rect 578432 643635 578496 643639
rect 578512 643695 578576 643699
rect 578512 643639 578516 643695
rect 578516 643639 578572 643695
rect 578572 643639 578576 643695
rect 578512 643635 578576 643639
rect 578592 643695 578656 643699
rect 578592 643639 578596 643695
rect 578596 643639 578652 643695
rect 578652 643639 578656 643695
rect 578592 643635 578656 643639
rect 578672 643695 578736 643699
rect 578672 643639 578676 643695
rect 578676 643639 578732 643695
rect 578732 643639 578736 643695
rect 578672 643635 578736 643639
rect 578752 643695 578816 643699
rect 578752 643639 578756 643695
rect 578756 643639 578812 643695
rect 578812 643639 578816 643695
rect 578752 643635 578816 643639
rect 577032 591690 577096 591694
rect 577032 591634 577036 591690
rect 577036 591634 577092 591690
rect 577092 591634 577096 591690
rect 577032 591630 577096 591634
rect 577112 591690 577176 591694
rect 577112 591634 577116 591690
rect 577116 591634 577172 591690
rect 577172 591634 577176 591690
rect 577112 591630 577176 591634
rect 577192 591690 577256 591694
rect 577192 591634 577196 591690
rect 577196 591634 577252 591690
rect 577252 591634 577256 591690
rect 577192 591630 577256 591634
rect 577272 591690 577336 591694
rect 577272 591634 577276 591690
rect 577276 591634 577332 591690
rect 577332 591634 577336 591690
rect 577272 591630 577336 591634
rect 577352 591690 577416 591694
rect 577352 591634 577356 591690
rect 577356 591634 577412 591690
rect 577412 591634 577416 591690
rect 577352 591630 577416 591634
rect 577432 591690 577496 591694
rect 577432 591634 577436 591690
rect 577436 591634 577492 591690
rect 577492 591634 577496 591690
rect 577432 591630 577496 591634
rect 577512 591690 577576 591694
rect 577512 591634 577516 591690
rect 577516 591634 577572 591690
rect 577572 591634 577576 591690
rect 577512 591630 577576 591634
rect 577032 591610 577096 591614
rect 577032 591554 577036 591610
rect 577036 591554 577092 591610
rect 577092 591554 577096 591610
rect 577032 591550 577096 591554
rect 577112 591610 577176 591614
rect 577112 591554 577116 591610
rect 577116 591554 577172 591610
rect 577172 591554 577176 591610
rect 577112 591550 577176 591554
rect 577192 591610 577256 591614
rect 577192 591554 577196 591610
rect 577196 591554 577252 591610
rect 577252 591554 577256 591610
rect 577192 591550 577256 591554
rect 577272 591610 577336 591614
rect 577272 591554 577276 591610
rect 577276 591554 577332 591610
rect 577332 591554 577336 591610
rect 577272 591550 577336 591554
rect 577352 591610 577416 591614
rect 577352 591554 577356 591610
rect 577356 591554 577412 591610
rect 577412 591554 577416 591610
rect 577352 591550 577416 591554
rect 577432 591610 577496 591614
rect 577432 591554 577436 591610
rect 577436 591554 577492 591610
rect 577492 591554 577496 591610
rect 577432 591550 577496 591554
rect 577512 591610 577576 591614
rect 577512 591554 577516 591610
rect 577516 591554 577572 591610
rect 577572 591554 577576 591610
rect 577512 591550 577576 591554
rect 577032 591530 577096 591534
rect 577032 591474 577036 591530
rect 577036 591474 577092 591530
rect 577092 591474 577096 591530
rect 577032 591470 577096 591474
rect 577112 591530 577176 591534
rect 577112 591474 577116 591530
rect 577116 591474 577172 591530
rect 577172 591474 577176 591530
rect 577112 591470 577176 591474
rect 577192 591530 577256 591534
rect 577192 591474 577196 591530
rect 577196 591474 577252 591530
rect 577252 591474 577256 591530
rect 577192 591470 577256 591474
rect 577272 591530 577336 591534
rect 577272 591474 577276 591530
rect 577276 591474 577332 591530
rect 577332 591474 577336 591530
rect 577272 591470 577336 591474
rect 577352 591530 577416 591534
rect 577352 591474 577356 591530
rect 577356 591474 577412 591530
rect 577412 591474 577416 591530
rect 577352 591470 577416 591474
rect 577432 591530 577496 591534
rect 577432 591474 577436 591530
rect 577436 591474 577492 591530
rect 577492 591474 577496 591530
rect 577432 591470 577496 591474
rect 577512 591530 577576 591534
rect 577512 591474 577516 591530
rect 577516 591474 577572 591530
rect 577572 591474 577576 591530
rect 577512 591470 577576 591474
rect 577032 591450 577096 591454
rect 577032 591394 577036 591450
rect 577036 591394 577092 591450
rect 577092 591394 577096 591450
rect 577032 591390 577096 591394
rect 577112 591450 577176 591454
rect 577112 591394 577116 591450
rect 577116 591394 577172 591450
rect 577172 591394 577176 591450
rect 577112 591390 577176 591394
rect 577192 591450 577256 591454
rect 577192 591394 577196 591450
rect 577196 591394 577252 591450
rect 577252 591394 577256 591450
rect 577192 591390 577256 591394
rect 577272 591450 577336 591454
rect 577272 591394 577276 591450
rect 577276 591394 577332 591450
rect 577332 591394 577336 591450
rect 577272 591390 577336 591394
rect 577352 591450 577416 591454
rect 577352 591394 577356 591450
rect 577356 591394 577412 591450
rect 577412 591394 577416 591450
rect 577352 591390 577416 591394
rect 577432 591450 577496 591454
rect 577432 591394 577436 591450
rect 577436 591394 577492 591450
rect 577492 591394 577496 591450
rect 577432 591390 577496 591394
rect 577512 591450 577576 591454
rect 577512 591394 577516 591450
rect 577516 591394 577572 591450
rect 577572 591394 577576 591450
rect 577512 591390 577576 591394
rect 578272 590895 578336 590899
rect 578272 590839 578276 590895
rect 578276 590839 578332 590895
rect 578332 590839 578336 590895
rect 578272 590835 578336 590839
rect 578352 590895 578416 590899
rect 578352 590839 578356 590895
rect 578356 590839 578412 590895
rect 578412 590839 578416 590895
rect 578352 590835 578416 590839
rect 578432 590895 578496 590899
rect 578432 590839 578436 590895
rect 578436 590839 578492 590895
rect 578492 590839 578496 590895
rect 578432 590835 578496 590839
rect 578512 590895 578576 590899
rect 578512 590839 578516 590895
rect 578516 590839 578572 590895
rect 578572 590839 578576 590895
rect 578512 590835 578576 590839
rect 578592 590895 578656 590899
rect 578592 590839 578596 590895
rect 578596 590839 578652 590895
rect 578652 590839 578656 590895
rect 578592 590835 578656 590839
rect 578672 590895 578736 590899
rect 578672 590839 578676 590895
rect 578676 590839 578732 590895
rect 578732 590839 578736 590895
rect 578672 590835 578736 590839
rect 578752 590895 578816 590899
rect 578752 590839 578756 590895
rect 578756 590839 578812 590895
rect 578812 590839 578816 590895
rect 578752 590835 578816 590839
rect 578272 590815 578336 590819
rect 578272 590759 578276 590815
rect 578276 590759 578332 590815
rect 578332 590759 578336 590815
rect 578272 590755 578336 590759
rect 578352 590815 578416 590819
rect 578352 590759 578356 590815
rect 578356 590759 578412 590815
rect 578412 590759 578416 590815
rect 578352 590755 578416 590759
rect 578432 590815 578496 590819
rect 578432 590759 578436 590815
rect 578436 590759 578492 590815
rect 578492 590759 578496 590815
rect 578432 590755 578496 590759
rect 578512 590815 578576 590819
rect 578512 590759 578516 590815
rect 578516 590759 578572 590815
rect 578572 590759 578576 590815
rect 578512 590755 578576 590759
rect 578592 590815 578656 590819
rect 578592 590759 578596 590815
rect 578596 590759 578652 590815
rect 578652 590759 578656 590815
rect 578592 590755 578656 590759
rect 578672 590815 578736 590819
rect 578672 590759 578676 590815
rect 578676 590759 578732 590815
rect 578732 590759 578736 590815
rect 578672 590755 578736 590759
rect 578752 590815 578816 590819
rect 578752 590759 578756 590815
rect 578756 590759 578812 590815
rect 578812 590759 578816 590815
rect 578752 590755 578816 590759
rect 578272 590735 578336 590739
rect 578272 590679 578276 590735
rect 578276 590679 578332 590735
rect 578332 590679 578336 590735
rect 578272 590675 578336 590679
rect 578352 590735 578416 590739
rect 578352 590679 578356 590735
rect 578356 590679 578412 590735
rect 578412 590679 578416 590735
rect 578352 590675 578416 590679
rect 578432 590735 578496 590739
rect 578432 590679 578436 590735
rect 578436 590679 578492 590735
rect 578492 590679 578496 590735
rect 578432 590675 578496 590679
rect 578512 590735 578576 590739
rect 578512 590679 578516 590735
rect 578516 590679 578572 590735
rect 578572 590679 578576 590735
rect 578512 590675 578576 590679
rect 578592 590735 578656 590739
rect 578592 590679 578596 590735
rect 578596 590679 578652 590735
rect 578652 590679 578656 590735
rect 578592 590675 578656 590679
rect 578672 590735 578736 590739
rect 578672 590679 578676 590735
rect 578676 590679 578732 590735
rect 578732 590679 578736 590735
rect 578672 590675 578736 590679
rect 578752 590735 578816 590739
rect 578752 590679 578756 590735
rect 578756 590679 578812 590735
rect 578812 590679 578816 590735
rect 578752 590675 578816 590679
rect 578272 590655 578336 590659
rect 578272 590599 578276 590655
rect 578276 590599 578332 590655
rect 578332 590599 578336 590655
rect 578272 590595 578336 590599
rect 578352 590655 578416 590659
rect 578352 590599 578356 590655
rect 578356 590599 578412 590655
rect 578412 590599 578416 590655
rect 578352 590595 578416 590599
rect 578432 590655 578496 590659
rect 578432 590599 578436 590655
rect 578436 590599 578492 590655
rect 578492 590599 578496 590655
rect 578432 590595 578496 590599
rect 578512 590655 578576 590659
rect 578512 590599 578516 590655
rect 578516 590599 578572 590655
rect 578572 590599 578576 590655
rect 578512 590595 578576 590599
rect 578592 590655 578656 590659
rect 578592 590599 578596 590655
rect 578596 590599 578652 590655
rect 578652 590599 578656 590655
rect 578592 590595 578656 590599
rect 578672 590655 578736 590659
rect 578672 590599 578676 590655
rect 578676 590599 578732 590655
rect 578732 590599 578736 590655
rect 578672 590595 578736 590599
rect 578752 590655 578816 590659
rect 578752 590599 578756 590655
rect 578756 590599 578812 590655
rect 578812 590599 578816 590655
rect 578752 590595 578816 590599
rect 505032 554598 505096 554602
rect 505032 554542 505036 554598
rect 505036 554542 505092 554598
rect 505092 554542 505096 554598
rect 505032 554538 505096 554542
rect 505112 554598 505176 554602
rect 505112 554542 505116 554598
rect 505116 554542 505172 554598
rect 505172 554542 505176 554598
rect 505112 554538 505176 554542
rect 505192 554598 505256 554602
rect 505192 554542 505196 554598
rect 505196 554542 505252 554598
rect 505252 554542 505256 554598
rect 505192 554538 505256 554542
rect 505272 554598 505336 554602
rect 505272 554542 505276 554598
rect 505276 554542 505332 554598
rect 505332 554542 505336 554598
rect 505272 554538 505336 554542
rect 505352 554598 505416 554602
rect 505352 554542 505356 554598
rect 505356 554542 505412 554598
rect 505412 554542 505416 554598
rect 505352 554538 505416 554542
rect 505432 554598 505496 554602
rect 505432 554542 505436 554598
rect 505436 554542 505492 554598
rect 505492 554542 505496 554598
rect 505432 554538 505496 554542
rect 505512 554598 505576 554602
rect 505512 554542 505516 554598
rect 505516 554542 505572 554598
rect 505572 554542 505576 554598
rect 505512 554538 505576 554542
rect 505032 554518 505096 554522
rect 505032 554462 505036 554518
rect 505036 554462 505092 554518
rect 505092 554462 505096 554518
rect 505032 554458 505096 554462
rect 505112 554518 505176 554522
rect 505112 554462 505116 554518
rect 505116 554462 505172 554518
rect 505172 554462 505176 554518
rect 505112 554458 505176 554462
rect 505192 554518 505256 554522
rect 505192 554462 505196 554518
rect 505196 554462 505252 554518
rect 505252 554462 505256 554518
rect 505192 554458 505256 554462
rect 505272 554518 505336 554522
rect 505272 554462 505276 554518
rect 505276 554462 505332 554518
rect 505332 554462 505336 554518
rect 505272 554458 505336 554462
rect 505352 554518 505416 554522
rect 505352 554462 505356 554518
rect 505356 554462 505412 554518
rect 505412 554462 505416 554518
rect 505352 554458 505416 554462
rect 505432 554518 505496 554522
rect 505432 554462 505436 554518
rect 505436 554462 505492 554518
rect 505492 554462 505496 554518
rect 505432 554458 505496 554462
rect 505512 554518 505576 554522
rect 505512 554462 505516 554518
rect 505516 554462 505572 554518
rect 505572 554462 505576 554518
rect 505512 554458 505576 554462
rect 505032 554438 505096 554442
rect 505032 554382 505036 554438
rect 505036 554382 505092 554438
rect 505092 554382 505096 554438
rect 505032 554378 505096 554382
rect 505112 554438 505176 554442
rect 505112 554382 505116 554438
rect 505116 554382 505172 554438
rect 505172 554382 505176 554438
rect 505112 554378 505176 554382
rect 505192 554438 505256 554442
rect 505192 554382 505196 554438
rect 505196 554382 505252 554438
rect 505252 554382 505256 554438
rect 505192 554378 505256 554382
rect 505272 554438 505336 554442
rect 505272 554382 505276 554438
rect 505276 554382 505332 554438
rect 505332 554382 505336 554438
rect 505272 554378 505336 554382
rect 505352 554438 505416 554442
rect 505352 554382 505356 554438
rect 505356 554382 505412 554438
rect 505412 554382 505416 554438
rect 505352 554378 505416 554382
rect 505432 554438 505496 554442
rect 505432 554382 505436 554438
rect 505436 554382 505492 554438
rect 505492 554382 505496 554438
rect 505432 554378 505496 554382
rect 505512 554438 505576 554442
rect 505512 554382 505516 554438
rect 505516 554382 505572 554438
rect 505572 554382 505576 554438
rect 505512 554378 505576 554382
rect 505032 554358 505096 554362
rect 505032 554302 505036 554358
rect 505036 554302 505092 554358
rect 505092 554302 505096 554358
rect 505032 554298 505096 554302
rect 505112 554358 505176 554362
rect 505112 554302 505116 554358
rect 505116 554302 505172 554358
rect 505172 554302 505176 554358
rect 505112 554298 505176 554302
rect 505192 554358 505256 554362
rect 505192 554302 505196 554358
rect 505196 554302 505252 554358
rect 505252 554302 505256 554358
rect 505192 554298 505256 554302
rect 505272 554358 505336 554362
rect 505272 554302 505276 554358
rect 505276 554302 505332 554358
rect 505332 554302 505336 554358
rect 505272 554298 505336 554302
rect 505352 554358 505416 554362
rect 505352 554302 505356 554358
rect 505356 554302 505412 554358
rect 505412 554302 505416 554358
rect 505352 554298 505416 554302
rect 505432 554358 505496 554362
rect 505432 554302 505436 554358
rect 505436 554302 505492 554358
rect 505492 554302 505496 554358
rect 505432 554298 505496 554302
rect 505512 554358 505576 554362
rect 505512 554302 505516 554358
rect 505516 554302 505572 554358
rect 505572 554302 505576 554358
rect 505512 554298 505576 554302
rect 506272 553803 506336 553807
rect 506272 553747 506276 553803
rect 506276 553747 506332 553803
rect 506332 553747 506336 553803
rect 506272 553743 506336 553747
rect 506352 553803 506416 553807
rect 506352 553747 506356 553803
rect 506356 553747 506412 553803
rect 506412 553747 506416 553803
rect 506352 553743 506416 553747
rect 506432 553803 506496 553807
rect 506432 553747 506436 553803
rect 506436 553747 506492 553803
rect 506492 553747 506496 553803
rect 506432 553743 506496 553747
rect 506512 553803 506576 553807
rect 506512 553747 506516 553803
rect 506516 553747 506572 553803
rect 506572 553747 506576 553803
rect 506512 553743 506576 553747
rect 506592 553803 506656 553807
rect 506592 553747 506596 553803
rect 506596 553747 506652 553803
rect 506652 553747 506656 553803
rect 506592 553743 506656 553747
rect 506672 553803 506736 553807
rect 506672 553747 506676 553803
rect 506676 553747 506732 553803
rect 506732 553747 506736 553803
rect 506672 553743 506736 553747
rect 506752 553803 506816 553807
rect 506752 553747 506756 553803
rect 506756 553747 506812 553803
rect 506812 553747 506816 553803
rect 506752 553743 506816 553747
rect 506272 553723 506336 553727
rect 506272 553667 506276 553723
rect 506276 553667 506332 553723
rect 506332 553667 506336 553723
rect 506272 553663 506336 553667
rect 506352 553723 506416 553727
rect 506352 553667 506356 553723
rect 506356 553667 506412 553723
rect 506412 553667 506416 553723
rect 506352 553663 506416 553667
rect 506432 553723 506496 553727
rect 506432 553667 506436 553723
rect 506436 553667 506492 553723
rect 506492 553667 506496 553723
rect 506432 553663 506496 553667
rect 506512 553723 506576 553727
rect 506512 553667 506516 553723
rect 506516 553667 506572 553723
rect 506572 553667 506576 553723
rect 506512 553663 506576 553667
rect 506592 553723 506656 553727
rect 506592 553667 506596 553723
rect 506596 553667 506652 553723
rect 506652 553667 506656 553723
rect 506592 553663 506656 553667
rect 506672 553723 506736 553727
rect 506672 553667 506676 553723
rect 506676 553667 506732 553723
rect 506732 553667 506736 553723
rect 506672 553663 506736 553667
rect 506752 553723 506816 553727
rect 506752 553667 506756 553723
rect 506756 553667 506812 553723
rect 506812 553667 506816 553723
rect 506752 553663 506816 553667
rect 506272 553643 506336 553647
rect 506272 553587 506276 553643
rect 506276 553587 506332 553643
rect 506332 553587 506336 553643
rect 506272 553583 506336 553587
rect 506352 553643 506416 553647
rect 506352 553587 506356 553643
rect 506356 553587 506412 553643
rect 506412 553587 506416 553643
rect 506352 553583 506416 553587
rect 506432 553643 506496 553647
rect 506432 553587 506436 553643
rect 506436 553587 506492 553643
rect 506492 553587 506496 553643
rect 506432 553583 506496 553587
rect 506512 553643 506576 553647
rect 506512 553587 506516 553643
rect 506516 553587 506572 553643
rect 506572 553587 506576 553643
rect 506512 553583 506576 553587
rect 506592 553643 506656 553647
rect 506592 553587 506596 553643
rect 506596 553587 506652 553643
rect 506652 553587 506656 553643
rect 506592 553583 506656 553587
rect 506672 553643 506736 553647
rect 506672 553587 506676 553643
rect 506676 553587 506732 553643
rect 506732 553587 506736 553643
rect 506672 553583 506736 553587
rect 506752 553643 506816 553647
rect 506752 553587 506756 553643
rect 506756 553587 506812 553643
rect 506812 553587 506816 553643
rect 506752 553583 506816 553587
rect 506272 553563 506336 553567
rect 506272 553507 506276 553563
rect 506276 553507 506332 553563
rect 506332 553507 506336 553563
rect 506272 553503 506336 553507
rect 506352 553563 506416 553567
rect 506352 553507 506356 553563
rect 506356 553507 506412 553563
rect 506412 553507 506416 553563
rect 506352 553503 506416 553507
rect 506432 553563 506496 553567
rect 506432 553507 506436 553563
rect 506436 553507 506492 553563
rect 506492 553507 506496 553563
rect 506432 553503 506496 553507
rect 506512 553563 506576 553567
rect 506512 553507 506516 553563
rect 506516 553507 506572 553563
rect 506572 553507 506576 553563
rect 506512 553503 506576 553507
rect 506592 553563 506656 553567
rect 506592 553507 506596 553563
rect 506596 553507 506652 553563
rect 506652 553507 506656 553563
rect 506592 553503 506656 553507
rect 506672 553563 506736 553567
rect 506672 553507 506676 553563
rect 506676 553507 506732 553563
rect 506732 553507 506736 553563
rect 506672 553503 506736 553507
rect 506752 553563 506816 553567
rect 506752 553507 506756 553563
rect 506756 553507 506812 553563
rect 506812 553507 506816 553563
rect 506752 553503 506816 553507
rect 577032 538514 577096 538518
rect 577032 538458 577036 538514
rect 577036 538458 577092 538514
rect 577092 538458 577096 538514
rect 577032 538454 577096 538458
rect 577112 538514 577176 538518
rect 577112 538458 577116 538514
rect 577116 538458 577172 538514
rect 577172 538458 577176 538514
rect 577112 538454 577176 538458
rect 577192 538514 577256 538518
rect 577192 538458 577196 538514
rect 577196 538458 577252 538514
rect 577252 538458 577256 538514
rect 577192 538454 577256 538458
rect 577272 538514 577336 538518
rect 577272 538458 577276 538514
rect 577276 538458 577332 538514
rect 577332 538458 577336 538514
rect 577272 538454 577336 538458
rect 577352 538514 577416 538518
rect 577352 538458 577356 538514
rect 577356 538458 577412 538514
rect 577412 538458 577416 538514
rect 577352 538454 577416 538458
rect 577432 538514 577496 538518
rect 577432 538458 577436 538514
rect 577436 538458 577492 538514
rect 577492 538458 577496 538514
rect 577432 538454 577496 538458
rect 577512 538514 577576 538518
rect 577512 538458 577516 538514
rect 577516 538458 577572 538514
rect 577572 538458 577576 538514
rect 577512 538454 577576 538458
rect 577032 538434 577096 538438
rect 577032 538378 577036 538434
rect 577036 538378 577092 538434
rect 577092 538378 577096 538434
rect 577032 538374 577096 538378
rect 577112 538434 577176 538438
rect 577112 538378 577116 538434
rect 577116 538378 577172 538434
rect 577172 538378 577176 538434
rect 577112 538374 577176 538378
rect 577192 538434 577256 538438
rect 577192 538378 577196 538434
rect 577196 538378 577252 538434
rect 577252 538378 577256 538434
rect 577192 538374 577256 538378
rect 577272 538434 577336 538438
rect 577272 538378 577276 538434
rect 577276 538378 577332 538434
rect 577332 538378 577336 538434
rect 577272 538374 577336 538378
rect 577352 538434 577416 538438
rect 577352 538378 577356 538434
rect 577356 538378 577412 538434
rect 577412 538378 577416 538434
rect 577352 538374 577416 538378
rect 577432 538434 577496 538438
rect 577432 538378 577436 538434
rect 577436 538378 577492 538434
rect 577492 538378 577496 538434
rect 577432 538374 577496 538378
rect 577512 538434 577576 538438
rect 577512 538378 577516 538434
rect 577516 538378 577572 538434
rect 577572 538378 577576 538434
rect 577512 538374 577576 538378
rect 577032 538354 577096 538358
rect 577032 538298 577036 538354
rect 577036 538298 577092 538354
rect 577092 538298 577096 538354
rect 577032 538294 577096 538298
rect 577112 538354 577176 538358
rect 577112 538298 577116 538354
rect 577116 538298 577172 538354
rect 577172 538298 577176 538354
rect 577112 538294 577176 538298
rect 577192 538354 577256 538358
rect 577192 538298 577196 538354
rect 577196 538298 577252 538354
rect 577252 538298 577256 538354
rect 577192 538294 577256 538298
rect 577272 538354 577336 538358
rect 577272 538298 577276 538354
rect 577276 538298 577332 538354
rect 577332 538298 577336 538354
rect 577272 538294 577336 538298
rect 577352 538354 577416 538358
rect 577352 538298 577356 538354
rect 577356 538298 577412 538354
rect 577412 538298 577416 538354
rect 577352 538294 577416 538298
rect 577432 538354 577496 538358
rect 577432 538298 577436 538354
rect 577436 538298 577492 538354
rect 577492 538298 577496 538354
rect 577432 538294 577496 538298
rect 577512 538354 577576 538358
rect 577512 538298 577516 538354
rect 577516 538298 577572 538354
rect 577572 538298 577576 538354
rect 577512 538294 577576 538298
rect 577032 538274 577096 538278
rect 577032 538218 577036 538274
rect 577036 538218 577092 538274
rect 577092 538218 577096 538274
rect 577032 538214 577096 538218
rect 577112 538274 577176 538278
rect 577112 538218 577116 538274
rect 577116 538218 577172 538274
rect 577172 538218 577176 538274
rect 577112 538214 577176 538218
rect 577192 538274 577256 538278
rect 577192 538218 577196 538274
rect 577196 538218 577252 538274
rect 577252 538218 577256 538274
rect 577192 538214 577256 538218
rect 577272 538274 577336 538278
rect 577272 538218 577276 538274
rect 577276 538218 577332 538274
rect 577332 538218 577336 538274
rect 577272 538214 577336 538218
rect 577352 538274 577416 538278
rect 577352 538218 577356 538274
rect 577356 538218 577412 538274
rect 577412 538218 577416 538274
rect 577352 538214 577416 538218
rect 577432 538274 577496 538278
rect 577432 538218 577436 538274
rect 577436 538218 577492 538274
rect 577492 538218 577496 538274
rect 577432 538214 577496 538218
rect 577512 538274 577576 538278
rect 577512 538218 577516 538274
rect 577516 538218 577572 538274
rect 577572 538218 577576 538274
rect 577512 538214 577576 538218
rect 578272 537719 578336 537723
rect 578272 537663 578276 537719
rect 578276 537663 578332 537719
rect 578332 537663 578336 537719
rect 578272 537659 578336 537663
rect 578352 537719 578416 537723
rect 578352 537663 578356 537719
rect 578356 537663 578412 537719
rect 578412 537663 578416 537719
rect 578352 537659 578416 537663
rect 578432 537719 578496 537723
rect 578432 537663 578436 537719
rect 578436 537663 578492 537719
rect 578492 537663 578496 537719
rect 578432 537659 578496 537663
rect 578512 537719 578576 537723
rect 578512 537663 578516 537719
rect 578516 537663 578572 537719
rect 578572 537663 578576 537719
rect 578512 537659 578576 537663
rect 578592 537719 578656 537723
rect 578592 537663 578596 537719
rect 578596 537663 578652 537719
rect 578652 537663 578656 537719
rect 578592 537659 578656 537663
rect 578672 537719 578736 537723
rect 578672 537663 578676 537719
rect 578676 537663 578732 537719
rect 578732 537663 578736 537719
rect 578672 537659 578736 537663
rect 578752 537719 578816 537723
rect 578752 537663 578756 537719
rect 578756 537663 578812 537719
rect 578812 537663 578816 537719
rect 578752 537659 578816 537663
rect 578272 537639 578336 537643
rect 578272 537583 578276 537639
rect 578276 537583 578332 537639
rect 578332 537583 578336 537639
rect 578272 537579 578336 537583
rect 578352 537639 578416 537643
rect 578352 537583 578356 537639
rect 578356 537583 578412 537639
rect 578412 537583 578416 537639
rect 578352 537579 578416 537583
rect 578432 537639 578496 537643
rect 578432 537583 578436 537639
rect 578436 537583 578492 537639
rect 578492 537583 578496 537639
rect 578432 537579 578496 537583
rect 578512 537639 578576 537643
rect 578512 537583 578516 537639
rect 578516 537583 578572 537639
rect 578572 537583 578576 537639
rect 578512 537579 578576 537583
rect 578592 537639 578656 537643
rect 578592 537583 578596 537639
rect 578596 537583 578652 537639
rect 578652 537583 578656 537639
rect 578592 537579 578656 537583
rect 578672 537639 578736 537643
rect 578672 537583 578676 537639
rect 578676 537583 578732 537639
rect 578732 537583 578736 537639
rect 578672 537579 578736 537583
rect 578752 537639 578816 537643
rect 578752 537583 578756 537639
rect 578756 537583 578812 537639
rect 578812 537583 578816 537639
rect 578752 537579 578816 537583
rect 578272 537559 578336 537563
rect 578272 537503 578276 537559
rect 578276 537503 578332 537559
rect 578332 537503 578336 537559
rect 578272 537499 578336 537503
rect 578352 537559 578416 537563
rect 578352 537503 578356 537559
rect 578356 537503 578412 537559
rect 578412 537503 578416 537559
rect 578352 537499 578416 537503
rect 578432 537559 578496 537563
rect 578432 537503 578436 537559
rect 578436 537503 578492 537559
rect 578492 537503 578496 537559
rect 578432 537499 578496 537503
rect 578512 537559 578576 537563
rect 578512 537503 578516 537559
rect 578516 537503 578572 537559
rect 578572 537503 578576 537559
rect 578512 537499 578576 537503
rect 578592 537559 578656 537563
rect 578592 537503 578596 537559
rect 578596 537503 578652 537559
rect 578652 537503 578656 537559
rect 578592 537499 578656 537503
rect 578672 537559 578736 537563
rect 578672 537503 578676 537559
rect 578676 537503 578732 537559
rect 578732 537503 578736 537559
rect 578672 537499 578736 537503
rect 578752 537559 578816 537563
rect 578752 537503 578756 537559
rect 578756 537503 578812 537559
rect 578812 537503 578816 537559
rect 578752 537499 578816 537503
rect 578272 537479 578336 537483
rect 578272 537423 578276 537479
rect 578276 537423 578332 537479
rect 578332 537423 578336 537479
rect 578272 537419 578336 537423
rect 578352 537479 578416 537483
rect 578352 537423 578356 537479
rect 578356 537423 578412 537479
rect 578412 537423 578416 537479
rect 578352 537419 578416 537423
rect 578432 537479 578496 537483
rect 578432 537423 578436 537479
rect 578436 537423 578492 537479
rect 578492 537423 578496 537479
rect 578432 537419 578496 537423
rect 578512 537479 578576 537483
rect 578512 537423 578516 537479
rect 578516 537423 578572 537479
rect 578572 537423 578576 537479
rect 578512 537419 578576 537423
rect 578592 537479 578656 537483
rect 578592 537423 578596 537479
rect 578596 537423 578652 537479
rect 578652 537423 578656 537479
rect 578592 537419 578656 537423
rect 578672 537479 578736 537483
rect 578672 537423 578676 537479
rect 578676 537423 578732 537479
rect 578732 537423 578736 537479
rect 578672 537419 578736 537423
rect 578752 537479 578816 537483
rect 578752 537423 578756 537479
rect 578756 537423 578812 537479
rect 578812 537423 578816 537479
rect 578752 537419 578816 537423
rect 577032 485338 577096 485342
rect 577032 485282 577036 485338
rect 577036 485282 577092 485338
rect 577092 485282 577096 485338
rect 577032 485278 577096 485282
rect 577112 485338 577176 485342
rect 577112 485282 577116 485338
rect 577116 485282 577172 485338
rect 577172 485282 577176 485338
rect 577112 485278 577176 485282
rect 577192 485338 577256 485342
rect 577192 485282 577196 485338
rect 577196 485282 577252 485338
rect 577252 485282 577256 485338
rect 577192 485278 577256 485282
rect 577272 485338 577336 485342
rect 577272 485282 577276 485338
rect 577276 485282 577332 485338
rect 577332 485282 577336 485338
rect 577272 485278 577336 485282
rect 577352 485338 577416 485342
rect 577352 485282 577356 485338
rect 577356 485282 577412 485338
rect 577412 485282 577416 485338
rect 577352 485278 577416 485282
rect 577432 485338 577496 485342
rect 577432 485282 577436 485338
rect 577436 485282 577492 485338
rect 577492 485282 577496 485338
rect 577432 485278 577496 485282
rect 577512 485338 577576 485342
rect 577512 485282 577516 485338
rect 577516 485282 577572 485338
rect 577572 485282 577576 485338
rect 577512 485278 577576 485282
rect 577032 485258 577096 485262
rect 577032 485202 577036 485258
rect 577036 485202 577092 485258
rect 577092 485202 577096 485258
rect 577032 485198 577096 485202
rect 577112 485258 577176 485262
rect 577112 485202 577116 485258
rect 577116 485202 577172 485258
rect 577172 485202 577176 485258
rect 577112 485198 577176 485202
rect 577192 485258 577256 485262
rect 577192 485202 577196 485258
rect 577196 485202 577252 485258
rect 577252 485202 577256 485258
rect 577192 485198 577256 485202
rect 577272 485258 577336 485262
rect 577272 485202 577276 485258
rect 577276 485202 577332 485258
rect 577332 485202 577336 485258
rect 577272 485198 577336 485202
rect 577352 485258 577416 485262
rect 577352 485202 577356 485258
rect 577356 485202 577412 485258
rect 577412 485202 577416 485258
rect 577352 485198 577416 485202
rect 577432 485258 577496 485262
rect 577432 485202 577436 485258
rect 577436 485202 577492 485258
rect 577492 485202 577496 485258
rect 577432 485198 577496 485202
rect 577512 485258 577576 485262
rect 577512 485202 577516 485258
rect 577516 485202 577572 485258
rect 577572 485202 577576 485258
rect 577512 485198 577576 485202
rect 577032 485178 577096 485182
rect 577032 485122 577036 485178
rect 577036 485122 577092 485178
rect 577092 485122 577096 485178
rect 577032 485118 577096 485122
rect 577112 485178 577176 485182
rect 577112 485122 577116 485178
rect 577116 485122 577172 485178
rect 577172 485122 577176 485178
rect 577112 485118 577176 485122
rect 577192 485178 577256 485182
rect 577192 485122 577196 485178
rect 577196 485122 577252 485178
rect 577252 485122 577256 485178
rect 577192 485118 577256 485122
rect 577272 485178 577336 485182
rect 577272 485122 577276 485178
rect 577276 485122 577332 485178
rect 577332 485122 577336 485178
rect 577272 485118 577336 485122
rect 577352 485178 577416 485182
rect 577352 485122 577356 485178
rect 577356 485122 577412 485178
rect 577412 485122 577416 485178
rect 577352 485118 577416 485122
rect 577432 485178 577496 485182
rect 577432 485122 577436 485178
rect 577436 485122 577492 485178
rect 577492 485122 577496 485178
rect 577432 485118 577496 485122
rect 577512 485178 577576 485182
rect 577512 485122 577516 485178
rect 577516 485122 577572 485178
rect 577572 485122 577576 485178
rect 577512 485118 577576 485122
rect 577032 485098 577096 485102
rect 577032 485042 577036 485098
rect 577036 485042 577092 485098
rect 577092 485042 577096 485098
rect 577032 485038 577096 485042
rect 577112 485098 577176 485102
rect 577112 485042 577116 485098
rect 577116 485042 577172 485098
rect 577172 485042 577176 485098
rect 577112 485038 577176 485042
rect 577192 485098 577256 485102
rect 577192 485042 577196 485098
rect 577196 485042 577252 485098
rect 577252 485042 577256 485098
rect 577192 485038 577256 485042
rect 577272 485098 577336 485102
rect 577272 485042 577276 485098
rect 577276 485042 577332 485098
rect 577332 485042 577336 485098
rect 577272 485038 577336 485042
rect 577352 485098 577416 485102
rect 577352 485042 577356 485098
rect 577356 485042 577412 485098
rect 577412 485042 577416 485098
rect 577352 485038 577416 485042
rect 577432 485098 577496 485102
rect 577432 485042 577436 485098
rect 577436 485042 577492 485098
rect 577492 485042 577496 485098
rect 577432 485038 577496 485042
rect 577512 485098 577576 485102
rect 577512 485042 577516 485098
rect 577516 485042 577572 485098
rect 577572 485042 577576 485098
rect 577512 485038 577576 485042
rect 578272 484543 578336 484547
rect 578272 484487 578276 484543
rect 578276 484487 578332 484543
rect 578332 484487 578336 484543
rect 578272 484483 578336 484487
rect 578352 484543 578416 484547
rect 578352 484487 578356 484543
rect 578356 484487 578412 484543
rect 578412 484487 578416 484543
rect 578352 484483 578416 484487
rect 578432 484543 578496 484547
rect 578432 484487 578436 484543
rect 578436 484487 578492 484543
rect 578492 484487 578496 484543
rect 578432 484483 578496 484487
rect 578512 484543 578576 484547
rect 578512 484487 578516 484543
rect 578516 484487 578572 484543
rect 578572 484487 578576 484543
rect 578512 484483 578576 484487
rect 578592 484543 578656 484547
rect 578592 484487 578596 484543
rect 578596 484487 578652 484543
rect 578652 484487 578656 484543
rect 578592 484483 578656 484487
rect 578672 484543 578736 484547
rect 578672 484487 578676 484543
rect 578676 484487 578732 484543
rect 578732 484487 578736 484543
rect 578672 484483 578736 484487
rect 578752 484543 578816 484547
rect 578752 484487 578756 484543
rect 578756 484487 578812 484543
rect 578812 484487 578816 484543
rect 578752 484483 578816 484487
rect 578272 484463 578336 484467
rect 578272 484407 578276 484463
rect 578276 484407 578332 484463
rect 578332 484407 578336 484463
rect 578272 484403 578336 484407
rect 578352 484463 578416 484467
rect 578352 484407 578356 484463
rect 578356 484407 578412 484463
rect 578412 484407 578416 484463
rect 578352 484403 578416 484407
rect 578432 484463 578496 484467
rect 578432 484407 578436 484463
rect 578436 484407 578492 484463
rect 578492 484407 578496 484463
rect 578432 484403 578496 484407
rect 578512 484463 578576 484467
rect 578512 484407 578516 484463
rect 578516 484407 578572 484463
rect 578572 484407 578576 484463
rect 578512 484403 578576 484407
rect 578592 484463 578656 484467
rect 578592 484407 578596 484463
rect 578596 484407 578652 484463
rect 578652 484407 578656 484463
rect 578592 484403 578656 484407
rect 578672 484463 578736 484467
rect 578672 484407 578676 484463
rect 578676 484407 578732 484463
rect 578732 484407 578736 484463
rect 578672 484403 578736 484407
rect 578752 484463 578816 484467
rect 578752 484407 578756 484463
rect 578756 484407 578812 484463
rect 578812 484407 578816 484463
rect 578752 484403 578816 484407
rect 578272 484383 578336 484387
rect 578272 484327 578276 484383
rect 578276 484327 578332 484383
rect 578332 484327 578336 484383
rect 578272 484323 578336 484327
rect 578352 484383 578416 484387
rect 578352 484327 578356 484383
rect 578356 484327 578412 484383
rect 578412 484327 578416 484383
rect 578352 484323 578416 484327
rect 578432 484383 578496 484387
rect 578432 484327 578436 484383
rect 578436 484327 578492 484383
rect 578492 484327 578496 484383
rect 578432 484323 578496 484327
rect 578512 484383 578576 484387
rect 578512 484327 578516 484383
rect 578516 484327 578572 484383
rect 578572 484327 578576 484383
rect 578512 484323 578576 484327
rect 578592 484383 578656 484387
rect 578592 484327 578596 484383
rect 578596 484327 578652 484383
rect 578652 484327 578656 484383
rect 578592 484323 578656 484327
rect 578672 484383 578736 484387
rect 578672 484327 578676 484383
rect 578676 484327 578732 484383
rect 578732 484327 578736 484383
rect 578672 484323 578736 484327
rect 578752 484383 578816 484387
rect 578752 484327 578756 484383
rect 578756 484327 578812 484383
rect 578812 484327 578816 484383
rect 578752 484323 578816 484327
rect 578272 484303 578336 484307
rect 578272 484247 578276 484303
rect 578276 484247 578332 484303
rect 578332 484247 578336 484303
rect 578272 484243 578336 484247
rect 578352 484303 578416 484307
rect 578352 484247 578356 484303
rect 578356 484247 578412 484303
rect 578412 484247 578416 484303
rect 578352 484243 578416 484247
rect 578432 484303 578496 484307
rect 578432 484247 578436 484303
rect 578436 484247 578492 484303
rect 578492 484247 578496 484303
rect 578432 484243 578496 484247
rect 578512 484303 578576 484307
rect 578512 484247 578516 484303
rect 578516 484247 578572 484303
rect 578572 484247 578576 484303
rect 578512 484243 578576 484247
rect 578592 484303 578656 484307
rect 578592 484247 578596 484303
rect 578596 484247 578652 484303
rect 578652 484247 578656 484303
rect 578592 484243 578656 484247
rect 578672 484303 578736 484307
rect 578672 484247 578676 484303
rect 578676 484247 578732 484303
rect 578732 484247 578736 484303
rect 578672 484243 578736 484247
rect 578752 484303 578816 484307
rect 578752 484247 578756 484303
rect 578756 484247 578812 484303
rect 578812 484247 578816 484303
rect 578752 484243 578816 484247
rect 470272 451481 470336 451485
rect 470272 451425 470276 451481
rect 470276 451425 470332 451481
rect 470332 451425 470336 451481
rect 470272 451421 470336 451425
rect 470352 451481 470416 451485
rect 470352 451425 470356 451481
rect 470356 451425 470412 451481
rect 470412 451425 470416 451481
rect 470352 451421 470416 451425
rect 470432 451481 470496 451485
rect 470432 451425 470436 451481
rect 470436 451425 470492 451481
rect 470492 451425 470496 451481
rect 470432 451421 470496 451425
rect 470512 451481 470576 451485
rect 470512 451425 470516 451481
rect 470516 451425 470572 451481
rect 470572 451425 470576 451481
rect 470512 451421 470576 451425
rect 470592 451481 470656 451485
rect 470592 451425 470596 451481
rect 470596 451425 470652 451481
rect 470652 451425 470656 451481
rect 470592 451421 470656 451425
rect 470672 451481 470736 451485
rect 470672 451425 470676 451481
rect 470676 451425 470732 451481
rect 470732 451425 470736 451481
rect 470672 451421 470736 451425
rect 470752 451481 470816 451485
rect 470752 451425 470756 451481
rect 470756 451425 470812 451481
rect 470812 451425 470816 451481
rect 470752 451421 470816 451425
rect 470272 451401 470336 451405
rect 470272 451345 470276 451401
rect 470276 451345 470332 451401
rect 470332 451345 470336 451401
rect 470272 451341 470336 451345
rect 470352 451401 470416 451405
rect 470352 451345 470356 451401
rect 470356 451345 470412 451401
rect 470412 451345 470416 451401
rect 470352 451341 470416 451345
rect 470432 451401 470496 451405
rect 470432 451345 470436 451401
rect 470436 451345 470492 451401
rect 470492 451345 470496 451401
rect 470432 451341 470496 451345
rect 470512 451401 470576 451405
rect 470512 451345 470516 451401
rect 470516 451345 470572 451401
rect 470572 451345 470576 451401
rect 470512 451341 470576 451345
rect 470592 451401 470656 451405
rect 470592 451345 470596 451401
rect 470596 451345 470652 451401
rect 470652 451345 470656 451401
rect 470592 451341 470656 451345
rect 470672 451401 470736 451405
rect 470672 451345 470676 451401
rect 470676 451345 470732 451401
rect 470732 451345 470736 451401
rect 470672 451341 470736 451345
rect 470752 451401 470816 451405
rect 470752 451345 470756 451401
rect 470756 451345 470812 451401
rect 470812 451345 470816 451401
rect 470752 451341 470816 451345
rect 470272 451321 470336 451325
rect 470272 451265 470276 451321
rect 470276 451265 470332 451321
rect 470332 451265 470336 451321
rect 470272 451261 470336 451265
rect 470352 451321 470416 451325
rect 470352 451265 470356 451321
rect 470356 451265 470412 451321
rect 470412 451265 470416 451321
rect 470352 451261 470416 451265
rect 470432 451321 470496 451325
rect 470432 451265 470436 451321
rect 470436 451265 470492 451321
rect 470492 451265 470496 451321
rect 470432 451261 470496 451265
rect 470512 451321 470576 451325
rect 470512 451265 470516 451321
rect 470516 451265 470572 451321
rect 470572 451265 470576 451321
rect 470512 451261 470576 451265
rect 470592 451321 470656 451325
rect 470592 451265 470596 451321
rect 470596 451265 470652 451321
rect 470652 451265 470656 451321
rect 470592 451261 470656 451265
rect 470672 451321 470736 451325
rect 470672 451265 470676 451321
rect 470676 451265 470732 451321
rect 470732 451265 470736 451321
rect 470672 451261 470736 451265
rect 470752 451321 470816 451325
rect 470752 451265 470756 451321
rect 470756 451265 470812 451321
rect 470812 451265 470816 451321
rect 470752 451261 470816 451265
rect 470272 451241 470336 451245
rect 470272 451185 470276 451241
rect 470276 451185 470332 451241
rect 470332 451185 470336 451241
rect 470272 451181 470336 451185
rect 470352 451241 470416 451245
rect 470352 451185 470356 451241
rect 470356 451185 470412 451241
rect 470412 451185 470416 451241
rect 470352 451181 470416 451185
rect 470432 451241 470496 451245
rect 470432 451185 470436 451241
rect 470436 451185 470492 451241
rect 470492 451185 470496 451241
rect 470432 451181 470496 451185
rect 470512 451241 470576 451245
rect 470512 451185 470516 451241
rect 470516 451185 470572 451241
rect 470572 451185 470576 451241
rect 470512 451181 470576 451185
rect 470592 451241 470656 451245
rect 470592 451185 470596 451241
rect 470596 451185 470652 451241
rect 470652 451185 470656 451241
rect 470592 451181 470656 451185
rect 470672 451241 470736 451245
rect 470672 451185 470676 451241
rect 470676 451185 470732 451241
rect 470732 451185 470736 451241
rect 470672 451181 470736 451185
rect 470752 451241 470816 451245
rect 470752 451185 470756 451241
rect 470756 451185 470812 451241
rect 470812 451185 470816 451241
rect 470752 451181 470816 451185
rect 469032 450395 469096 450399
rect 469032 450339 469036 450395
rect 469036 450339 469092 450395
rect 469092 450339 469096 450395
rect 469032 450335 469096 450339
rect 469112 450395 469176 450399
rect 469112 450339 469116 450395
rect 469116 450339 469172 450395
rect 469172 450339 469176 450395
rect 469112 450335 469176 450339
rect 469192 450395 469256 450399
rect 469192 450339 469196 450395
rect 469196 450339 469252 450395
rect 469252 450339 469256 450395
rect 469192 450335 469256 450339
rect 469272 450395 469336 450399
rect 469272 450339 469276 450395
rect 469276 450339 469332 450395
rect 469332 450339 469336 450395
rect 469272 450335 469336 450339
rect 469352 450395 469416 450399
rect 469352 450339 469356 450395
rect 469356 450339 469412 450395
rect 469412 450339 469416 450395
rect 469352 450335 469416 450339
rect 469432 450395 469496 450399
rect 469432 450339 469436 450395
rect 469436 450339 469492 450395
rect 469492 450339 469496 450395
rect 469432 450335 469496 450339
rect 469512 450395 469576 450399
rect 469512 450339 469516 450395
rect 469516 450339 469572 450395
rect 469572 450339 469576 450395
rect 469512 450335 469576 450339
rect 469032 450315 469096 450319
rect 469032 450259 469036 450315
rect 469036 450259 469092 450315
rect 469092 450259 469096 450315
rect 469032 450255 469096 450259
rect 469112 450315 469176 450319
rect 469112 450259 469116 450315
rect 469116 450259 469172 450315
rect 469172 450259 469176 450315
rect 469112 450255 469176 450259
rect 469192 450315 469256 450319
rect 469192 450259 469196 450315
rect 469196 450259 469252 450315
rect 469252 450259 469256 450315
rect 469192 450255 469256 450259
rect 469272 450315 469336 450319
rect 469272 450259 469276 450315
rect 469276 450259 469332 450315
rect 469332 450259 469336 450315
rect 469272 450255 469336 450259
rect 469352 450315 469416 450319
rect 469352 450259 469356 450315
rect 469356 450259 469412 450315
rect 469412 450259 469416 450315
rect 469352 450255 469416 450259
rect 469432 450315 469496 450319
rect 469432 450259 469436 450315
rect 469436 450259 469492 450315
rect 469492 450259 469496 450315
rect 469432 450255 469496 450259
rect 469512 450315 469576 450319
rect 469512 450259 469516 450315
rect 469516 450259 469572 450315
rect 469572 450259 469576 450315
rect 469512 450255 469576 450259
rect 469032 450235 469096 450239
rect 469032 450179 469036 450235
rect 469036 450179 469092 450235
rect 469092 450179 469096 450235
rect 469032 450175 469096 450179
rect 469112 450235 469176 450239
rect 469112 450179 469116 450235
rect 469116 450179 469172 450235
rect 469172 450179 469176 450235
rect 469112 450175 469176 450179
rect 469192 450235 469256 450239
rect 469192 450179 469196 450235
rect 469196 450179 469252 450235
rect 469252 450179 469256 450235
rect 469192 450175 469256 450179
rect 469272 450235 469336 450239
rect 469272 450179 469276 450235
rect 469276 450179 469332 450235
rect 469332 450179 469336 450235
rect 469272 450175 469336 450179
rect 469352 450235 469416 450239
rect 469352 450179 469356 450235
rect 469356 450179 469412 450235
rect 469412 450179 469416 450235
rect 469352 450175 469416 450179
rect 469432 450235 469496 450239
rect 469432 450179 469436 450235
rect 469436 450179 469492 450235
rect 469492 450179 469496 450235
rect 469432 450175 469496 450179
rect 469512 450235 469576 450239
rect 469512 450179 469516 450235
rect 469516 450179 469572 450235
rect 469572 450179 469576 450235
rect 469512 450175 469576 450179
rect 478460 450198 478524 450262
rect 481220 450198 481284 450262
rect 487844 450258 487908 450262
rect 487844 450202 487849 450258
rect 487849 450202 487908 450258
rect 487844 450198 487908 450202
rect 469032 450155 469096 450159
rect 469032 450099 469036 450155
rect 469036 450099 469092 450155
rect 469092 450099 469096 450155
rect 469032 450095 469096 450099
rect 469112 450155 469176 450159
rect 469112 450099 469116 450155
rect 469116 450099 469172 450155
rect 469172 450099 469176 450155
rect 469112 450095 469176 450099
rect 469192 450155 469256 450159
rect 469192 450099 469196 450155
rect 469196 450099 469252 450155
rect 469252 450099 469256 450155
rect 469192 450095 469256 450099
rect 469272 450155 469336 450159
rect 469272 450099 469276 450155
rect 469276 450099 469332 450155
rect 469332 450099 469336 450155
rect 469272 450095 469336 450099
rect 469352 450155 469416 450159
rect 469352 450099 469356 450155
rect 469356 450099 469412 450155
rect 469412 450099 469416 450155
rect 469352 450095 469416 450099
rect 469432 450155 469496 450159
rect 469432 450099 469436 450155
rect 469436 450099 469492 450155
rect 469492 450099 469496 450155
rect 469432 450095 469496 450099
rect 469512 450155 469576 450159
rect 469512 450099 469516 450155
rect 469516 450099 469572 450155
rect 469572 450099 469576 450155
rect 469512 450095 469576 450099
rect 473676 449654 473740 449718
rect 470272 449310 470336 449314
rect 470272 449254 470276 449310
rect 470276 449254 470332 449310
rect 470332 449254 470336 449310
rect 470272 449250 470336 449254
rect 470352 449310 470416 449314
rect 470352 449254 470356 449310
rect 470356 449254 470412 449310
rect 470412 449254 470416 449310
rect 470352 449250 470416 449254
rect 470432 449310 470496 449314
rect 470432 449254 470436 449310
rect 470436 449254 470492 449310
rect 470492 449254 470496 449310
rect 470432 449250 470496 449254
rect 470512 449310 470576 449314
rect 470512 449254 470516 449310
rect 470516 449254 470572 449310
rect 470572 449254 470576 449310
rect 470512 449250 470576 449254
rect 470592 449310 470656 449314
rect 470592 449254 470596 449310
rect 470596 449254 470652 449310
rect 470652 449254 470656 449310
rect 470592 449250 470656 449254
rect 470672 449310 470736 449314
rect 470672 449254 470676 449310
rect 470676 449254 470732 449310
rect 470732 449254 470736 449310
rect 470672 449250 470736 449254
rect 470752 449310 470816 449314
rect 470752 449254 470756 449310
rect 470756 449254 470812 449310
rect 470812 449254 470816 449310
rect 470752 449250 470816 449254
rect 470272 449230 470336 449234
rect 470272 449174 470276 449230
rect 470276 449174 470332 449230
rect 470332 449174 470336 449230
rect 470272 449170 470336 449174
rect 470352 449230 470416 449234
rect 470352 449174 470356 449230
rect 470356 449174 470412 449230
rect 470412 449174 470416 449230
rect 470352 449170 470416 449174
rect 470432 449230 470496 449234
rect 470432 449174 470436 449230
rect 470436 449174 470492 449230
rect 470492 449174 470496 449230
rect 470432 449170 470496 449174
rect 470512 449230 470576 449234
rect 470512 449174 470516 449230
rect 470516 449174 470572 449230
rect 470572 449174 470576 449230
rect 470512 449170 470576 449174
rect 470592 449230 470656 449234
rect 470592 449174 470596 449230
rect 470596 449174 470652 449230
rect 470652 449174 470656 449230
rect 470592 449170 470656 449174
rect 470672 449230 470736 449234
rect 470672 449174 470676 449230
rect 470676 449174 470732 449230
rect 470732 449174 470736 449230
rect 470672 449170 470736 449174
rect 470752 449230 470816 449234
rect 470752 449174 470756 449230
rect 470756 449174 470812 449230
rect 470812 449174 470816 449230
rect 470752 449170 470816 449174
rect 470272 449150 470336 449154
rect 470272 449094 470276 449150
rect 470276 449094 470332 449150
rect 470332 449094 470336 449150
rect 470272 449090 470336 449094
rect 470352 449150 470416 449154
rect 470352 449094 470356 449150
rect 470356 449094 470412 449150
rect 470412 449094 470416 449150
rect 470352 449090 470416 449094
rect 470432 449150 470496 449154
rect 470432 449094 470436 449150
rect 470436 449094 470492 449150
rect 470492 449094 470496 449150
rect 470432 449090 470496 449094
rect 470512 449150 470576 449154
rect 470512 449094 470516 449150
rect 470516 449094 470572 449150
rect 470572 449094 470576 449150
rect 470512 449090 470576 449094
rect 470592 449150 470656 449154
rect 470592 449094 470596 449150
rect 470596 449094 470652 449150
rect 470652 449094 470656 449150
rect 470592 449090 470656 449094
rect 470672 449150 470736 449154
rect 470672 449094 470676 449150
rect 470676 449094 470732 449150
rect 470732 449094 470736 449150
rect 470672 449090 470736 449094
rect 470752 449150 470816 449154
rect 470752 449094 470756 449150
rect 470756 449094 470812 449150
rect 470812 449094 470816 449150
rect 470752 449090 470816 449094
rect 470272 449070 470336 449074
rect 470272 449014 470276 449070
rect 470276 449014 470332 449070
rect 470332 449014 470336 449070
rect 470272 449010 470336 449014
rect 470352 449070 470416 449074
rect 470352 449014 470356 449070
rect 470356 449014 470412 449070
rect 470412 449014 470416 449070
rect 470352 449010 470416 449014
rect 470432 449070 470496 449074
rect 470432 449014 470436 449070
rect 470436 449014 470492 449070
rect 470492 449014 470496 449070
rect 470432 449010 470496 449014
rect 470512 449070 470576 449074
rect 470512 449014 470516 449070
rect 470516 449014 470572 449070
rect 470572 449014 470576 449070
rect 470512 449010 470576 449014
rect 470592 449070 470656 449074
rect 470592 449014 470596 449070
rect 470596 449014 470652 449070
rect 470652 449014 470656 449070
rect 470592 449010 470656 449014
rect 470672 449070 470736 449074
rect 470672 449014 470676 449070
rect 470676 449014 470732 449070
rect 470732 449014 470736 449070
rect 470672 449010 470736 449014
rect 470752 449070 470816 449074
rect 470752 449014 470756 449070
rect 470756 449014 470812 449070
rect 470812 449014 470816 449070
rect 470752 449010 470816 449014
rect 544332 445710 544396 445774
rect 541572 445302 541636 445366
rect 470272 433082 470336 433086
rect 470272 433026 470276 433082
rect 470276 433026 470332 433082
rect 470332 433026 470336 433082
rect 470272 433022 470336 433026
rect 470352 433082 470416 433086
rect 470352 433026 470356 433082
rect 470356 433026 470412 433082
rect 470412 433026 470416 433082
rect 470352 433022 470416 433026
rect 470432 433082 470496 433086
rect 470432 433026 470436 433082
rect 470436 433026 470492 433082
rect 470492 433026 470496 433082
rect 470432 433022 470496 433026
rect 470512 433082 470576 433086
rect 470512 433026 470516 433082
rect 470516 433026 470572 433082
rect 470572 433026 470576 433082
rect 470512 433022 470576 433026
rect 470592 433082 470656 433086
rect 470592 433026 470596 433082
rect 470596 433026 470652 433082
rect 470652 433026 470656 433082
rect 470592 433022 470656 433026
rect 470672 433082 470736 433086
rect 470672 433026 470676 433082
rect 470676 433026 470732 433082
rect 470732 433026 470736 433082
rect 470672 433022 470736 433026
rect 470752 433082 470816 433086
rect 470752 433026 470756 433082
rect 470756 433026 470812 433082
rect 470812 433026 470816 433082
rect 470752 433022 470816 433026
rect 470272 433002 470336 433006
rect 470272 432946 470276 433002
rect 470276 432946 470332 433002
rect 470332 432946 470336 433002
rect 470272 432942 470336 432946
rect 470352 433002 470416 433006
rect 470352 432946 470356 433002
rect 470356 432946 470412 433002
rect 470412 432946 470416 433002
rect 470352 432942 470416 432946
rect 470432 433002 470496 433006
rect 470432 432946 470436 433002
rect 470436 432946 470492 433002
rect 470492 432946 470496 433002
rect 470432 432942 470496 432946
rect 470512 433002 470576 433006
rect 470512 432946 470516 433002
rect 470516 432946 470572 433002
rect 470572 432946 470576 433002
rect 470512 432942 470576 432946
rect 470592 433002 470656 433006
rect 470592 432946 470596 433002
rect 470596 432946 470652 433002
rect 470652 432946 470656 433002
rect 470592 432942 470656 432946
rect 470672 433002 470736 433006
rect 470672 432946 470676 433002
rect 470676 432946 470732 433002
rect 470732 432946 470736 433002
rect 470672 432942 470736 432946
rect 470752 433002 470816 433006
rect 470752 432946 470756 433002
rect 470756 432946 470812 433002
rect 470812 432946 470816 433002
rect 470752 432942 470816 432946
rect 470272 432922 470336 432926
rect 470272 432866 470276 432922
rect 470276 432866 470332 432922
rect 470332 432866 470336 432922
rect 470272 432862 470336 432866
rect 470352 432922 470416 432926
rect 470352 432866 470356 432922
rect 470356 432866 470412 432922
rect 470412 432866 470416 432922
rect 470352 432862 470416 432866
rect 470432 432922 470496 432926
rect 470432 432866 470436 432922
rect 470436 432866 470492 432922
rect 470492 432866 470496 432922
rect 470432 432862 470496 432866
rect 470512 432922 470576 432926
rect 470512 432866 470516 432922
rect 470516 432866 470572 432922
rect 470572 432866 470576 432922
rect 470512 432862 470576 432866
rect 470592 432922 470656 432926
rect 470592 432866 470596 432922
rect 470596 432866 470652 432922
rect 470652 432866 470656 432922
rect 470592 432862 470656 432866
rect 470672 432922 470736 432926
rect 470672 432866 470676 432922
rect 470676 432866 470732 432922
rect 470732 432866 470736 432922
rect 470672 432862 470736 432866
rect 470752 432922 470816 432926
rect 470752 432866 470756 432922
rect 470756 432866 470812 432922
rect 470812 432866 470816 432922
rect 470752 432862 470816 432866
rect 470272 432842 470336 432846
rect 470272 432786 470276 432842
rect 470276 432786 470332 432842
rect 470332 432786 470336 432842
rect 470272 432782 470336 432786
rect 470352 432842 470416 432846
rect 470352 432786 470356 432842
rect 470356 432786 470412 432842
rect 470412 432786 470416 432842
rect 470352 432782 470416 432786
rect 470432 432842 470496 432846
rect 470432 432786 470436 432842
rect 470436 432786 470492 432842
rect 470492 432786 470496 432842
rect 470432 432782 470496 432786
rect 470512 432842 470576 432846
rect 470512 432786 470516 432842
rect 470516 432786 470572 432842
rect 470572 432786 470576 432842
rect 470512 432782 470576 432786
rect 470592 432842 470656 432846
rect 470592 432786 470596 432842
rect 470596 432786 470652 432842
rect 470652 432786 470656 432842
rect 470592 432782 470656 432786
rect 470672 432842 470736 432846
rect 470672 432786 470676 432842
rect 470676 432786 470732 432842
rect 470732 432786 470736 432842
rect 470672 432782 470736 432786
rect 470752 432842 470816 432846
rect 470752 432786 470756 432842
rect 470756 432786 470812 432842
rect 470812 432786 470816 432842
rect 470752 432782 470816 432786
rect 483612 432850 483676 432854
rect 483612 432794 483662 432850
rect 483662 432794 483676 432850
rect 483612 432790 483676 432794
rect 483612 432306 483676 432310
rect 483612 432250 483626 432306
rect 483626 432250 483676 432306
rect 483612 432246 483676 432250
rect 577032 432298 577096 432302
rect 577032 432242 577036 432298
rect 577036 432242 577092 432298
rect 577092 432242 577096 432298
rect 577032 432238 577096 432242
rect 577112 432298 577176 432302
rect 577112 432242 577116 432298
rect 577116 432242 577172 432298
rect 577172 432242 577176 432298
rect 577112 432238 577176 432242
rect 577192 432298 577256 432302
rect 577192 432242 577196 432298
rect 577196 432242 577252 432298
rect 577252 432242 577256 432298
rect 577192 432238 577256 432242
rect 577272 432298 577336 432302
rect 577272 432242 577276 432298
rect 577276 432242 577332 432298
rect 577332 432242 577336 432298
rect 577272 432238 577336 432242
rect 577352 432298 577416 432302
rect 577352 432242 577356 432298
rect 577356 432242 577412 432298
rect 577412 432242 577416 432298
rect 577352 432238 577416 432242
rect 577432 432298 577496 432302
rect 577432 432242 577436 432298
rect 577436 432242 577492 432298
rect 577492 432242 577496 432298
rect 577432 432238 577496 432242
rect 577512 432298 577576 432302
rect 577512 432242 577516 432298
rect 577516 432242 577572 432298
rect 577572 432242 577576 432298
rect 577512 432238 577576 432242
rect 481220 432170 481284 432174
rect 481220 432114 481270 432170
rect 481270 432114 481284 432170
rect 481220 432110 481284 432114
rect 577032 432218 577096 432222
rect 577032 432162 577036 432218
rect 577036 432162 577092 432218
rect 577092 432162 577096 432218
rect 577032 432158 577096 432162
rect 577112 432218 577176 432222
rect 577112 432162 577116 432218
rect 577116 432162 577172 432218
rect 577172 432162 577176 432218
rect 577112 432158 577176 432162
rect 577192 432218 577256 432222
rect 577192 432162 577196 432218
rect 577196 432162 577252 432218
rect 577252 432162 577256 432218
rect 577192 432158 577256 432162
rect 577272 432218 577336 432222
rect 577272 432162 577276 432218
rect 577276 432162 577332 432218
rect 577332 432162 577336 432218
rect 577272 432158 577336 432162
rect 577352 432218 577416 432222
rect 577352 432162 577356 432218
rect 577356 432162 577412 432218
rect 577412 432162 577416 432218
rect 577352 432158 577416 432162
rect 577432 432218 577496 432222
rect 577432 432162 577436 432218
rect 577436 432162 577492 432218
rect 577492 432162 577496 432218
rect 577432 432158 577496 432162
rect 577512 432218 577576 432222
rect 577512 432162 577516 432218
rect 577516 432162 577572 432218
rect 577572 432162 577576 432218
rect 577512 432158 577576 432162
rect 577032 432138 577096 432142
rect 577032 432082 577036 432138
rect 577036 432082 577092 432138
rect 577092 432082 577096 432138
rect 577032 432078 577096 432082
rect 577112 432138 577176 432142
rect 577112 432082 577116 432138
rect 577116 432082 577172 432138
rect 577172 432082 577176 432138
rect 577112 432078 577176 432082
rect 577192 432138 577256 432142
rect 577192 432082 577196 432138
rect 577196 432082 577252 432138
rect 577252 432082 577256 432138
rect 577192 432078 577256 432082
rect 577272 432138 577336 432142
rect 577272 432082 577276 432138
rect 577276 432082 577332 432138
rect 577332 432082 577336 432138
rect 577272 432078 577336 432082
rect 577352 432138 577416 432142
rect 577352 432082 577356 432138
rect 577356 432082 577412 432138
rect 577412 432082 577416 432138
rect 577352 432078 577416 432082
rect 577432 432138 577496 432142
rect 577432 432082 577436 432138
rect 577436 432082 577492 432138
rect 577492 432082 577496 432138
rect 577432 432078 577496 432082
rect 577512 432138 577576 432142
rect 577512 432082 577516 432138
rect 577516 432082 577572 432138
rect 577572 432082 577576 432138
rect 577512 432078 577576 432082
rect 469032 431995 469096 431999
rect 469032 431939 469036 431995
rect 469036 431939 469092 431995
rect 469092 431939 469096 431995
rect 469032 431935 469096 431939
rect 469112 431995 469176 431999
rect 469112 431939 469116 431995
rect 469116 431939 469172 431995
rect 469172 431939 469176 431995
rect 469112 431935 469176 431939
rect 469192 431995 469256 431999
rect 469192 431939 469196 431995
rect 469196 431939 469252 431995
rect 469252 431939 469256 431995
rect 469192 431935 469256 431939
rect 469272 431995 469336 431999
rect 469272 431939 469276 431995
rect 469276 431939 469332 431995
rect 469332 431939 469336 431995
rect 469272 431935 469336 431939
rect 469352 431995 469416 431999
rect 469352 431939 469356 431995
rect 469356 431939 469412 431995
rect 469412 431939 469416 431995
rect 469352 431935 469416 431939
rect 469432 431995 469496 431999
rect 469432 431939 469436 431995
rect 469436 431939 469492 431995
rect 469492 431939 469496 431995
rect 469432 431935 469496 431939
rect 469512 431995 469576 431999
rect 469512 431939 469516 431995
rect 469516 431939 469572 431995
rect 469572 431939 469576 431995
rect 469512 431935 469576 431939
rect 577032 432058 577096 432062
rect 577032 432002 577036 432058
rect 577036 432002 577092 432058
rect 577092 432002 577096 432058
rect 577032 431998 577096 432002
rect 577112 432058 577176 432062
rect 577112 432002 577116 432058
rect 577116 432002 577172 432058
rect 577172 432002 577176 432058
rect 577112 431998 577176 432002
rect 577192 432058 577256 432062
rect 577192 432002 577196 432058
rect 577196 432002 577252 432058
rect 577252 432002 577256 432058
rect 577192 431998 577256 432002
rect 577272 432058 577336 432062
rect 577272 432002 577276 432058
rect 577276 432002 577332 432058
rect 577332 432002 577336 432058
rect 577272 431998 577336 432002
rect 577352 432058 577416 432062
rect 577352 432002 577356 432058
rect 577356 432002 577412 432058
rect 577412 432002 577416 432058
rect 577352 431998 577416 432002
rect 577432 432058 577496 432062
rect 577432 432002 577436 432058
rect 577436 432002 577492 432058
rect 577492 432002 577496 432058
rect 577432 431998 577496 432002
rect 577512 432058 577576 432062
rect 577512 432002 577516 432058
rect 577516 432002 577572 432058
rect 577572 432002 577576 432058
rect 577512 431998 577576 432002
rect 469032 431915 469096 431919
rect 469032 431859 469036 431915
rect 469036 431859 469092 431915
rect 469092 431859 469096 431915
rect 469032 431855 469096 431859
rect 469112 431915 469176 431919
rect 469112 431859 469116 431915
rect 469116 431859 469172 431915
rect 469172 431859 469176 431915
rect 469112 431855 469176 431859
rect 469192 431915 469256 431919
rect 469192 431859 469196 431915
rect 469196 431859 469252 431915
rect 469252 431859 469256 431915
rect 469192 431855 469256 431859
rect 469272 431915 469336 431919
rect 469272 431859 469276 431915
rect 469276 431859 469332 431915
rect 469332 431859 469336 431915
rect 469272 431855 469336 431859
rect 469352 431915 469416 431919
rect 469352 431859 469356 431915
rect 469356 431859 469412 431915
rect 469412 431859 469416 431915
rect 469352 431855 469416 431859
rect 469432 431915 469496 431919
rect 469432 431859 469436 431915
rect 469436 431859 469492 431915
rect 469492 431859 469496 431915
rect 469432 431855 469496 431859
rect 469512 431915 469576 431919
rect 469512 431859 469516 431915
rect 469516 431859 469572 431915
rect 469572 431859 469576 431915
rect 469512 431855 469576 431859
rect 469032 431835 469096 431839
rect 469032 431779 469036 431835
rect 469036 431779 469092 431835
rect 469092 431779 469096 431835
rect 469032 431775 469096 431779
rect 469112 431835 469176 431839
rect 469112 431779 469116 431835
rect 469116 431779 469172 431835
rect 469172 431779 469176 431835
rect 469112 431775 469176 431779
rect 469192 431835 469256 431839
rect 469192 431779 469196 431835
rect 469196 431779 469252 431835
rect 469252 431779 469256 431835
rect 469192 431775 469256 431779
rect 469272 431835 469336 431839
rect 469272 431779 469276 431835
rect 469276 431779 469332 431835
rect 469332 431779 469336 431835
rect 469272 431775 469336 431779
rect 469352 431835 469416 431839
rect 469352 431779 469356 431835
rect 469356 431779 469412 431835
rect 469412 431779 469416 431835
rect 469352 431775 469416 431779
rect 469432 431835 469496 431839
rect 469432 431779 469436 431835
rect 469436 431779 469492 431835
rect 469492 431779 469496 431835
rect 469432 431775 469496 431779
rect 469512 431835 469576 431839
rect 469512 431779 469516 431835
rect 469516 431779 469572 431835
rect 469572 431779 469576 431835
rect 469512 431775 469576 431779
rect 473676 431838 473740 431902
rect 469032 431755 469096 431759
rect 469032 431699 469036 431755
rect 469036 431699 469092 431755
rect 469092 431699 469096 431755
rect 469032 431695 469096 431699
rect 469112 431755 469176 431759
rect 469112 431699 469116 431755
rect 469116 431699 469172 431755
rect 469172 431699 469176 431755
rect 469112 431695 469176 431699
rect 469192 431755 469256 431759
rect 469192 431699 469196 431755
rect 469196 431699 469252 431755
rect 469252 431699 469256 431755
rect 469192 431695 469256 431699
rect 469272 431755 469336 431759
rect 469272 431699 469276 431755
rect 469276 431699 469332 431755
rect 469332 431699 469336 431755
rect 469272 431695 469336 431699
rect 469352 431755 469416 431759
rect 469352 431699 469356 431755
rect 469356 431699 469412 431755
rect 469412 431699 469416 431755
rect 469352 431695 469416 431699
rect 469432 431755 469496 431759
rect 469432 431699 469436 431755
rect 469436 431699 469492 431755
rect 469492 431699 469496 431755
rect 469432 431695 469496 431699
rect 469512 431755 469576 431759
rect 469512 431699 469516 431755
rect 469516 431699 469572 431755
rect 469572 431699 469576 431755
rect 469512 431695 469576 431699
rect 478460 431566 478524 431630
rect 488396 431626 488460 431630
rect 488396 431570 488433 431626
rect 488433 431570 488460 431626
rect 488396 431566 488460 431570
rect 578272 431503 578336 431507
rect 578272 431447 578276 431503
rect 578276 431447 578332 431503
rect 578332 431447 578336 431503
rect 578272 431443 578336 431447
rect 578352 431503 578416 431507
rect 578352 431447 578356 431503
rect 578356 431447 578412 431503
rect 578412 431447 578416 431503
rect 578352 431443 578416 431447
rect 578432 431503 578496 431507
rect 578432 431447 578436 431503
rect 578436 431447 578492 431503
rect 578492 431447 578496 431503
rect 578432 431443 578496 431447
rect 578512 431503 578576 431507
rect 578512 431447 578516 431503
rect 578516 431447 578572 431503
rect 578572 431447 578576 431503
rect 578512 431443 578576 431447
rect 578592 431503 578656 431507
rect 578592 431447 578596 431503
rect 578596 431447 578652 431503
rect 578652 431447 578656 431503
rect 578592 431443 578656 431447
rect 578672 431503 578736 431507
rect 578672 431447 578676 431503
rect 578676 431447 578732 431503
rect 578732 431447 578736 431503
rect 578672 431443 578736 431447
rect 578752 431503 578816 431507
rect 578752 431447 578756 431503
rect 578756 431447 578812 431503
rect 578812 431447 578816 431503
rect 578752 431443 578816 431447
rect 578272 431423 578336 431427
rect 578272 431367 578276 431423
rect 578276 431367 578332 431423
rect 578332 431367 578336 431423
rect 578272 431363 578336 431367
rect 578352 431423 578416 431427
rect 578352 431367 578356 431423
rect 578356 431367 578412 431423
rect 578412 431367 578416 431423
rect 578352 431363 578416 431367
rect 578432 431423 578496 431427
rect 578432 431367 578436 431423
rect 578436 431367 578492 431423
rect 578492 431367 578496 431423
rect 578432 431363 578496 431367
rect 578512 431423 578576 431427
rect 578512 431367 578516 431423
rect 578516 431367 578572 431423
rect 578572 431367 578576 431423
rect 578512 431363 578576 431367
rect 578592 431423 578656 431427
rect 578592 431367 578596 431423
rect 578596 431367 578652 431423
rect 578652 431367 578656 431423
rect 578592 431363 578656 431367
rect 578672 431423 578736 431427
rect 578672 431367 578676 431423
rect 578676 431367 578732 431423
rect 578732 431367 578736 431423
rect 578672 431363 578736 431367
rect 578752 431423 578816 431427
rect 578752 431367 578756 431423
rect 578756 431367 578812 431423
rect 578812 431367 578816 431423
rect 578752 431363 578816 431367
rect 578272 431343 578336 431347
rect 578272 431287 578276 431343
rect 578276 431287 578332 431343
rect 578332 431287 578336 431343
rect 578272 431283 578336 431287
rect 578352 431343 578416 431347
rect 578352 431287 578356 431343
rect 578356 431287 578412 431343
rect 578412 431287 578416 431343
rect 578352 431283 578416 431287
rect 578432 431343 578496 431347
rect 578432 431287 578436 431343
rect 578436 431287 578492 431343
rect 578492 431287 578496 431343
rect 578432 431283 578496 431287
rect 578512 431343 578576 431347
rect 578512 431287 578516 431343
rect 578516 431287 578572 431343
rect 578572 431287 578576 431343
rect 578512 431283 578576 431287
rect 578592 431343 578656 431347
rect 578592 431287 578596 431343
rect 578596 431287 578652 431343
rect 578652 431287 578656 431343
rect 578592 431283 578656 431287
rect 578672 431343 578736 431347
rect 578672 431287 578676 431343
rect 578676 431287 578732 431343
rect 578732 431287 578736 431343
rect 578672 431283 578736 431287
rect 578752 431343 578816 431347
rect 578752 431287 578756 431343
rect 578756 431287 578812 431343
rect 578812 431287 578816 431343
rect 578752 431283 578816 431287
rect 578272 431263 578336 431267
rect 578272 431207 578276 431263
rect 578276 431207 578332 431263
rect 578332 431207 578336 431263
rect 578272 431203 578336 431207
rect 578352 431263 578416 431267
rect 578352 431207 578356 431263
rect 578356 431207 578412 431263
rect 578412 431207 578416 431263
rect 578352 431203 578416 431207
rect 578432 431263 578496 431267
rect 578432 431207 578436 431263
rect 578436 431207 578492 431263
rect 578492 431207 578496 431263
rect 578432 431203 578496 431207
rect 578512 431263 578576 431267
rect 578512 431207 578516 431263
rect 578516 431207 578572 431263
rect 578572 431207 578576 431263
rect 578512 431203 578576 431207
rect 578592 431263 578656 431267
rect 578592 431207 578596 431263
rect 578596 431207 578652 431263
rect 578652 431207 578656 431263
rect 578592 431203 578656 431207
rect 578672 431263 578736 431267
rect 578672 431207 578676 431263
rect 578676 431207 578732 431263
rect 578732 431207 578736 431263
rect 578672 431203 578736 431207
rect 578752 431263 578816 431267
rect 578752 431207 578756 431263
rect 578756 431207 578812 431263
rect 578812 431207 578816 431263
rect 578752 431203 578816 431207
rect 470272 430910 470336 430914
rect 470272 430854 470276 430910
rect 470276 430854 470332 430910
rect 470332 430854 470336 430910
rect 470272 430850 470336 430854
rect 470352 430910 470416 430914
rect 470352 430854 470356 430910
rect 470356 430854 470412 430910
rect 470412 430854 470416 430910
rect 470352 430850 470416 430854
rect 470432 430910 470496 430914
rect 470432 430854 470436 430910
rect 470436 430854 470492 430910
rect 470492 430854 470496 430910
rect 470432 430850 470496 430854
rect 470512 430910 470576 430914
rect 470512 430854 470516 430910
rect 470516 430854 470572 430910
rect 470572 430854 470576 430910
rect 470512 430850 470576 430854
rect 470592 430910 470656 430914
rect 470592 430854 470596 430910
rect 470596 430854 470652 430910
rect 470652 430854 470656 430910
rect 470592 430850 470656 430854
rect 470672 430910 470736 430914
rect 470672 430854 470676 430910
rect 470676 430854 470732 430910
rect 470732 430854 470736 430910
rect 470672 430850 470736 430854
rect 470752 430910 470816 430914
rect 470752 430854 470756 430910
rect 470756 430854 470812 430910
rect 470812 430854 470816 430910
rect 470752 430850 470816 430854
rect 470272 430830 470336 430834
rect 470272 430774 470276 430830
rect 470276 430774 470332 430830
rect 470332 430774 470336 430830
rect 470272 430770 470336 430774
rect 470352 430830 470416 430834
rect 470352 430774 470356 430830
rect 470356 430774 470412 430830
rect 470412 430774 470416 430830
rect 470352 430770 470416 430774
rect 470432 430830 470496 430834
rect 470432 430774 470436 430830
rect 470436 430774 470492 430830
rect 470492 430774 470496 430830
rect 470432 430770 470496 430774
rect 470512 430830 470576 430834
rect 470512 430774 470516 430830
rect 470516 430774 470572 430830
rect 470572 430774 470576 430830
rect 470512 430770 470576 430774
rect 470592 430830 470656 430834
rect 470592 430774 470596 430830
rect 470596 430774 470652 430830
rect 470652 430774 470656 430830
rect 470592 430770 470656 430774
rect 470672 430830 470736 430834
rect 470672 430774 470676 430830
rect 470676 430774 470732 430830
rect 470732 430774 470736 430830
rect 470672 430770 470736 430774
rect 470752 430830 470816 430834
rect 470752 430774 470756 430830
rect 470756 430774 470812 430830
rect 470812 430774 470816 430830
rect 470752 430770 470816 430774
rect 470272 430750 470336 430754
rect 470272 430694 470276 430750
rect 470276 430694 470332 430750
rect 470332 430694 470336 430750
rect 470272 430690 470336 430694
rect 470352 430750 470416 430754
rect 470352 430694 470356 430750
rect 470356 430694 470412 430750
rect 470412 430694 470416 430750
rect 470352 430690 470416 430694
rect 470432 430750 470496 430754
rect 470432 430694 470436 430750
rect 470436 430694 470492 430750
rect 470492 430694 470496 430750
rect 470432 430690 470496 430694
rect 470512 430750 470576 430754
rect 470512 430694 470516 430750
rect 470516 430694 470572 430750
rect 470572 430694 470576 430750
rect 470512 430690 470576 430694
rect 470592 430750 470656 430754
rect 470592 430694 470596 430750
rect 470596 430694 470652 430750
rect 470652 430694 470656 430750
rect 470592 430690 470656 430694
rect 470672 430750 470736 430754
rect 470672 430694 470676 430750
rect 470676 430694 470732 430750
rect 470732 430694 470736 430750
rect 470672 430690 470736 430694
rect 470752 430750 470816 430754
rect 470752 430694 470756 430750
rect 470756 430694 470812 430750
rect 470812 430694 470816 430750
rect 470752 430690 470816 430694
rect 470272 430670 470336 430674
rect 470272 430614 470276 430670
rect 470276 430614 470332 430670
rect 470332 430614 470336 430670
rect 470272 430610 470336 430614
rect 470352 430670 470416 430674
rect 470352 430614 470356 430670
rect 470356 430614 470412 430670
rect 470412 430614 470416 430670
rect 470352 430610 470416 430614
rect 470432 430670 470496 430674
rect 470432 430614 470436 430670
rect 470436 430614 470492 430670
rect 470492 430614 470496 430670
rect 470432 430610 470496 430614
rect 470512 430670 470576 430674
rect 470512 430614 470516 430670
rect 470516 430614 470572 430670
rect 470572 430614 470576 430670
rect 470512 430610 470576 430614
rect 470592 430670 470656 430674
rect 470592 430614 470596 430670
rect 470596 430614 470652 430670
rect 470652 430614 470656 430670
rect 470592 430610 470656 430614
rect 470672 430670 470736 430674
rect 470672 430614 470676 430670
rect 470676 430614 470732 430670
rect 470732 430614 470736 430670
rect 470672 430610 470736 430614
rect 470752 430670 470816 430674
rect 470752 430614 470756 430670
rect 470756 430614 470812 430670
rect 470812 430614 470816 430670
rect 470752 430610 470816 430614
rect 480116 427894 480180 427958
rect 486556 427894 486620 427958
rect 488396 413886 488460 413950
rect 470272 412082 470336 412086
rect 470272 412026 470276 412082
rect 470276 412026 470332 412082
rect 470332 412026 470336 412082
rect 470272 412022 470336 412026
rect 470352 412082 470416 412086
rect 470352 412026 470356 412082
rect 470356 412026 470412 412082
rect 470412 412026 470416 412082
rect 470352 412022 470416 412026
rect 470432 412082 470496 412086
rect 470432 412026 470436 412082
rect 470436 412026 470492 412082
rect 470492 412026 470496 412082
rect 470432 412022 470496 412026
rect 470512 412082 470576 412086
rect 470512 412026 470516 412082
rect 470516 412026 470572 412082
rect 470572 412026 470576 412082
rect 470512 412022 470576 412026
rect 470592 412082 470656 412086
rect 470592 412026 470596 412082
rect 470596 412026 470652 412082
rect 470652 412026 470656 412082
rect 470592 412022 470656 412026
rect 470672 412082 470736 412086
rect 470672 412026 470676 412082
rect 470676 412026 470732 412082
rect 470732 412026 470736 412082
rect 470672 412022 470736 412026
rect 470752 412082 470816 412086
rect 470752 412026 470756 412082
rect 470756 412026 470812 412082
rect 470812 412026 470816 412082
rect 470752 412022 470816 412026
rect 470272 412002 470336 412006
rect 470272 411946 470276 412002
rect 470276 411946 470332 412002
rect 470332 411946 470336 412002
rect 470272 411942 470336 411946
rect 470352 412002 470416 412006
rect 470352 411946 470356 412002
rect 470356 411946 470412 412002
rect 470412 411946 470416 412002
rect 470352 411942 470416 411946
rect 470432 412002 470496 412006
rect 470432 411946 470436 412002
rect 470436 411946 470492 412002
rect 470492 411946 470496 412002
rect 470432 411942 470496 411946
rect 470512 412002 470576 412006
rect 470512 411946 470516 412002
rect 470516 411946 470572 412002
rect 470572 411946 470576 412002
rect 470512 411942 470576 411946
rect 470592 412002 470656 412006
rect 470592 411946 470596 412002
rect 470596 411946 470652 412002
rect 470652 411946 470656 412002
rect 470592 411942 470656 411946
rect 470672 412002 470736 412006
rect 470672 411946 470676 412002
rect 470676 411946 470732 412002
rect 470732 411946 470736 412002
rect 470672 411942 470736 411946
rect 470752 412002 470816 412006
rect 470752 411946 470756 412002
rect 470756 411946 470812 412002
rect 470812 411946 470816 412002
rect 470752 411942 470816 411946
rect 470272 411922 470336 411926
rect 470272 411866 470276 411922
rect 470276 411866 470332 411922
rect 470332 411866 470336 411922
rect 470272 411862 470336 411866
rect 470352 411922 470416 411926
rect 470352 411866 470356 411922
rect 470356 411866 470412 411922
rect 470412 411866 470416 411922
rect 470352 411862 470416 411866
rect 470432 411922 470496 411926
rect 470432 411866 470436 411922
rect 470436 411866 470492 411922
rect 470492 411866 470496 411922
rect 470432 411862 470496 411866
rect 470512 411922 470576 411926
rect 470512 411866 470516 411922
rect 470516 411866 470572 411922
rect 470572 411866 470576 411922
rect 470512 411862 470576 411866
rect 470592 411922 470656 411926
rect 470592 411866 470596 411922
rect 470596 411866 470652 411922
rect 470652 411866 470656 411922
rect 470592 411862 470656 411866
rect 470672 411922 470736 411926
rect 470672 411866 470676 411922
rect 470676 411866 470732 411922
rect 470732 411866 470736 411922
rect 470672 411862 470736 411866
rect 470752 411922 470816 411926
rect 470752 411866 470756 411922
rect 470756 411866 470812 411922
rect 470812 411866 470816 411922
rect 470752 411862 470816 411866
rect 470272 411842 470336 411846
rect 470272 411786 470276 411842
rect 470276 411786 470332 411842
rect 470332 411786 470336 411842
rect 470272 411782 470336 411786
rect 470352 411842 470416 411846
rect 470352 411786 470356 411842
rect 470356 411786 470412 411842
rect 470412 411786 470416 411842
rect 470352 411782 470416 411786
rect 470432 411842 470496 411846
rect 470432 411786 470436 411842
rect 470436 411786 470492 411842
rect 470492 411786 470496 411842
rect 470432 411782 470496 411786
rect 470512 411842 470576 411846
rect 470512 411786 470516 411842
rect 470516 411786 470572 411842
rect 470572 411786 470576 411842
rect 470512 411782 470576 411786
rect 470592 411842 470656 411846
rect 470592 411786 470596 411842
rect 470596 411786 470652 411842
rect 470652 411786 470656 411842
rect 470592 411782 470656 411786
rect 470672 411842 470736 411846
rect 470672 411786 470676 411842
rect 470676 411786 470732 411842
rect 470732 411786 470736 411842
rect 470672 411782 470736 411786
rect 470752 411842 470816 411846
rect 470752 411786 470756 411842
rect 470756 411786 470812 411842
rect 470812 411786 470816 411842
rect 470752 411782 470816 411786
rect 469032 410996 469096 411000
rect 469032 410940 469036 410996
rect 469036 410940 469092 410996
rect 469092 410940 469096 410996
rect 469032 410936 469096 410940
rect 469112 410996 469176 411000
rect 469112 410940 469116 410996
rect 469116 410940 469172 410996
rect 469172 410940 469176 410996
rect 469112 410936 469176 410940
rect 469192 410996 469256 411000
rect 469192 410940 469196 410996
rect 469196 410940 469252 410996
rect 469252 410940 469256 410996
rect 469192 410936 469256 410940
rect 469272 410996 469336 411000
rect 469272 410940 469276 410996
rect 469276 410940 469332 410996
rect 469332 410940 469336 410996
rect 469272 410936 469336 410940
rect 469352 410996 469416 411000
rect 469352 410940 469356 410996
rect 469356 410940 469412 410996
rect 469412 410940 469416 410996
rect 469352 410936 469416 410940
rect 469432 410996 469496 411000
rect 469432 410940 469436 410996
rect 469436 410940 469492 410996
rect 469492 410940 469496 410996
rect 469432 410936 469496 410940
rect 469512 410996 469576 411000
rect 469512 410940 469516 410996
rect 469516 410940 469572 410996
rect 469572 410940 469576 410996
rect 469512 410936 469576 410940
rect 469032 410916 469096 410920
rect 469032 410860 469036 410916
rect 469036 410860 469092 410916
rect 469092 410860 469096 410916
rect 469032 410856 469096 410860
rect 469112 410916 469176 410920
rect 469112 410860 469116 410916
rect 469116 410860 469172 410916
rect 469172 410860 469176 410916
rect 469112 410856 469176 410860
rect 469192 410916 469256 410920
rect 469192 410860 469196 410916
rect 469196 410860 469252 410916
rect 469252 410860 469256 410916
rect 469192 410856 469256 410860
rect 469272 410916 469336 410920
rect 469272 410860 469276 410916
rect 469276 410860 469332 410916
rect 469332 410860 469336 410916
rect 469272 410856 469336 410860
rect 469352 410916 469416 410920
rect 469352 410860 469356 410916
rect 469356 410860 469412 410916
rect 469412 410860 469416 410916
rect 469352 410856 469416 410860
rect 469432 410916 469496 410920
rect 469432 410860 469436 410916
rect 469436 410860 469492 410916
rect 469492 410860 469496 410916
rect 469432 410856 469496 410860
rect 469512 410916 469576 410920
rect 469512 410860 469516 410916
rect 469516 410860 469572 410916
rect 469572 410860 469576 410916
rect 469512 410856 469576 410860
rect 473676 410954 473740 410958
rect 473676 410898 473726 410954
rect 473726 410898 473740 410954
rect 473676 410894 473740 410898
rect 469032 410836 469096 410840
rect 469032 410780 469036 410836
rect 469036 410780 469092 410836
rect 469092 410780 469096 410836
rect 469032 410776 469096 410780
rect 469112 410836 469176 410840
rect 469112 410780 469116 410836
rect 469116 410780 469172 410836
rect 469172 410780 469176 410836
rect 469112 410776 469176 410780
rect 469192 410836 469256 410840
rect 469192 410780 469196 410836
rect 469196 410780 469252 410836
rect 469252 410780 469256 410836
rect 469192 410776 469256 410780
rect 469272 410836 469336 410840
rect 469272 410780 469276 410836
rect 469276 410780 469332 410836
rect 469332 410780 469336 410836
rect 469272 410776 469336 410780
rect 469352 410836 469416 410840
rect 469352 410780 469356 410836
rect 469356 410780 469412 410836
rect 469412 410780 469416 410836
rect 469352 410776 469416 410780
rect 469432 410836 469496 410840
rect 469432 410780 469436 410836
rect 469436 410780 469492 410836
rect 469492 410780 469496 410836
rect 469432 410776 469496 410780
rect 469512 410836 469576 410840
rect 469512 410780 469516 410836
rect 469516 410780 469572 410836
rect 469572 410780 469576 410836
rect 469512 410776 469576 410780
rect 469032 410756 469096 410760
rect 469032 410700 469036 410756
rect 469036 410700 469092 410756
rect 469092 410700 469096 410756
rect 469032 410696 469096 410700
rect 469112 410756 469176 410760
rect 469112 410700 469116 410756
rect 469116 410700 469172 410756
rect 469172 410700 469176 410756
rect 469112 410696 469176 410700
rect 469192 410756 469256 410760
rect 469192 410700 469196 410756
rect 469196 410700 469252 410756
rect 469252 410700 469256 410756
rect 469192 410696 469256 410700
rect 469272 410756 469336 410760
rect 469272 410700 469276 410756
rect 469276 410700 469332 410756
rect 469332 410700 469336 410756
rect 469272 410696 469336 410700
rect 469352 410756 469416 410760
rect 469352 410700 469356 410756
rect 469356 410700 469412 410756
rect 469412 410700 469416 410756
rect 469352 410696 469416 410700
rect 469432 410756 469496 410760
rect 469432 410700 469436 410756
rect 469436 410700 469492 410756
rect 469492 410700 469496 410756
rect 469432 410696 469496 410700
rect 469512 410756 469576 410760
rect 469512 410700 469516 410756
rect 469516 410700 469572 410756
rect 469572 410700 469576 410756
rect 469512 410696 469576 410700
rect 484164 410410 484228 410414
rect 484164 410354 484178 410410
rect 484178 410354 484228 410410
rect 484164 410350 484228 410354
rect 478460 410138 478524 410142
rect 478460 410082 478474 410138
rect 478474 410082 478524 410138
rect 478460 410078 478524 410082
rect 481404 410138 481468 410142
rect 481404 410082 481418 410138
rect 481418 410082 481468 410138
rect 481404 410078 481468 410082
rect 470272 409910 470336 409914
rect 470272 409854 470276 409910
rect 470276 409854 470332 409910
rect 470332 409854 470336 409910
rect 470272 409850 470336 409854
rect 470352 409910 470416 409914
rect 470352 409854 470356 409910
rect 470356 409854 470412 409910
rect 470412 409854 470416 409910
rect 470352 409850 470416 409854
rect 470432 409910 470496 409914
rect 470432 409854 470436 409910
rect 470436 409854 470492 409910
rect 470492 409854 470496 409910
rect 470432 409850 470496 409854
rect 470512 409910 470576 409914
rect 470512 409854 470516 409910
rect 470516 409854 470572 409910
rect 470572 409854 470576 409910
rect 470512 409850 470576 409854
rect 470592 409910 470656 409914
rect 470592 409854 470596 409910
rect 470596 409854 470652 409910
rect 470652 409854 470656 409910
rect 470592 409850 470656 409854
rect 470672 409910 470736 409914
rect 470672 409854 470676 409910
rect 470676 409854 470732 409910
rect 470732 409854 470736 409910
rect 470672 409850 470736 409854
rect 470752 409910 470816 409914
rect 470752 409854 470756 409910
rect 470756 409854 470812 409910
rect 470812 409854 470816 409910
rect 470752 409850 470816 409854
rect 470272 409830 470336 409834
rect 470272 409774 470276 409830
rect 470276 409774 470332 409830
rect 470332 409774 470336 409830
rect 470272 409770 470336 409774
rect 470352 409830 470416 409834
rect 470352 409774 470356 409830
rect 470356 409774 470412 409830
rect 470412 409774 470416 409830
rect 470352 409770 470416 409774
rect 470432 409830 470496 409834
rect 470432 409774 470436 409830
rect 470436 409774 470492 409830
rect 470492 409774 470496 409830
rect 470432 409770 470496 409774
rect 470512 409830 470576 409834
rect 470512 409774 470516 409830
rect 470516 409774 470572 409830
rect 470572 409774 470576 409830
rect 470512 409770 470576 409774
rect 470592 409830 470656 409834
rect 470592 409774 470596 409830
rect 470596 409774 470652 409830
rect 470652 409774 470656 409830
rect 470592 409770 470656 409774
rect 470672 409830 470736 409834
rect 470672 409774 470676 409830
rect 470676 409774 470732 409830
rect 470732 409774 470736 409830
rect 470672 409770 470736 409774
rect 470752 409830 470816 409834
rect 470752 409774 470756 409830
rect 470756 409774 470812 409830
rect 470812 409774 470816 409830
rect 470752 409770 470816 409774
rect 470272 409750 470336 409754
rect 470272 409694 470276 409750
rect 470276 409694 470332 409750
rect 470332 409694 470336 409750
rect 470272 409690 470336 409694
rect 470352 409750 470416 409754
rect 470352 409694 470356 409750
rect 470356 409694 470412 409750
rect 470412 409694 470416 409750
rect 470352 409690 470416 409694
rect 470432 409750 470496 409754
rect 470432 409694 470436 409750
rect 470436 409694 470492 409750
rect 470492 409694 470496 409750
rect 470432 409690 470496 409694
rect 470512 409750 470576 409754
rect 470512 409694 470516 409750
rect 470516 409694 470572 409750
rect 470572 409694 470576 409750
rect 470512 409690 470576 409694
rect 470592 409750 470656 409754
rect 470592 409694 470596 409750
rect 470596 409694 470652 409750
rect 470652 409694 470656 409750
rect 470592 409690 470656 409694
rect 470672 409750 470736 409754
rect 470672 409694 470676 409750
rect 470676 409694 470732 409750
rect 470732 409694 470736 409750
rect 470672 409690 470736 409694
rect 470752 409750 470816 409754
rect 470752 409694 470756 409750
rect 470756 409694 470812 409750
rect 470812 409694 470816 409750
rect 470752 409690 470816 409694
rect 470272 409670 470336 409674
rect 470272 409614 470276 409670
rect 470276 409614 470332 409670
rect 470332 409614 470336 409670
rect 470272 409610 470336 409614
rect 470352 409670 470416 409674
rect 470352 409614 470356 409670
rect 470356 409614 470412 409670
rect 470412 409614 470416 409670
rect 470352 409610 470416 409614
rect 470432 409670 470496 409674
rect 470432 409614 470436 409670
rect 470436 409614 470492 409670
rect 470492 409614 470496 409670
rect 470432 409610 470496 409614
rect 470512 409670 470576 409674
rect 470512 409614 470516 409670
rect 470516 409614 470572 409670
rect 470572 409614 470576 409670
rect 470512 409610 470576 409614
rect 470592 409670 470656 409674
rect 470592 409614 470596 409670
rect 470596 409614 470652 409670
rect 470652 409614 470656 409670
rect 470592 409610 470656 409614
rect 470672 409670 470736 409674
rect 470672 409614 470676 409670
rect 470676 409614 470732 409670
rect 470732 409614 470736 409670
rect 470672 409610 470736 409614
rect 470752 409670 470816 409674
rect 470752 409614 470756 409670
rect 470756 409614 470812 409670
rect 470812 409614 470816 409670
rect 470752 409610 470816 409614
rect 541572 409262 541636 409326
rect 544332 409322 544396 409326
rect 544332 409266 544346 409322
rect 544346 409266 544396 409322
rect 544332 409262 544396 409266
rect 480116 407494 480180 407558
rect 482876 407086 482940 407150
rect 485636 407086 485700 407150
rect 473676 391990 473740 392054
rect 474964 391990 475028 392054
rect 489316 391990 489380 392054
rect 470272 391083 470336 391087
rect 470272 391027 470276 391083
rect 470276 391027 470332 391083
rect 470332 391027 470336 391083
rect 470272 391023 470336 391027
rect 470352 391083 470416 391087
rect 470352 391027 470356 391083
rect 470356 391027 470412 391083
rect 470412 391027 470416 391083
rect 470352 391023 470416 391027
rect 470432 391083 470496 391087
rect 470432 391027 470436 391083
rect 470436 391027 470492 391083
rect 470492 391027 470496 391083
rect 470432 391023 470496 391027
rect 470512 391083 470576 391087
rect 470512 391027 470516 391083
rect 470516 391027 470572 391083
rect 470572 391027 470576 391083
rect 470512 391023 470576 391027
rect 470592 391083 470656 391087
rect 470592 391027 470596 391083
rect 470596 391027 470652 391083
rect 470652 391027 470656 391083
rect 470592 391023 470656 391027
rect 470672 391083 470736 391087
rect 470672 391027 470676 391083
rect 470676 391027 470732 391083
rect 470732 391027 470736 391083
rect 470672 391023 470736 391027
rect 470752 391083 470816 391087
rect 470752 391027 470756 391083
rect 470756 391027 470812 391083
rect 470812 391027 470816 391083
rect 470752 391023 470816 391027
rect 470272 391003 470336 391007
rect 470272 390947 470276 391003
rect 470276 390947 470332 391003
rect 470332 390947 470336 391003
rect 470272 390943 470336 390947
rect 470352 391003 470416 391007
rect 470352 390947 470356 391003
rect 470356 390947 470412 391003
rect 470412 390947 470416 391003
rect 470352 390943 470416 390947
rect 470432 391003 470496 391007
rect 470432 390947 470436 391003
rect 470436 390947 470492 391003
rect 470492 390947 470496 391003
rect 470432 390943 470496 390947
rect 470512 391003 470576 391007
rect 470512 390947 470516 391003
rect 470516 390947 470572 391003
rect 470572 390947 470576 391003
rect 470512 390943 470576 390947
rect 470592 391003 470656 391007
rect 470592 390947 470596 391003
rect 470596 390947 470652 391003
rect 470652 390947 470656 391003
rect 470592 390943 470656 390947
rect 470672 391003 470736 391007
rect 470672 390947 470676 391003
rect 470676 390947 470732 391003
rect 470732 390947 470736 391003
rect 470672 390943 470736 390947
rect 470752 391003 470816 391007
rect 470752 390947 470756 391003
rect 470756 390947 470812 391003
rect 470812 390947 470816 391003
rect 470752 390943 470816 390947
rect 470272 390923 470336 390927
rect 470272 390867 470276 390923
rect 470276 390867 470332 390923
rect 470332 390867 470336 390923
rect 470272 390863 470336 390867
rect 470352 390923 470416 390927
rect 470352 390867 470356 390923
rect 470356 390867 470412 390923
rect 470412 390867 470416 390923
rect 470352 390863 470416 390867
rect 470432 390923 470496 390927
rect 470432 390867 470436 390923
rect 470436 390867 470492 390923
rect 470492 390867 470496 390923
rect 470432 390863 470496 390867
rect 470512 390923 470576 390927
rect 470512 390867 470516 390923
rect 470516 390867 470572 390923
rect 470572 390867 470576 390923
rect 470512 390863 470576 390867
rect 470592 390923 470656 390927
rect 470592 390867 470596 390923
rect 470596 390867 470652 390923
rect 470652 390867 470656 390923
rect 470592 390863 470656 390867
rect 470672 390923 470736 390927
rect 470672 390867 470676 390923
rect 470676 390867 470732 390923
rect 470732 390867 470736 390923
rect 470672 390863 470736 390867
rect 470752 390923 470816 390927
rect 470752 390867 470756 390923
rect 470756 390867 470812 390923
rect 470812 390867 470816 390923
rect 470752 390863 470816 390867
rect 470272 390843 470336 390847
rect 470272 390787 470276 390843
rect 470276 390787 470332 390843
rect 470332 390787 470336 390843
rect 470272 390783 470336 390787
rect 470352 390843 470416 390847
rect 470352 390787 470356 390843
rect 470356 390787 470412 390843
rect 470412 390787 470416 390843
rect 470352 390783 470416 390787
rect 470432 390843 470496 390847
rect 470432 390787 470436 390843
rect 470436 390787 470492 390843
rect 470492 390787 470496 390843
rect 470432 390783 470496 390787
rect 470512 390843 470576 390847
rect 470512 390787 470516 390843
rect 470516 390787 470572 390843
rect 470572 390787 470576 390843
rect 470512 390783 470576 390787
rect 470592 390843 470656 390847
rect 470592 390787 470596 390843
rect 470596 390787 470652 390843
rect 470652 390787 470656 390843
rect 470592 390783 470656 390787
rect 470672 390843 470736 390847
rect 470672 390787 470676 390843
rect 470676 390787 470732 390843
rect 470732 390787 470736 390843
rect 470672 390783 470736 390787
rect 470752 390843 470816 390847
rect 470752 390787 470756 390843
rect 470756 390787 470812 390843
rect 470812 390787 470816 390843
rect 470752 390783 470816 390787
rect 484900 390235 484964 390299
rect 469032 390000 469096 390004
rect 469032 389944 469036 390000
rect 469036 389944 469092 390000
rect 469092 389944 469096 390000
rect 469032 389940 469096 389944
rect 469112 390000 469176 390004
rect 469112 389944 469116 390000
rect 469116 389944 469172 390000
rect 469172 389944 469176 390000
rect 469112 389940 469176 389944
rect 469192 390000 469256 390004
rect 469192 389944 469196 390000
rect 469196 389944 469252 390000
rect 469252 389944 469256 390000
rect 469192 389940 469256 389944
rect 469272 390000 469336 390004
rect 469272 389944 469276 390000
rect 469276 389944 469332 390000
rect 469332 389944 469336 390000
rect 469272 389940 469336 389944
rect 469352 390000 469416 390004
rect 469352 389944 469356 390000
rect 469356 389944 469412 390000
rect 469412 389944 469416 390000
rect 469352 389940 469416 389944
rect 469432 390000 469496 390004
rect 469432 389944 469436 390000
rect 469436 389944 469492 390000
rect 469492 389944 469496 390000
rect 469432 389940 469496 389944
rect 469512 390000 469576 390004
rect 469512 389944 469516 390000
rect 469516 389944 469572 390000
rect 469572 389944 469576 390000
rect 469512 389940 469576 389944
rect 469032 389920 469096 389924
rect 469032 389864 469036 389920
rect 469036 389864 469092 389920
rect 469092 389864 469096 389920
rect 469032 389860 469096 389864
rect 469112 389920 469176 389924
rect 469112 389864 469116 389920
rect 469116 389864 469172 389920
rect 469172 389864 469176 389920
rect 469112 389860 469176 389864
rect 469192 389920 469256 389924
rect 469192 389864 469196 389920
rect 469196 389864 469252 389920
rect 469252 389864 469256 389920
rect 469192 389860 469256 389864
rect 469272 389920 469336 389924
rect 469272 389864 469276 389920
rect 469276 389864 469332 389920
rect 469332 389864 469336 389920
rect 469272 389860 469336 389864
rect 469352 389920 469416 389924
rect 469352 389864 469356 389920
rect 469356 389864 469412 389920
rect 469412 389864 469416 389920
rect 469352 389860 469416 389864
rect 469432 389920 469496 389924
rect 469432 389864 469436 389920
rect 469436 389864 469492 389920
rect 469492 389864 469496 389920
rect 469432 389860 469496 389864
rect 469512 389920 469576 389924
rect 469512 389864 469516 389920
rect 469516 389864 469572 389920
rect 469572 389864 469576 389920
rect 469512 389860 469576 389864
rect 469032 389840 469096 389844
rect 469032 389784 469036 389840
rect 469036 389784 469092 389840
rect 469092 389784 469096 389840
rect 469032 389780 469096 389784
rect 469112 389840 469176 389844
rect 469112 389784 469116 389840
rect 469116 389784 469172 389840
rect 469172 389784 469176 389840
rect 469112 389780 469176 389784
rect 469192 389840 469256 389844
rect 469192 389784 469196 389840
rect 469196 389784 469252 389840
rect 469252 389784 469256 389840
rect 469192 389780 469256 389784
rect 469272 389840 469336 389844
rect 469272 389784 469276 389840
rect 469276 389784 469332 389840
rect 469332 389784 469336 389840
rect 469272 389780 469336 389784
rect 469352 389840 469416 389844
rect 469352 389784 469356 389840
rect 469356 389784 469412 389840
rect 469412 389784 469416 389840
rect 469352 389780 469416 389784
rect 469432 389840 469496 389844
rect 469432 389784 469436 389840
rect 469436 389784 469492 389840
rect 469492 389784 469496 389840
rect 469432 389780 469496 389784
rect 469512 389840 469576 389844
rect 469512 389784 469516 389840
rect 469516 389784 469572 389840
rect 469572 389784 469576 389840
rect 469512 389780 469576 389784
rect 469032 389760 469096 389764
rect 469032 389704 469036 389760
rect 469036 389704 469092 389760
rect 469092 389704 469096 389760
rect 469032 389700 469096 389704
rect 469112 389760 469176 389764
rect 469112 389704 469116 389760
rect 469116 389704 469172 389760
rect 469172 389704 469176 389760
rect 469112 389700 469176 389704
rect 469192 389760 469256 389764
rect 469192 389704 469196 389760
rect 469196 389704 469252 389760
rect 469252 389704 469256 389760
rect 469192 389700 469256 389704
rect 469272 389760 469336 389764
rect 469272 389704 469276 389760
rect 469276 389704 469332 389760
rect 469332 389704 469336 389760
rect 469272 389700 469336 389704
rect 469352 389760 469416 389764
rect 469352 389704 469356 389760
rect 469356 389704 469412 389760
rect 469412 389704 469416 389760
rect 469352 389700 469416 389704
rect 469432 389760 469496 389764
rect 469432 389704 469436 389760
rect 469436 389704 469492 389760
rect 469492 389704 469496 389760
rect 469432 389700 469496 389704
rect 469512 389760 469576 389764
rect 469512 389704 469516 389760
rect 469516 389704 469572 389760
rect 469572 389704 469576 389760
rect 469512 389700 469576 389704
rect 481772 389406 481836 389470
rect 489316 389466 489380 389470
rect 489316 389410 489366 389466
rect 489366 389410 489380 389466
rect 489316 389406 489380 389410
rect 474964 389330 475028 389334
rect 474964 389274 474978 389330
rect 474978 389274 475028 389330
rect 474964 389270 475028 389274
rect 478644 389330 478708 389334
rect 478644 389274 478690 389330
rect 478690 389274 478708 389330
rect 478644 389270 478708 389274
rect 470272 388910 470336 388914
rect 470272 388854 470276 388910
rect 470276 388854 470332 388910
rect 470332 388854 470336 388910
rect 470272 388850 470336 388854
rect 470352 388910 470416 388914
rect 470352 388854 470356 388910
rect 470356 388854 470412 388910
rect 470412 388854 470416 388910
rect 470352 388850 470416 388854
rect 470432 388910 470496 388914
rect 470432 388854 470436 388910
rect 470436 388854 470492 388910
rect 470492 388854 470496 388910
rect 470432 388850 470496 388854
rect 470512 388910 470576 388914
rect 470512 388854 470516 388910
rect 470516 388854 470572 388910
rect 470572 388854 470576 388910
rect 470512 388850 470576 388854
rect 470592 388910 470656 388914
rect 470592 388854 470596 388910
rect 470596 388854 470652 388910
rect 470652 388854 470656 388910
rect 470592 388850 470656 388854
rect 470672 388910 470736 388914
rect 470672 388854 470676 388910
rect 470676 388854 470732 388910
rect 470732 388854 470736 388910
rect 470672 388850 470736 388854
rect 470752 388910 470816 388914
rect 470752 388854 470756 388910
rect 470756 388854 470812 388910
rect 470812 388854 470816 388910
rect 470752 388850 470816 388854
rect 470272 388830 470336 388834
rect 470272 388774 470276 388830
rect 470276 388774 470332 388830
rect 470332 388774 470336 388830
rect 470272 388770 470336 388774
rect 470352 388830 470416 388834
rect 470352 388774 470356 388830
rect 470356 388774 470412 388830
rect 470412 388774 470416 388830
rect 470352 388770 470416 388774
rect 470432 388830 470496 388834
rect 470432 388774 470436 388830
rect 470436 388774 470492 388830
rect 470492 388774 470496 388830
rect 470432 388770 470496 388774
rect 470512 388830 470576 388834
rect 470512 388774 470516 388830
rect 470516 388774 470572 388830
rect 470572 388774 470576 388830
rect 470512 388770 470576 388774
rect 470592 388830 470656 388834
rect 470592 388774 470596 388830
rect 470596 388774 470652 388830
rect 470652 388774 470656 388830
rect 470592 388770 470656 388774
rect 470672 388830 470736 388834
rect 470672 388774 470676 388830
rect 470676 388774 470732 388830
rect 470732 388774 470736 388830
rect 470672 388770 470736 388774
rect 470752 388830 470816 388834
rect 470752 388774 470756 388830
rect 470756 388774 470812 388830
rect 470812 388774 470816 388830
rect 470752 388770 470816 388774
rect 470272 388750 470336 388754
rect 470272 388694 470276 388750
rect 470276 388694 470332 388750
rect 470332 388694 470336 388750
rect 470272 388690 470336 388694
rect 470352 388750 470416 388754
rect 470352 388694 470356 388750
rect 470356 388694 470412 388750
rect 470412 388694 470416 388750
rect 470352 388690 470416 388694
rect 470432 388750 470496 388754
rect 470432 388694 470436 388750
rect 470436 388694 470492 388750
rect 470492 388694 470496 388750
rect 470432 388690 470496 388694
rect 470512 388750 470576 388754
rect 470512 388694 470516 388750
rect 470516 388694 470572 388750
rect 470572 388694 470576 388750
rect 470512 388690 470576 388694
rect 470592 388750 470656 388754
rect 470592 388694 470596 388750
rect 470596 388694 470652 388750
rect 470652 388694 470656 388750
rect 470592 388690 470656 388694
rect 470672 388750 470736 388754
rect 470672 388694 470676 388750
rect 470676 388694 470732 388750
rect 470732 388694 470736 388750
rect 470672 388690 470736 388694
rect 470752 388750 470816 388754
rect 470752 388694 470756 388750
rect 470756 388694 470812 388750
rect 470812 388694 470816 388750
rect 470752 388690 470816 388694
rect 470272 388670 470336 388674
rect 470272 388614 470276 388670
rect 470276 388614 470332 388670
rect 470332 388614 470336 388670
rect 470272 388610 470336 388614
rect 470352 388670 470416 388674
rect 470352 388614 470356 388670
rect 470356 388614 470412 388670
rect 470412 388614 470416 388670
rect 470352 388610 470416 388614
rect 470432 388670 470496 388674
rect 470432 388614 470436 388670
rect 470436 388614 470492 388670
rect 470492 388614 470496 388670
rect 470432 388610 470496 388614
rect 470512 388670 470576 388674
rect 470512 388614 470516 388670
rect 470516 388614 470572 388670
rect 470572 388614 470576 388670
rect 470512 388610 470576 388614
rect 470592 388670 470656 388674
rect 470592 388614 470596 388670
rect 470596 388614 470652 388670
rect 470652 388614 470656 388670
rect 470592 388610 470656 388614
rect 470672 388670 470736 388674
rect 470672 388614 470676 388670
rect 470676 388614 470732 388670
rect 470732 388614 470736 388670
rect 470672 388610 470736 388614
rect 470752 388670 470816 388674
rect 470752 388614 470756 388670
rect 470756 388614 470812 388670
rect 470812 388614 470816 388670
rect 470752 388610 470816 388614
rect 486740 386414 486804 386478
rect 577032 379122 577096 379126
rect 577032 379066 577036 379122
rect 577036 379066 577092 379122
rect 577092 379066 577096 379122
rect 577032 379062 577096 379066
rect 577112 379122 577176 379126
rect 577112 379066 577116 379122
rect 577116 379066 577172 379122
rect 577172 379066 577176 379122
rect 577112 379062 577176 379066
rect 577192 379122 577256 379126
rect 577192 379066 577196 379122
rect 577196 379066 577252 379122
rect 577252 379066 577256 379122
rect 577192 379062 577256 379066
rect 577272 379122 577336 379126
rect 577272 379066 577276 379122
rect 577276 379066 577332 379122
rect 577332 379066 577336 379122
rect 577272 379062 577336 379066
rect 577352 379122 577416 379126
rect 577352 379066 577356 379122
rect 577356 379066 577412 379122
rect 577412 379066 577416 379122
rect 577352 379062 577416 379066
rect 577432 379122 577496 379126
rect 577432 379066 577436 379122
rect 577436 379066 577492 379122
rect 577492 379066 577496 379122
rect 577432 379062 577496 379066
rect 577512 379122 577576 379126
rect 577512 379066 577516 379122
rect 577516 379066 577572 379122
rect 577572 379066 577576 379122
rect 577512 379062 577576 379066
rect 577032 379042 577096 379046
rect 577032 378986 577036 379042
rect 577036 378986 577092 379042
rect 577092 378986 577096 379042
rect 577032 378982 577096 378986
rect 577112 379042 577176 379046
rect 577112 378986 577116 379042
rect 577116 378986 577172 379042
rect 577172 378986 577176 379042
rect 577112 378982 577176 378986
rect 577192 379042 577256 379046
rect 577192 378986 577196 379042
rect 577196 378986 577252 379042
rect 577252 378986 577256 379042
rect 577192 378982 577256 378986
rect 577272 379042 577336 379046
rect 577272 378986 577276 379042
rect 577276 378986 577332 379042
rect 577332 378986 577336 379042
rect 577272 378982 577336 378986
rect 577352 379042 577416 379046
rect 577352 378986 577356 379042
rect 577356 378986 577412 379042
rect 577412 378986 577416 379042
rect 577352 378982 577416 378986
rect 577432 379042 577496 379046
rect 577432 378986 577436 379042
rect 577436 378986 577492 379042
rect 577492 378986 577496 379042
rect 577432 378982 577496 378986
rect 577512 379042 577576 379046
rect 577512 378986 577516 379042
rect 577516 378986 577572 379042
rect 577572 378986 577576 379042
rect 577512 378982 577576 378986
rect 577032 378962 577096 378966
rect 577032 378906 577036 378962
rect 577036 378906 577092 378962
rect 577092 378906 577096 378962
rect 577032 378902 577096 378906
rect 577112 378962 577176 378966
rect 577112 378906 577116 378962
rect 577116 378906 577172 378962
rect 577172 378906 577176 378962
rect 577112 378902 577176 378906
rect 577192 378962 577256 378966
rect 577192 378906 577196 378962
rect 577196 378906 577252 378962
rect 577252 378906 577256 378962
rect 577192 378902 577256 378906
rect 577272 378962 577336 378966
rect 577272 378906 577276 378962
rect 577276 378906 577332 378962
rect 577332 378906 577336 378962
rect 577272 378902 577336 378906
rect 577352 378962 577416 378966
rect 577352 378906 577356 378962
rect 577356 378906 577412 378962
rect 577412 378906 577416 378962
rect 577352 378902 577416 378906
rect 577432 378962 577496 378966
rect 577432 378906 577436 378962
rect 577436 378906 577492 378962
rect 577492 378906 577496 378962
rect 577432 378902 577496 378906
rect 577512 378962 577576 378966
rect 577512 378906 577516 378962
rect 577516 378906 577572 378962
rect 577572 378906 577576 378962
rect 577512 378902 577576 378906
rect 577032 378882 577096 378886
rect 577032 378826 577036 378882
rect 577036 378826 577092 378882
rect 577092 378826 577096 378882
rect 577032 378822 577096 378826
rect 577112 378882 577176 378886
rect 577112 378826 577116 378882
rect 577116 378826 577172 378882
rect 577172 378826 577176 378882
rect 577112 378822 577176 378826
rect 577192 378882 577256 378886
rect 577192 378826 577196 378882
rect 577196 378826 577252 378882
rect 577252 378826 577256 378882
rect 577192 378822 577256 378826
rect 577272 378882 577336 378886
rect 577272 378826 577276 378882
rect 577276 378826 577332 378882
rect 577332 378826 577336 378882
rect 577272 378822 577336 378826
rect 577352 378882 577416 378886
rect 577352 378826 577356 378882
rect 577356 378826 577412 378882
rect 577412 378826 577416 378882
rect 577352 378822 577416 378826
rect 577432 378882 577496 378886
rect 577432 378826 577436 378882
rect 577436 378826 577492 378882
rect 577492 378826 577496 378882
rect 577432 378822 577496 378826
rect 577512 378882 577576 378886
rect 577512 378826 577516 378882
rect 577516 378826 577572 378882
rect 577572 378826 577576 378882
rect 577512 378822 577576 378826
rect 578272 378327 578336 378331
rect 578272 378271 578276 378327
rect 578276 378271 578332 378327
rect 578332 378271 578336 378327
rect 578272 378267 578336 378271
rect 578352 378327 578416 378331
rect 578352 378271 578356 378327
rect 578356 378271 578412 378327
rect 578412 378271 578416 378327
rect 578352 378267 578416 378271
rect 578432 378327 578496 378331
rect 578432 378271 578436 378327
rect 578436 378271 578492 378327
rect 578492 378271 578496 378327
rect 578432 378267 578496 378271
rect 578512 378327 578576 378331
rect 578512 378271 578516 378327
rect 578516 378271 578572 378327
rect 578572 378271 578576 378327
rect 578512 378267 578576 378271
rect 578592 378327 578656 378331
rect 578592 378271 578596 378327
rect 578596 378271 578652 378327
rect 578652 378271 578656 378327
rect 578592 378267 578656 378271
rect 578672 378327 578736 378331
rect 578672 378271 578676 378327
rect 578676 378271 578732 378327
rect 578732 378271 578736 378327
rect 578672 378267 578736 378271
rect 578752 378327 578816 378331
rect 578752 378271 578756 378327
rect 578756 378271 578812 378327
rect 578812 378271 578816 378327
rect 578752 378267 578816 378271
rect 578272 378247 578336 378251
rect 578272 378191 578276 378247
rect 578276 378191 578332 378247
rect 578332 378191 578336 378247
rect 578272 378187 578336 378191
rect 578352 378247 578416 378251
rect 578352 378191 578356 378247
rect 578356 378191 578412 378247
rect 578412 378191 578416 378247
rect 578352 378187 578416 378191
rect 578432 378247 578496 378251
rect 578432 378191 578436 378247
rect 578436 378191 578492 378247
rect 578492 378191 578496 378247
rect 578432 378187 578496 378191
rect 578512 378247 578576 378251
rect 578512 378191 578516 378247
rect 578516 378191 578572 378247
rect 578572 378191 578576 378247
rect 578512 378187 578576 378191
rect 578592 378247 578656 378251
rect 578592 378191 578596 378247
rect 578596 378191 578652 378247
rect 578652 378191 578656 378247
rect 578592 378187 578656 378191
rect 578672 378247 578736 378251
rect 578672 378191 578676 378247
rect 578676 378191 578732 378247
rect 578732 378191 578736 378247
rect 578672 378187 578736 378191
rect 578752 378247 578816 378251
rect 578752 378191 578756 378247
rect 578756 378191 578812 378247
rect 578812 378191 578816 378247
rect 578752 378187 578816 378191
rect 578272 378167 578336 378171
rect 578272 378111 578276 378167
rect 578276 378111 578332 378167
rect 578332 378111 578336 378167
rect 578272 378107 578336 378111
rect 578352 378167 578416 378171
rect 578352 378111 578356 378167
rect 578356 378111 578412 378167
rect 578412 378111 578416 378167
rect 578352 378107 578416 378111
rect 578432 378167 578496 378171
rect 578432 378111 578436 378167
rect 578436 378111 578492 378167
rect 578492 378111 578496 378167
rect 578432 378107 578496 378111
rect 578512 378167 578576 378171
rect 578512 378111 578516 378167
rect 578516 378111 578572 378167
rect 578572 378111 578576 378167
rect 578512 378107 578576 378111
rect 578592 378167 578656 378171
rect 578592 378111 578596 378167
rect 578596 378111 578652 378167
rect 578652 378111 578656 378167
rect 578592 378107 578656 378111
rect 578672 378167 578736 378171
rect 578672 378111 578676 378167
rect 578676 378111 578732 378167
rect 578732 378111 578736 378167
rect 578672 378107 578736 378111
rect 578752 378167 578816 378171
rect 578752 378111 578756 378167
rect 578756 378111 578812 378167
rect 578812 378111 578816 378167
rect 578752 378107 578816 378111
rect 578272 378087 578336 378091
rect 578272 378031 578276 378087
rect 578276 378031 578332 378087
rect 578332 378031 578336 378087
rect 578272 378027 578336 378031
rect 578352 378087 578416 378091
rect 578352 378031 578356 378087
rect 578356 378031 578412 378087
rect 578412 378031 578416 378087
rect 578352 378027 578416 378031
rect 578432 378087 578496 378091
rect 578432 378031 578436 378087
rect 578436 378031 578492 378087
rect 578492 378031 578496 378087
rect 578432 378027 578496 378031
rect 578512 378087 578576 378091
rect 578512 378031 578516 378087
rect 578516 378031 578572 378087
rect 578572 378031 578576 378087
rect 578512 378027 578576 378031
rect 578592 378087 578656 378091
rect 578592 378031 578596 378087
rect 578596 378031 578652 378087
rect 578652 378031 578656 378087
rect 578592 378027 578656 378031
rect 578672 378087 578736 378091
rect 578672 378031 578676 378087
rect 578676 378031 578732 378087
rect 578732 378031 578736 378087
rect 578672 378027 578736 378031
rect 578752 378087 578816 378091
rect 578752 378031 578756 378087
rect 578756 378031 578812 378087
rect 578812 378031 578816 378087
rect 578752 378027 578816 378031
rect 541572 373086 541636 373150
rect 544332 373086 544396 373150
rect 482876 370094 482940 370158
rect 470272 358483 470336 358487
rect 470272 358427 470276 358483
rect 470276 358427 470332 358483
rect 470332 358427 470336 358483
rect 470272 358423 470336 358427
rect 470352 358483 470416 358487
rect 470352 358427 470356 358483
rect 470356 358427 470412 358483
rect 470412 358427 470416 358483
rect 470352 358423 470416 358427
rect 470432 358483 470496 358487
rect 470432 358427 470436 358483
rect 470436 358427 470492 358483
rect 470492 358427 470496 358483
rect 470432 358423 470496 358427
rect 470512 358483 470576 358487
rect 470512 358427 470516 358483
rect 470516 358427 470572 358483
rect 470572 358427 470576 358483
rect 470512 358423 470576 358427
rect 470592 358483 470656 358487
rect 470592 358427 470596 358483
rect 470596 358427 470652 358483
rect 470652 358427 470656 358483
rect 470592 358423 470656 358427
rect 470672 358483 470736 358487
rect 470672 358427 470676 358483
rect 470676 358427 470732 358483
rect 470732 358427 470736 358483
rect 470672 358423 470736 358427
rect 470752 358483 470816 358487
rect 470752 358427 470756 358483
rect 470756 358427 470812 358483
rect 470812 358427 470816 358483
rect 470752 358423 470816 358427
rect 470272 358403 470336 358407
rect 470272 358347 470276 358403
rect 470276 358347 470332 358403
rect 470332 358347 470336 358403
rect 470272 358343 470336 358347
rect 470352 358403 470416 358407
rect 470352 358347 470356 358403
rect 470356 358347 470412 358403
rect 470412 358347 470416 358403
rect 470352 358343 470416 358347
rect 470432 358403 470496 358407
rect 470432 358347 470436 358403
rect 470436 358347 470492 358403
rect 470492 358347 470496 358403
rect 470432 358343 470496 358347
rect 470512 358403 470576 358407
rect 470512 358347 470516 358403
rect 470516 358347 470572 358403
rect 470572 358347 470576 358403
rect 470512 358343 470576 358347
rect 470592 358403 470656 358407
rect 470592 358347 470596 358403
rect 470596 358347 470652 358403
rect 470652 358347 470656 358403
rect 470592 358343 470656 358347
rect 470672 358403 470736 358407
rect 470672 358347 470676 358403
rect 470676 358347 470732 358403
rect 470732 358347 470736 358403
rect 470672 358343 470736 358347
rect 470752 358403 470816 358407
rect 470752 358347 470756 358403
rect 470756 358347 470812 358403
rect 470812 358347 470816 358403
rect 470752 358343 470816 358347
rect 470272 358323 470336 358327
rect 470272 358267 470276 358323
rect 470276 358267 470332 358323
rect 470332 358267 470336 358323
rect 470272 358263 470336 358267
rect 470352 358323 470416 358327
rect 470352 358267 470356 358323
rect 470356 358267 470412 358323
rect 470412 358267 470416 358323
rect 470352 358263 470416 358267
rect 470432 358323 470496 358327
rect 470432 358267 470436 358323
rect 470436 358267 470492 358323
rect 470492 358267 470496 358323
rect 470432 358263 470496 358267
rect 470512 358323 470576 358327
rect 470512 358267 470516 358323
rect 470516 358267 470572 358323
rect 470572 358267 470576 358323
rect 470512 358263 470576 358267
rect 470592 358323 470656 358327
rect 470592 358267 470596 358323
rect 470596 358267 470652 358323
rect 470652 358267 470656 358323
rect 470592 358263 470656 358267
rect 470672 358323 470736 358327
rect 470672 358267 470676 358323
rect 470676 358267 470732 358323
rect 470732 358267 470736 358323
rect 470672 358263 470736 358267
rect 470752 358323 470816 358327
rect 470752 358267 470756 358323
rect 470756 358267 470812 358323
rect 470812 358267 470816 358323
rect 470752 358263 470816 358267
rect 470272 358243 470336 358247
rect 470272 358187 470276 358243
rect 470276 358187 470332 358243
rect 470332 358187 470336 358243
rect 470272 358183 470336 358187
rect 470352 358243 470416 358247
rect 470352 358187 470356 358243
rect 470356 358187 470412 358243
rect 470412 358187 470416 358243
rect 470352 358183 470416 358187
rect 470432 358243 470496 358247
rect 470432 358187 470436 358243
rect 470436 358187 470492 358243
rect 470492 358187 470496 358243
rect 470432 358183 470496 358187
rect 470512 358243 470576 358247
rect 470512 358187 470516 358243
rect 470516 358187 470572 358243
rect 470572 358187 470576 358243
rect 470512 358183 470576 358187
rect 470592 358243 470656 358247
rect 470592 358187 470596 358243
rect 470596 358187 470652 358243
rect 470652 358187 470656 358243
rect 470592 358183 470656 358187
rect 470672 358243 470736 358247
rect 470672 358187 470676 358243
rect 470676 358187 470732 358243
rect 470732 358187 470736 358243
rect 470672 358183 470736 358187
rect 470752 358243 470816 358247
rect 470752 358187 470756 358243
rect 470756 358187 470812 358243
rect 470812 358187 470816 358243
rect 470752 358183 470816 358187
rect 478644 357990 478708 358054
rect 481772 358050 481836 358054
rect 481772 357994 481822 358050
rect 481822 357994 481836 358050
rect 481772 357990 481836 357994
rect 484900 358050 484964 358054
rect 484900 357994 484950 358050
rect 484950 357994 484964 358050
rect 484900 357990 484964 357994
rect 488396 358050 488460 358054
rect 488396 357994 488446 358050
rect 488446 357994 488460 358050
rect 488396 357990 488460 357994
rect 489316 357990 489380 358054
rect 474964 357506 475028 357510
rect 474964 357450 475014 357506
rect 475014 357450 475028 357506
rect 474964 357446 475028 357450
rect 469032 357397 469096 357401
rect 469032 357341 469036 357397
rect 469036 357341 469092 357397
rect 469092 357341 469096 357397
rect 469032 357337 469096 357341
rect 469112 357397 469176 357401
rect 469112 357341 469116 357397
rect 469116 357341 469172 357397
rect 469172 357341 469176 357397
rect 469112 357337 469176 357341
rect 469192 357397 469256 357401
rect 469192 357341 469196 357397
rect 469196 357341 469252 357397
rect 469252 357341 469256 357397
rect 469192 357337 469256 357341
rect 469272 357397 469336 357401
rect 469272 357341 469276 357397
rect 469276 357341 469332 357397
rect 469332 357341 469336 357397
rect 469272 357337 469336 357341
rect 469352 357397 469416 357401
rect 469352 357341 469356 357397
rect 469356 357341 469412 357397
rect 469412 357341 469416 357397
rect 469352 357337 469416 357341
rect 469432 357397 469496 357401
rect 469432 357341 469436 357397
rect 469436 357341 469492 357397
rect 469492 357341 469496 357397
rect 469432 357337 469496 357341
rect 469512 357397 469576 357401
rect 469512 357341 469516 357397
rect 469516 357341 469572 357397
rect 469572 357341 469576 357397
rect 469512 357337 469576 357341
rect 469032 357317 469096 357321
rect 469032 357261 469036 357317
rect 469036 357261 469092 357317
rect 469092 357261 469096 357317
rect 469032 357257 469096 357261
rect 469112 357317 469176 357321
rect 469112 357261 469116 357317
rect 469116 357261 469172 357317
rect 469172 357261 469176 357317
rect 469112 357257 469176 357261
rect 469192 357317 469256 357321
rect 469192 357261 469196 357317
rect 469196 357261 469252 357317
rect 469252 357261 469256 357317
rect 469192 357257 469256 357261
rect 469272 357317 469336 357321
rect 469272 357261 469276 357317
rect 469276 357261 469332 357317
rect 469332 357261 469336 357317
rect 469272 357257 469336 357261
rect 469352 357317 469416 357321
rect 469352 357261 469356 357317
rect 469356 357261 469412 357317
rect 469412 357261 469416 357317
rect 469352 357257 469416 357261
rect 469432 357317 469496 357321
rect 469432 357261 469436 357317
rect 469436 357261 469492 357317
rect 469492 357261 469496 357317
rect 469432 357257 469496 357261
rect 469512 357317 469576 357321
rect 469512 357261 469516 357317
rect 469516 357261 469572 357317
rect 469572 357261 469576 357317
rect 469512 357257 469576 357261
rect 469032 357237 469096 357241
rect 469032 357181 469036 357237
rect 469036 357181 469092 357237
rect 469092 357181 469096 357237
rect 469032 357177 469096 357181
rect 469112 357237 469176 357241
rect 469112 357181 469116 357237
rect 469116 357181 469172 357237
rect 469172 357181 469176 357237
rect 469112 357177 469176 357181
rect 469192 357237 469256 357241
rect 469192 357181 469196 357237
rect 469196 357181 469252 357237
rect 469252 357181 469256 357237
rect 469192 357177 469256 357181
rect 469272 357237 469336 357241
rect 469272 357181 469276 357237
rect 469276 357181 469332 357237
rect 469332 357181 469336 357237
rect 469272 357177 469336 357181
rect 469352 357237 469416 357241
rect 469352 357181 469356 357237
rect 469356 357181 469412 357237
rect 469412 357181 469416 357237
rect 469352 357177 469416 357181
rect 469432 357237 469496 357241
rect 469432 357181 469436 357237
rect 469436 357181 469492 357237
rect 469492 357181 469496 357237
rect 469432 357177 469496 357181
rect 469512 357237 469576 357241
rect 469512 357181 469516 357237
rect 469516 357181 469572 357237
rect 469572 357181 469576 357237
rect 469512 357177 469576 357181
rect 469032 357157 469096 357161
rect 469032 357101 469036 357157
rect 469036 357101 469092 357157
rect 469092 357101 469096 357157
rect 469032 357097 469096 357101
rect 469112 357157 469176 357161
rect 469112 357101 469116 357157
rect 469116 357101 469172 357157
rect 469172 357101 469176 357157
rect 469112 357097 469176 357101
rect 469192 357157 469256 357161
rect 469192 357101 469196 357157
rect 469196 357101 469252 357157
rect 469252 357101 469256 357157
rect 469192 357097 469256 357101
rect 469272 357157 469336 357161
rect 469272 357101 469276 357157
rect 469276 357101 469332 357157
rect 469332 357101 469336 357157
rect 469272 357097 469336 357101
rect 469352 357157 469416 357161
rect 469352 357101 469356 357157
rect 469356 357101 469412 357157
rect 469412 357101 469416 357157
rect 469352 357097 469416 357101
rect 469432 357157 469496 357161
rect 469432 357101 469436 357157
rect 469436 357101 469492 357157
rect 469492 357101 469496 357157
rect 469432 357097 469496 357101
rect 469512 357157 469576 357161
rect 469512 357101 469516 357157
rect 469516 357101 469572 357157
rect 469572 357101 469576 357157
rect 469512 357097 469576 357101
rect 470272 356310 470336 356314
rect 470272 356254 470276 356310
rect 470276 356254 470332 356310
rect 470332 356254 470336 356310
rect 470272 356250 470336 356254
rect 470352 356310 470416 356314
rect 470352 356254 470356 356310
rect 470356 356254 470412 356310
rect 470412 356254 470416 356310
rect 470352 356250 470416 356254
rect 470432 356310 470496 356314
rect 470432 356254 470436 356310
rect 470436 356254 470492 356310
rect 470492 356254 470496 356310
rect 470432 356250 470496 356254
rect 470512 356310 470576 356314
rect 470512 356254 470516 356310
rect 470516 356254 470572 356310
rect 470572 356254 470576 356310
rect 470512 356250 470576 356254
rect 470592 356310 470656 356314
rect 470592 356254 470596 356310
rect 470596 356254 470652 356310
rect 470652 356254 470656 356310
rect 470592 356250 470656 356254
rect 470672 356310 470736 356314
rect 470672 356254 470676 356310
rect 470676 356254 470732 356310
rect 470732 356254 470736 356310
rect 470672 356250 470736 356254
rect 470752 356310 470816 356314
rect 470752 356254 470756 356310
rect 470756 356254 470812 356310
rect 470812 356254 470816 356310
rect 470752 356250 470816 356254
rect 470272 356230 470336 356234
rect 470272 356174 470276 356230
rect 470276 356174 470332 356230
rect 470332 356174 470336 356230
rect 470272 356170 470336 356174
rect 470352 356230 470416 356234
rect 470352 356174 470356 356230
rect 470356 356174 470412 356230
rect 470412 356174 470416 356230
rect 470352 356170 470416 356174
rect 470432 356230 470496 356234
rect 470432 356174 470436 356230
rect 470436 356174 470492 356230
rect 470492 356174 470496 356230
rect 470432 356170 470496 356174
rect 470512 356230 470576 356234
rect 470512 356174 470516 356230
rect 470516 356174 470572 356230
rect 470572 356174 470576 356230
rect 470512 356170 470576 356174
rect 470592 356230 470656 356234
rect 470592 356174 470596 356230
rect 470596 356174 470652 356230
rect 470652 356174 470656 356230
rect 470592 356170 470656 356174
rect 470672 356230 470736 356234
rect 470672 356174 470676 356230
rect 470676 356174 470732 356230
rect 470732 356174 470736 356230
rect 470672 356170 470736 356174
rect 470752 356230 470816 356234
rect 470752 356174 470756 356230
rect 470756 356174 470812 356230
rect 470812 356174 470816 356230
rect 470752 356170 470816 356174
rect 470272 356150 470336 356154
rect 470272 356094 470276 356150
rect 470276 356094 470332 356150
rect 470332 356094 470336 356150
rect 470272 356090 470336 356094
rect 470352 356150 470416 356154
rect 470352 356094 470356 356150
rect 470356 356094 470412 356150
rect 470412 356094 470416 356150
rect 470352 356090 470416 356094
rect 470432 356150 470496 356154
rect 470432 356094 470436 356150
rect 470436 356094 470492 356150
rect 470492 356094 470496 356150
rect 470432 356090 470496 356094
rect 470512 356150 470576 356154
rect 470512 356094 470516 356150
rect 470516 356094 470572 356150
rect 470572 356094 470576 356150
rect 470512 356090 470576 356094
rect 470592 356150 470656 356154
rect 470592 356094 470596 356150
rect 470596 356094 470652 356150
rect 470652 356094 470656 356150
rect 470592 356090 470656 356094
rect 470672 356150 470736 356154
rect 470672 356094 470676 356150
rect 470676 356094 470732 356150
rect 470732 356094 470736 356150
rect 470672 356090 470736 356094
rect 470752 356150 470816 356154
rect 470752 356094 470756 356150
rect 470756 356094 470812 356150
rect 470812 356094 470816 356150
rect 470752 356090 470816 356094
rect 470272 356070 470336 356074
rect 470272 356014 470276 356070
rect 470276 356014 470332 356070
rect 470332 356014 470336 356070
rect 470272 356010 470336 356014
rect 470352 356070 470416 356074
rect 470352 356014 470356 356070
rect 470356 356014 470412 356070
rect 470412 356014 470416 356070
rect 470352 356010 470416 356014
rect 470432 356070 470496 356074
rect 470432 356014 470436 356070
rect 470436 356014 470492 356070
rect 470492 356014 470496 356070
rect 470432 356010 470496 356014
rect 470512 356070 470576 356074
rect 470512 356014 470516 356070
rect 470516 356014 470572 356070
rect 470572 356014 470576 356070
rect 470512 356010 470576 356014
rect 470592 356070 470656 356074
rect 470592 356014 470596 356070
rect 470596 356014 470652 356070
rect 470652 356014 470656 356070
rect 470592 356010 470656 356014
rect 470672 356070 470736 356074
rect 470672 356014 470676 356070
rect 470676 356014 470732 356070
rect 470732 356014 470736 356070
rect 470672 356010 470736 356014
rect 470752 356070 470816 356074
rect 470752 356014 470756 356070
rect 470756 356014 470812 356070
rect 470812 356014 470816 356070
rect 470752 356010 470816 356014
rect 485452 351870 485516 351934
rect 473676 343710 473740 343774
rect 474964 343710 475028 343774
rect 470272 342482 470336 342486
rect 470272 342426 470276 342482
rect 470276 342426 470332 342482
rect 470332 342426 470336 342482
rect 470272 342422 470336 342426
rect 470352 342482 470416 342486
rect 470352 342426 470356 342482
rect 470356 342426 470412 342482
rect 470412 342426 470416 342482
rect 470352 342422 470416 342426
rect 470432 342482 470496 342486
rect 470432 342426 470436 342482
rect 470436 342426 470492 342482
rect 470492 342426 470496 342482
rect 470432 342422 470496 342426
rect 470512 342482 470576 342486
rect 470512 342426 470516 342482
rect 470516 342426 470572 342482
rect 470572 342426 470576 342482
rect 470512 342422 470576 342426
rect 470592 342482 470656 342486
rect 470592 342426 470596 342482
rect 470596 342426 470652 342482
rect 470652 342426 470656 342482
rect 470592 342422 470656 342426
rect 470672 342482 470736 342486
rect 470672 342426 470676 342482
rect 470676 342426 470732 342482
rect 470732 342426 470736 342482
rect 470672 342422 470736 342426
rect 470752 342482 470816 342486
rect 470752 342426 470756 342482
rect 470756 342426 470812 342482
rect 470812 342426 470816 342482
rect 470752 342422 470816 342426
rect 470272 342402 470336 342406
rect 470272 342346 470276 342402
rect 470276 342346 470332 342402
rect 470332 342346 470336 342402
rect 470272 342342 470336 342346
rect 470352 342402 470416 342406
rect 470352 342346 470356 342402
rect 470356 342346 470412 342402
rect 470412 342346 470416 342402
rect 470352 342342 470416 342346
rect 470432 342402 470496 342406
rect 470432 342346 470436 342402
rect 470436 342346 470492 342402
rect 470492 342346 470496 342402
rect 470432 342342 470496 342346
rect 470512 342402 470576 342406
rect 470512 342346 470516 342402
rect 470516 342346 470572 342402
rect 470572 342346 470576 342402
rect 470512 342342 470576 342346
rect 470592 342402 470656 342406
rect 470592 342346 470596 342402
rect 470596 342346 470652 342402
rect 470652 342346 470656 342402
rect 470592 342342 470656 342346
rect 470672 342402 470736 342406
rect 470672 342346 470676 342402
rect 470676 342346 470732 342402
rect 470732 342346 470736 342402
rect 470672 342342 470736 342346
rect 470752 342402 470816 342406
rect 470752 342346 470756 342402
rect 470756 342346 470812 342402
rect 470812 342346 470816 342402
rect 470752 342342 470816 342346
rect 470272 342322 470336 342326
rect 470272 342266 470276 342322
rect 470276 342266 470332 342322
rect 470332 342266 470336 342322
rect 470272 342262 470336 342266
rect 470352 342322 470416 342326
rect 470352 342266 470356 342322
rect 470356 342266 470412 342322
rect 470412 342266 470416 342322
rect 470352 342262 470416 342266
rect 470432 342322 470496 342326
rect 470432 342266 470436 342322
rect 470436 342266 470492 342322
rect 470492 342266 470496 342322
rect 470432 342262 470496 342266
rect 470512 342322 470576 342326
rect 470512 342266 470516 342322
rect 470516 342266 470572 342322
rect 470572 342266 470576 342322
rect 470512 342262 470576 342266
rect 470592 342322 470656 342326
rect 470592 342266 470596 342322
rect 470596 342266 470652 342322
rect 470652 342266 470656 342322
rect 470592 342262 470656 342266
rect 470672 342322 470736 342326
rect 470672 342266 470676 342322
rect 470676 342266 470732 342322
rect 470732 342266 470736 342322
rect 470672 342262 470736 342266
rect 470752 342322 470816 342326
rect 470752 342266 470756 342322
rect 470756 342266 470812 342322
rect 470812 342266 470816 342322
rect 470752 342262 470816 342266
rect 470272 342242 470336 342246
rect 470272 342186 470276 342242
rect 470276 342186 470332 342242
rect 470332 342186 470336 342242
rect 470272 342182 470336 342186
rect 470352 342242 470416 342246
rect 470352 342186 470356 342242
rect 470356 342186 470412 342242
rect 470412 342186 470416 342242
rect 470352 342182 470416 342186
rect 470432 342242 470496 342246
rect 470432 342186 470436 342242
rect 470436 342186 470492 342242
rect 470492 342186 470496 342242
rect 470432 342182 470496 342186
rect 470512 342242 470576 342246
rect 470512 342186 470516 342242
rect 470516 342186 470572 342242
rect 470572 342186 470576 342242
rect 470512 342182 470576 342186
rect 470592 342242 470656 342246
rect 470592 342186 470596 342242
rect 470596 342186 470652 342242
rect 470652 342186 470656 342242
rect 470592 342182 470656 342186
rect 470672 342242 470736 342246
rect 470672 342186 470676 342242
rect 470676 342186 470732 342242
rect 470732 342186 470736 342242
rect 470672 342182 470736 342186
rect 470752 342242 470816 342246
rect 470752 342186 470756 342242
rect 470756 342186 470812 342242
rect 470812 342186 470816 342242
rect 470752 342182 470816 342186
rect 469032 341395 469096 341399
rect 469032 341339 469036 341395
rect 469036 341339 469092 341395
rect 469092 341339 469096 341395
rect 469032 341335 469096 341339
rect 469112 341395 469176 341399
rect 469112 341339 469116 341395
rect 469116 341339 469172 341395
rect 469172 341339 469176 341395
rect 469112 341335 469176 341339
rect 469192 341395 469256 341399
rect 469192 341339 469196 341395
rect 469196 341339 469252 341395
rect 469252 341339 469256 341395
rect 469192 341335 469256 341339
rect 469272 341395 469336 341399
rect 469272 341339 469276 341395
rect 469276 341339 469332 341395
rect 469332 341339 469336 341395
rect 469272 341335 469336 341339
rect 469352 341395 469416 341399
rect 469352 341339 469356 341395
rect 469356 341339 469412 341395
rect 469412 341339 469416 341395
rect 469352 341335 469416 341339
rect 469432 341395 469496 341399
rect 469432 341339 469436 341395
rect 469436 341339 469492 341395
rect 469492 341339 469496 341395
rect 469432 341335 469496 341339
rect 469512 341395 469576 341399
rect 469512 341339 469516 341395
rect 469516 341339 469572 341395
rect 469572 341339 469576 341395
rect 469512 341335 469576 341339
rect 469032 341315 469096 341319
rect 469032 341259 469036 341315
rect 469036 341259 469092 341315
rect 469092 341259 469096 341315
rect 469032 341255 469096 341259
rect 469112 341315 469176 341319
rect 469112 341259 469116 341315
rect 469116 341259 469172 341315
rect 469172 341259 469176 341315
rect 469112 341255 469176 341259
rect 469192 341315 469256 341319
rect 469192 341259 469196 341315
rect 469196 341259 469252 341315
rect 469252 341259 469256 341315
rect 469192 341255 469256 341259
rect 469272 341315 469336 341319
rect 469272 341259 469276 341315
rect 469276 341259 469332 341315
rect 469332 341259 469336 341315
rect 469272 341255 469336 341259
rect 469352 341315 469416 341319
rect 469352 341259 469356 341315
rect 469356 341259 469412 341315
rect 469412 341259 469416 341315
rect 469352 341255 469416 341259
rect 469432 341315 469496 341319
rect 469432 341259 469436 341315
rect 469436 341259 469492 341315
rect 469492 341259 469496 341315
rect 469432 341255 469496 341259
rect 469512 341315 469576 341319
rect 469512 341259 469516 341315
rect 469516 341259 469572 341315
rect 469572 341259 469576 341315
rect 469512 341255 469576 341259
rect 469032 341235 469096 341239
rect 469032 341179 469036 341235
rect 469036 341179 469092 341235
rect 469092 341179 469096 341235
rect 469032 341175 469096 341179
rect 469112 341235 469176 341239
rect 469112 341179 469116 341235
rect 469116 341179 469172 341235
rect 469172 341179 469176 341235
rect 469112 341175 469176 341179
rect 469192 341235 469256 341239
rect 469192 341179 469196 341235
rect 469196 341179 469252 341235
rect 469252 341179 469256 341235
rect 469192 341175 469256 341179
rect 469272 341235 469336 341239
rect 469272 341179 469276 341235
rect 469276 341179 469332 341235
rect 469332 341179 469336 341235
rect 469272 341175 469336 341179
rect 469352 341235 469416 341239
rect 469352 341179 469356 341235
rect 469356 341179 469412 341235
rect 469412 341179 469416 341235
rect 469352 341175 469416 341179
rect 469432 341235 469496 341239
rect 469432 341179 469436 341235
rect 469436 341179 469492 341235
rect 469492 341179 469496 341235
rect 469432 341175 469496 341179
rect 469512 341235 469576 341239
rect 469512 341179 469516 341235
rect 469516 341179 469572 341235
rect 469572 341179 469576 341235
rect 469512 341175 469576 341179
rect 469032 341155 469096 341159
rect 469032 341099 469036 341155
rect 469036 341099 469092 341155
rect 469092 341099 469096 341155
rect 469032 341095 469096 341099
rect 469112 341155 469176 341159
rect 469112 341099 469116 341155
rect 469116 341099 469172 341155
rect 469172 341099 469176 341155
rect 469112 341095 469176 341099
rect 469192 341155 469256 341159
rect 469192 341099 469196 341155
rect 469196 341099 469252 341155
rect 469252 341099 469256 341155
rect 469192 341095 469256 341099
rect 469272 341155 469336 341159
rect 469272 341099 469276 341155
rect 469276 341099 469332 341155
rect 469332 341099 469336 341155
rect 469272 341095 469336 341099
rect 469352 341155 469416 341159
rect 469352 341099 469356 341155
rect 469356 341099 469412 341155
rect 469412 341099 469416 341155
rect 469352 341095 469416 341099
rect 469432 341155 469496 341159
rect 469432 341099 469436 341155
rect 469436 341099 469492 341155
rect 469492 341099 469496 341155
rect 469432 341095 469496 341099
rect 469512 341155 469576 341159
rect 469512 341099 469516 341155
rect 469516 341099 469572 341155
rect 469572 341099 469576 341155
rect 469512 341095 469576 341099
rect 478460 340990 478524 341054
rect 481404 340990 481468 341054
rect 488028 340990 488092 341054
rect 473676 340446 473740 340510
rect 470272 340310 470336 340314
rect 470272 340254 470276 340310
rect 470276 340254 470332 340310
rect 470332 340254 470336 340310
rect 470272 340250 470336 340254
rect 470352 340310 470416 340314
rect 470352 340254 470356 340310
rect 470356 340254 470412 340310
rect 470412 340254 470416 340310
rect 470352 340250 470416 340254
rect 470432 340310 470496 340314
rect 470432 340254 470436 340310
rect 470436 340254 470492 340310
rect 470492 340254 470496 340310
rect 470432 340250 470496 340254
rect 470512 340310 470576 340314
rect 470512 340254 470516 340310
rect 470516 340254 470572 340310
rect 470572 340254 470576 340310
rect 470512 340250 470576 340254
rect 470592 340310 470656 340314
rect 470592 340254 470596 340310
rect 470596 340254 470652 340310
rect 470652 340254 470656 340310
rect 470592 340250 470656 340254
rect 470672 340310 470736 340314
rect 470672 340254 470676 340310
rect 470676 340254 470732 340310
rect 470732 340254 470736 340310
rect 470672 340250 470736 340254
rect 470752 340310 470816 340314
rect 470752 340254 470756 340310
rect 470756 340254 470812 340310
rect 470812 340254 470816 340310
rect 470752 340250 470816 340254
rect 470272 340230 470336 340234
rect 470272 340174 470276 340230
rect 470276 340174 470332 340230
rect 470332 340174 470336 340230
rect 470272 340170 470336 340174
rect 470352 340230 470416 340234
rect 470352 340174 470356 340230
rect 470356 340174 470412 340230
rect 470412 340174 470416 340230
rect 470352 340170 470416 340174
rect 470432 340230 470496 340234
rect 470432 340174 470436 340230
rect 470436 340174 470492 340230
rect 470492 340174 470496 340230
rect 470432 340170 470496 340174
rect 470512 340230 470576 340234
rect 470512 340174 470516 340230
rect 470516 340174 470572 340230
rect 470572 340174 470576 340230
rect 470512 340170 470576 340174
rect 470592 340230 470656 340234
rect 470592 340174 470596 340230
rect 470596 340174 470652 340230
rect 470652 340174 470656 340230
rect 470592 340170 470656 340174
rect 470672 340230 470736 340234
rect 470672 340174 470676 340230
rect 470676 340174 470732 340230
rect 470732 340174 470736 340230
rect 470672 340170 470736 340174
rect 470752 340230 470816 340234
rect 470752 340174 470756 340230
rect 470756 340174 470812 340230
rect 470812 340174 470816 340230
rect 470752 340170 470816 340174
rect 470272 340150 470336 340154
rect 470272 340094 470276 340150
rect 470276 340094 470332 340150
rect 470332 340094 470336 340150
rect 470272 340090 470336 340094
rect 470352 340150 470416 340154
rect 470352 340094 470356 340150
rect 470356 340094 470412 340150
rect 470412 340094 470416 340150
rect 470352 340090 470416 340094
rect 470432 340150 470496 340154
rect 470432 340094 470436 340150
rect 470436 340094 470492 340150
rect 470492 340094 470496 340150
rect 470432 340090 470496 340094
rect 470512 340150 470576 340154
rect 470512 340094 470516 340150
rect 470516 340094 470572 340150
rect 470572 340094 470576 340150
rect 470512 340090 470576 340094
rect 470592 340150 470656 340154
rect 470592 340094 470596 340150
rect 470596 340094 470652 340150
rect 470652 340094 470656 340150
rect 470592 340090 470656 340094
rect 470672 340150 470736 340154
rect 470672 340094 470676 340150
rect 470676 340094 470732 340150
rect 470732 340094 470736 340150
rect 470672 340090 470736 340094
rect 470752 340150 470816 340154
rect 470752 340094 470756 340150
rect 470756 340094 470812 340150
rect 470812 340094 470816 340150
rect 470752 340090 470816 340094
rect 470272 340070 470336 340074
rect 470272 340014 470276 340070
rect 470276 340014 470332 340070
rect 470332 340014 470336 340070
rect 470272 340010 470336 340014
rect 470352 340070 470416 340074
rect 470352 340014 470356 340070
rect 470356 340014 470412 340070
rect 470412 340014 470416 340070
rect 470352 340010 470416 340014
rect 470432 340070 470496 340074
rect 470432 340014 470436 340070
rect 470436 340014 470492 340070
rect 470492 340014 470496 340070
rect 470432 340010 470496 340014
rect 470512 340070 470576 340074
rect 470512 340014 470516 340070
rect 470516 340014 470572 340070
rect 470572 340014 470576 340070
rect 470512 340010 470576 340014
rect 470592 340070 470656 340074
rect 470592 340014 470596 340070
rect 470596 340014 470652 340070
rect 470652 340014 470656 340070
rect 470592 340010 470656 340014
rect 470672 340070 470736 340074
rect 470672 340014 470676 340070
rect 470676 340014 470732 340070
rect 470732 340014 470736 340070
rect 470672 340010 470736 340014
rect 470752 340070 470816 340074
rect 470752 340014 470756 340070
rect 470756 340014 470812 340070
rect 470812 340014 470816 340070
rect 470752 340010 470816 340014
rect 541572 339494 541636 339558
rect 544332 339494 544396 339558
rect 486556 335414 486620 335478
rect 485636 334054 485700 334118
rect 486740 332694 486804 332758
rect 577032 325946 577096 325950
rect 577032 325890 577036 325946
rect 577036 325890 577092 325946
rect 577092 325890 577096 325946
rect 577032 325886 577096 325890
rect 577112 325946 577176 325950
rect 577112 325890 577116 325946
rect 577116 325890 577172 325946
rect 577172 325890 577176 325946
rect 577112 325886 577176 325890
rect 577192 325946 577256 325950
rect 577192 325890 577196 325946
rect 577196 325890 577252 325946
rect 577252 325890 577256 325946
rect 577192 325886 577256 325890
rect 577272 325946 577336 325950
rect 577272 325890 577276 325946
rect 577276 325890 577332 325946
rect 577332 325890 577336 325946
rect 577272 325886 577336 325890
rect 577352 325946 577416 325950
rect 577352 325890 577356 325946
rect 577356 325890 577412 325946
rect 577412 325890 577416 325946
rect 577352 325886 577416 325890
rect 577432 325946 577496 325950
rect 577432 325890 577436 325946
rect 577436 325890 577492 325946
rect 577492 325890 577496 325946
rect 577432 325886 577496 325890
rect 577512 325946 577576 325950
rect 577512 325890 577516 325946
rect 577516 325890 577572 325946
rect 577572 325890 577576 325946
rect 577512 325886 577576 325890
rect 577032 325866 577096 325870
rect 577032 325810 577036 325866
rect 577036 325810 577092 325866
rect 577092 325810 577096 325866
rect 577032 325806 577096 325810
rect 577112 325866 577176 325870
rect 577112 325810 577116 325866
rect 577116 325810 577172 325866
rect 577172 325810 577176 325866
rect 577112 325806 577176 325810
rect 577192 325866 577256 325870
rect 577192 325810 577196 325866
rect 577196 325810 577252 325866
rect 577252 325810 577256 325866
rect 577192 325806 577256 325810
rect 577272 325866 577336 325870
rect 577272 325810 577276 325866
rect 577276 325810 577332 325866
rect 577332 325810 577336 325866
rect 577272 325806 577336 325810
rect 577352 325866 577416 325870
rect 577352 325810 577356 325866
rect 577356 325810 577412 325866
rect 577412 325810 577416 325866
rect 577352 325806 577416 325810
rect 577432 325866 577496 325870
rect 577432 325810 577436 325866
rect 577436 325810 577492 325866
rect 577492 325810 577496 325866
rect 577432 325806 577496 325810
rect 577512 325866 577576 325870
rect 577512 325810 577516 325866
rect 577516 325810 577572 325866
rect 577572 325810 577576 325866
rect 577512 325806 577576 325810
rect 577032 325786 577096 325790
rect 577032 325730 577036 325786
rect 577036 325730 577092 325786
rect 577092 325730 577096 325786
rect 577032 325726 577096 325730
rect 577112 325786 577176 325790
rect 577112 325730 577116 325786
rect 577116 325730 577172 325786
rect 577172 325730 577176 325786
rect 577112 325726 577176 325730
rect 577192 325786 577256 325790
rect 577192 325730 577196 325786
rect 577196 325730 577252 325786
rect 577252 325730 577256 325786
rect 577192 325726 577256 325730
rect 577272 325786 577336 325790
rect 577272 325730 577276 325786
rect 577276 325730 577332 325786
rect 577332 325730 577336 325786
rect 577272 325726 577336 325730
rect 577352 325786 577416 325790
rect 577352 325730 577356 325786
rect 577356 325730 577412 325786
rect 577412 325730 577416 325786
rect 577352 325726 577416 325730
rect 577432 325786 577496 325790
rect 577432 325730 577436 325786
rect 577436 325730 577492 325786
rect 577492 325730 577496 325786
rect 577432 325726 577496 325730
rect 577512 325786 577576 325790
rect 577512 325730 577516 325786
rect 577516 325730 577572 325786
rect 577572 325730 577576 325786
rect 577512 325726 577576 325730
rect 577032 325706 577096 325710
rect 577032 325650 577036 325706
rect 577036 325650 577092 325706
rect 577092 325650 577096 325706
rect 577032 325646 577096 325650
rect 577112 325706 577176 325710
rect 577112 325650 577116 325706
rect 577116 325650 577172 325706
rect 577172 325650 577176 325706
rect 577112 325646 577176 325650
rect 577192 325706 577256 325710
rect 577192 325650 577196 325706
rect 577196 325650 577252 325706
rect 577252 325650 577256 325706
rect 577192 325646 577256 325650
rect 577272 325706 577336 325710
rect 577272 325650 577276 325706
rect 577276 325650 577332 325706
rect 577332 325650 577336 325706
rect 577272 325646 577336 325650
rect 577352 325706 577416 325710
rect 577352 325650 577356 325706
rect 577356 325650 577412 325706
rect 577412 325650 577416 325706
rect 577352 325646 577416 325650
rect 577432 325706 577496 325710
rect 577432 325650 577436 325706
rect 577436 325650 577492 325706
rect 577492 325650 577496 325706
rect 577432 325646 577496 325650
rect 577512 325706 577576 325710
rect 577512 325650 577516 325706
rect 577516 325650 577572 325706
rect 577572 325650 577576 325706
rect 577512 325646 577576 325650
rect 578272 325151 578336 325155
rect 578272 325095 578276 325151
rect 578276 325095 578332 325151
rect 578332 325095 578336 325151
rect 578272 325091 578336 325095
rect 578352 325151 578416 325155
rect 578352 325095 578356 325151
rect 578356 325095 578412 325151
rect 578412 325095 578416 325151
rect 578352 325091 578416 325095
rect 578432 325151 578496 325155
rect 578432 325095 578436 325151
rect 578436 325095 578492 325151
rect 578492 325095 578496 325151
rect 578432 325091 578496 325095
rect 578512 325151 578576 325155
rect 578512 325095 578516 325151
rect 578516 325095 578572 325151
rect 578572 325095 578576 325151
rect 578512 325091 578576 325095
rect 578592 325151 578656 325155
rect 578592 325095 578596 325151
rect 578596 325095 578652 325151
rect 578652 325095 578656 325151
rect 578592 325091 578656 325095
rect 578672 325151 578736 325155
rect 578672 325095 578676 325151
rect 578676 325095 578732 325151
rect 578732 325095 578736 325151
rect 578672 325091 578736 325095
rect 578752 325151 578816 325155
rect 578752 325095 578756 325151
rect 578756 325095 578812 325151
rect 578812 325095 578816 325151
rect 578752 325091 578816 325095
rect 578272 325071 578336 325075
rect 578272 325015 578276 325071
rect 578276 325015 578332 325071
rect 578332 325015 578336 325071
rect 578272 325011 578336 325015
rect 578352 325071 578416 325075
rect 578352 325015 578356 325071
rect 578356 325015 578412 325071
rect 578412 325015 578416 325071
rect 578352 325011 578416 325015
rect 578432 325071 578496 325075
rect 578432 325015 578436 325071
rect 578436 325015 578492 325071
rect 578492 325015 578496 325071
rect 578432 325011 578496 325015
rect 578512 325071 578576 325075
rect 578512 325015 578516 325071
rect 578516 325015 578572 325071
rect 578572 325015 578576 325071
rect 578512 325011 578576 325015
rect 578592 325071 578656 325075
rect 578592 325015 578596 325071
rect 578596 325015 578652 325071
rect 578652 325015 578656 325071
rect 578592 325011 578656 325015
rect 578672 325071 578736 325075
rect 578672 325015 578676 325071
rect 578676 325015 578732 325071
rect 578732 325015 578736 325071
rect 578672 325011 578736 325015
rect 578752 325071 578816 325075
rect 578752 325015 578756 325071
rect 578756 325015 578812 325071
rect 578812 325015 578816 325071
rect 578752 325011 578816 325015
rect 578272 324991 578336 324995
rect 578272 324935 578276 324991
rect 578276 324935 578332 324991
rect 578332 324935 578336 324991
rect 578272 324931 578336 324935
rect 578352 324991 578416 324995
rect 578352 324935 578356 324991
rect 578356 324935 578412 324991
rect 578412 324935 578416 324991
rect 578352 324931 578416 324935
rect 578432 324991 578496 324995
rect 578432 324935 578436 324991
rect 578436 324935 578492 324991
rect 578492 324935 578496 324991
rect 578432 324931 578496 324935
rect 578512 324991 578576 324995
rect 578512 324935 578516 324991
rect 578516 324935 578572 324991
rect 578572 324935 578576 324991
rect 578512 324931 578576 324935
rect 578592 324991 578656 324995
rect 578592 324935 578596 324991
rect 578596 324935 578652 324991
rect 578652 324935 578656 324991
rect 578592 324931 578656 324935
rect 578672 324991 578736 324995
rect 578672 324935 578676 324991
rect 578676 324935 578732 324991
rect 578732 324935 578736 324991
rect 578672 324931 578736 324935
rect 578752 324991 578816 324995
rect 578752 324935 578756 324991
rect 578756 324935 578812 324991
rect 578812 324935 578816 324991
rect 578752 324931 578816 324935
rect 578272 324911 578336 324915
rect 578272 324855 578276 324911
rect 578276 324855 578332 324911
rect 578332 324855 578336 324911
rect 578272 324851 578336 324855
rect 578352 324911 578416 324915
rect 578352 324855 578356 324911
rect 578356 324855 578412 324911
rect 578412 324855 578416 324911
rect 578352 324851 578416 324855
rect 578432 324911 578496 324915
rect 578432 324855 578436 324911
rect 578436 324855 578492 324911
rect 578492 324855 578496 324911
rect 578432 324851 578496 324855
rect 578512 324911 578576 324915
rect 578512 324855 578516 324911
rect 578516 324855 578572 324911
rect 578572 324855 578576 324911
rect 578512 324851 578576 324855
rect 578592 324911 578656 324915
rect 578592 324855 578596 324911
rect 578596 324855 578652 324911
rect 578652 324855 578656 324911
rect 578592 324851 578656 324855
rect 578672 324911 578736 324915
rect 578672 324855 578676 324911
rect 578676 324855 578732 324911
rect 578732 324855 578736 324911
rect 578672 324851 578736 324855
rect 578752 324911 578816 324915
rect 578752 324855 578756 324911
rect 578756 324855 578812 324911
rect 578812 324855 578816 324911
rect 578752 324851 578816 324855
rect 470272 322482 470336 322486
rect 470272 322426 470276 322482
rect 470276 322426 470332 322482
rect 470332 322426 470336 322482
rect 470272 322422 470336 322426
rect 470352 322482 470416 322486
rect 470352 322426 470356 322482
rect 470356 322426 470412 322482
rect 470412 322426 470416 322482
rect 470352 322422 470416 322426
rect 470432 322482 470496 322486
rect 470432 322426 470436 322482
rect 470436 322426 470492 322482
rect 470492 322426 470496 322482
rect 470432 322422 470496 322426
rect 470512 322482 470576 322486
rect 470512 322426 470516 322482
rect 470516 322426 470572 322482
rect 470572 322426 470576 322482
rect 470512 322422 470576 322426
rect 470592 322482 470656 322486
rect 470592 322426 470596 322482
rect 470596 322426 470652 322482
rect 470652 322426 470656 322482
rect 470592 322422 470656 322426
rect 470672 322482 470736 322486
rect 470672 322426 470676 322482
rect 470676 322426 470732 322482
rect 470732 322426 470736 322482
rect 470672 322422 470736 322426
rect 470752 322482 470816 322486
rect 470752 322426 470756 322482
rect 470756 322426 470812 322482
rect 470812 322426 470816 322482
rect 470752 322422 470816 322426
rect 470272 322402 470336 322406
rect 470272 322346 470276 322402
rect 470276 322346 470332 322402
rect 470332 322346 470336 322402
rect 470272 322342 470336 322346
rect 470352 322402 470416 322406
rect 470352 322346 470356 322402
rect 470356 322346 470412 322402
rect 470412 322346 470416 322402
rect 470352 322342 470416 322346
rect 470432 322402 470496 322406
rect 470432 322346 470436 322402
rect 470436 322346 470492 322402
rect 470492 322346 470496 322402
rect 470432 322342 470496 322346
rect 470512 322402 470576 322406
rect 470512 322346 470516 322402
rect 470516 322346 470572 322402
rect 470572 322346 470576 322402
rect 470512 322342 470576 322346
rect 470592 322402 470656 322406
rect 470592 322346 470596 322402
rect 470596 322346 470652 322402
rect 470652 322346 470656 322402
rect 470592 322342 470656 322346
rect 470672 322402 470736 322406
rect 470672 322346 470676 322402
rect 470676 322346 470732 322402
rect 470732 322346 470736 322402
rect 470672 322342 470736 322346
rect 470752 322402 470816 322406
rect 470752 322346 470756 322402
rect 470756 322346 470812 322402
rect 470812 322346 470816 322402
rect 470752 322342 470816 322346
rect 470272 322322 470336 322326
rect 470272 322266 470276 322322
rect 470276 322266 470332 322322
rect 470332 322266 470336 322322
rect 470272 322262 470336 322266
rect 470352 322322 470416 322326
rect 470352 322266 470356 322322
rect 470356 322266 470412 322322
rect 470412 322266 470416 322322
rect 470352 322262 470416 322266
rect 470432 322322 470496 322326
rect 470432 322266 470436 322322
rect 470436 322266 470492 322322
rect 470492 322266 470496 322322
rect 470432 322262 470496 322266
rect 470512 322322 470576 322326
rect 470512 322266 470516 322322
rect 470516 322266 470572 322322
rect 470572 322266 470576 322322
rect 470512 322262 470576 322266
rect 470592 322322 470656 322326
rect 470592 322266 470596 322322
rect 470596 322266 470652 322322
rect 470652 322266 470656 322322
rect 470592 322262 470656 322266
rect 470672 322322 470736 322326
rect 470672 322266 470676 322322
rect 470676 322266 470732 322322
rect 470732 322266 470736 322322
rect 470672 322262 470736 322266
rect 470752 322322 470816 322326
rect 470752 322266 470756 322322
rect 470756 322266 470812 322322
rect 470812 322266 470816 322322
rect 470752 322262 470816 322266
rect 470272 322242 470336 322246
rect 470272 322186 470276 322242
rect 470276 322186 470332 322242
rect 470332 322186 470336 322242
rect 470272 322182 470336 322186
rect 470352 322242 470416 322246
rect 470352 322186 470356 322242
rect 470356 322186 470412 322242
rect 470412 322186 470416 322242
rect 470352 322182 470416 322186
rect 470432 322242 470496 322246
rect 470432 322186 470436 322242
rect 470436 322186 470492 322242
rect 470492 322186 470496 322242
rect 470432 322182 470496 322186
rect 470512 322242 470576 322246
rect 470512 322186 470516 322242
rect 470516 322186 470572 322242
rect 470572 322186 470576 322242
rect 470512 322182 470576 322186
rect 470592 322242 470656 322246
rect 470592 322186 470596 322242
rect 470596 322186 470652 322242
rect 470652 322186 470656 322242
rect 470592 322182 470656 322186
rect 470672 322242 470736 322246
rect 470672 322186 470676 322242
rect 470676 322186 470732 322242
rect 470732 322186 470736 322242
rect 470672 322182 470736 322186
rect 470752 322242 470816 322246
rect 470752 322186 470756 322242
rect 470756 322186 470812 322242
rect 470812 322186 470816 322242
rect 470752 322182 470816 322186
rect 483612 322086 483676 322150
rect 483612 321542 483676 321606
rect 469032 321395 469096 321399
rect 469032 321339 469036 321395
rect 469036 321339 469092 321395
rect 469092 321339 469096 321395
rect 469032 321335 469096 321339
rect 469112 321395 469176 321399
rect 469112 321339 469116 321395
rect 469116 321339 469172 321395
rect 469172 321339 469176 321395
rect 469112 321335 469176 321339
rect 469192 321395 469256 321399
rect 469192 321339 469196 321395
rect 469196 321339 469252 321395
rect 469252 321339 469256 321395
rect 469192 321335 469256 321339
rect 469272 321395 469336 321399
rect 469272 321339 469276 321395
rect 469276 321339 469332 321395
rect 469332 321339 469336 321395
rect 469272 321335 469336 321339
rect 469352 321395 469416 321399
rect 469352 321339 469356 321395
rect 469356 321339 469412 321395
rect 469412 321339 469416 321395
rect 469352 321335 469416 321339
rect 469432 321395 469496 321399
rect 469432 321339 469436 321395
rect 469436 321339 469492 321395
rect 469492 321339 469496 321395
rect 469432 321335 469496 321339
rect 469512 321395 469576 321399
rect 469512 321339 469516 321395
rect 469516 321339 469572 321395
rect 469572 321339 469576 321395
rect 469512 321335 469576 321339
rect 469032 321315 469096 321319
rect 469032 321259 469036 321315
rect 469036 321259 469092 321315
rect 469092 321259 469096 321315
rect 469032 321255 469096 321259
rect 469112 321315 469176 321319
rect 469112 321259 469116 321315
rect 469116 321259 469172 321315
rect 469172 321259 469176 321315
rect 469112 321255 469176 321259
rect 469192 321315 469256 321319
rect 469192 321259 469196 321315
rect 469196 321259 469252 321315
rect 469252 321259 469256 321315
rect 469192 321255 469256 321259
rect 469272 321315 469336 321319
rect 469272 321259 469276 321315
rect 469276 321259 469332 321315
rect 469332 321259 469336 321315
rect 469272 321255 469336 321259
rect 469352 321315 469416 321319
rect 469352 321259 469356 321315
rect 469356 321259 469412 321315
rect 469412 321259 469416 321315
rect 469352 321255 469416 321259
rect 469432 321315 469496 321319
rect 469432 321259 469436 321315
rect 469436 321259 469492 321315
rect 469492 321259 469496 321315
rect 469432 321255 469496 321259
rect 469512 321315 469576 321319
rect 469512 321259 469516 321315
rect 469516 321259 469572 321315
rect 469572 321259 469576 321315
rect 469512 321255 469576 321259
rect 473676 321270 473740 321334
rect 469032 321235 469096 321239
rect 469032 321179 469036 321235
rect 469036 321179 469092 321235
rect 469092 321179 469096 321235
rect 469032 321175 469096 321179
rect 469112 321235 469176 321239
rect 469112 321179 469116 321235
rect 469116 321179 469172 321235
rect 469172 321179 469176 321235
rect 469112 321175 469176 321179
rect 469192 321235 469256 321239
rect 469192 321179 469196 321235
rect 469196 321179 469252 321235
rect 469252 321179 469256 321235
rect 469192 321175 469256 321179
rect 469272 321235 469336 321239
rect 469272 321179 469276 321235
rect 469276 321179 469332 321235
rect 469332 321179 469336 321235
rect 469272 321175 469336 321179
rect 469352 321235 469416 321239
rect 469352 321179 469356 321235
rect 469356 321179 469412 321235
rect 469412 321179 469416 321235
rect 469352 321175 469416 321179
rect 469432 321235 469496 321239
rect 469432 321179 469436 321235
rect 469436 321179 469492 321235
rect 469492 321179 469496 321235
rect 469432 321175 469496 321179
rect 469512 321235 469576 321239
rect 469512 321179 469516 321235
rect 469516 321179 469572 321235
rect 469572 321179 469576 321235
rect 469512 321175 469576 321179
rect 469032 321155 469096 321159
rect 469032 321099 469036 321155
rect 469036 321099 469092 321155
rect 469092 321099 469096 321155
rect 469032 321095 469096 321099
rect 469112 321155 469176 321159
rect 469112 321099 469116 321155
rect 469116 321099 469172 321155
rect 469172 321099 469176 321155
rect 469112 321095 469176 321099
rect 469192 321155 469256 321159
rect 469192 321099 469196 321155
rect 469196 321099 469252 321155
rect 469252 321099 469256 321155
rect 469192 321095 469256 321099
rect 469272 321155 469336 321159
rect 469272 321099 469276 321155
rect 469276 321099 469332 321155
rect 469332 321099 469336 321155
rect 469272 321095 469336 321099
rect 469352 321155 469416 321159
rect 469352 321099 469356 321155
rect 469356 321099 469412 321155
rect 469412 321099 469416 321155
rect 469352 321095 469416 321099
rect 469432 321155 469496 321159
rect 469432 321099 469436 321155
rect 469436 321099 469492 321155
rect 469492 321099 469496 321155
rect 469432 321095 469496 321099
rect 469512 321155 469576 321159
rect 469512 321099 469516 321155
rect 469516 321099 469572 321155
rect 469572 321099 469576 321155
rect 469512 321095 469576 321099
rect 481036 320998 481100 321062
rect 488028 320998 488092 321062
rect 478644 320862 478708 320926
rect 470272 320310 470336 320314
rect 470272 320254 470276 320310
rect 470276 320254 470332 320310
rect 470332 320254 470336 320310
rect 470272 320250 470336 320254
rect 470352 320310 470416 320314
rect 470352 320254 470356 320310
rect 470356 320254 470412 320310
rect 470412 320254 470416 320310
rect 470352 320250 470416 320254
rect 470432 320310 470496 320314
rect 470432 320254 470436 320310
rect 470436 320254 470492 320310
rect 470492 320254 470496 320310
rect 470432 320250 470496 320254
rect 470512 320310 470576 320314
rect 470512 320254 470516 320310
rect 470516 320254 470572 320310
rect 470572 320254 470576 320310
rect 470512 320250 470576 320254
rect 470592 320310 470656 320314
rect 470592 320254 470596 320310
rect 470596 320254 470652 320310
rect 470652 320254 470656 320310
rect 470592 320250 470656 320254
rect 470672 320310 470736 320314
rect 470672 320254 470676 320310
rect 470676 320254 470732 320310
rect 470732 320254 470736 320310
rect 470672 320250 470736 320254
rect 470752 320310 470816 320314
rect 470752 320254 470756 320310
rect 470756 320254 470812 320310
rect 470812 320254 470816 320310
rect 470752 320250 470816 320254
rect 470272 320230 470336 320234
rect 470272 320174 470276 320230
rect 470276 320174 470332 320230
rect 470332 320174 470336 320230
rect 470272 320170 470336 320174
rect 470352 320230 470416 320234
rect 470352 320174 470356 320230
rect 470356 320174 470412 320230
rect 470412 320174 470416 320230
rect 470352 320170 470416 320174
rect 470432 320230 470496 320234
rect 470432 320174 470436 320230
rect 470436 320174 470492 320230
rect 470492 320174 470496 320230
rect 470432 320170 470496 320174
rect 470512 320230 470576 320234
rect 470512 320174 470516 320230
rect 470516 320174 470572 320230
rect 470572 320174 470576 320230
rect 470512 320170 470576 320174
rect 470592 320230 470656 320234
rect 470592 320174 470596 320230
rect 470596 320174 470652 320230
rect 470652 320174 470656 320230
rect 470592 320170 470656 320174
rect 470672 320230 470736 320234
rect 470672 320174 470676 320230
rect 470676 320174 470732 320230
rect 470732 320174 470736 320230
rect 470672 320170 470736 320174
rect 470752 320230 470816 320234
rect 470752 320174 470756 320230
rect 470756 320174 470812 320230
rect 470812 320174 470816 320230
rect 470752 320170 470816 320174
rect 470272 320150 470336 320154
rect 470272 320094 470276 320150
rect 470276 320094 470332 320150
rect 470332 320094 470336 320150
rect 470272 320090 470336 320094
rect 470352 320150 470416 320154
rect 470352 320094 470356 320150
rect 470356 320094 470412 320150
rect 470412 320094 470416 320150
rect 470352 320090 470416 320094
rect 470432 320150 470496 320154
rect 470432 320094 470436 320150
rect 470436 320094 470492 320150
rect 470492 320094 470496 320150
rect 470432 320090 470496 320094
rect 470512 320150 470576 320154
rect 470512 320094 470516 320150
rect 470516 320094 470572 320150
rect 470572 320094 470576 320150
rect 470512 320090 470576 320094
rect 470592 320150 470656 320154
rect 470592 320094 470596 320150
rect 470596 320094 470652 320150
rect 470652 320094 470656 320150
rect 470592 320090 470656 320094
rect 470672 320150 470736 320154
rect 470672 320094 470676 320150
rect 470676 320094 470732 320150
rect 470732 320094 470736 320150
rect 470672 320090 470736 320094
rect 470752 320150 470816 320154
rect 470752 320094 470756 320150
rect 470756 320094 470812 320150
rect 470812 320094 470816 320150
rect 470752 320090 470816 320094
rect 470272 320070 470336 320074
rect 470272 320014 470276 320070
rect 470276 320014 470332 320070
rect 470332 320014 470336 320070
rect 470272 320010 470336 320014
rect 470352 320070 470416 320074
rect 470352 320014 470356 320070
rect 470356 320014 470412 320070
rect 470412 320014 470416 320070
rect 470352 320010 470416 320014
rect 470432 320070 470496 320074
rect 470432 320014 470436 320070
rect 470436 320014 470492 320070
rect 470492 320014 470496 320070
rect 470432 320010 470496 320014
rect 470512 320070 470576 320074
rect 470512 320014 470516 320070
rect 470516 320014 470572 320070
rect 470572 320014 470576 320070
rect 470512 320010 470576 320014
rect 470592 320070 470656 320074
rect 470592 320014 470596 320070
rect 470596 320014 470652 320070
rect 470652 320014 470656 320070
rect 470592 320010 470656 320014
rect 470672 320070 470736 320074
rect 470672 320014 470676 320070
rect 470676 320014 470732 320070
rect 470732 320014 470736 320070
rect 470672 320010 470736 320014
rect 470752 320070 470816 320074
rect 470752 320014 470756 320070
rect 470756 320014 470812 320070
rect 470812 320014 470816 320070
rect 470752 320010 470816 320014
rect 470272 307082 470336 307086
rect 470272 307026 470276 307082
rect 470276 307026 470332 307082
rect 470332 307026 470336 307082
rect 470272 307022 470336 307026
rect 470352 307082 470416 307086
rect 470352 307026 470356 307082
rect 470356 307026 470412 307082
rect 470412 307026 470416 307082
rect 470352 307022 470416 307026
rect 470432 307082 470496 307086
rect 470432 307026 470436 307082
rect 470436 307026 470492 307082
rect 470492 307026 470496 307082
rect 470432 307022 470496 307026
rect 470512 307082 470576 307086
rect 470512 307026 470516 307082
rect 470516 307026 470572 307082
rect 470572 307026 470576 307082
rect 470512 307022 470576 307026
rect 470592 307082 470656 307086
rect 470592 307026 470596 307082
rect 470596 307026 470652 307082
rect 470652 307026 470656 307082
rect 470592 307022 470656 307026
rect 470672 307082 470736 307086
rect 470672 307026 470676 307082
rect 470676 307026 470732 307082
rect 470732 307026 470736 307082
rect 470672 307022 470736 307026
rect 470752 307082 470816 307086
rect 470752 307026 470756 307082
rect 470756 307026 470812 307082
rect 470812 307026 470816 307082
rect 470752 307022 470816 307026
rect 470272 307002 470336 307006
rect 470272 306946 470276 307002
rect 470276 306946 470332 307002
rect 470332 306946 470336 307002
rect 470272 306942 470336 306946
rect 470352 307002 470416 307006
rect 470352 306946 470356 307002
rect 470356 306946 470412 307002
rect 470412 306946 470416 307002
rect 470352 306942 470416 306946
rect 470432 307002 470496 307006
rect 470432 306946 470436 307002
rect 470436 306946 470492 307002
rect 470492 306946 470496 307002
rect 470432 306942 470496 306946
rect 470512 307002 470576 307006
rect 470512 306946 470516 307002
rect 470516 306946 470572 307002
rect 470572 306946 470576 307002
rect 470512 306942 470576 306946
rect 470592 307002 470656 307006
rect 470592 306946 470596 307002
rect 470596 306946 470652 307002
rect 470652 306946 470656 307002
rect 470592 306942 470656 306946
rect 470672 307002 470736 307006
rect 470672 306946 470676 307002
rect 470676 306946 470732 307002
rect 470732 306946 470736 307002
rect 470672 306942 470736 306946
rect 470752 307002 470816 307006
rect 470752 306946 470756 307002
rect 470756 306946 470812 307002
rect 470812 306946 470816 307002
rect 470752 306942 470816 306946
rect 470272 306922 470336 306926
rect 470272 306866 470276 306922
rect 470276 306866 470332 306922
rect 470332 306866 470336 306922
rect 470272 306862 470336 306866
rect 470352 306922 470416 306926
rect 470352 306866 470356 306922
rect 470356 306866 470412 306922
rect 470412 306866 470416 306922
rect 470352 306862 470416 306866
rect 470432 306922 470496 306926
rect 470432 306866 470436 306922
rect 470436 306866 470492 306922
rect 470492 306866 470496 306922
rect 470432 306862 470496 306866
rect 470512 306922 470576 306926
rect 470512 306866 470516 306922
rect 470516 306866 470572 306922
rect 470572 306866 470576 306922
rect 470512 306862 470576 306866
rect 470592 306922 470656 306926
rect 470592 306866 470596 306922
rect 470596 306866 470652 306922
rect 470652 306866 470656 306922
rect 470592 306862 470656 306866
rect 470672 306922 470736 306926
rect 470672 306866 470676 306922
rect 470676 306866 470732 306922
rect 470732 306866 470736 306922
rect 470672 306862 470736 306866
rect 470752 306922 470816 306926
rect 470752 306866 470756 306922
rect 470756 306866 470812 306922
rect 470812 306866 470816 306922
rect 470752 306862 470816 306866
rect 470272 306842 470336 306846
rect 470272 306786 470276 306842
rect 470276 306786 470332 306842
rect 470332 306786 470336 306842
rect 470272 306782 470336 306786
rect 470352 306842 470416 306846
rect 470352 306786 470356 306842
rect 470356 306786 470412 306842
rect 470412 306786 470416 306842
rect 470352 306782 470416 306786
rect 470432 306842 470496 306846
rect 470432 306786 470436 306842
rect 470436 306786 470492 306842
rect 470492 306786 470496 306842
rect 470432 306782 470496 306786
rect 470512 306842 470576 306846
rect 470512 306786 470516 306842
rect 470516 306786 470572 306842
rect 470572 306786 470576 306842
rect 470512 306782 470576 306786
rect 470592 306842 470656 306846
rect 470592 306786 470596 306842
rect 470596 306786 470652 306842
rect 470652 306786 470656 306842
rect 470592 306782 470656 306786
rect 470672 306842 470736 306846
rect 470672 306786 470676 306842
rect 470676 306786 470732 306842
rect 470732 306786 470736 306842
rect 470672 306782 470736 306786
rect 470752 306842 470816 306846
rect 470752 306786 470756 306842
rect 470756 306786 470812 306842
rect 470812 306786 470816 306842
rect 470752 306782 470816 306786
rect 480852 306506 480916 306510
rect 480852 306450 480902 306506
rect 480902 306450 480916 306506
rect 480852 306446 480916 306450
rect 487660 306310 487724 306374
rect 469032 305997 469096 306001
rect 469032 305941 469036 305997
rect 469036 305941 469092 305997
rect 469092 305941 469096 305997
rect 469032 305937 469096 305941
rect 469112 305997 469176 306001
rect 469112 305941 469116 305997
rect 469116 305941 469172 305997
rect 469172 305941 469176 305997
rect 469112 305937 469176 305941
rect 469192 305997 469256 306001
rect 469192 305941 469196 305997
rect 469196 305941 469252 305997
rect 469252 305941 469256 305997
rect 469192 305937 469256 305941
rect 469272 305997 469336 306001
rect 469272 305941 469276 305997
rect 469276 305941 469332 305997
rect 469332 305941 469336 305997
rect 469272 305937 469336 305941
rect 469352 305997 469416 306001
rect 469352 305941 469356 305997
rect 469356 305941 469412 305997
rect 469412 305941 469416 305997
rect 469352 305937 469416 305941
rect 469432 305997 469496 306001
rect 469432 305941 469436 305997
rect 469436 305941 469492 305997
rect 469492 305941 469496 305997
rect 469432 305937 469496 305941
rect 469512 305997 469576 306001
rect 469512 305941 469516 305997
rect 469516 305941 469572 305997
rect 469572 305941 469576 305997
rect 469512 305937 469576 305941
rect 469032 305917 469096 305921
rect 469032 305861 469036 305917
rect 469036 305861 469092 305917
rect 469092 305861 469096 305917
rect 469032 305857 469096 305861
rect 469112 305917 469176 305921
rect 469112 305861 469116 305917
rect 469116 305861 469172 305917
rect 469172 305861 469176 305917
rect 469112 305857 469176 305861
rect 469192 305917 469256 305921
rect 469192 305861 469196 305917
rect 469196 305861 469252 305917
rect 469252 305861 469256 305917
rect 469192 305857 469256 305861
rect 469272 305917 469336 305921
rect 469272 305861 469276 305917
rect 469276 305861 469332 305917
rect 469332 305861 469336 305917
rect 469272 305857 469336 305861
rect 469352 305917 469416 305921
rect 469352 305861 469356 305917
rect 469356 305861 469412 305917
rect 469412 305861 469416 305917
rect 469352 305857 469416 305861
rect 469432 305917 469496 305921
rect 469432 305861 469436 305917
rect 469436 305861 469492 305917
rect 469492 305861 469496 305917
rect 469432 305857 469496 305861
rect 469512 305917 469576 305921
rect 469512 305861 469516 305917
rect 469516 305861 469572 305917
rect 469572 305861 469576 305917
rect 469512 305857 469576 305861
rect 473676 305962 473740 305966
rect 473676 305906 473726 305962
rect 473726 305906 473740 305962
rect 473676 305902 473740 305906
rect 469032 305837 469096 305841
rect 469032 305781 469036 305837
rect 469036 305781 469092 305837
rect 469092 305781 469096 305837
rect 469032 305777 469096 305781
rect 469112 305837 469176 305841
rect 469112 305781 469116 305837
rect 469116 305781 469172 305837
rect 469172 305781 469176 305837
rect 469112 305777 469176 305781
rect 469192 305837 469256 305841
rect 469192 305781 469196 305837
rect 469196 305781 469252 305837
rect 469252 305781 469256 305837
rect 469192 305777 469256 305781
rect 469272 305837 469336 305841
rect 469272 305781 469276 305837
rect 469276 305781 469332 305837
rect 469332 305781 469336 305837
rect 469272 305777 469336 305781
rect 469352 305837 469416 305841
rect 469352 305781 469356 305837
rect 469356 305781 469412 305837
rect 469412 305781 469416 305837
rect 469352 305777 469416 305781
rect 469432 305837 469496 305841
rect 469432 305781 469436 305837
rect 469436 305781 469492 305837
rect 469492 305781 469496 305837
rect 469432 305777 469496 305781
rect 469512 305837 469576 305841
rect 469512 305781 469516 305837
rect 469516 305781 469572 305837
rect 469572 305781 469576 305837
rect 469512 305777 469576 305781
rect 469032 305757 469096 305761
rect 469032 305701 469036 305757
rect 469036 305701 469092 305757
rect 469092 305701 469096 305757
rect 469032 305697 469096 305701
rect 469112 305757 469176 305761
rect 469112 305701 469116 305757
rect 469116 305701 469172 305757
rect 469172 305701 469176 305757
rect 469112 305697 469176 305701
rect 469192 305757 469256 305761
rect 469192 305701 469196 305757
rect 469196 305701 469252 305757
rect 469252 305701 469256 305757
rect 469192 305697 469256 305701
rect 469272 305757 469336 305761
rect 469272 305701 469276 305757
rect 469276 305701 469332 305757
rect 469332 305701 469336 305757
rect 469272 305697 469336 305701
rect 469352 305757 469416 305761
rect 469352 305701 469356 305757
rect 469356 305701 469412 305757
rect 469412 305701 469416 305757
rect 469352 305697 469416 305701
rect 469432 305757 469496 305761
rect 469432 305701 469436 305757
rect 469436 305701 469492 305757
rect 469492 305701 469496 305757
rect 469432 305697 469496 305701
rect 469512 305757 469576 305761
rect 469512 305701 469516 305757
rect 469516 305701 469572 305757
rect 469572 305701 469576 305757
rect 469512 305697 469576 305701
rect 478828 305630 478892 305694
rect 484164 305554 484228 305558
rect 484164 305498 484178 305554
rect 484178 305498 484228 305554
rect 484164 305494 484228 305498
rect 470272 304910 470336 304914
rect 470272 304854 470276 304910
rect 470276 304854 470332 304910
rect 470332 304854 470336 304910
rect 470272 304850 470336 304854
rect 470352 304910 470416 304914
rect 470352 304854 470356 304910
rect 470356 304854 470412 304910
rect 470412 304854 470416 304910
rect 470352 304850 470416 304854
rect 470432 304910 470496 304914
rect 470432 304854 470436 304910
rect 470436 304854 470492 304910
rect 470492 304854 470496 304910
rect 470432 304850 470496 304854
rect 470512 304910 470576 304914
rect 470512 304854 470516 304910
rect 470516 304854 470572 304910
rect 470572 304854 470576 304910
rect 470512 304850 470576 304854
rect 470592 304910 470656 304914
rect 470592 304854 470596 304910
rect 470596 304854 470652 304910
rect 470652 304854 470656 304910
rect 470592 304850 470656 304854
rect 470672 304910 470736 304914
rect 470672 304854 470676 304910
rect 470676 304854 470732 304910
rect 470732 304854 470736 304910
rect 470672 304850 470736 304854
rect 470752 304910 470816 304914
rect 470752 304854 470756 304910
rect 470756 304854 470812 304910
rect 470812 304854 470816 304910
rect 470752 304850 470816 304854
rect 470272 304830 470336 304834
rect 470272 304774 470276 304830
rect 470276 304774 470332 304830
rect 470332 304774 470336 304830
rect 470272 304770 470336 304774
rect 470352 304830 470416 304834
rect 470352 304774 470356 304830
rect 470356 304774 470412 304830
rect 470412 304774 470416 304830
rect 470352 304770 470416 304774
rect 470432 304830 470496 304834
rect 470432 304774 470436 304830
rect 470436 304774 470492 304830
rect 470492 304774 470496 304830
rect 470432 304770 470496 304774
rect 470512 304830 470576 304834
rect 470512 304774 470516 304830
rect 470516 304774 470572 304830
rect 470572 304774 470576 304830
rect 470512 304770 470576 304774
rect 470592 304830 470656 304834
rect 470592 304774 470596 304830
rect 470596 304774 470652 304830
rect 470652 304774 470656 304830
rect 470592 304770 470656 304774
rect 470672 304830 470736 304834
rect 470672 304774 470676 304830
rect 470676 304774 470732 304830
rect 470732 304774 470736 304830
rect 470672 304770 470736 304774
rect 470752 304830 470816 304834
rect 470752 304774 470756 304830
rect 470756 304774 470812 304830
rect 470812 304774 470816 304830
rect 470752 304770 470816 304774
rect 470272 304750 470336 304754
rect 470272 304694 470276 304750
rect 470276 304694 470332 304750
rect 470332 304694 470336 304750
rect 470272 304690 470336 304694
rect 470352 304750 470416 304754
rect 470352 304694 470356 304750
rect 470356 304694 470412 304750
rect 470412 304694 470416 304750
rect 470352 304690 470416 304694
rect 470432 304750 470496 304754
rect 470432 304694 470436 304750
rect 470436 304694 470492 304750
rect 470492 304694 470496 304750
rect 470432 304690 470496 304694
rect 470512 304750 470576 304754
rect 470512 304694 470516 304750
rect 470516 304694 470572 304750
rect 470572 304694 470576 304750
rect 470512 304690 470576 304694
rect 470592 304750 470656 304754
rect 470592 304694 470596 304750
rect 470596 304694 470652 304750
rect 470652 304694 470656 304750
rect 470592 304690 470656 304694
rect 470672 304750 470736 304754
rect 470672 304694 470676 304750
rect 470676 304694 470732 304750
rect 470732 304694 470736 304750
rect 470672 304690 470736 304694
rect 470752 304750 470816 304754
rect 470752 304694 470756 304750
rect 470756 304694 470812 304750
rect 470812 304694 470816 304750
rect 470752 304690 470816 304694
rect 470272 304670 470336 304674
rect 470272 304614 470276 304670
rect 470276 304614 470332 304670
rect 470332 304614 470336 304670
rect 470272 304610 470336 304614
rect 470352 304670 470416 304674
rect 470352 304614 470356 304670
rect 470356 304614 470412 304670
rect 470412 304614 470416 304670
rect 470352 304610 470416 304614
rect 470432 304670 470496 304674
rect 470432 304614 470436 304670
rect 470436 304614 470492 304670
rect 470492 304614 470496 304670
rect 470432 304610 470496 304614
rect 470512 304670 470576 304674
rect 470512 304614 470516 304670
rect 470516 304614 470572 304670
rect 470572 304614 470576 304670
rect 470512 304610 470576 304614
rect 470592 304670 470656 304674
rect 470592 304614 470596 304670
rect 470596 304614 470652 304670
rect 470652 304614 470656 304670
rect 470592 304610 470656 304614
rect 470672 304670 470736 304674
rect 470672 304614 470676 304670
rect 470676 304614 470732 304670
rect 470732 304614 470736 304670
rect 470672 304610 470736 304614
rect 470752 304670 470816 304674
rect 470752 304614 470756 304670
rect 470756 304614 470812 304670
rect 470812 304614 470816 304670
rect 470752 304610 470816 304614
rect 541572 303726 541636 303790
rect 544332 303726 544396 303790
rect 480852 302230 480916 302294
rect 473676 289718 473740 289782
rect 476068 289718 476132 289782
rect 482140 288358 482204 288422
rect 470272 287483 470336 287487
rect 470272 287427 470276 287483
rect 470276 287427 470332 287483
rect 470332 287427 470336 287483
rect 470272 287423 470336 287427
rect 470352 287483 470416 287487
rect 470352 287427 470356 287483
rect 470356 287427 470412 287483
rect 470412 287427 470416 287483
rect 470352 287423 470416 287427
rect 470432 287483 470496 287487
rect 470432 287427 470436 287483
rect 470436 287427 470492 287483
rect 470492 287427 470496 287483
rect 470432 287423 470496 287427
rect 470512 287483 470576 287487
rect 470512 287427 470516 287483
rect 470516 287427 470572 287483
rect 470572 287427 470576 287483
rect 470512 287423 470576 287427
rect 470592 287483 470656 287487
rect 470592 287427 470596 287483
rect 470596 287427 470652 287483
rect 470652 287427 470656 287483
rect 470592 287423 470656 287427
rect 470672 287483 470736 287487
rect 470672 287427 470676 287483
rect 470676 287427 470732 287483
rect 470732 287427 470736 287483
rect 470672 287423 470736 287427
rect 470752 287483 470816 287487
rect 470752 287427 470756 287483
rect 470756 287427 470812 287483
rect 470812 287427 470816 287483
rect 470752 287423 470816 287427
rect 470272 287403 470336 287407
rect 470272 287347 470276 287403
rect 470276 287347 470332 287403
rect 470332 287347 470336 287403
rect 470272 287343 470336 287347
rect 470352 287403 470416 287407
rect 470352 287347 470356 287403
rect 470356 287347 470412 287403
rect 470412 287347 470416 287403
rect 470352 287343 470416 287347
rect 470432 287403 470496 287407
rect 470432 287347 470436 287403
rect 470436 287347 470492 287403
rect 470492 287347 470496 287403
rect 470432 287343 470496 287347
rect 470512 287403 470576 287407
rect 470512 287347 470516 287403
rect 470516 287347 470572 287403
rect 470572 287347 470576 287403
rect 470512 287343 470576 287347
rect 470592 287403 470656 287407
rect 470592 287347 470596 287403
rect 470596 287347 470652 287403
rect 470652 287347 470656 287403
rect 470592 287343 470656 287347
rect 470672 287403 470736 287407
rect 470672 287347 470676 287403
rect 470676 287347 470732 287403
rect 470732 287347 470736 287403
rect 470672 287343 470736 287347
rect 470752 287403 470816 287407
rect 470752 287347 470756 287403
rect 470756 287347 470812 287403
rect 470812 287347 470816 287403
rect 470752 287343 470816 287347
rect 470272 287323 470336 287327
rect 470272 287267 470276 287323
rect 470276 287267 470332 287323
rect 470332 287267 470336 287323
rect 470272 287263 470336 287267
rect 470352 287323 470416 287327
rect 470352 287267 470356 287323
rect 470356 287267 470412 287323
rect 470412 287267 470416 287323
rect 470352 287263 470416 287267
rect 470432 287323 470496 287327
rect 470432 287267 470436 287323
rect 470436 287267 470492 287323
rect 470492 287267 470496 287323
rect 470432 287263 470496 287267
rect 470512 287323 470576 287327
rect 470512 287267 470516 287323
rect 470516 287267 470572 287323
rect 470572 287267 470576 287323
rect 470512 287263 470576 287267
rect 470592 287323 470656 287327
rect 470592 287267 470596 287323
rect 470596 287267 470652 287323
rect 470652 287267 470656 287323
rect 470592 287263 470656 287267
rect 470672 287323 470736 287327
rect 470672 287267 470676 287323
rect 470676 287267 470732 287323
rect 470732 287267 470736 287323
rect 470672 287263 470736 287267
rect 470752 287323 470816 287327
rect 470752 287267 470756 287323
rect 470756 287267 470812 287323
rect 470812 287267 470816 287323
rect 470752 287263 470816 287267
rect 470272 287243 470336 287247
rect 470272 287187 470276 287243
rect 470276 287187 470332 287243
rect 470332 287187 470336 287243
rect 470272 287183 470336 287187
rect 470352 287243 470416 287247
rect 470352 287187 470356 287243
rect 470356 287187 470412 287243
rect 470412 287187 470416 287243
rect 470352 287183 470416 287187
rect 470432 287243 470496 287247
rect 470432 287187 470436 287243
rect 470436 287187 470492 287243
rect 470492 287187 470496 287243
rect 470432 287183 470496 287187
rect 470512 287243 470576 287247
rect 470512 287187 470516 287243
rect 470516 287187 470572 287243
rect 470572 287187 470576 287243
rect 470512 287183 470576 287187
rect 470592 287243 470656 287247
rect 470592 287187 470596 287243
rect 470596 287187 470652 287243
rect 470652 287187 470656 287243
rect 470592 287183 470656 287187
rect 470672 287243 470736 287247
rect 470672 287187 470676 287243
rect 470676 287187 470732 287243
rect 470732 287187 470736 287243
rect 470672 287183 470736 287187
rect 470752 287243 470816 287247
rect 470752 287187 470756 287243
rect 470756 287187 470812 287243
rect 470812 287187 470816 287243
rect 470752 287183 470816 287187
rect 478828 286862 478892 286926
rect 488396 286726 488460 286790
rect 476068 286590 476132 286654
rect 484164 286590 484228 286654
rect 469032 286398 469096 286402
rect 469032 286342 469036 286398
rect 469036 286342 469092 286398
rect 469092 286342 469096 286398
rect 469032 286338 469096 286342
rect 469112 286398 469176 286402
rect 469112 286342 469116 286398
rect 469116 286342 469172 286398
rect 469172 286342 469176 286398
rect 469112 286338 469176 286342
rect 469192 286398 469256 286402
rect 469192 286342 469196 286398
rect 469196 286342 469252 286398
rect 469252 286342 469256 286398
rect 469192 286338 469256 286342
rect 469272 286398 469336 286402
rect 469272 286342 469276 286398
rect 469276 286342 469332 286398
rect 469332 286342 469336 286398
rect 469272 286338 469336 286342
rect 469352 286398 469416 286402
rect 469352 286342 469356 286398
rect 469356 286342 469412 286398
rect 469412 286342 469416 286398
rect 469352 286338 469416 286342
rect 469432 286398 469496 286402
rect 469432 286342 469436 286398
rect 469436 286342 469492 286398
rect 469492 286342 469496 286398
rect 469432 286338 469496 286342
rect 469512 286398 469576 286402
rect 469512 286342 469516 286398
rect 469516 286342 469572 286398
rect 469572 286342 469576 286398
rect 469512 286338 469576 286342
rect 469032 286318 469096 286322
rect 469032 286262 469036 286318
rect 469036 286262 469092 286318
rect 469092 286262 469096 286318
rect 469032 286258 469096 286262
rect 469112 286318 469176 286322
rect 469112 286262 469116 286318
rect 469116 286262 469172 286318
rect 469172 286262 469176 286318
rect 469112 286258 469176 286262
rect 469192 286318 469256 286322
rect 469192 286262 469196 286318
rect 469196 286262 469252 286318
rect 469252 286262 469256 286318
rect 469192 286258 469256 286262
rect 469272 286318 469336 286322
rect 469272 286262 469276 286318
rect 469276 286262 469332 286318
rect 469332 286262 469336 286318
rect 469272 286258 469336 286262
rect 469352 286318 469416 286322
rect 469352 286262 469356 286318
rect 469356 286262 469412 286318
rect 469412 286262 469416 286318
rect 469352 286258 469416 286262
rect 469432 286318 469496 286322
rect 469432 286262 469436 286318
rect 469436 286262 469492 286318
rect 469492 286262 469496 286318
rect 469432 286258 469496 286262
rect 469512 286318 469576 286322
rect 469512 286262 469516 286318
rect 469516 286262 469572 286318
rect 469572 286262 469576 286318
rect 469512 286258 469576 286262
rect 469032 286238 469096 286242
rect 469032 286182 469036 286238
rect 469036 286182 469092 286238
rect 469092 286182 469096 286238
rect 469032 286178 469096 286182
rect 469112 286238 469176 286242
rect 469112 286182 469116 286238
rect 469116 286182 469172 286238
rect 469172 286182 469176 286238
rect 469112 286178 469176 286182
rect 469192 286238 469256 286242
rect 469192 286182 469196 286238
rect 469196 286182 469252 286238
rect 469252 286182 469256 286238
rect 469192 286178 469256 286182
rect 469272 286238 469336 286242
rect 469272 286182 469276 286238
rect 469276 286182 469332 286238
rect 469332 286182 469336 286238
rect 469272 286178 469336 286182
rect 469352 286238 469416 286242
rect 469352 286182 469356 286238
rect 469356 286182 469412 286238
rect 469412 286182 469416 286238
rect 469352 286178 469416 286182
rect 469432 286238 469496 286242
rect 469432 286182 469436 286238
rect 469436 286182 469492 286238
rect 469492 286182 469496 286238
rect 469432 286178 469496 286182
rect 469512 286238 469576 286242
rect 469512 286182 469516 286238
rect 469516 286182 469572 286238
rect 469572 286182 469576 286238
rect 469512 286178 469576 286182
rect 469032 286158 469096 286162
rect 469032 286102 469036 286158
rect 469036 286102 469092 286158
rect 469092 286102 469096 286158
rect 469032 286098 469096 286102
rect 469112 286158 469176 286162
rect 469112 286102 469116 286158
rect 469116 286102 469172 286158
rect 469172 286102 469176 286158
rect 469112 286098 469176 286102
rect 469192 286158 469256 286162
rect 469192 286102 469196 286158
rect 469196 286102 469252 286158
rect 469252 286102 469256 286158
rect 469192 286098 469256 286102
rect 469272 286158 469336 286162
rect 469272 286102 469276 286158
rect 469276 286102 469332 286158
rect 469332 286102 469336 286158
rect 469272 286098 469336 286102
rect 469352 286158 469416 286162
rect 469352 286102 469356 286158
rect 469356 286102 469412 286158
rect 469412 286102 469416 286158
rect 469352 286098 469416 286102
rect 469432 286158 469496 286162
rect 469432 286102 469436 286158
rect 469436 286102 469492 286158
rect 469492 286102 469496 286158
rect 469432 286098 469496 286102
rect 469512 286158 469576 286162
rect 469512 286102 469516 286158
rect 469516 286102 469572 286158
rect 469572 286102 469576 286158
rect 469512 286098 469576 286102
rect 482140 285698 482204 285702
rect 482140 285642 482190 285698
rect 482190 285642 482204 285698
rect 482140 285638 482204 285642
rect 470272 285310 470336 285314
rect 470272 285254 470276 285310
rect 470276 285254 470332 285310
rect 470332 285254 470336 285310
rect 470272 285250 470336 285254
rect 470352 285310 470416 285314
rect 470352 285254 470356 285310
rect 470356 285254 470412 285310
rect 470412 285254 470416 285310
rect 470352 285250 470416 285254
rect 470432 285310 470496 285314
rect 470432 285254 470436 285310
rect 470436 285254 470492 285310
rect 470492 285254 470496 285310
rect 470432 285250 470496 285254
rect 470512 285310 470576 285314
rect 470512 285254 470516 285310
rect 470516 285254 470572 285310
rect 470572 285254 470576 285310
rect 470512 285250 470576 285254
rect 470592 285310 470656 285314
rect 470592 285254 470596 285310
rect 470596 285254 470652 285310
rect 470652 285254 470656 285310
rect 470592 285250 470656 285254
rect 470672 285310 470736 285314
rect 470672 285254 470676 285310
rect 470676 285254 470732 285310
rect 470732 285254 470736 285310
rect 470672 285250 470736 285254
rect 470752 285310 470816 285314
rect 470752 285254 470756 285310
rect 470756 285254 470812 285310
rect 470812 285254 470816 285310
rect 470752 285250 470816 285254
rect 470272 285230 470336 285234
rect 470272 285174 470276 285230
rect 470276 285174 470332 285230
rect 470332 285174 470336 285230
rect 470272 285170 470336 285174
rect 470352 285230 470416 285234
rect 470352 285174 470356 285230
rect 470356 285174 470412 285230
rect 470412 285174 470416 285230
rect 470352 285170 470416 285174
rect 470432 285230 470496 285234
rect 470432 285174 470436 285230
rect 470436 285174 470492 285230
rect 470492 285174 470496 285230
rect 470432 285170 470496 285174
rect 470512 285230 470576 285234
rect 470512 285174 470516 285230
rect 470516 285174 470572 285230
rect 470572 285174 470576 285230
rect 470512 285170 470576 285174
rect 470592 285230 470656 285234
rect 470592 285174 470596 285230
rect 470596 285174 470652 285230
rect 470652 285174 470656 285230
rect 470592 285170 470656 285174
rect 470672 285230 470736 285234
rect 470672 285174 470676 285230
rect 470676 285174 470732 285230
rect 470732 285174 470736 285230
rect 470672 285170 470736 285174
rect 470752 285230 470816 285234
rect 470752 285174 470756 285230
rect 470756 285174 470812 285230
rect 470812 285174 470816 285230
rect 470752 285170 470816 285174
rect 470272 285150 470336 285154
rect 470272 285094 470276 285150
rect 470276 285094 470332 285150
rect 470332 285094 470336 285150
rect 470272 285090 470336 285094
rect 470352 285150 470416 285154
rect 470352 285094 470356 285150
rect 470356 285094 470412 285150
rect 470412 285094 470416 285150
rect 470352 285090 470416 285094
rect 470432 285150 470496 285154
rect 470432 285094 470436 285150
rect 470436 285094 470492 285150
rect 470492 285094 470496 285150
rect 470432 285090 470496 285094
rect 470512 285150 470576 285154
rect 470512 285094 470516 285150
rect 470516 285094 470572 285150
rect 470572 285094 470576 285150
rect 470512 285090 470576 285094
rect 470592 285150 470656 285154
rect 470592 285094 470596 285150
rect 470596 285094 470652 285150
rect 470652 285094 470656 285150
rect 470592 285090 470656 285094
rect 470672 285150 470736 285154
rect 470672 285094 470676 285150
rect 470676 285094 470732 285150
rect 470732 285094 470736 285150
rect 470672 285090 470736 285094
rect 470752 285150 470816 285154
rect 470752 285094 470756 285150
rect 470756 285094 470812 285150
rect 470812 285094 470816 285150
rect 470752 285090 470816 285094
rect 470272 285070 470336 285074
rect 470272 285014 470276 285070
rect 470276 285014 470332 285070
rect 470332 285014 470336 285070
rect 470272 285010 470336 285014
rect 470352 285070 470416 285074
rect 470352 285014 470356 285070
rect 470356 285014 470412 285070
rect 470412 285014 470416 285070
rect 470352 285010 470416 285014
rect 470432 285070 470496 285074
rect 470432 285014 470436 285070
rect 470436 285014 470492 285070
rect 470492 285014 470496 285070
rect 470432 285010 470496 285014
rect 470512 285070 470576 285074
rect 470512 285014 470516 285070
rect 470516 285014 470572 285070
rect 470572 285014 470576 285070
rect 470512 285010 470576 285014
rect 470592 285070 470656 285074
rect 470592 285014 470596 285070
rect 470596 285014 470652 285070
rect 470652 285014 470656 285070
rect 470592 285010 470656 285014
rect 470672 285070 470736 285074
rect 470672 285014 470676 285070
rect 470676 285014 470732 285070
rect 470732 285014 470736 285070
rect 470672 285010 470736 285014
rect 470752 285070 470816 285074
rect 470752 285014 470756 285070
rect 470756 285014 470812 285070
rect 470812 285014 470816 285070
rect 470752 285010 470816 285014
rect 482140 273262 482204 273326
rect 577032 272906 577096 272910
rect 577032 272850 577036 272906
rect 577036 272850 577092 272906
rect 577092 272850 577096 272906
rect 577032 272846 577096 272850
rect 577112 272906 577176 272910
rect 577112 272850 577116 272906
rect 577116 272850 577172 272906
rect 577172 272850 577176 272906
rect 577112 272846 577176 272850
rect 577192 272906 577256 272910
rect 577192 272850 577196 272906
rect 577196 272850 577252 272906
rect 577252 272850 577256 272906
rect 577192 272846 577256 272850
rect 577272 272906 577336 272910
rect 577272 272850 577276 272906
rect 577276 272850 577332 272906
rect 577332 272850 577336 272906
rect 577272 272846 577336 272850
rect 577352 272906 577416 272910
rect 577352 272850 577356 272906
rect 577356 272850 577412 272906
rect 577412 272850 577416 272906
rect 577352 272846 577416 272850
rect 577432 272906 577496 272910
rect 577432 272850 577436 272906
rect 577436 272850 577492 272906
rect 577492 272850 577496 272906
rect 577432 272846 577496 272850
rect 577512 272906 577576 272910
rect 577512 272850 577516 272906
rect 577516 272850 577572 272906
rect 577572 272850 577576 272906
rect 577512 272846 577576 272850
rect 577032 272826 577096 272830
rect 577032 272770 577036 272826
rect 577036 272770 577092 272826
rect 577092 272770 577096 272826
rect 577032 272766 577096 272770
rect 577112 272826 577176 272830
rect 577112 272770 577116 272826
rect 577116 272770 577172 272826
rect 577172 272770 577176 272826
rect 577112 272766 577176 272770
rect 577192 272826 577256 272830
rect 577192 272770 577196 272826
rect 577196 272770 577252 272826
rect 577252 272770 577256 272826
rect 577192 272766 577256 272770
rect 577272 272826 577336 272830
rect 577272 272770 577276 272826
rect 577276 272770 577332 272826
rect 577332 272770 577336 272826
rect 577272 272766 577336 272770
rect 577352 272826 577416 272830
rect 577352 272770 577356 272826
rect 577356 272770 577412 272826
rect 577412 272770 577416 272826
rect 577352 272766 577416 272770
rect 577432 272826 577496 272830
rect 577432 272770 577436 272826
rect 577436 272770 577492 272826
rect 577492 272770 577496 272826
rect 577432 272766 577496 272770
rect 577512 272826 577576 272830
rect 577512 272770 577516 272826
rect 577516 272770 577572 272826
rect 577572 272770 577576 272826
rect 577512 272766 577576 272770
rect 577032 272746 577096 272750
rect 577032 272690 577036 272746
rect 577036 272690 577092 272746
rect 577092 272690 577096 272746
rect 577032 272686 577096 272690
rect 577112 272746 577176 272750
rect 577112 272690 577116 272746
rect 577116 272690 577172 272746
rect 577172 272690 577176 272746
rect 577112 272686 577176 272690
rect 577192 272746 577256 272750
rect 577192 272690 577196 272746
rect 577196 272690 577252 272746
rect 577252 272690 577256 272746
rect 577192 272686 577256 272690
rect 577272 272746 577336 272750
rect 577272 272690 577276 272746
rect 577276 272690 577332 272746
rect 577332 272690 577336 272746
rect 577272 272686 577336 272690
rect 577352 272746 577416 272750
rect 577352 272690 577356 272746
rect 577356 272690 577412 272746
rect 577412 272690 577416 272746
rect 577352 272686 577416 272690
rect 577432 272746 577496 272750
rect 577432 272690 577436 272746
rect 577436 272690 577492 272746
rect 577492 272690 577496 272746
rect 577432 272686 577496 272690
rect 577512 272746 577576 272750
rect 577512 272690 577516 272746
rect 577516 272690 577572 272746
rect 577572 272690 577576 272746
rect 577512 272686 577576 272690
rect 484164 272582 484228 272646
rect 577032 272666 577096 272670
rect 577032 272610 577036 272666
rect 577036 272610 577092 272666
rect 577092 272610 577096 272666
rect 577032 272606 577096 272610
rect 577112 272666 577176 272670
rect 577112 272610 577116 272666
rect 577116 272610 577172 272666
rect 577172 272610 577176 272666
rect 577112 272606 577176 272610
rect 577192 272666 577256 272670
rect 577192 272610 577196 272666
rect 577196 272610 577252 272666
rect 577252 272610 577256 272666
rect 577192 272606 577256 272610
rect 577272 272666 577336 272670
rect 577272 272610 577276 272666
rect 577276 272610 577332 272666
rect 577332 272610 577336 272666
rect 577272 272606 577336 272610
rect 577352 272666 577416 272670
rect 577352 272610 577356 272666
rect 577356 272610 577412 272666
rect 577412 272610 577416 272666
rect 577352 272606 577416 272610
rect 577432 272666 577496 272670
rect 577432 272610 577436 272666
rect 577436 272610 577492 272666
rect 577492 272610 577496 272666
rect 577432 272606 577496 272610
rect 577512 272666 577576 272670
rect 577512 272610 577516 272666
rect 577516 272610 577572 272666
rect 577572 272610 577576 272666
rect 577512 272606 577576 272610
rect 578272 272111 578336 272115
rect 578272 272055 578276 272111
rect 578276 272055 578332 272111
rect 578332 272055 578336 272111
rect 578272 272051 578336 272055
rect 578352 272111 578416 272115
rect 578352 272055 578356 272111
rect 578356 272055 578412 272111
rect 578412 272055 578416 272111
rect 578352 272051 578416 272055
rect 578432 272111 578496 272115
rect 578432 272055 578436 272111
rect 578436 272055 578492 272111
rect 578492 272055 578496 272111
rect 578432 272051 578496 272055
rect 578512 272111 578576 272115
rect 578512 272055 578516 272111
rect 578516 272055 578572 272111
rect 578572 272055 578576 272111
rect 578512 272051 578576 272055
rect 578592 272111 578656 272115
rect 578592 272055 578596 272111
rect 578596 272055 578652 272111
rect 578652 272055 578656 272111
rect 578592 272051 578656 272055
rect 578672 272111 578736 272115
rect 578672 272055 578676 272111
rect 578676 272055 578732 272111
rect 578732 272055 578736 272111
rect 578672 272051 578736 272055
rect 578752 272111 578816 272115
rect 578752 272055 578756 272111
rect 578756 272055 578812 272111
rect 578812 272055 578816 272111
rect 578752 272051 578816 272055
rect 578272 272031 578336 272035
rect 578272 271975 578276 272031
rect 578276 271975 578332 272031
rect 578332 271975 578336 272031
rect 578272 271971 578336 271975
rect 578352 272031 578416 272035
rect 578352 271975 578356 272031
rect 578356 271975 578412 272031
rect 578412 271975 578416 272031
rect 578352 271971 578416 271975
rect 578432 272031 578496 272035
rect 578432 271975 578436 272031
rect 578436 271975 578492 272031
rect 578492 271975 578496 272031
rect 578432 271971 578496 271975
rect 578512 272031 578576 272035
rect 578512 271975 578516 272031
rect 578516 271975 578572 272031
rect 578572 271975 578576 272031
rect 578512 271971 578576 271975
rect 578592 272031 578656 272035
rect 578592 271975 578596 272031
rect 578596 271975 578652 272031
rect 578652 271975 578656 272031
rect 578592 271971 578656 271975
rect 578672 272031 578736 272035
rect 578672 271975 578676 272031
rect 578676 271975 578732 272031
rect 578732 271975 578736 272031
rect 578672 271971 578736 271975
rect 578752 272031 578816 272035
rect 578752 271975 578756 272031
rect 578756 271975 578812 272031
rect 578812 271975 578816 272031
rect 578752 271971 578816 271975
rect 578272 271951 578336 271955
rect 578272 271895 578276 271951
rect 578276 271895 578332 271951
rect 578332 271895 578336 271951
rect 578272 271891 578336 271895
rect 578352 271951 578416 271955
rect 578352 271895 578356 271951
rect 578356 271895 578412 271951
rect 578412 271895 578416 271951
rect 578352 271891 578416 271895
rect 578432 271951 578496 271955
rect 578432 271895 578436 271951
rect 578436 271895 578492 271951
rect 578492 271895 578496 271951
rect 578432 271891 578496 271895
rect 578512 271951 578576 271955
rect 578512 271895 578516 271951
rect 578516 271895 578572 271951
rect 578572 271895 578576 271951
rect 578512 271891 578576 271895
rect 578592 271951 578656 271955
rect 578592 271895 578596 271951
rect 578596 271895 578652 271951
rect 578652 271895 578656 271951
rect 578592 271891 578656 271895
rect 578672 271951 578736 271955
rect 578672 271895 578676 271951
rect 578676 271895 578732 271951
rect 578732 271895 578736 271951
rect 578672 271891 578736 271895
rect 578752 271951 578816 271955
rect 578752 271895 578756 271951
rect 578756 271895 578812 271951
rect 578812 271895 578816 271951
rect 578752 271891 578816 271895
rect 578272 271871 578336 271875
rect 578272 271815 578276 271871
rect 578276 271815 578332 271871
rect 578332 271815 578336 271871
rect 578272 271811 578336 271815
rect 578352 271871 578416 271875
rect 578352 271815 578356 271871
rect 578356 271815 578412 271871
rect 578412 271815 578416 271871
rect 578352 271811 578416 271815
rect 578432 271871 578496 271875
rect 578432 271815 578436 271871
rect 578436 271815 578492 271871
rect 578492 271815 578496 271871
rect 578432 271811 578496 271815
rect 578512 271871 578576 271875
rect 578512 271815 578516 271871
rect 578516 271815 578572 271871
rect 578572 271815 578576 271871
rect 578512 271811 578576 271815
rect 578592 271871 578656 271875
rect 578592 271815 578596 271871
rect 578596 271815 578652 271871
rect 578652 271815 578656 271871
rect 578592 271811 578656 271815
rect 578672 271871 578736 271875
rect 578672 271815 578676 271871
rect 578676 271815 578732 271871
rect 578732 271815 578736 271871
rect 578672 271811 578736 271815
rect 578752 271871 578816 271875
rect 578752 271815 578756 271871
rect 578756 271815 578812 271871
rect 578812 271815 578816 271871
rect 578752 271811 578816 271815
rect 470272 267483 470336 267487
rect 470272 267427 470276 267483
rect 470276 267427 470332 267483
rect 470332 267427 470336 267483
rect 470272 267423 470336 267427
rect 470352 267483 470416 267487
rect 470352 267427 470356 267483
rect 470356 267427 470412 267483
rect 470412 267427 470416 267483
rect 470352 267423 470416 267427
rect 470432 267483 470496 267487
rect 470432 267427 470436 267483
rect 470436 267427 470492 267483
rect 470492 267427 470496 267483
rect 470432 267423 470496 267427
rect 470512 267483 470576 267487
rect 470512 267427 470516 267483
rect 470516 267427 470572 267483
rect 470572 267427 470576 267483
rect 470512 267423 470576 267427
rect 470592 267483 470656 267487
rect 470592 267427 470596 267483
rect 470596 267427 470652 267483
rect 470652 267427 470656 267483
rect 470592 267423 470656 267427
rect 470672 267483 470736 267487
rect 470672 267427 470676 267483
rect 470676 267427 470732 267483
rect 470732 267427 470736 267483
rect 470672 267423 470736 267427
rect 470752 267483 470816 267487
rect 470752 267427 470756 267483
rect 470756 267427 470812 267483
rect 470812 267427 470816 267483
rect 470752 267423 470816 267427
rect 470272 267403 470336 267407
rect 470272 267347 470276 267403
rect 470276 267347 470332 267403
rect 470332 267347 470336 267403
rect 470272 267343 470336 267347
rect 470352 267403 470416 267407
rect 470352 267347 470356 267403
rect 470356 267347 470412 267403
rect 470412 267347 470416 267403
rect 470352 267343 470416 267347
rect 470432 267403 470496 267407
rect 470432 267347 470436 267403
rect 470436 267347 470492 267403
rect 470492 267347 470496 267403
rect 470432 267343 470496 267347
rect 470512 267403 470576 267407
rect 470512 267347 470516 267403
rect 470516 267347 470572 267403
rect 470572 267347 470576 267403
rect 470512 267343 470576 267347
rect 470592 267403 470656 267407
rect 470592 267347 470596 267403
rect 470596 267347 470652 267403
rect 470652 267347 470656 267403
rect 470592 267343 470656 267347
rect 470672 267403 470736 267407
rect 470672 267347 470676 267403
rect 470676 267347 470732 267403
rect 470732 267347 470736 267403
rect 470672 267343 470736 267347
rect 470752 267403 470816 267407
rect 470752 267347 470756 267403
rect 470756 267347 470812 267403
rect 470812 267347 470816 267403
rect 470752 267343 470816 267347
rect 470272 267323 470336 267327
rect 470272 267267 470276 267323
rect 470276 267267 470332 267323
rect 470332 267267 470336 267323
rect 470272 267263 470336 267267
rect 470352 267323 470416 267327
rect 470352 267267 470356 267323
rect 470356 267267 470412 267323
rect 470412 267267 470416 267323
rect 470352 267263 470416 267267
rect 470432 267323 470496 267327
rect 470432 267267 470436 267323
rect 470436 267267 470492 267323
rect 470492 267267 470496 267323
rect 470432 267263 470496 267267
rect 470512 267323 470576 267327
rect 470512 267267 470516 267323
rect 470516 267267 470572 267323
rect 470572 267267 470576 267323
rect 470512 267263 470576 267267
rect 470592 267323 470656 267327
rect 470592 267267 470596 267323
rect 470596 267267 470652 267323
rect 470652 267267 470656 267323
rect 470592 267263 470656 267267
rect 470672 267323 470736 267327
rect 470672 267267 470676 267323
rect 470676 267267 470732 267323
rect 470732 267267 470736 267323
rect 470672 267263 470736 267267
rect 470752 267323 470816 267327
rect 470752 267267 470756 267323
rect 470756 267267 470812 267323
rect 470812 267267 470816 267323
rect 470752 267263 470816 267267
rect 470272 267243 470336 267247
rect 470272 267187 470276 267243
rect 470276 267187 470332 267243
rect 470332 267187 470336 267243
rect 470272 267183 470336 267187
rect 470352 267243 470416 267247
rect 470352 267187 470356 267243
rect 470356 267187 470412 267243
rect 470412 267187 470416 267243
rect 470352 267183 470416 267187
rect 470432 267243 470496 267247
rect 470432 267187 470436 267243
rect 470436 267187 470492 267243
rect 470492 267187 470496 267243
rect 470432 267183 470496 267187
rect 470512 267243 470576 267247
rect 470512 267187 470516 267243
rect 470516 267187 470572 267243
rect 470572 267187 470576 267243
rect 470512 267183 470576 267187
rect 470592 267243 470656 267247
rect 470592 267187 470596 267243
rect 470596 267187 470652 267243
rect 470652 267187 470656 267243
rect 470592 267183 470656 267187
rect 470672 267243 470736 267247
rect 470672 267187 470676 267243
rect 470676 267187 470732 267243
rect 470732 267187 470736 267243
rect 470672 267183 470736 267187
rect 470752 267243 470816 267247
rect 470752 267187 470756 267243
rect 470756 267187 470812 267243
rect 470812 267187 470816 267243
rect 470752 267183 470816 267187
rect 488396 267066 488460 267070
rect 488396 267010 488446 267066
rect 488446 267010 488460 267066
rect 488396 267006 488460 267010
rect 469032 266397 469096 266401
rect 469032 266341 469036 266397
rect 469036 266341 469092 266397
rect 469092 266341 469096 266397
rect 469032 266337 469096 266341
rect 469112 266397 469176 266401
rect 469112 266341 469116 266397
rect 469116 266341 469172 266397
rect 469172 266341 469176 266397
rect 469112 266337 469176 266341
rect 469192 266397 469256 266401
rect 469192 266341 469196 266397
rect 469196 266341 469252 266397
rect 469252 266341 469256 266397
rect 469192 266337 469256 266341
rect 469272 266397 469336 266401
rect 469272 266341 469276 266397
rect 469276 266341 469332 266397
rect 469332 266341 469336 266397
rect 469272 266337 469336 266341
rect 469352 266397 469416 266401
rect 469352 266341 469356 266397
rect 469356 266341 469412 266397
rect 469412 266341 469416 266397
rect 469352 266337 469416 266341
rect 469432 266397 469496 266401
rect 469432 266341 469436 266397
rect 469436 266341 469492 266397
rect 469492 266341 469496 266397
rect 469432 266337 469496 266341
rect 469512 266397 469576 266401
rect 469512 266341 469516 266397
rect 469516 266341 469572 266397
rect 469572 266341 469576 266397
rect 469512 266337 469576 266341
rect 469032 266317 469096 266321
rect 469032 266261 469036 266317
rect 469036 266261 469092 266317
rect 469092 266261 469096 266317
rect 469032 266257 469096 266261
rect 469112 266317 469176 266321
rect 469112 266261 469116 266317
rect 469116 266261 469172 266317
rect 469172 266261 469176 266317
rect 469112 266257 469176 266261
rect 469192 266317 469256 266321
rect 469192 266261 469196 266317
rect 469196 266261 469252 266317
rect 469252 266261 469256 266317
rect 469192 266257 469256 266261
rect 469272 266317 469336 266321
rect 469272 266261 469276 266317
rect 469276 266261 469332 266317
rect 469332 266261 469336 266317
rect 469272 266257 469336 266261
rect 469352 266317 469416 266321
rect 469352 266261 469356 266317
rect 469356 266261 469412 266317
rect 469412 266261 469416 266317
rect 469352 266257 469416 266261
rect 469432 266317 469496 266321
rect 469432 266261 469436 266317
rect 469436 266261 469492 266317
rect 469492 266261 469496 266317
rect 469432 266257 469496 266261
rect 469512 266317 469576 266321
rect 469512 266261 469516 266317
rect 469516 266261 469572 266317
rect 469572 266261 469576 266317
rect 469512 266257 469576 266261
rect 469032 266237 469096 266241
rect 469032 266181 469036 266237
rect 469036 266181 469092 266237
rect 469092 266181 469096 266237
rect 469032 266177 469096 266181
rect 469112 266237 469176 266241
rect 469112 266181 469116 266237
rect 469116 266181 469172 266237
rect 469172 266181 469176 266237
rect 469112 266177 469176 266181
rect 469192 266237 469256 266241
rect 469192 266181 469196 266237
rect 469196 266181 469252 266237
rect 469252 266181 469256 266237
rect 469192 266177 469256 266181
rect 469272 266237 469336 266241
rect 469272 266181 469276 266237
rect 469276 266181 469332 266237
rect 469332 266181 469336 266237
rect 469272 266177 469336 266181
rect 469352 266237 469416 266241
rect 469352 266181 469356 266237
rect 469356 266181 469412 266237
rect 469412 266181 469416 266237
rect 469352 266177 469416 266181
rect 469432 266237 469496 266241
rect 469432 266181 469436 266237
rect 469436 266181 469492 266237
rect 469492 266181 469496 266237
rect 469432 266177 469496 266181
rect 469512 266237 469576 266241
rect 469512 266181 469516 266237
rect 469516 266181 469572 266237
rect 469572 266181 469576 266237
rect 469512 266177 469576 266181
rect 469032 266157 469096 266161
rect 469032 266101 469036 266157
rect 469036 266101 469092 266157
rect 469092 266101 469096 266157
rect 469032 266097 469096 266101
rect 469112 266157 469176 266161
rect 469112 266101 469116 266157
rect 469116 266101 469172 266157
rect 469172 266101 469176 266157
rect 469112 266097 469176 266101
rect 469192 266157 469256 266161
rect 469192 266101 469196 266157
rect 469196 266101 469252 266157
rect 469252 266101 469256 266157
rect 469192 266097 469256 266101
rect 469272 266157 469336 266161
rect 469272 266101 469276 266157
rect 469276 266101 469332 266157
rect 469332 266101 469336 266157
rect 469272 266097 469336 266101
rect 469352 266157 469416 266161
rect 469352 266101 469356 266157
rect 469356 266101 469412 266157
rect 469412 266101 469416 266157
rect 469352 266097 469416 266101
rect 469432 266157 469496 266161
rect 469432 266101 469436 266157
rect 469436 266101 469492 266157
rect 469492 266101 469496 266157
rect 469432 266097 469496 266101
rect 469512 266157 469576 266161
rect 469512 266101 469516 266157
rect 469516 266101 469572 266157
rect 469572 266101 469576 266157
rect 469512 266097 469576 266101
rect 479012 265978 479076 265982
rect 479012 265922 479062 265978
rect 479062 265922 479076 265978
rect 479012 265918 479076 265922
rect 470272 265310 470336 265314
rect 470272 265254 470276 265310
rect 470276 265254 470332 265310
rect 470332 265254 470336 265310
rect 470272 265250 470336 265254
rect 470352 265310 470416 265314
rect 470352 265254 470356 265310
rect 470356 265254 470412 265310
rect 470412 265254 470416 265310
rect 470352 265250 470416 265254
rect 470432 265310 470496 265314
rect 470432 265254 470436 265310
rect 470436 265254 470492 265310
rect 470492 265254 470496 265310
rect 470432 265250 470496 265254
rect 470512 265310 470576 265314
rect 470512 265254 470516 265310
rect 470516 265254 470572 265310
rect 470572 265254 470576 265310
rect 470512 265250 470576 265254
rect 470592 265310 470656 265314
rect 470592 265254 470596 265310
rect 470596 265254 470652 265310
rect 470652 265254 470656 265310
rect 470592 265250 470656 265254
rect 470672 265310 470736 265314
rect 470672 265254 470676 265310
rect 470676 265254 470732 265310
rect 470732 265254 470736 265310
rect 470672 265250 470736 265254
rect 470752 265310 470816 265314
rect 470752 265254 470756 265310
rect 470756 265254 470812 265310
rect 470812 265254 470816 265310
rect 470752 265250 470816 265254
rect 470272 265230 470336 265234
rect 470272 265174 470276 265230
rect 470276 265174 470332 265230
rect 470332 265174 470336 265230
rect 470272 265170 470336 265174
rect 470352 265230 470416 265234
rect 470352 265174 470356 265230
rect 470356 265174 470412 265230
rect 470412 265174 470416 265230
rect 470352 265170 470416 265174
rect 470432 265230 470496 265234
rect 470432 265174 470436 265230
rect 470436 265174 470492 265230
rect 470492 265174 470496 265230
rect 470432 265170 470496 265174
rect 470512 265230 470576 265234
rect 470512 265174 470516 265230
rect 470516 265174 470572 265230
rect 470572 265174 470576 265230
rect 470512 265170 470576 265174
rect 470592 265230 470656 265234
rect 470592 265174 470596 265230
rect 470596 265174 470652 265230
rect 470652 265174 470656 265230
rect 470592 265170 470656 265174
rect 470672 265230 470736 265234
rect 470672 265174 470676 265230
rect 470676 265174 470732 265230
rect 470732 265174 470736 265230
rect 470672 265170 470736 265174
rect 470752 265230 470816 265234
rect 470752 265174 470756 265230
rect 470756 265174 470812 265230
rect 470812 265174 470816 265230
rect 470752 265170 470816 265174
rect 470272 265150 470336 265154
rect 470272 265094 470276 265150
rect 470276 265094 470332 265150
rect 470332 265094 470336 265150
rect 470272 265090 470336 265094
rect 470352 265150 470416 265154
rect 470352 265094 470356 265150
rect 470356 265094 470412 265150
rect 470412 265094 470416 265150
rect 470352 265090 470416 265094
rect 470432 265150 470496 265154
rect 470432 265094 470436 265150
rect 470436 265094 470492 265150
rect 470492 265094 470496 265150
rect 470432 265090 470496 265094
rect 470512 265150 470576 265154
rect 470512 265094 470516 265150
rect 470516 265094 470572 265150
rect 470572 265094 470576 265150
rect 470512 265090 470576 265094
rect 470592 265150 470656 265154
rect 470592 265094 470596 265150
rect 470596 265094 470652 265150
rect 470652 265094 470656 265150
rect 470592 265090 470656 265094
rect 470672 265150 470736 265154
rect 470672 265094 470676 265150
rect 470676 265094 470732 265150
rect 470732 265094 470736 265150
rect 470672 265090 470736 265094
rect 470752 265150 470816 265154
rect 470752 265094 470756 265150
rect 470756 265094 470812 265150
rect 470812 265094 470816 265150
rect 470752 265090 470816 265094
rect 470272 265070 470336 265074
rect 470272 265014 470276 265070
rect 470276 265014 470332 265070
rect 470332 265014 470336 265070
rect 470272 265010 470336 265014
rect 470352 265070 470416 265074
rect 470352 265014 470356 265070
rect 470356 265014 470412 265070
rect 470412 265014 470416 265070
rect 470352 265010 470416 265014
rect 470432 265070 470496 265074
rect 470432 265014 470436 265070
rect 470436 265014 470492 265070
rect 470492 265014 470496 265070
rect 470432 265010 470496 265014
rect 470512 265070 470576 265074
rect 470512 265014 470516 265070
rect 470516 265014 470572 265070
rect 470572 265014 470576 265070
rect 470512 265010 470576 265014
rect 470592 265070 470656 265074
rect 470592 265014 470596 265070
rect 470596 265014 470652 265070
rect 470652 265014 470656 265070
rect 470592 265010 470656 265014
rect 470672 265070 470736 265074
rect 470672 265014 470676 265070
rect 470676 265014 470732 265070
rect 470732 265014 470736 265070
rect 470672 265010 470736 265014
rect 470752 265070 470816 265074
rect 470752 265014 470756 265070
rect 470756 265014 470812 265070
rect 470812 265014 470816 265070
rect 470752 265010 470816 265014
rect 476436 265026 476500 265030
rect 476436 264970 476486 265026
rect 476486 264970 476500 265026
rect 476436 264966 476500 264970
rect 477356 264966 477420 265030
rect 480116 264966 480180 265030
rect 480116 245518 480180 245582
rect 577032 233059 577096 233063
rect 577032 233003 577036 233059
rect 577036 233003 577092 233059
rect 577092 233003 577096 233059
rect 577032 232999 577096 233003
rect 577112 233059 577176 233063
rect 577112 233003 577116 233059
rect 577116 233003 577172 233059
rect 577172 233003 577176 233059
rect 577112 232999 577176 233003
rect 577192 233059 577256 233063
rect 577192 233003 577196 233059
rect 577196 233003 577252 233059
rect 577252 233003 577256 233059
rect 577192 232999 577256 233003
rect 577272 233059 577336 233063
rect 577272 233003 577276 233059
rect 577276 233003 577332 233059
rect 577332 233003 577336 233059
rect 577272 232999 577336 233003
rect 577352 233059 577416 233063
rect 577352 233003 577356 233059
rect 577356 233003 577412 233059
rect 577412 233003 577416 233059
rect 577352 232999 577416 233003
rect 577432 233059 577496 233063
rect 577432 233003 577436 233059
rect 577436 233003 577492 233059
rect 577492 233003 577496 233059
rect 577432 232999 577496 233003
rect 577512 233059 577576 233063
rect 577512 233003 577516 233059
rect 577516 233003 577572 233059
rect 577572 233003 577576 233059
rect 577512 232999 577576 233003
rect 577032 232979 577096 232983
rect 577032 232923 577036 232979
rect 577036 232923 577092 232979
rect 577092 232923 577096 232979
rect 577032 232919 577096 232923
rect 577112 232979 577176 232983
rect 577112 232923 577116 232979
rect 577116 232923 577172 232979
rect 577172 232923 577176 232979
rect 577112 232919 577176 232923
rect 577192 232979 577256 232983
rect 577192 232923 577196 232979
rect 577196 232923 577252 232979
rect 577252 232923 577256 232979
rect 577192 232919 577256 232923
rect 577272 232979 577336 232983
rect 577272 232923 577276 232979
rect 577276 232923 577332 232979
rect 577332 232923 577336 232979
rect 577272 232919 577336 232923
rect 577352 232979 577416 232983
rect 577352 232923 577356 232979
rect 577356 232923 577412 232979
rect 577412 232923 577416 232979
rect 577352 232919 577416 232923
rect 577432 232979 577496 232983
rect 577432 232923 577436 232979
rect 577436 232923 577492 232979
rect 577492 232923 577496 232979
rect 577432 232919 577496 232923
rect 577512 232979 577576 232983
rect 577512 232923 577516 232979
rect 577516 232923 577572 232979
rect 577572 232923 577576 232979
rect 577512 232919 577576 232923
rect 577032 232899 577096 232903
rect 577032 232843 577036 232899
rect 577036 232843 577092 232899
rect 577092 232843 577096 232899
rect 577032 232839 577096 232843
rect 577112 232899 577176 232903
rect 577112 232843 577116 232899
rect 577116 232843 577172 232899
rect 577172 232843 577176 232899
rect 577112 232839 577176 232843
rect 577192 232899 577256 232903
rect 577192 232843 577196 232899
rect 577196 232843 577252 232899
rect 577252 232843 577256 232899
rect 577192 232839 577256 232843
rect 577272 232899 577336 232903
rect 577272 232843 577276 232899
rect 577276 232843 577332 232899
rect 577332 232843 577336 232899
rect 577272 232839 577336 232843
rect 577352 232899 577416 232903
rect 577352 232843 577356 232899
rect 577356 232843 577412 232899
rect 577412 232843 577416 232899
rect 577352 232839 577416 232843
rect 577432 232899 577496 232903
rect 577432 232843 577436 232899
rect 577436 232843 577492 232899
rect 577492 232843 577496 232899
rect 577432 232839 577496 232843
rect 577512 232899 577576 232903
rect 577512 232843 577516 232899
rect 577516 232843 577572 232899
rect 577572 232843 577576 232899
rect 577512 232839 577576 232843
rect 577032 232819 577096 232823
rect 577032 232763 577036 232819
rect 577036 232763 577092 232819
rect 577092 232763 577096 232819
rect 577032 232759 577096 232763
rect 577112 232819 577176 232823
rect 577112 232763 577116 232819
rect 577116 232763 577172 232819
rect 577172 232763 577176 232819
rect 577112 232759 577176 232763
rect 577192 232819 577256 232823
rect 577192 232763 577196 232819
rect 577196 232763 577252 232819
rect 577252 232763 577256 232819
rect 577192 232759 577256 232763
rect 577272 232819 577336 232823
rect 577272 232763 577276 232819
rect 577276 232763 577332 232819
rect 577332 232763 577336 232819
rect 577272 232759 577336 232763
rect 577352 232819 577416 232823
rect 577352 232763 577356 232819
rect 577356 232763 577412 232819
rect 577412 232763 577416 232819
rect 577352 232759 577416 232763
rect 577432 232819 577496 232823
rect 577432 232763 577436 232819
rect 577436 232763 577492 232819
rect 577492 232763 577496 232819
rect 577432 232759 577496 232763
rect 577512 232819 577576 232823
rect 577512 232763 577516 232819
rect 577516 232763 577572 232819
rect 577572 232763 577576 232819
rect 577512 232759 577576 232763
rect 578272 232264 578336 232268
rect 578272 232208 578276 232264
rect 578276 232208 578332 232264
rect 578332 232208 578336 232264
rect 578272 232204 578336 232208
rect 578352 232264 578416 232268
rect 578352 232208 578356 232264
rect 578356 232208 578412 232264
rect 578412 232208 578416 232264
rect 578352 232204 578416 232208
rect 578432 232264 578496 232268
rect 578432 232208 578436 232264
rect 578436 232208 578492 232264
rect 578492 232208 578496 232264
rect 578432 232204 578496 232208
rect 578512 232264 578576 232268
rect 578512 232208 578516 232264
rect 578516 232208 578572 232264
rect 578572 232208 578576 232264
rect 578512 232204 578576 232208
rect 578592 232264 578656 232268
rect 578592 232208 578596 232264
rect 578596 232208 578652 232264
rect 578652 232208 578656 232264
rect 578592 232204 578656 232208
rect 578672 232264 578736 232268
rect 578672 232208 578676 232264
rect 578676 232208 578732 232264
rect 578732 232208 578736 232264
rect 578672 232204 578736 232208
rect 578752 232264 578816 232268
rect 578752 232208 578756 232264
rect 578756 232208 578812 232264
rect 578812 232208 578816 232264
rect 578752 232204 578816 232208
rect 578272 232184 578336 232188
rect 578272 232128 578276 232184
rect 578276 232128 578332 232184
rect 578332 232128 578336 232184
rect 578272 232124 578336 232128
rect 578352 232184 578416 232188
rect 578352 232128 578356 232184
rect 578356 232128 578412 232184
rect 578412 232128 578416 232184
rect 578352 232124 578416 232128
rect 578432 232184 578496 232188
rect 578432 232128 578436 232184
rect 578436 232128 578492 232184
rect 578492 232128 578496 232184
rect 578432 232124 578496 232128
rect 578512 232184 578576 232188
rect 578512 232128 578516 232184
rect 578516 232128 578572 232184
rect 578572 232128 578576 232184
rect 578512 232124 578576 232128
rect 578592 232184 578656 232188
rect 578592 232128 578596 232184
rect 578596 232128 578652 232184
rect 578652 232128 578656 232184
rect 578592 232124 578656 232128
rect 578672 232184 578736 232188
rect 578672 232128 578676 232184
rect 578676 232128 578732 232184
rect 578732 232128 578736 232184
rect 578672 232124 578736 232128
rect 578752 232184 578816 232188
rect 578752 232128 578756 232184
rect 578756 232128 578812 232184
rect 578812 232128 578816 232184
rect 578752 232124 578816 232128
rect 578272 232104 578336 232108
rect 578272 232048 578276 232104
rect 578276 232048 578332 232104
rect 578332 232048 578336 232104
rect 578272 232044 578336 232048
rect 578352 232104 578416 232108
rect 578352 232048 578356 232104
rect 578356 232048 578412 232104
rect 578412 232048 578416 232104
rect 578352 232044 578416 232048
rect 578432 232104 578496 232108
rect 578432 232048 578436 232104
rect 578436 232048 578492 232104
rect 578492 232048 578496 232104
rect 578432 232044 578496 232048
rect 578512 232104 578576 232108
rect 578512 232048 578516 232104
rect 578516 232048 578572 232104
rect 578572 232048 578576 232104
rect 578512 232044 578576 232048
rect 578592 232104 578656 232108
rect 578592 232048 578596 232104
rect 578596 232048 578652 232104
rect 578652 232048 578656 232104
rect 578592 232044 578656 232048
rect 578672 232104 578736 232108
rect 578672 232048 578676 232104
rect 578676 232048 578732 232104
rect 578732 232048 578736 232104
rect 578672 232044 578736 232048
rect 578752 232104 578816 232108
rect 578752 232048 578756 232104
rect 578756 232048 578812 232104
rect 578812 232048 578816 232104
rect 578752 232044 578816 232048
rect 578272 232024 578336 232028
rect 578272 231968 578276 232024
rect 578276 231968 578332 232024
rect 578332 231968 578336 232024
rect 578272 231964 578336 231968
rect 578352 232024 578416 232028
rect 578352 231968 578356 232024
rect 578356 231968 578412 232024
rect 578412 231968 578416 232024
rect 578352 231964 578416 231968
rect 578432 232024 578496 232028
rect 578432 231968 578436 232024
rect 578436 231968 578492 232024
rect 578492 231968 578496 232024
rect 578432 231964 578496 231968
rect 578512 232024 578576 232028
rect 578512 231968 578516 232024
rect 578516 231968 578572 232024
rect 578572 231968 578576 232024
rect 578512 231964 578576 231968
rect 578592 232024 578656 232028
rect 578592 231968 578596 232024
rect 578596 231968 578652 232024
rect 578652 231968 578656 232024
rect 578592 231964 578656 231968
rect 578672 232024 578736 232028
rect 578672 231968 578676 232024
rect 578676 231968 578732 232024
rect 578732 231968 578736 232024
rect 578672 231964 578736 231968
rect 578752 232024 578816 232028
rect 578752 231968 578756 232024
rect 578756 231968 578812 232024
rect 578812 231968 578816 232024
rect 578752 231964 578816 231968
rect 477356 205670 477420 205734
<< metal4 >>
rect -8726 711560 -8106 711592
rect -8726 711324 -8694 711560
rect -8458 711324 -8374 711560
rect -8138 711324 -8106 711560
rect -8726 711240 -8106 711324
rect -8726 711004 -8694 711240
rect -8458 711004 -8374 711240
rect -8138 711004 -8106 711240
rect -8726 695336 -8106 711004
rect -8726 695100 -8694 695336
rect -8458 695100 -8374 695336
rect -8138 695100 -8106 695336
rect -8726 695016 -8106 695100
rect -8726 694780 -8694 695016
rect -8458 694780 -8374 695016
rect -8138 694780 -8106 695016
rect -8726 659336 -8106 694780
rect -8726 659100 -8694 659336
rect -8458 659100 -8374 659336
rect -8138 659100 -8106 659336
rect -8726 659016 -8106 659100
rect -8726 658780 -8694 659016
rect -8458 658780 -8374 659016
rect -8138 658780 -8106 659016
rect -8726 623336 -8106 658780
rect -8726 623100 -8694 623336
rect -8458 623100 -8374 623336
rect -8138 623100 -8106 623336
rect -8726 623016 -8106 623100
rect -8726 622780 -8694 623016
rect -8458 622780 -8374 623016
rect -8138 622780 -8106 623016
rect -8726 587336 -8106 622780
rect -8726 587100 -8694 587336
rect -8458 587100 -8374 587336
rect -8138 587100 -8106 587336
rect -8726 587016 -8106 587100
rect -8726 586780 -8694 587016
rect -8458 586780 -8374 587016
rect -8138 586780 -8106 587016
rect -8726 551336 -8106 586780
rect -8726 551100 -8694 551336
rect -8458 551100 -8374 551336
rect -8138 551100 -8106 551336
rect -8726 551016 -8106 551100
rect -8726 550780 -8694 551016
rect -8458 550780 -8374 551016
rect -8138 550780 -8106 551016
rect -8726 515336 -8106 550780
rect -8726 515100 -8694 515336
rect -8458 515100 -8374 515336
rect -8138 515100 -8106 515336
rect -8726 515016 -8106 515100
rect -8726 514780 -8694 515016
rect -8458 514780 -8374 515016
rect -8138 514780 -8106 515016
rect -8726 479336 -8106 514780
rect -8726 479100 -8694 479336
rect -8458 479100 -8374 479336
rect -8138 479100 -8106 479336
rect -8726 479016 -8106 479100
rect -8726 478780 -8694 479016
rect -8458 478780 -8374 479016
rect -8138 478780 -8106 479016
rect -8726 443336 -8106 478780
rect -8726 443100 -8694 443336
rect -8458 443100 -8374 443336
rect -8138 443100 -8106 443336
rect -8726 443016 -8106 443100
rect -8726 442780 -8694 443016
rect -8458 442780 -8374 443016
rect -8138 442780 -8106 443016
rect -8726 407336 -8106 442780
rect -8726 407100 -8694 407336
rect -8458 407100 -8374 407336
rect -8138 407100 -8106 407336
rect -8726 407016 -8106 407100
rect -8726 406780 -8694 407016
rect -8458 406780 -8374 407016
rect -8138 406780 -8106 407016
rect -8726 371336 -8106 406780
rect -8726 371100 -8694 371336
rect -8458 371100 -8374 371336
rect -8138 371100 -8106 371336
rect -8726 371016 -8106 371100
rect -8726 370780 -8694 371016
rect -8458 370780 -8374 371016
rect -8138 370780 -8106 371016
rect -8726 335336 -8106 370780
rect -8726 335100 -8694 335336
rect -8458 335100 -8374 335336
rect -8138 335100 -8106 335336
rect -8726 335016 -8106 335100
rect -8726 334780 -8694 335016
rect -8458 334780 -8374 335016
rect -8138 334780 -8106 335016
rect -8726 299336 -8106 334780
rect -8726 299100 -8694 299336
rect -8458 299100 -8374 299336
rect -8138 299100 -8106 299336
rect -8726 299016 -8106 299100
rect -8726 298780 -8694 299016
rect -8458 298780 -8374 299016
rect -8138 298780 -8106 299016
rect -8726 263336 -8106 298780
rect -8726 263100 -8694 263336
rect -8458 263100 -8374 263336
rect -8138 263100 -8106 263336
rect -8726 263016 -8106 263100
rect -8726 262780 -8694 263016
rect -8458 262780 -8374 263016
rect -8138 262780 -8106 263016
rect -8726 227336 -8106 262780
rect -8726 227100 -8694 227336
rect -8458 227100 -8374 227336
rect -8138 227100 -8106 227336
rect -8726 227016 -8106 227100
rect -8726 226780 -8694 227016
rect -8458 226780 -8374 227016
rect -8138 226780 -8106 227016
rect -8726 191336 -8106 226780
rect -8726 191100 -8694 191336
rect -8458 191100 -8374 191336
rect -8138 191100 -8106 191336
rect -8726 191016 -8106 191100
rect -8726 190780 -8694 191016
rect -8458 190780 -8374 191016
rect -8138 190780 -8106 191016
rect -8726 155336 -8106 190780
rect -8726 155100 -8694 155336
rect -8458 155100 -8374 155336
rect -8138 155100 -8106 155336
rect -8726 155016 -8106 155100
rect -8726 154780 -8694 155016
rect -8458 154780 -8374 155016
rect -8138 154780 -8106 155016
rect -8726 119336 -8106 154780
rect -8726 119100 -8694 119336
rect -8458 119100 -8374 119336
rect -8138 119100 -8106 119336
rect -8726 119016 -8106 119100
rect -8726 118780 -8694 119016
rect -8458 118780 -8374 119016
rect -8138 118780 -8106 119016
rect -8726 83336 -8106 118780
rect -8726 83100 -8694 83336
rect -8458 83100 -8374 83336
rect -8138 83100 -8106 83336
rect -8726 83016 -8106 83100
rect -8726 82780 -8694 83016
rect -8458 82780 -8374 83016
rect -8138 82780 -8106 83016
rect -8726 47336 -8106 82780
rect -8726 47100 -8694 47336
rect -8458 47100 -8374 47336
rect -8138 47100 -8106 47336
rect -8726 47016 -8106 47100
rect -8726 46780 -8694 47016
rect -8458 46780 -8374 47016
rect -8138 46780 -8106 47016
rect -8726 11336 -8106 46780
rect -8726 11100 -8694 11336
rect -8458 11100 -8374 11336
rect -8138 11100 -8106 11336
rect -8726 11016 -8106 11100
rect -8726 10780 -8694 11016
rect -8458 10780 -8374 11016
rect -8138 10780 -8106 11016
rect -8726 -7064 -8106 10780
rect -7766 710600 -7146 710632
rect -7766 710364 -7734 710600
rect -7498 710364 -7414 710600
rect -7178 710364 -7146 710600
rect -7766 710280 -7146 710364
rect -7766 710044 -7734 710280
rect -7498 710044 -7414 710280
rect -7178 710044 -7146 710280
rect -7766 694096 -7146 710044
rect -7766 693860 -7734 694096
rect -7498 693860 -7414 694096
rect -7178 693860 -7146 694096
rect -7766 693776 -7146 693860
rect -7766 693540 -7734 693776
rect -7498 693540 -7414 693776
rect -7178 693540 -7146 693776
rect -7766 658096 -7146 693540
rect -7766 657860 -7734 658096
rect -7498 657860 -7414 658096
rect -7178 657860 -7146 658096
rect -7766 657776 -7146 657860
rect -7766 657540 -7734 657776
rect -7498 657540 -7414 657776
rect -7178 657540 -7146 657776
rect -7766 622096 -7146 657540
rect -7766 621860 -7734 622096
rect -7498 621860 -7414 622096
rect -7178 621860 -7146 622096
rect -7766 621776 -7146 621860
rect -7766 621540 -7734 621776
rect -7498 621540 -7414 621776
rect -7178 621540 -7146 621776
rect -7766 586096 -7146 621540
rect -7766 585860 -7734 586096
rect -7498 585860 -7414 586096
rect -7178 585860 -7146 586096
rect -7766 585776 -7146 585860
rect -7766 585540 -7734 585776
rect -7498 585540 -7414 585776
rect -7178 585540 -7146 585776
rect -7766 550096 -7146 585540
rect -7766 549860 -7734 550096
rect -7498 549860 -7414 550096
rect -7178 549860 -7146 550096
rect -7766 549776 -7146 549860
rect -7766 549540 -7734 549776
rect -7498 549540 -7414 549776
rect -7178 549540 -7146 549776
rect -7766 514096 -7146 549540
rect -7766 513860 -7734 514096
rect -7498 513860 -7414 514096
rect -7178 513860 -7146 514096
rect -7766 513776 -7146 513860
rect -7766 513540 -7734 513776
rect -7498 513540 -7414 513776
rect -7178 513540 -7146 513776
rect -7766 478096 -7146 513540
rect -7766 477860 -7734 478096
rect -7498 477860 -7414 478096
rect -7178 477860 -7146 478096
rect -7766 477776 -7146 477860
rect -7766 477540 -7734 477776
rect -7498 477540 -7414 477776
rect -7178 477540 -7146 477776
rect -7766 442096 -7146 477540
rect -7766 441860 -7734 442096
rect -7498 441860 -7414 442096
rect -7178 441860 -7146 442096
rect -7766 441776 -7146 441860
rect -7766 441540 -7734 441776
rect -7498 441540 -7414 441776
rect -7178 441540 -7146 441776
rect -7766 406096 -7146 441540
rect -7766 405860 -7734 406096
rect -7498 405860 -7414 406096
rect -7178 405860 -7146 406096
rect -7766 405776 -7146 405860
rect -7766 405540 -7734 405776
rect -7498 405540 -7414 405776
rect -7178 405540 -7146 405776
rect -7766 370096 -7146 405540
rect -7766 369860 -7734 370096
rect -7498 369860 -7414 370096
rect -7178 369860 -7146 370096
rect -7766 369776 -7146 369860
rect -7766 369540 -7734 369776
rect -7498 369540 -7414 369776
rect -7178 369540 -7146 369776
rect -7766 334096 -7146 369540
rect -7766 333860 -7734 334096
rect -7498 333860 -7414 334096
rect -7178 333860 -7146 334096
rect -7766 333776 -7146 333860
rect -7766 333540 -7734 333776
rect -7498 333540 -7414 333776
rect -7178 333540 -7146 333776
rect -7766 298096 -7146 333540
rect -7766 297860 -7734 298096
rect -7498 297860 -7414 298096
rect -7178 297860 -7146 298096
rect -7766 297776 -7146 297860
rect -7766 297540 -7734 297776
rect -7498 297540 -7414 297776
rect -7178 297540 -7146 297776
rect -7766 262096 -7146 297540
rect -7766 261860 -7734 262096
rect -7498 261860 -7414 262096
rect -7178 261860 -7146 262096
rect -7766 261776 -7146 261860
rect -7766 261540 -7734 261776
rect -7498 261540 -7414 261776
rect -7178 261540 -7146 261776
rect -7766 226096 -7146 261540
rect -7766 225860 -7734 226096
rect -7498 225860 -7414 226096
rect -7178 225860 -7146 226096
rect -7766 225776 -7146 225860
rect -7766 225540 -7734 225776
rect -7498 225540 -7414 225776
rect -7178 225540 -7146 225776
rect -7766 190096 -7146 225540
rect -7766 189860 -7734 190096
rect -7498 189860 -7414 190096
rect -7178 189860 -7146 190096
rect -7766 189776 -7146 189860
rect -7766 189540 -7734 189776
rect -7498 189540 -7414 189776
rect -7178 189540 -7146 189776
rect -7766 154096 -7146 189540
rect -7766 153860 -7734 154096
rect -7498 153860 -7414 154096
rect -7178 153860 -7146 154096
rect -7766 153776 -7146 153860
rect -7766 153540 -7734 153776
rect -7498 153540 -7414 153776
rect -7178 153540 -7146 153776
rect -7766 118096 -7146 153540
rect -7766 117860 -7734 118096
rect -7498 117860 -7414 118096
rect -7178 117860 -7146 118096
rect -7766 117776 -7146 117860
rect -7766 117540 -7734 117776
rect -7498 117540 -7414 117776
rect -7178 117540 -7146 117776
rect -7766 82096 -7146 117540
rect -7766 81860 -7734 82096
rect -7498 81860 -7414 82096
rect -7178 81860 -7146 82096
rect -7766 81776 -7146 81860
rect -7766 81540 -7734 81776
rect -7498 81540 -7414 81776
rect -7178 81540 -7146 81776
rect -7766 46096 -7146 81540
rect -7766 45860 -7734 46096
rect -7498 45860 -7414 46096
rect -7178 45860 -7146 46096
rect -7766 45776 -7146 45860
rect -7766 45540 -7734 45776
rect -7498 45540 -7414 45776
rect -7178 45540 -7146 45776
rect -7766 10096 -7146 45540
rect -7766 9860 -7734 10096
rect -7498 9860 -7414 10096
rect -7178 9860 -7146 10096
rect -7766 9776 -7146 9860
rect -7766 9540 -7734 9776
rect -7498 9540 -7414 9776
rect -7178 9540 -7146 9776
rect -7766 -6104 -7146 9540
rect -6806 709640 -6186 709672
rect -6806 709404 -6774 709640
rect -6538 709404 -6454 709640
rect -6218 709404 -6186 709640
rect -6806 709320 -6186 709404
rect -6806 709084 -6774 709320
rect -6538 709084 -6454 709320
rect -6218 709084 -6186 709320
rect -6806 692856 -6186 709084
rect -6806 692620 -6774 692856
rect -6538 692620 -6454 692856
rect -6218 692620 -6186 692856
rect -6806 692536 -6186 692620
rect -6806 692300 -6774 692536
rect -6538 692300 -6454 692536
rect -6218 692300 -6186 692536
rect -6806 656856 -6186 692300
rect -6806 656620 -6774 656856
rect -6538 656620 -6454 656856
rect -6218 656620 -6186 656856
rect -6806 656536 -6186 656620
rect -6806 656300 -6774 656536
rect -6538 656300 -6454 656536
rect -6218 656300 -6186 656536
rect -6806 620856 -6186 656300
rect -6806 620620 -6774 620856
rect -6538 620620 -6454 620856
rect -6218 620620 -6186 620856
rect -6806 620536 -6186 620620
rect -6806 620300 -6774 620536
rect -6538 620300 -6454 620536
rect -6218 620300 -6186 620536
rect -6806 584856 -6186 620300
rect -6806 584620 -6774 584856
rect -6538 584620 -6454 584856
rect -6218 584620 -6186 584856
rect -6806 584536 -6186 584620
rect -6806 584300 -6774 584536
rect -6538 584300 -6454 584536
rect -6218 584300 -6186 584536
rect -6806 548856 -6186 584300
rect -6806 548620 -6774 548856
rect -6538 548620 -6454 548856
rect -6218 548620 -6186 548856
rect -6806 548536 -6186 548620
rect -6806 548300 -6774 548536
rect -6538 548300 -6454 548536
rect -6218 548300 -6186 548536
rect -6806 512856 -6186 548300
rect -6806 512620 -6774 512856
rect -6538 512620 -6454 512856
rect -6218 512620 -6186 512856
rect -6806 512536 -6186 512620
rect -6806 512300 -6774 512536
rect -6538 512300 -6454 512536
rect -6218 512300 -6186 512536
rect -6806 476856 -6186 512300
rect -6806 476620 -6774 476856
rect -6538 476620 -6454 476856
rect -6218 476620 -6186 476856
rect -6806 476536 -6186 476620
rect -6806 476300 -6774 476536
rect -6538 476300 -6454 476536
rect -6218 476300 -6186 476536
rect -6806 440856 -6186 476300
rect -6806 440620 -6774 440856
rect -6538 440620 -6454 440856
rect -6218 440620 -6186 440856
rect -6806 440536 -6186 440620
rect -6806 440300 -6774 440536
rect -6538 440300 -6454 440536
rect -6218 440300 -6186 440536
rect -6806 404856 -6186 440300
rect -6806 404620 -6774 404856
rect -6538 404620 -6454 404856
rect -6218 404620 -6186 404856
rect -6806 404536 -6186 404620
rect -6806 404300 -6774 404536
rect -6538 404300 -6454 404536
rect -6218 404300 -6186 404536
rect -6806 368856 -6186 404300
rect -6806 368620 -6774 368856
rect -6538 368620 -6454 368856
rect -6218 368620 -6186 368856
rect -6806 368536 -6186 368620
rect -6806 368300 -6774 368536
rect -6538 368300 -6454 368536
rect -6218 368300 -6186 368536
rect -6806 332856 -6186 368300
rect -6806 332620 -6774 332856
rect -6538 332620 -6454 332856
rect -6218 332620 -6186 332856
rect -6806 332536 -6186 332620
rect -6806 332300 -6774 332536
rect -6538 332300 -6454 332536
rect -6218 332300 -6186 332536
rect -6806 296856 -6186 332300
rect -6806 296620 -6774 296856
rect -6538 296620 -6454 296856
rect -6218 296620 -6186 296856
rect -6806 296536 -6186 296620
rect -6806 296300 -6774 296536
rect -6538 296300 -6454 296536
rect -6218 296300 -6186 296536
rect -6806 260856 -6186 296300
rect -6806 260620 -6774 260856
rect -6538 260620 -6454 260856
rect -6218 260620 -6186 260856
rect -6806 260536 -6186 260620
rect -6806 260300 -6774 260536
rect -6538 260300 -6454 260536
rect -6218 260300 -6186 260536
rect -6806 224856 -6186 260300
rect -6806 224620 -6774 224856
rect -6538 224620 -6454 224856
rect -6218 224620 -6186 224856
rect -6806 224536 -6186 224620
rect -6806 224300 -6774 224536
rect -6538 224300 -6454 224536
rect -6218 224300 -6186 224536
rect -6806 188856 -6186 224300
rect -6806 188620 -6774 188856
rect -6538 188620 -6454 188856
rect -6218 188620 -6186 188856
rect -6806 188536 -6186 188620
rect -6806 188300 -6774 188536
rect -6538 188300 -6454 188536
rect -6218 188300 -6186 188536
rect -6806 152856 -6186 188300
rect -6806 152620 -6774 152856
rect -6538 152620 -6454 152856
rect -6218 152620 -6186 152856
rect -6806 152536 -6186 152620
rect -6806 152300 -6774 152536
rect -6538 152300 -6454 152536
rect -6218 152300 -6186 152536
rect -6806 116856 -6186 152300
rect -6806 116620 -6774 116856
rect -6538 116620 -6454 116856
rect -6218 116620 -6186 116856
rect -6806 116536 -6186 116620
rect -6806 116300 -6774 116536
rect -6538 116300 -6454 116536
rect -6218 116300 -6186 116536
rect -6806 80856 -6186 116300
rect -6806 80620 -6774 80856
rect -6538 80620 -6454 80856
rect -6218 80620 -6186 80856
rect -6806 80536 -6186 80620
rect -6806 80300 -6774 80536
rect -6538 80300 -6454 80536
rect -6218 80300 -6186 80536
rect -6806 44856 -6186 80300
rect -6806 44620 -6774 44856
rect -6538 44620 -6454 44856
rect -6218 44620 -6186 44856
rect -6806 44536 -6186 44620
rect -6806 44300 -6774 44536
rect -6538 44300 -6454 44536
rect -6218 44300 -6186 44536
rect -6806 8856 -6186 44300
rect -6806 8620 -6774 8856
rect -6538 8620 -6454 8856
rect -6218 8620 -6186 8856
rect -6806 8536 -6186 8620
rect -6806 8300 -6774 8536
rect -6538 8300 -6454 8536
rect -6218 8300 -6186 8536
rect -6806 -5144 -6186 8300
rect -5846 708680 -5226 708712
rect -5846 708444 -5814 708680
rect -5578 708444 -5494 708680
rect -5258 708444 -5226 708680
rect -5846 708360 -5226 708444
rect -5846 708124 -5814 708360
rect -5578 708124 -5494 708360
rect -5258 708124 -5226 708360
rect -5846 691616 -5226 708124
rect -5846 691380 -5814 691616
rect -5578 691380 -5494 691616
rect -5258 691380 -5226 691616
rect -5846 691296 -5226 691380
rect -5846 691060 -5814 691296
rect -5578 691060 -5494 691296
rect -5258 691060 -5226 691296
rect -5846 655616 -5226 691060
rect -5846 655380 -5814 655616
rect -5578 655380 -5494 655616
rect -5258 655380 -5226 655616
rect -5846 655296 -5226 655380
rect -5846 655060 -5814 655296
rect -5578 655060 -5494 655296
rect -5258 655060 -5226 655296
rect -5846 619616 -5226 655060
rect -5846 619380 -5814 619616
rect -5578 619380 -5494 619616
rect -5258 619380 -5226 619616
rect -5846 619296 -5226 619380
rect -5846 619060 -5814 619296
rect -5578 619060 -5494 619296
rect -5258 619060 -5226 619296
rect -5846 583616 -5226 619060
rect -5846 583380 -5814 583616
rect -5578 583380 -5494 583616
rect -5258 583380 -5226 583616
rect -5846 583296 -5226 583380
rect -5846 583060 -5814 583296
rect -5578 583060 -5494 583296
rect -5258 583060 -5226 583296
rect -5846 547616 -5226 583060
rect -5846 547380 -5814 547616
rect -5578 547380 -5494 547616
rect -5258 547380 -5226 547616
rect -5846 547296 -5226 547380
rect -5846 547060 -5814 547296
rect -5578 547060 -5494 547296
rect -5258 547060 -5226 547296
rect -5846 511616 -5226 547060
rect -5846 511380 -5814 511616
rect -5578 511380 -5494 511616
rect -5258 511380 -5226 511616
rect -5846 511296 -5226 511380
rect -5846 511060 -5814 511296
rect -5578 511060 -5494 511296
rect -5258 511060 -5226 511296
rect -5846 475616 -5226 511060
rect -5846 475380 -5814 475616
rect -5578 475380 -5494 475616
rect -5258 475380 -5226 475616
rect -5846 475296 -5226 475380
rect -5846 475060 -5814 475296
rect -5578 475060 -5494 475296
rect -5258 475060 -5226 475296
rect -5846 439616 -5226 475060
rect -5846 439380 -5814 439616
rect -5578 439380 -5494 439616
rect -5258 439380 -5226 439616
rect -5846 439296 -5226 439380
rect -5846 439060 -5814 439296
rect -5578 439060 -5494 439296
rect -5258 439060 -5226 439296
rect -5846 403616 -5226 439060
rect -5846 403380 -5814 403616
rect -5578 403380 -5494 403616
rect -5258 403380 -5226 403616
rect -5846 403296 -5226 403380
rect -5846 403060 -5814 403296
rect -5578 403060 -5494 403296
rect -5258 403060 -5226 403296
rect -5846 367616 -5226 403060
rect -5846 367380 -5814 367616
rect -5578 367380 -5494 367616
rect -5258 367380 -5226 367616
rect -5846 367296 -5226 367380
rect -5846 367060 -5814 367296
rect -5578 367060 -5494 367296
rect -5258 367060 -5226 367296
rect -5846 331616 -5226 367060
rect -5846 331380 -5814 331616
rect -5578 331380 -5494 331616
rect -5258 331380 -5226 331616
rect -5846 331296 -5226 331380
rect -5846 331060 -5814 331296
rect -5578 331060 -5494 331296
rect -5258 331060 -5226 331296
rect -5846 295616 -5226 331060
rect -5846 295380 -5814 295616
rect -5578 295380 -5494 295616
rect -5258 295380 -5226 295616
rect -5846 295296 -5226 295380
rect -5846 295060 -5814 295296
rect -5578 295060 -5494 295296
rect -5258 295060 -5226 295296
rect -5846 259616 -5226 295060
rect -5846 259380 -5814 259616
rect -5578 259380 -5494 259616
rect -5258 259380 -5226 259616
rect -5846 259296 -5226 259380
rect -5846 259060 -5814 259296
rect -5578 259060 -5494 259296
rect -5258 259060 -5226 259296
rect -5846 223616 -5226 259060
rect -5846 223380 -5814 223616
rect -5578 223380 -5494 223616
rect -5258 223380 -5226 223616
rect -5846 223296 -5226 223380
rect -5846 223060 -5814 223296
rect -5578 223060 -5494 223296
rect -5258 223060 -5226 223296
rect -5846 187616 -5226 223060
rect -5846 187380 -5814 187616
rect -5578 187380 -5494 187616
rect -5258 187380 -5226 187616
rect -5846 187296 -5226 187380
rect -5846 187060 -5814 187296
rect -5578 187060 -5494 187296
rect -5258 187060 -5226 187296
rect -5846 151616 -5226 187060
rect -5846 151380 -5814 151616
rect -5578 151380 -5494 151616
rect -5258 151380 -5226 151616
rect -5846 151296 -5226 151380
rect -5846 151060 -5814 151296
rect -5578 151060 -5494 151296
rect -5258 151060 -5226 151296
rect -5846 115616 -5226 151060
rect -5846 115380 -5814 115616
rect -5578 115380 -5494 115616
rect -5258 115380 -5226 115616
rect -5846 115296 -5226 115380
rect -5846 115060 -5814 115296
rect -5578 115060 -5494 115296
rect -5258 115060 -5226 115296
rect -5846 79616 -5226 115060
rect -5846 79380 -5814 79616
rect -5578 79380 -5494 79616
rect -5258 79380 -5226 79616
rect -5846 79296 -5226 79380
rect -5846 79060 -5814 79296
rect -5578 79060 -5494 79296
rect -5258 79060 -5226 79296
rect -5846 43616 -5226 79060
rect -5846 43380 -5814 43616
rect -5578 43380 -5494 43616
rect -5258 43380 -5226 43616
rect -5846 43296 -5226 43380
rect -5846 43060 -5814 43296
rect -5578 43060 -5494 43296
rect -5258 43060 -5226 43296
rect -5846 7616 -5226 43060
rect -5846 7380 -5814 7616
rect -5578 7380 -5494 7616
rect -5258 7380 -5226 7616
rect -5846 7296 -5226 7380
rect -5846 7060 -5814 7296
rect -5578 7060 -5494 7296
rect -5258 7060 -5226 7296
rect -5846 -4184 -5226 7060
rect -4886 707720 -4266 707752
rect -4886 707484 -4854 707720
rect -4618 707484 -4534 707720
rect -4298 707484 -4266 707720
rect -4886 707400 -4266 707484
rect -4886 707164 -4854 707400
rect -4618 707164 -4534 707400
rect -4298 707164 -4266 707400
rect -4886 690376 -4266 707164
rect -4886 690140 -4854 690376
rect -4618 690140 -4534 690376
rect -4298 690140 -4266 690376
rect -4886 690056 -4266 690140
rect -4886 689820 -4854 690056
rect -4618 689820 -4534 690056
rect -4298 689820 -4266 690056
rect -4886 654376 -4266 689820
rect -4886 654140 -4854 654376
rect -4618 654140 -4534 654376
rect -4298 654140 -4266 654376
rect -4886 654056 -4266 654140
rect -4886 653820 -4854 654056
rect -4618 653820 -4534 654056
rect -4298 653820 -4266 654056
rect -4886 618376 -4266 653820
rect -4886 618140 -4854 618376
rect -4618 618140 -4534 618376
rect -4298 618140 -4266 618376
rect -4886 618056 -4266 618140
rect -4886 617820 -4854 618056
rect -4618 617820 -4534 618056
rect -4298 617820 -4266 618056
rect -4886 582376 -4266 617820
rect -4886 582140 -4854 582376
rect -4618 582140 -4534 582376
rect -4298 582140 -4266 582376
rect -4886 582056 -4266 582140
rect -4886 581820 -4854 582056
rect -4618 581820 -4534 582056
rect -4298 581820 -4266 582056
rect -4886 546376 -4266 581820
rect -4886 546140 -4854 546376
rect -4618 546140 -4534 546376
rect -4298 546140 -4266 546376
rect -4886 546056 -4266 546140
rect -4886 545820 -4854 546056
rect -4618 545820 -4534 546056
rect -4298 545820 -4266 546056
rect -4886 510376 -4266 545820
rect -4886 510140 -4854 510376
rect -4618 510140 -4534 510376
rect -4298 510140 -4266 510376
rect -4886 510056 -4266 510140
rect -4886 509820 -4854 510056
rect -4618 509820 -4534 510056
rect -4298 509820 -4266 510056
rect -4886 474376 -4266 509820
rect -4886 474140 -4854 474376
rect -4618 474140 -4534 474376
rect -4298 474140 -4266 474376
rect -4886 474056 -4266 474140
rect -4886 473820 -4854 474056
rect -4618 473820 -4534 474056
rect -4298 473820 -4266 474056
rect -4886 438376 -4266 473820
rect -4886 438140 -4854 438376
rect -4618 438140 -4534 438376
rect -4298 438140 -4266 438376
rect -4886 438056 -4266 438140
rect -4886 437820 -4854 438056
rect -4618 437820 -4534 438056
rect -4298 437820 -4266 438056
rect -4886 402376 -4266 437820
rect -4886 402140 -4854 402376
rect -4618 402140 -4534 402376
rect -4298 402140 -4266 402376
rect -4886 402056 -4266 402140
rect -4886 401820 -4854 402056
rect -4618 401820 -4534 402056
rect -4298 401820 -4266 402056
rect -4886 366376 -4266 401820
rect -4886 366140 -4854 366376
rect -4618 366140 -4534 366376
rect -4298 366140 -4266 366376
rect -4886 366056 -4266 366140
rect -4886 365820 -4854 366056
rect -4618 365820 -4534 366056
rect -4298 365820 -4266 366056
rect -4886 330376 -4266 365820
rect -4886 330140 -4854 330376
rect -4618 330140 -4534 330376
rect -4298 330140 -4266 330376
rect -4886 330056 -4266 330140
rect -4886 329820 -4854 330056
rect -4618 329820 -4534 330056
rect -4298 329820 -4266 330056
rect -4886 294376 -4266 329820
rect -4886 294140 -4854 294376
rect -4618 294140 -4534 294376
rect -4298 294140 -4266 294376
rect -4886 294056 -4266 294140
rect -4886 293820 -4854 294056
rect -4618 293820 -4534 294056
rect -4298 293820 -4266 294056
rect -4886 258376 -4266 293820
rect -4886 258140 -4854 258376
rect -4618 258140 -4534 258376
rect -4298 258140 -4266 258376
rect -4886 258056 -4266 258140
rect -4886 257820 -4854 258056
rect -4618 257820 -4534 258056
rect -4298 257820 -4266 258056
rect -4886 222376 -4266 257820
rect -4886 222140 -4854 222376
rect -4618 222140 -4534 222376
rect -4298 222140 -4266 222376
rect -4886 222056 -4266 222140
rect -4886 221820 -4854 222056
rect -4618 221820 -4534 222056
rect -4298 221820 -4266 222056
rect -4886 186376 -4266 221820
rect -4886 186140 -4854 186376
rect -4618 186140 -4534 186376
rect -4298 186140 -4266 186376
rect -4886 186056 -4266 186140
rect -4886 185820 -4854 186056
rect -4618 185820 -4534 186056
rect -4298 185820 -4266 186056
rect -4886 150376 -4266 185820
rect -4886 150140 -4854 150376
rect -4618 150140 -4534 150376
rect -4298 150140 -4266 150376
rect -4886 150056 -4266 150140
rect -4886 149820 -4854 150056
rect -4618 149820 -4534 150056
rect -4298 149820 -4266 150056
rect -4886 114376 -4266 149820
rect -4886 114140 -4854 114376
rect -4618 114140 -4534 114376
rect -4298 114140 -4266 114376
rect -4886 114056 -4266 114140
rect -4886 113820 -4854 114056
rect -4618 113820 -4534 114056
rect -4298 113820 -4266 114056
rect -4886 78376 -4266 113820
rect -4886 78140 -4854 78376
rect -4618 78140 -4534 78376
rect -4298 78140 -4266 78376
rect -4886 78056 -4266 78140
rect -4886 77820 -4854 78056
rect -4618 77820 -4534 78056
rect -4298 77820 -4266 78056
rect -4886 42376 -4266 77820
rect -4886 42140 -4854 42376
rect -4618 42140 -4534 42376
rect -4298 42140 -4266 42376
rect -4886 42056 -4266 42140
rect -4886 41820 -4854 42056
rect -4618 41820 -4534 42056
rect -4298 41820 -4266 42056
rect -4886 6376 -4266 41820
rect -4886 6140 -4854 6376
rect -4618 6140 -4534 6376
rect -4298 6140 -4266 6376
rect -4886 6056 -4266 6140
rect -4886 5820 -4854 6056
rect -4618 5820 -4534 6056
rect -4298 5820 -4266 6056
rect -4886 -3224 -4266 5820
rect -3926 706760 -3306 706792
rect -3926 706524 -3894 706760
rect -3658 706524 -3574 706760
rect -3338 706524 -3306 706760
rect -3926 706440 -3306 706524
rect -3926 706204 -3894 706440
rect -3658 706204 -3574 706440
rect -3338 706204 -3306 706440
rect -3926 689136 -3306 706204
rect -3926 688900 -3894 689136
rect -3658 688900 -3574 689136
rect -3338 688900 -3306 689136
rect -3926 688816 -3306 688900
rect -3926 688580 -3894 688816
rect -3658 688580 -3574 688816
rect -3338 688580 -3306 688816
rect -3926 653136 -3306 688580
rect -3926 652900 -3894 653136
rect -3658 652900 -3574 653136
rect -3338 652900 -3306 653136
rect -3926 652816 -3306 652900
rect -3926 652580 -3894 652816
rect -3658 652580 -3574 652816
rect -3338 652580 -3306 652816
rect -3926 617136 -3306 652580
rect -3926 616900 -3894 617136
rect -3658 616900 -3574 617136
rect -3338 616900 -3306 617136
rect -3926 616816 -3306 616900
rect -3926 616580 -3894 616816
rect -3658 616580 -3574 616816
rect -3338 616580 -3306 616816
rect -3926 581136 -3306 616580
rect -3926 580900 -3894 581136
rect -3658 580900 -3574 581136
rect -3338 580900 -3306 581136
rect -3926 580816 -3306 580900
rect -3926 580580 -3894 580816
rect -3658 580580 -3574 580816
rect -3338 580580 -3306 580816
rect -3926 545136 -3306 580580
rect -3926 544900 -3894 545136
rect -3658 544900 -3574 545136
rect -3338 544900 -3306 545136
rect -3926 544816 -3306 544900
rect -3926 544580 -3894 544816
rect -3658 544580 -3574 544816
rect -3338 544580 -3306 544816
rect -3926 509136 -3306 544580
rect -3926 508900 -3894 509136
rect -3658 508900 -3574 509136
rect -3338 508900 -3306 509136
rect -3926 508816 -3306 508900
rect -3926 508580 -3894 508816
rect -3658 508580 -3574 508816
rect -3338 508580 -3306 508816
rect -3926 473136 -3306 508580
rect -3926 472900 -3894 473136
rect -3658 472900 -3574 473136
rect -3338 472900 -3306 473136
rect -3926 472816 -3306 472900
rect -3926 472580 -3894 472816
rect -3658 472580 -3574 472816
rect -3338 472580 -3306 472816
rect -3926 437136 -3306 472580
rect -3926 436900 -3894 437136
rect -3658 436900 -3574 437136
rect -3338 436900 -3306 437136
rect -3926 436816 -3306 436900
rect -3926 436580 -3894 436816
rect -3658 436580 -3574 436816
rect -3338 436580 -3306 436816
rect -3926 401136 -3306 436580
rect -3926 400900 -3894 401136
rect -3658 400900 -3574 401136
rect -3338 400900 -3306 401136
rect -3926 400816 -3306 400900
rect -3926 400580 -3894 400816
rect -3658 400580 -3574 400816
rect -3338 400580 -3306 400816
rect -3926 365136 -3306 400580
rect -3926 364900 -3894 365136
rect -3658 364900 -3574 365136
rect -3338 364900 -3306 365136
rect -3926 364816 -3306 364900
rect -3926 364580 -3894 364816
rect -3658 364580 -3574 364816
rect -3338 364580 -3306 364816
rect -3926 329136 -3306 364580
rect -3926 328900 -3894 329136
rect -3658 328900 -3574 329136
rect -3338 328900 -3306 329136
rect -3926 328816 -3306 328900
rect -3926 328580 -3894 328816
rect -3658 328580 -3574 328816
rect -3338 328580 -3306 328816
rect -3926 293136 -3306 328580
rect -3926 292900 -3894 293136
rect -3658 292900 -3574 293136
rect -3338 292900 -3306 293136
rect -3926 292816 -3306 292900
rect -3926 292580 -3894 292816
rect -3658 292580 -3574 292816
rect -3338 292580 -3306 292816
rect -3926 257136 -3306 292580
rect -3926 256900 -3894 257136
rect -3658 256900 -3574 257136
rect -3338 256900 -3306 257136
rect -3926 256816 -3306 256900
rect -3926 256580 -3894 256816
rect -3658 256580 -3574 256816
rect -3338 256580 -3306 256816
rect -3926 221136 -3306 256580
rect -3926 220900 -3894 221136
rect -3658 220900 -3574 221136
rect -3338 220900 -3306 221136
rect -3926 220816 -3306 220900
rect -3926 220580 -3894 220816
rect -3658 220580 -3574 220816
rect -3338 220580 -3306 220816
rect -3926 185136 -3306 220580
rect -3926 184900 -3894 185136
rect -3658 184900 -3574 185136
rect -3338 184900 -3306 185136
rect -3926 184816 -3306 184900
rect -3926 184580 -3894 184816
rect -3658 184580 -3574 184816
rect -3338 184580 -3306 184816
rect -3926 149136 -3306 184580
rect -3926 148900 -3894 149136
rect -3658 148900 -3574 149136
rect -3338 148900 -3306 149136
rect -3926 148816 -3306 148900
rect -3926 148580 -3894 148816
rect -3658 148580 -3574 148816
rect -3338 148580 -3306 148816
rect -3926 113136 -3306 148580
rect -3926 112900 -3894 113136
rect -3658 112900 -3574 113136
rect -3338 112900 -3306 113136
rect -3926 112816 -3306 112900
rect -3926 112580 -3894 112816
rect -3658 112580 -3574 112816
rect -3338 112580 -3306 112816
rect -3926 77136 -3306 112580
rect -3926 76900 -3894 77136
rect -3658 76900 -3574 77136
rect -3338 76900 -3306 77136
rect -3926 76816 -3306 76900
rect -3926 76580 -3894 76816
rect -3658 76580 -3574 76816
rect -3338 76580 -3306 76816
rect -3926 41136 -3306 76580
rect -3926 40900 -3894 41136
rect -3658 40900 -3574 41136
rect -3338 40900 -3306 41136
rect -3926 40816 -3306 40900
rect -3926 40580 -3894 40816
rect -3658 40580 -3574 40816
rect -3338 40580 -3306 40816
rect -3926 5136 -3306 40580
rect -3926 4900 -3894 5136
rect -3658 4900 -3574 5136
rect -3338 4900 -3306 5136
rect -3926 4816 -3306 4900
rect -3926 4580 -3894 4816
rect -3658 4580 -3574 4816
rect -3338 4580 -3306 4816
rect -3926 -2264 -3306 4580
rect -2966 705800 -2346 705832
rect -2966 705564 -2934 705800
rect -2698 705564 -2614 705800
rect -2378 705564 -2346 705800
rect -2966 705480 -2346 705564
rect -2966 705244 -2934 705480
rect -2698 705244 -2614 705480
rect -2378 705244 -2346 705480
rect -2966 687896 -2346 705244
rect -2966 687660 -2934 687896
rect -2698 687660 -2614 687896
rect -2378 687660 -2346 687896
rect -2966 687576 -2346 687660
rect -2966 687340 -2934 687576
rect -2698 687340 -2614 687576
rect -2378 687340 -2346 687576
rect -2966 651896 -2346 687340
rect -2966 651660 -2934 651896
rect -2698 651660 -2614 651896
rect -2378 651660 -2346 651896
rect -2966 651576 -2346 651660
rect -2966 651340 -2934 651576
rect -2698 651340 -2614 651576
rect -2378 651340 -2346 651576
rect -2966 615896 -2346 651340
rect -2966 615660 -2934 615896
rect -2698 615660 -2614 615896
rect -2378 615660 -2346 615896
rect -2966 615576 -2346 615660
rect -2966 615340 -2934 615576
rect -2698 615340 -2614 615576
rect -2378 615340 -2346 615576
rect -2966 579896 -2346 615340
rect -2966 579660 -2934 579896
rect -2698 579660 -2614 579896
rect -2378 579660 -2346 579896
rect -2966 579576 -2346 579660
rect -2966 579340 -2934 579576
rect -2698 579340 -2614 579576
rect -2378 579340 -2346 579576
rect -2966 543896 -2346 579340
rect -2966 543660 -2934 543896
rect -2698 543660 -2614 543896
rect -2378 543660 -2346 543896
rect -2966 543576 -2346 543660
rect -2966 543340 -2934 543576
rect -2698 543340 -2614 543576
rect -2378 543340 -2346 543576
rect -2966 507896 -2346 543340
rect -2966 507660 -2934 507896
rect -2698 507660 -2614 507896
rect -2378 507660 -2346 507896
rect -2966 507576 -2346 507660
rect -2966 507340 -2934 507576
rect -2698 507340 -2614 507576
rect -2378 507340 -2346 507576
rect -2966 471896 -2346 507340
rect -2966 471660 -2934 471896
rect -2698 471660 -2614 471896
rect -2378 471660 -2346 471896
rect -2966 471576 -2346 471660
rect -2966 471340 -2934 471576
rect -2698 471340 -2614 471576
rect -2378 471340 -2346 471576
rect -2966 435896 -2346 471340
rect -2966 435660 -2934 435896
rect -2698 435660 -2614 435896
rect -2378 435660 -2346 435896
rect -2966 435576 -2346 435660
rect -2966 435340 -2934 435576
rect -2698 435340 -2614 435576
rect -2378 435340 -2346 435576
rect -2966 399896 -2346 435340
rect -2966 399660 -2934 399896
rect -2698 399660 -2614 399896
rect -2378 399660 -2346 399896
rect -2966 399576 -2346 399660
rect -2966 399340 -2934 399576
rect -2698 399340 -2614 399576
rect -2378 399340 -2346 399576
rect -2966 363896 -2346 399340
rect -2966 363660 -2934 363896
rect -2698 363660 -2614 363896
rect -2378 363660 -2346 363896
rect -2966 363576 -2346 363660
rect -2966 363340 -2934 363576
rect -2698 363340 -2614 363576
rect -2378 363340 -2346 363576
rect -2966 327896 -2346 363340
rect -2966 327660 -2934 327896
rect -2698 327660 -2614 327896
rect -2378 327660 -2346 327896
rect -2966 327576 -2346 327660
rect -2966 327340 -2934 327576
rect -2698 327340 -2614 327576
rect -2378 327340 -2346 327576
rect -2966 291896 -2346 327340
rect -2966 291660 -2934 291896
rect -2698 291660 -2614 291896
rect -2378 291660 -2346 291896
rect -2966 291576 -2346 291660
rect -2966 291340 -2934 291576
rect -2698 291340 -2614 291576
rect -2378 291340 -2346 291576
rect -2966 255896 -2346 291340
rect -2966 255660 -2934 255896
rect -2698 255660 -2614 255896
rect -2378 255660 -2346 255896
rect -2966 255576 -2346 255660
rect -2966 255340 -2934 255576
rect -2698 255340 -2614 255576
rect -2378 255340 -2346 255576
rect -2966 219896 -2346 255340
rect -2966 219660 -2934 219896
rect -2698 219660 -2614 219896
rect -2378 219660 -2346 219896
rect -2966 219576 -2346 219660
rect -2966 219340 -2934 219576
rect -2698 219340 -2614 219576
rect -2378 219340 -2346 219576
rect -2966 183896 -2346 219340
rect -2966 183660 -2934 183896
rect -2698 183660 -2614 183896
rect -2378 183660 -2346 183896
rect -2966 183576 -2346 183660
rect -2966 183340 -2934 183576
rect -2698 183340 -2614 183576
rect -2378 183340 -2346 183576
rect -2966 147896 -2346 183340
rect -2966 147660 -2934 147896
rect -2698 147660 -2614 147896
rect -2378 147660 -2346 147896
rect -2966 147576 -2346 147660
rect -2966 147340 -2934 147576
rect -2698 147340 -2614 147576
rect -2378 147340 -2346 147576
rect -2966 111896 -2346 147340
rect -2966 111660 -2934 111896
rect -2698 111660 -2614 111896
rect -2378 111660 -2346 111896
rect -2966 111576 -2346 111660
rect -2966 111340 -2934 111576
rect -2698 111340 -2614 111576
rect -2378 111340 -2346 111576
rect -2966 75896 -2346 111340
rect -2966 75660 -2934 75896
rect -2698 75660 -2614 75896
rect -2378 75660 -2346 75896
rect -2966 75576 -2346 75660
rect -2966 75340 -2934 75576
rect -2698 75340 -2614 75576
rect -2378 75340 -2346 75576
rect -2966 39896 -2346 75340
rect -2966 39660 -2934 39896
rect -2698 39660 -2614 39896
rect -2378 39660 -2346 39896
rect -2966 39576 -2346 39660
rect -2966 39340 -2934 39576
rect -2698 39340 -2614 39576
rect -2378 39340 -2346 39576
rect -2966 3896 -2346 39340
rect -2966 3660 -2934 3896
rect -2698 3660 -2614 3896
rect -2378 3660 -2346 3896
rect -2966 3576 -2346 3660
rect -2966 3340 -2934 3576
rect -2698 3340 -2614 3576
rect -2378 3340 -2346 3576
rect -2966 -1304 -2346 3340
rect -2006 704840 -1386 704872
rect -2006 704604 -1974 704840
rect -1738 704604 -1654 704840
rect -1418 704604 -1386 704840
rect -2006 704520 -1386 704604
rect -2006 704284 -1974 704520
rect -1738 704284 -1654 704520
rect -1418 704284 -1386 704520
rect -2006 686656 -1386 704284
rect -2006 686420 -1974 686656
rect -1738 686420 -1654 686656
rect -1418 686420 -1386 686656
rect -2006 686336 -1386 686420
rect -2006 686100 -1974 686336
rect -1738 686100 -1654 686336
rect -1418 686100 -1386 686336
rect -2006 650656 -1386 686100
rect -2006 650420 -1974 650656
rect -1738 650420 -1654 650656
rect -1418 650420 -1386 650656
rect -2006 650336 -1386 650420
rect -2006 650100 -1974 650336
rect -1738 650100 -1654 650336
rect -1418 650100 -1386 650336
rect -2006 614656 -1386 650100
rect -2006 614420 -1974 614656
rect -1738 614420 -1654 614656
rect -1418 614420 -1386 614656
rect -2006 614336 -1386 614420
rect -2006 614100 -1974 614336
rect -1738 614100 -1654 614336
rect -1418 614100 -1386 614336
rect -2006 578656 -1386 614100
rect -2006 578420 -1974 578656
rect -1738 578420 -1654 578656
rect -1418 578420 -1386 578656
rect -2006 578336 -1386 578420
rect -2006 578100 -1974 578336
rect -1738 578100 -1654 578336
rect -1418 578100 -1386 578336
rect -2006 542656 -1386 578100
rect -2006 542420 -1974 542656
rect -1738 542420 -1654 542656
rect -1418 542420 -1386 542656
rect -2006 542336 -1386 542420
rect -2006 542100 -1974 542336
rect -1738 542100 -1654 542336
rect -1418 542100 -1386 542336
rect -2006 506656 -1386 542100
rect -2006 506420 -1974 506656
rect -1738 506420 -1654 506656
rect -1418 506420 -1386 506656
rect -2006 506336 -1386 506420
rect -2006 506100 -1974 506336
rect -1738 506100 -1654 506336
rect -1418 506100 -1386 506336
rect -2006 470656 -1386 506100
rect -2006 470420 -1974 470656
rect -1738 470420 -1654 470656
rect -1418 470420 -1386 470656
rect -2006 470336 -1386 470420
rect -2006 470100 -1974 470336
rect -1738 470100 -1654 470336
rect -1418 470100 -1386 470336
rect -2006 434656 -1386 470100
rect -2006 434420 -1974 434656
rect -1738 434420 -1654 434656
rect -1418 434420 -1386 434656
rect -2006 434336 -1386 434420
rect -2006 434100 -1974 434336
rect -1738 434100 -1654 434336
rect -1418 434100 -1386 434336
rect -2006 398656 -1386 434100
rect -2006 398420 -1974 398656
rect -1738 398420 -1654 398656
rect -1418 398420 -1386 398656
rect -2006 398336 -1386 398420
rect -2006 398100 -1974 398336
rect -1738 398100 -1654 398336
rect -1418 398100 -1386 398336
rect -2006 362656 -1386 398100
rect -2006 362420 -1974 362656
rect -1738 362420 -1654 362656
rect -1418 362420 -1386 362656
rect -2006 362336 -1386 362420
rect -2006 362100 -1974 362336
rect -1738 362100 -1654 362336
rect -1418 362100 -1386 362336
rect -2006 326656 -1386 362100
rect -2006 326420 -1974 326656
rect -1738 326420 -1654 326656
rect -1418 326420 -1386 326656
rect -2006 326336 -1386 326420
rect -2006 326100 -1974 326336
rect -1738 326100 -1654 326336
rect -1418 326100 -1386 326336
rect -2006 290656 -1386 326100
rect -2006 290420 -1974 290656
rect -1738 290420 -1654 290656
rect -1418 290420 -1386 290656
rect -2006 290336 -1386 290420
rect -2006 290100 -1974 290336
rect -1738 290100 -1654 290336
rect -1418 290100 -1386 290336
rect -2006 254656 -1386 290100
rect -2006 254420 -1974 254656
rect -1738 254420 -1654 254656
rect -1418 254420 -1386 254656
rect -2006 254336 -1386 254420
rect -2006 254100 -1974 254336
rect -1738 254100 -1654 254336
rect -1418 254100 -1386 254336
rect -2006 218656 -1386 254100
rect -2006 218420 -1974 218656
rect -1738 218420 -1654 218656
rect -1418 218420 -1386 218656
rect -2006 218336 -1386 218420
rect -2006 218100 -1974 218336
rect -1738 218100 -1654 218336
rect -1418 218100 -1386 218336
rect -2006 182656 -1386 218100
rect -2006 182420 -1974 182656
rect -1738 182420 -1654 182656
rect -1418 182420 -1386 182656
rect -2006 182336 -1386 182420
rect -2006 182100 -1974 182336
rect -1738 182100 -1654 182336
rect -1418 182100 -1386 182336
rect -2006 146656 -1386 182100
rect -2006 146420 -1974 146656
rect -1738 146420 -1654 146656
rect -1418 146420 -1386 146656
rect -2006 146336 -1386 146420
rect -2006 146100 -1974 146336
rect -1738 146100 -1654 146336
rect -1418 146100 -1386 146336
rect -2006 110656 -1386 146100
rect -2006 110420 -1974 110656
rect -1738 110420 -1654 110656
rect -1418 110420 -1386 110656
rect -2006 110336 -1386 110420
rect -2006 110100 -1974 110336
rect -1738 110100 -1654 110336
rect -1418 110100 -1386 110336
rect -2006 74656 -1386 110100
rect -2006 74420 -1974 74656
rect -1738 74420 -1654 74656
rect -1418 74420 -1386 74656
rect -2006 74336 -1386 74420
rect -2006 74100 -1974 74336
rect -1738 74100 -1654 74336
rect -1418 74100 -1386 74336
rect -2006 38656 -1386 74100
rect -2006 38420 -1974 38656
rect -1738 38420 -1654 38656
rect -1418 38420 -1386 38656
rect -2006 38336 -1386 38420
rect -2006 38100 -1974 38336
rect -1738 38100 -1654 38336
rect -1418 38100 -1386 38336
rect -2006 2656 -1386 38100
rect -2006 2420 -1974 2656
rect -1738 2420 -1654 2656
rect -1418 2420 -1386 2656
rect -2006 2336 -1386 2420
rect -2006 2100 -1974 2336
rect -1738 2100 -1654 2336
rect -1418 2100 -1386 2336
rect -2006 -344 -1386 2100
rect -2006 -580 -1974 -344
rect -1738 -580 -1654 -344
rect -1418 -580 -1386 -344
rect -2006 -664 -1386 -580
rect -2006 -900 -1974 -664
rect -1738 -900 -1654 -664
rect -1418 -900 -1386 -664
rect -2006 -932 -1386 -900
rect 994 704840 1614 711592
rect 994 704604 1026 704840
rect 1262 704604 1346 704840
rect 1582 704604 1614 704840
rect 994 704520 1614 704604
rect 994 704284 1026 704520
rect 1262 704284 1346 704520
rect 1582 704284 1614 704520
rect 994 686656 1614 704284
rect 994 686420 1026 686656
rect 1262 686420 1346 686656
rect 1582 686420 1614 686656
rect 994 686336 1614 686420
rect 994 686100 1026 686336
rect 1262 686100 1346 686336
rect 1582 686100 1614 686336
rect 994 650656 1614 686100
rect 994 650420 1026 650656
rect 1262 650420 1346 650656
rect 1582 650420 1614 650656
rect 994 650336 1614 650420
rect 994 650100 1026 650336
rect 1262 650100 1346 650336
rect 1582 650100 1614 650336
rect 994 614656 1614 650100
rect 994 614420 1026 614656
rect 1262 614420 1346 614656
rect 1582 614420 1614 614656
rect 994 614336 1614 614420
rect 994 614100 1026 614336
rect 1262 614100 1346 614336
rect 1582 614100 1614 614336
rect 994 578656 1614 614100
rect 994 578420 1026 578656
rect 1262 578420 1346 578656
rect 1582 578420 1614 578656
rect 994 578336 1614 578420
rect 994 578100 1026 578336
rect 1262 578100 1346 578336
rect 1582 578100 1614 578336
rect 994 542656 1614 578100
rect 994 542420 1026 542656
rect 1262 542420 1346 542656
rect 1582 542420 1614 542656
rect 994 542336 1614 542420
rect 994 542100 1026 542336
rect 1262 542100 1346 542336
rect 1582 542100 1614 542336
rect 994 506656 1614 542100
rect 994 506420 1026 506656
rect 1262 506420 1346 506656
rect 1582 506420 1614 506656
rect 994 506336 1614 506420
rect 994 506100 1026 506336
rect 1262 506100 1346 506336
rect 1582 506100 1614 506336
rect 994 470656 1614 506100
rect 994 470420 1026 470656
rect 1262 470420 1346 470656
rect 1582 470420 1614 470656
rect 994 470336 1614 470420
rect 994 470100 1026 470336
rect 1262 470100 1346 470336
rect 1582 470100 1614 470336
rect 994 434656 1614 470100
rect 994 434420 1026 434656
rect 1262 434420 1346 434656
rect 1582 434420 1614 434656
rect 994 434336 1614 434420
rect 994 434100 1026 434336
rect 1262 434100 1346 434336
rect 1582 434100 1614 434336
rect 994 398656 1614 434100
rect 994 398420 1026 398656
rect 1262 398420 1346 398656
rect 1582 398420 1614 398656
rect 994 398336 1614 398420
rect 994 398100 1026 398336
rect 1262 398100 1346 398336
rect 1582 398100 1614 398336
rect 994 362656 1614 398100
rect 994 362420 1026 362656
rect 1262 362420 1346 362656
rect 1582 362420 1614 362656
rect 994 362336 1614 362420
rect 994 362100 1026 362336
rect 1262 362100 1346 362336
rect 1582 362100 1614 362336
rect 994 326656 1614 362100
rect 994 326420 1026 326656
rect 1262 326420 1346 326656
rect 1582 326420 1614 326656
rect 994 326336 1614 326420
rect 994 326100 1026 326336
rect 1262 326100 1346 326336
rect 1582 326100 1614 326336
rect 994 290656 1614 326100
rect 994 290420 1026 290656
rect 1262 290420 1346 290656
rect 1582 290420 1614 290656
rect 994 290336 1614 290420
rect 994 290100 1026 290336
rect 1262 290100 1346 290336
rect 1582 290100 1614 290336
rect 994 254656 1614 290100
rect 994 254420 1026 254656
rect 1262 254420 1346 254656
rect 1582 254420 1614 254656
rect 994 254336 1614 254420
rect 994 254100 1026 254336
rect 1262 254100 1346 254336
rect 1582 254100 1614 254336
rect 994 218656 1614 254100
rect 994 218420 1026 218656
rect 1262 218420 1346 218656
rect 1582 218420 1614 218656
rect 994 218336 1614 218420
rect 994 218100 1026 218336
rect 1262 218100 1346 218336
rect 1582 218100 1614 218336
rect 994 182656 1614 218100
rect 994 182420 1026 182656
rect 1262 182420 1346 182656
rect 1582 182420 1614 182656
rect 994 182336 1614 182420
rect 994 182100 1026 182336
rect 1262 182100 1346 182336
rect 1582 182100 1614 182336
rect 994 146656 1614 182100
rect 994 146420 1026 146656
rect 1262 146420 1346 146656
rect 1582 146420 1614 146656
rect 994 146336 1614 146420
rect 994 146100 1026 146336
rect 1262 146100 1346 146336
rect 1582 146100 1614 146336
rect 994 110656 1614 146100
rect 994 110420 1026 110656
rect 1262 110420 1346 110656
rect 1582 110420 1614 110656
rect 994 110336 1614 110420
rect 994 110100 1026 110336
rect 1262 110100 1346 110336
rect 1582 110100 1614 110336
rect 994 74656 1614 110100
rect 994 74420 1026 74656
rect 1262 74420 1346 74656
rect 1582 74420 1614 74656
rect 994 74336 1614 74420
rect 994 74100 1026 74336
rect 1262 74100 1346 74336
rect 1582 74100 1614 74336
rect 994 38656 1614 74100
rect 994 38420 1026 38656
rect 1262 38420 1346 38656
rect 1582 38420 1614 38656
rect 994 38336 1614 38420
rect 994 38100 1026 38336
rect 1262 38100 1346 38336
rect 1582 38100 1614 38336
rect 994 2656 1614 38100
rect 994 2420 1026 2656
rect 1262 2420 1346 2656
rect 1582 2420 1614 2656
rect 994 2336 1614 2420
rect 994 2100 1026 2336
rect 1262 2100 1346 2336
rect 1582 2100 1614 2336
rect 994 -344 1614 2100
rect 994 -580 1026 -344
rect 1262 -580 1346 -344
rect 1582 -580 1614 -344
rect 994 -664 1614 -580
rect 994 -900 1026 -664
rect 1262 -900 1346 -664
rect 1582 -900 1614 -664
rect -2966 -1540 -2934 -1304
rect -2698 -1540 -2614 -1304
rect -2378 -1540 -2346 -1304
rect -2966 -1624 -2346 -1540
rect -2966 -1860 -2934 -1624
rect -2698 -1860 -2614 -1624
rect -2378 -1860 -2346 -1624
rect -2966 -1892 -2346 -1860
rect -3926 -2500 -3894 -2264
rect -3658 -2500 -3574 -2264
rect -3338 -2500 -3306 -2264
rect -3926 -2584 -3306 -2500
rect -3926 -2820 -3894 -2584
rect -3658 -2820 -3574 -2584
rect -3338 -2820 -3306 -2584
rect -3926 -2852 -3306 -2820
rect -4886 -3460 -4854 -3224
rect -4618 -3460 -4534 -3224
rect -4298 -3460 -4266 -3224
rect -4886 -3544 -4266 -3460
rect -4886 -3780 -4854 -3544
rect -4618 -3780 -4534 -3544
rect -4298 -3780 -4266 -3544
rect -4886 -3812 -4266 -3780
rect -5846 -4420 -5814 -4184
rect -5578 -4420 -5494 -4184
rect -5258 -4420 -5226 -4184
rect -5846 -4504 -5226 -4420
rect -5846 -4740 -5814 -4504
rect -5578 -4740 -5494 -4504
rect -5258 -4740 -5226 -4504
rect -5846 -4772 -5226 -4740
rect -6806 -5380 -6774 -5144
rect -6538 -5380 -6454 -5144
rect -6218 -5380 -6186 -5144
rect -6806 -5464 -6186 -5380
rect -6806 -5700 -6774 -5464
rect -6538 -5700 -6454 -5464
rect -6218 -5700 -6186 -5464
rect -6806 -5732 -6186 -5700
rect -7766 -6340 -7734 -6104
rect -7498 -6340 -7414 -6104
rect -7178 -6340 -7146 -6104
rect -7766 -6424 -7146 -6340
rect -7766 -6660 -7734 -6424
rect -7498 -6660 -7414 -6424
rect -7178 -6660 -7146 -6424
rect -7766 -6692 -7146 -6660
rect -8726 -7300 -8694 -7064
rect -8458 -7300 -8374 -7064
rect -8138 -7300 -8106 -7064
rect -8726 -7384 -8106 -7300
rect -8726 -7620 -8694 -7384
rect -8458 -7620 -8374 -7384
rect -8138 -7620 -8106 -7384
rect -8726 -7652 -8106 -7620
rect 994 -7652 1614 -900
rect 2234 705800 2854 711592
rect 2234 705564 2266 705800
rect 2502 705564 2586 705800
rect 2822 705564 2854 705800
rect 2234 705480 2854 705564
rect 2234 705244 2266 705480
rect 2502 705244 2586 705480
rect 2822 705244 2854 705480
rect 2234 687896 2854 705244
rect 2234 687660 2266 687896
rect 2502 687660 2586 687896
rect 2822 687660 2854 687896
rect 2234 687576 2854 687660
rect 2234 687340 2266 687576
rect 2502 687340 2586 687576
rect 2822 687340 2854 687576
rect 2234 651896 2854 687340
rect 2234 651660 2266 651896
rect 2502 651660 2586 651896
rect 2822 651660 2854 651896
rect 2234 651576 2854 651660
rect 2234 651340 2266 651576
rect 2502 651340 2586 651576
rect 2822 651340 2854 651576
rect 2234 615896 2854 651340
rect 2234 615660 2266 615896
rect 2502 615660 2586 615896
rect 2822 615660 2854 615896
rect 2234 615576 2854 615660
rect 2234 615340 2266 615576
rect 2502 615340 2586 615576
rect 2822 615340 2854 615576
rect 2234 579896 2854 615340
rect 2234 579660 2266 579896
rect 2502 579660 2586 579896
rect 2822 579660 2854 579896
rect 2234 579576 2854 579660
rect 2234 579340 2266 579576
rect 2502 579340 2586 579576
rect 2822 579340 2854 579576
rect 2234 543896 2854 579340
rect 2234 543660 2266 543896
rect 2502 543660 2586 543896
rect 2822 543660 2854 543896
rect 2234 543576 2854 543660
rect 2234 543340 2266 543576
rect 2502 543340 2586 543576
rect 2822 543340 2854 543576
rect 2234 507896 2854 543340
rect 2234 507660 2266 507896
rect 2502 507660 2586 507896
rect 2822 507660 2854 507896
rect 2234 507576 2854 507660
rect 2234 507340 2266 507576
rect 2502 507340 2586 507576
rect 2822 507340 2854 507576
rect 2234 471896 2854 507340
rect 2234 471660 2266 471896
rect 2502 471660 2586 471896
rect 2822 471660 2854 471896
rect 2234 471576 2854 471660
rect 2234 471340 2266 471576
rect 2502 471340 2586 471576
rect 2822 471340 2854 471576
rect 2234 435896 2854 471340
rect 2234 435660 2266 435896
rect 2502 435660 2586 435896
rect 2822 435660 2854 435896
rect 2234 435576 2854 435660
rect 2234 435340 2266 435576
rect 2502 435340 2586 435576
rect 2822 435340 2854 435576
rect 2234 399896 2854 435340
rect 2234 399660 2266 399896
rect 2502 399660 2586 399896
rect 2822 399660 2854 399896
rect 2234 399576 2854 399660
rect 2234 399340 2266 399576
rect 2502 399340 2586 399576
rect 2822 399340 2854 399576
rect 2234 363896 2854 399340
rect 2234 363660 2266 363896
rect 2502 363660 2586 363896
rect 2822 363660 2854 363896
rect 2234 363576 2854 363660
rect 2234 363340 2266 363576
rect 2502 363340 2586 363576
rect 2822 363340 2854 363576
rect 2234 327896 2854 363340
rect 2234 327660 2266 327896
rect 2502 327660 2586 327896
rect 2822 327660 2854 327896
rect 2234 327576 2854 327660
rect 2234 327340 2266 327576
rect 2502 327340 2586 327576
rect 2822 327340 2854 327576
rect 2234 291896 2854 327340
rect 2234 291660 2266 291896
rect 2502 291660 2586 291896
rect 2822 291660 2854 291896
rect 2234 291576 2854 291660
rect 2234 291340 2266 291576
rect 2502 291340 2586 291576
rect 2822 291340 2854 291576
rect 2234 255896 2854 291340
rect 2234 255660 2266 255896
rect 2502 255660 2586 255896
rect 2822 255660 2854 255896
rect 2234 255576 2854 255660
rect 2234 255340 2266 255576
rect 2502 255340 2586 255576
rect 2822 255340 2854 255576
rect 2234 219896 2854 255340
rect 2234 219660 2266 219896
rect 2502 219660 2586 219896
rect 2822 219660 2854 219896
rect 2234 219576 2854 219660
rect 2234 219340 2266 219576
rect 2502 219340 2586 219576
rect 2822 219340 2854 219576
rect 2234 183896 2854 219340
rect 2234 183660 2266 183896
rect 2502 183660 2586 183896
rect 2822 183660 2854 183896
rect 2234 183576 2854 183660
rect 2234 183340 2266 183576
rect 2502 183340 2586 183576
rect 2822 183340 2854 183576
rect 2234 147896 2854 183340
rect 2234 147660 2266 147896
rect 2502 147660 2586 147896
rect 2822 147660 2854 147896
rect 2234 147576 2854 147660
rect 2234 147340 2266 147576
rect 2502 147340 2586 147576
rect 2822 147340 2854 147576
rect 2234 111896 2854 147340
rect 2234 111660 2266 111896
rect 2502 111660 2586 111896
rect 2822 111660 2854 111896
rect 2234 111576 2854 111660
rect 2234 111340 2266 111576
rect 2502 111340 2586 111576
rect 2822 111340 2854 111576
rect 2234 75896 2854 111340
rect 2234 75660 2266 75896
rect 2502 75660 2586 75896
rect 2822 75660 2854 75896
rect 2234 75576 2854 75660
rect 2234 75340 2266 75576
rect 2502 75340 2586 75576
rect 2822 75340 2854 75576
rect 2234 39896 2854 75340
rect 2234 39660 2266 39896
rect 2502 39660 2586 39896
rect 2822 39660 2854 39896
rect 2234 39576 2854 39660
rect 2234 39340 2266 39576
rect 2502 39340 2586 39576
rect 2822 39340 2854 39576
rect 2234 3896 2854 39340
rect 2234 3660 2266 3896
rect 2502 3660 2586 3896
rect 2822 3660 2854 3896
rect 2234 3576 2854 3660
rect 2234 3340 2266 3576
rect 2502 3340 2586 3576
rect 2822 3340 2854 3576
rect 2234 -1304 2854 3340
rect 2234 -1540 2266 -1304
rect 2502 -1540 2586 -1304
rect 2822 -1540 2854 -1304
rect 2234 -1624 2854 -1540
rect 2234 -1860 2266 -1624
rect 2502 -1860 2586 -1624
rect 2822 -1860 2854 -1624
rect 2234 -7652 2854 -1860
rect 3474 706760 4094 711592
rect 3474 706524 3506 706760
rect 3742 706524 3826 706760
rect 4062 706524 4094 706760
rect 3474 706440 4094 706524
rect 3474 706204 3506 706440
rect 3742 706204 3826 706440
rect 4062 706204 4094 706440
rect 3474 689136 4094 706204
rect 3474 688900 3506 689136
rect 3742 688900 3826 689136
rect 4062 688900 4094 689136
rect 3474 688816 4094 688900
rect 3474 688580 3506 688816
rect 3742 688580 3826 688816
rect 4062 688580 4094 688816
rect 3474 653136 4094 688580
rect 3474 652900 3506 653136
rect 3742 652900 3826 653136
rect 4062 652900 4094 653136
rect 3474 652816 4094 652900
rect 3474 652580 3506 652816
rect 3742 652580 3826 652816
rect 4062 652580 4094 652816
rect 3474 617136 4094 652580
rect 3474 616900 3506 617136
rect 3742 616900 3826 617136
rect 4062 616900 4094 617136
rect 3474 616816 4094 616900
rect 3474 616580 3506 616816
rect 3742 616580 3826 616816
rect 4062 616580 4094 616816
rect 3474 581136 4094 616580
rect 3474 580900 3506 581136
rect 3742 580900 3826 581136
rect 4062 580900 4094 581136
rect 3474 580816 4094 580900
rect 3474 580580 3506 580816
rect 3742 580580 3826 580816
rect 4062 580580 4094 580816
rect 3474 545136 4094 580580
rect 3474 544900 3506 545136
rect 3742 544900 3826 545136
rect 4062 544900 4094 545136
rect 3474 544816 4094 544900
rect 3474 544580 3506 544816
rect 3742 544580 3826 544816
rect 4062 544580 4094 544816
rect 3474 509136 4094 544580
rect 3474 508900 3506 509136
rect 3742 508900 3826 509136
rect 4062 508900 4094 509136
rect 3474 508816 4094 508900
rect 3474 508580 3506 508816
rect 3742 508580 3826 508816
rect 4062 508580 4094 508816
rect 3474 473136 4094 508580
rect 3474 472900 3506 473136
rect 3742 472900 3826 473136
rect 4062 472900 4094 473136
rect 3474 472816 4094 472900
rect 3474 472580 3506 472816
rect 3742 472580 3826 472816
rect 4062 472580 4094 472816
rect 3474 437136 4094 472580
rect 3474 436900 3506 437136
rect 3742 436900 3826 437136
rect 4062 436900 4094 437136
rect 3474 436816 4094 436900
rect 3474 436580 3506 436816
rect 3742 436580 3826 436816
rect 4062 436580 4094 436816
rect 3474 401136 4094 436580
rect 3474 400900 3506 401136
rect 3742 400900 3826 401136
rect 4062 400900 4094 401136
rect 3474 400816 4094 400900
rect 3474 400580 3506 400816
rect 3742 400580 3826 400816
rect 4062 400580 4094 400816
rect 3474 365136 4094 400580
rect 3474 364900 3506 365136
rect 3742 364900 3826 365136
rect 4062 364900 4094 365136
rect 3474 364816 4094 364900
rect 3474 364580 3506 364816
rect 3742 364580 3826 364816
rect 4062 364580 4094 364816
rect 3474 329136 4094 364580
rect 3474 328900 3506 329136
rect 3742 328900 3826 329136
rect 4062 328900 4094 329136
rect 3474 328816 4094 328900
rect 3474 328580 3506 328816
rect 3742 328580 3826 328816
rect 4062 328580 4094 328816
rect 3474 293136 4094 328580
rect 3474 292900 3506 293136
rect 3742 292900 3826 293136
rect 4062 292900 4094 293136
rect 3474 292816 4094 292900
rect 3474 292580 3506 292816
rect 3742 292580 3826 292816
rect 4062 292580 4094 292816
rect 3474 257136 4094 292580
rect 3474 256900 3506 257136
rect 3742 256900 3826 257136
rect 4062 256900 4094 257136
rect 3474 256816 4094 256900
rect 3474 256580 3506 256816
rect 3742 256580 3826 256816
rect 4062 256580 4094 256816
rect 3474 221136 4094 256580
rect 3474 220900 3506 221136
rect 3742 220900 3826 221136
rect 4062 220900 4094 221136
rect 3474 220816 4094 220900
rect 3474 220580 3506 220816
rect 3742 220580 3826 220816
rect 4062 220580 4094 220816
rect 3474 185136 4094 220580
rect 3474 184900 3506 185136
rect 3742 184900 3826 185136
rect 4062 184900 4094 185136
rect 3474 184816 4094 184900
rect 3474 184580 3506 184816
rect 3742 184580 3826 184816
rect 4062 184580 4094 184816
rect 3474 149136 4094 184580
rect 3474 148900 3506 149136
rect 3742 148900 3826 149136
rect 4062 148900 4094 149136
rect 3474 148816 4094 148900
rect 3474 148580 3506 148816
rect 3742 148580 3826 148816
rect 4062 148580 4094 148816
rect 3474 113136 4094 148580
rect 3474 112900 3506 113136
rect 3742 112900 3826 113136
rect 4062 112900 4094 113136
rect 3474 112816 4094 112900
rect 3474 112580 3506 112816
rect 3742 112580 3826 112816
rect 4062 112580 4094 112816
rect 3474 77136 4094 112580
rect 3474 76900 3506 77136
rect 3742 76900 3826 77136
rect 4062 76900 4094 77136
rect 3474 76816 4094 76900
rect 3474 76580 3506 76816
rect 3742 76580 3826 76816
rect 4062 76580 4094 76816
rect 3474 41136 4094 76580
rect 3474 40900 3506 41136
rect 3742 40900 3826 41136
rect 4062 40900 4094 41136
rect 3474 40816 4094 40900
rect 3474 40580 3506 40816
rect 3742 40580 3826 40816
rect 4062 40580 4094 40816
rect 3474 5136 4094 40580
rect 3474 4900 3506 5136
rect 3742 4900 3826 5136
rect 4062 4900 4094 5136
rect 3474 4816 4094 4900
rect 3474 4580 3506 4816
rect 3742 4580 3826 4816
rect 4062 4580 4094 4816
rect 3474 -2264 4094 4580
rect 3474 -2500 3506 -2264
rect 3742 -2500 3826 -2264
rect 4062 -2500 4094 -2264
rect 3474 -2584 4094 -2500
rect 3474 -2820 3506 -2584
rect 3742 -2820 3826 -2584
rect 4062 -2820 4094 -2584
rect 3474 -7652 4094 -2820
rect 4714 707720 5334 711592
rect 4714 707484 4746 707720
rect 4982 707484 5066 707720
rect 5302 707484 5334 707720
rect 4714 707400 5334 707484
rect 4714 707164 4746 707400
rect 4982 707164 5066 707400
rect 5302 707164 5334 707400
rect 4714 690376 5334 707164
rect 4714 690140 4746 690376
rect 4982 690140 5066 690376
rect 5302 690140 5334 690376
rect 4714 690056 5334 690140
rect 4714 689820 4746 690056
rect 4982 689820 5066 690056
rect 5302 689820 5334 690056
rect 4714 654376 5334 689820
rect 4714 654140 4746 654376
rect 4982 654140 5066 654376
rect 5302 654140 5334 654376
rect 4714 654056 5334 654140
rect 4714 653820 4746 654056
rect 4982 653820 5066 654056
rect 5302 653820 5334 654056
rect 4714 618376 5334 653820
rect 4714 618140 4746 618376
rect 4982 618140 5066 618376
rect 5302 618140 5334 618376
rect 4714 618056 5334 618140
rect 4714 617820 4746 618056
rect 4982 617820 5066 618056
rect 5302 617820 5334 618056
rect 4714 582376 5334 617820
rect 4714 582140 4746 582376
rect 4982 582140 5066 582376
rect 5302 582140 5334 582376
rect 4714 582056 5334 582140
rect 4714 581820 4746 582056
rect 4982 581820 5066 582056
rect 5302 581820 5334 582056
rect 4714 546376 5334 581820
rect 4714 546140 4746 546376
rect 4982 546140 5066 546376
rect 5302 546140 5334 546376
rect 4714 546056 5334 546140
rect 4714 545820 4746 546056
rect 4982 545820 5066 546056
rect 5302 545820 5334 546056
rect 4714 510376 5334 545820
rect 4714 510140 4746 510376
rect 4982 510140 5066 510376
rect 5302 510140 5334 510376
rect 4714 510056 5334 510140
rect 4714 509820 4746 510056
rect 4982 509820 5066 510056
rect 5302 509820 5334 510056
rect 4714 474376 5334 509820
rect 4714 474140 4746 474376
rect 4982 474140 5066 474376
rect 5302 474140 5334 474376
rect 4714 474056 5334 474140
rect 4714 473820 4746 474056
rect 4982 473820 5066 474056
rect 5302 473820 5334 474056
rect 4714 438376 5334 473820
rect 4714 438140 4746 438376
rect 4982 438140 5066 438376
rect 5302 438140 5334 438376
rect 4714 438056 5334 438140
rect 4714 437820 4746 438056
rect 4982 437820 5066 438056
rect 5302 437820 5334 438056
rect 4714 402376 5334 437820
rect 4714 402140 4746 402376
rect 4982 402140 5066 402376
rect 5302 402140 5334 402376
rect 4714 402056 5334 402140
rect 4714 401820 4746 402056
rect 4982 401820 5066 402056
rect 5302 401820 5334 402056
rect 4714 366376 5334 401820
rect 4714 366140 4746 366376
rect 4982 366140 5066 366376
rect 5302 366140 5334 366376
rect 4714 366056 5334 366140
rect 4714 365820 4746 366056
rect 4982 365820 5066 366056
rect 5302 365820 5334 366056
rect 4714 330376 5334 365820
rect 4714 330140 4746 330376
rect 4982 330140 5066 330376
rect 5302 330140 5334 330376
rect 4714 330056 5334 330140
rect 4714 329820 4746 330056
rect 4982 329820 5066 330056
rect 5302 329820 5334 330056
rect 4714 294376 5334 329820
rect 4714 294140 4746 294376
rect 4982 294140 5066 294376
rect 5302 294140 5334 294376
rect 4714 294056 5334 294140
rect 4714 293820 4746 294056
rect 4982 293820 5066 294056
rect 5302 293820 5334 294056
rect 4714 258376 5334 293820
rect 4714 258140 4746 258376
rect 4982 258140 5066 258376
rect 5302 258140 5334 258376
rect 4714 258056 5334 258140
rect 4714 257820 4746 258056
rect 4982 257820 5066 258056
rect 5302 257820 5334 258056
rect 4714 222376 5334 257820
rect 4714 222140 4746 222376
rect 4982 222140 5066 222376
rect 5302 222140 5334 222376
rect 4714 222056 5334 222140
rect 4714 221820 4746 222056
rect 4982 221820 5066 222056
rect 5302 221820 5334 222056
rect 4714 186376 5334 221820
rect 4714 186140 4746 186376
rect 4982 186140 5066 186376
rect 5302 186140 5334 186376
rect 4714 186056 5334 186140
rect 4714 185820 4746 186056
rect 4982 185820 5066 186056
rect 5302 185820 5334 186056
rect 4714 150376 5334 185820
rect 4714 150140 4746 150376
rect 4982 150140 5066 150376
rect 5302 150140 5334 150376
rect 4714 150056 5334 150140
rect 4714 149820 4746 150056
rect 4982 149820 5066 150056
rect 5302 149820 5334 150056
rect 4714 114376 5334 149820
rect 4714 114140 4746 114376
rect 4982 114140 5066 114376
rect 5302 114140 5334 114376
rect 4714 114056 5334 114140
rect 4714 113820 4746 114056
rect 4982 113820 5066 114056
rect 5302 113820 5334 114056
rect 4714 78376 5334 113820
rect 4714 78140 4746 78376
rect 4982 78140 5066 78376
rect 5302 78140 5334 78376
rect 4714 78056 5334 78140
rect 4714 77820 4746 78056
rect 4982 77820 5066 78056
rect 5302 77820 5334 78056
rect 4714 42376 5334 77820
rect 4714 42140 4746 42376
rect 4982 42140 5066 42376
rect 5302 42140 5334 42376
rect 4714 42056 5334 42140
rect 4714 41820 4746 42056
rect 4982 41820 5066 42056
rect 5302 41820 5334 42056
rect 4714 6376 5334 41820
rect 4714 6140 4746 6376
rect 4982 6140 5066 6376
rect 5302 6140 5334 6376
rect 4714 6056 5334 6140
rect 4714 5820 4746 6056
rect 4982 5820 5066 6056
rect 5302 5820 5334 6056
rect 4714 -3224 5334 5820
rect 4714 -3460 4746 -3224
rect 4982 -3460 5066 -3224
rect 5302 -3460 5334 -3224
rect 4714 -3544 5334 -3460
rect 4714 -3780 4746 -3544
rect 4982 -3780 5066 -3544
rect 5302 -3780 5334 -3544
rect 4714 -7652 5334 -3780
rect 5954 708680 6574 711592
rect 5954 708444 5986 708680
rect 6222 708444 6306 708680
rect 6542 708444 6574 708680
rect 5954 708360 6574 708444
rect 5954 708124 5986 708360
rect 6222 708124 6306 708360
rect 6542 708124 6574 708360
rect 5954 691616 6574 708124
rect 5954 691380 5986 691616
rect 6222 691380 6306 691616
rect 6542 691380 6574 691616
rect 5954 691296 6574 691380
rect 5954 691060 5986 691296
rect 6222 691060 6306 691296
rect 6542 691060 6574 691296
rect 5954 655616 6574 691060
rect 5954 655380 5986 655616
rect 6222 655380 6306 655616
rect 6542 655380 6574 655616
rect 5954 655296 6574 655380
rect 5954 655060 5986 655296
rect 6222 655060 6306 655296
rect 6542 655060 6574 655296
rect 5954 619616 6574 655060
rect 5954 619380 5986 619616
rect 6222 619380 6306 619616
rect 6542 619380 6574 619616
rect 5954 619296 6574 619380
rect 5954 619060 5986 619296
rect 6222 619060 6306 619296
rect 6542 619060 6574 619296
rect 5954 583616 6574 619060
rect 5954 583380 5986 583616
rect 6222 583380 6306 583616
rect 6542 583380 6574 583616
rect 5954 583296 6574 583380
rect 5954 583060 5986 583296
rect 6222 583060 6306 583296
rect 6542 583060 6574 583296
rect 5954 547616 6574 583060
rect 5954 547380 5986 547616
rect 6222 547380 6306 547616
rect 6542 547380 6574 547616
rect 5954 547296 6574 547380
rect 5954 547060 5986 547296
rect 6222 547060 6306 547296
rect 6542 547060 6574 547296
rect 5954 511616 6574 547060
rect 5954 511380 5986 511616
rect 6222 511380 6306 511616
rect 6542 511380 6574 511616
rect 5954 511296 6574 511380
rect 5954 511060 5986 511296
rect 6222 511060 6306 511296
rect 6542 511060 6574 511296
rect 5954 475616 6574 511060
rect 5954 475380 5986 475616
rect 6222 475380 6306 475616
rect 6542 475380 6574 475616
rect 5954 475296 6574 475380
rect 5954 475060 5986 475296
rect 6222 475060 6306 475296
rect 6542 475060 6574 475296
rect 5954 439616 6574 475060
rect 5954 439380 5986 439616
rect 6222 439380 6306 439616
rect 6542 439380 6574 439616
rect 5954 439296 6574 439380
rect 5954 439060 5986 439296
rect 6222 439060 6306 439296
rect 6542 439060 6574 439296
rect 5954 403616 6574 439060
rect 5954 403380 5986 403616
rect 6222 403380 6306 403616
rect 6542 403380 6574 403616
rect 5954 403296 6574 403380
rect 5954 403060 5986 403296
rect 6222 403060 6306 403296
rect 6542 403060 6574 403296
rect 5954 367616 6574 403060
rect 5954 367380 5986 367616
rect 6222 367380 6306 367616
rect 6542 367380 6574 367616
rect 5954 367296 6574 367380
rect 5954 367060 5986 367296
rect 6222 367060 6306 367296
rect 6542 367060 6574 367296
rect 5954 331616 6574 367060
rect 5954 331380 5986 331616
rect 6222 331380 6306 331616
rect 6542 331380 6574 331616
rect 5954 331296 6574 331380
rect 5954 331060 5986 331296
rect 6222 331060 6306 331296
rect 6542 331060 6574 331296
rect 5954 295616 6574 331060
rect 5954 295380 5986 295616
rect 6222 295380 6306 295616
rect 6542 295380 6574 295616
rect 5954 295296 6574 295380
rect 5954 295060 5986 295296
rect 6222 295060 6306 295296
rect 6542 295060 6574 295296
rect 5954 259616 6574 295060
rect 5954 259380 5986 259616
rect 6222 259380 6306 259616
rect 6542 259380 6574 259616
rect 5954 259296 6574 259380
rect 5954 259060 5986 259296
rect 6222 259060 6306 259296
rect 6542 259060 6574 259296
rect 5954 223616 6574 259060
rect 5954 223380 5986 223616
rect 6222 223380 6306 223616
rect 6542 223380 6574 223616
rect 5954 223296 6574 223380
rect 5954 223060 5986 223296
rect 6222 223060 6306 223296
rect 6542 223060 6574 223296
rect 5954 187616 6574 223060
rect 5954 187380 5986 187616
rect 6222 187380 6306 187616
rect 6542 187380 6574 187616
rect 5954 187296 6574 187380
rect 5954 187060 5986 187296
rect 6222 187060 6306 187296
rect 6542 187060 6574 187296
rect 5954 151616 6574 187060
rect 5954 151380 5986 151616
rect 6222 151380 6306 151616
rect 6542 151380 6574 151616
rect 5954 151296 6574 151380
rect 5954 151060 5986 151296
rect 6222 151060 6306 151296
rect 6542 151060 6574 151296
rect 5954 115616 6574 151060
rect 5954 115380 5986 115616
rect 6222 115380 6306 115616
rect 6542 115380 6574 115616
rect 5954 115296 6574 115380
rect 5954 115060 5986 115296
rect 6222 115060 6306 115296
rect 6542 115060 6574 115296
rect 5954 79616 6574 115060
rect 5954 79380 5986 79616
rect 6222 79380 6306 79616
rect 6542 79380 6574 79616
rect 5954 79296 6574 79380
rect 5954 79060 5986 79296
rect 6222 79060 6306 79296
rect 6542 79060 6574 79296
rect 5954 43616 6574 79060
rect 5954 43380 5986 43616
rect 6222 43380 6306 43616
rect 6542 43380 6574 43616
rect 5954 43296 6574 43380
rect 5954 43060 5986 43296
rect 6222 43060 6306 43296
rect 6542 43060 6574 43296
rect 5954 7616 6574 43060
rect 5954 7380 5986 7616
rect 6222 7380 6306 7616
rect 6542 7380 6574 7616
rect 5954 7296 6574 7380
rect 5954 7060 5986 7296
rect 6222 7060 6306 7296
rect 6542 7060 6574 7296
rect 5954 -4184 6574 7060
rect 5954 -4420 5986 -4184
rect 6222 -4420 6306 -4184
rect 6542 -4420 6574 -4184
rect 5954 -4504 6574 -4420
rect 5954 -4740 5986 -4504
rect 6222 -4740 6306 -4504
rect 6542 -4740 6574 -4504
rect 5954 -7652 6574 -4740
rect 7194 709640 7814 711592
rect 7194 709404 7226 709640
rect 7462 709404 7546 709640
rect 7782 709404 7814 709640
rect 7194 709320 7814 709404
rect 7194 709084 7226 709320
rect 7462 709084 7546 709320
rect 7782 709084 7814 709320
rect 7194 692856 7814 709084
rect 7194 692620 7226 692856
rect 7462 692620 7546 692856
rect 7782 692620 7814 692856
rect 7194 692536 7814 692620
rect 7194 692300 7226 692536
rect 7462 692300 7546 692536
rect 7782 692300 7814 692536
rect 7194 656856 7814 692300
rect 7194 656620 7226 656856
rect 7462 656620 7546 656856
rect 7782 656620 7814 656856
rect 7194 656536 7814 656620
rect 7194 656300 7226 656536
rect 7462 656300 7546 656536
rect 7782 656300 7814 656536
rect 7194 620856 7814 656300
rect 7194 620620 7226 620856
rect 7462 620620 7546 620856
rect 7782 620620 7814 620856
rect 7194 620536 7814 620620
rect 7194 620300 7226 620536
rect 7462 620300 7546 620536
rect 7782 620300 7814 620536
rect 7194 584856 7814 620300
rect 7194 584620 7226 584856
rect 7462 584620 7546 584856
rect 7782 584620 7814 584856
rect 7194 584536 7814 584620
rect 7194 584300 7226 584536
rect 7462 584300 7546 584536
rect 7782 584300 7814 584536
rect 7194 548856 7814 584300
rect 7194 548620 7226 548856
rect 7462 548620 7546 548856
rect 7782 548620 7814 548856
rect 7194 548536 7814 548620
rect 7194 548300 7226 548536
rect 7462 548300 7546 548536
rect 7782 548300 7814 548536
rect 7194 512856 7814 548300
rect 7194 512620 7226 512856
rect 7462 512620 7546 512856
rect 7782 512620 7814 512856
rect 7194 512536 7814 512620
rect 7194 512300 7226 512536
rect 7462 512300 7546 512536
rect 7782 512300 7814 512536
rect 7194 476856 7814 512300
rect 7194 476620 7226 476856
rect 7462 476620 7546 476856
rect 7782 476620 7814 476856
rect 7194 476536 7814 476620
rect 7194 476300 7226 476536
rect 7462 476300 7546 476536
rect 7782 476300 7814 476536
rect 7194 440856 7814 476300
rect 7194 440620 7226 440856
rect 7462 440620 7546 440856
rect 7782 440620 7814 440856
rect 7194 440536 7814 440620
rect 7194 440300 7226 440536
rect 7462 440300 7546 440536
rect 7782 440300 7814 440536
rect 7194 404856 7814 440300
rect 7194 404620 7226 404856
rect 7462 404620 7546 404856
rect 7782 404620 7814 404856
rect 7194 404536 7814 404620
rect 7194 404300 7226 404536
rect 7462 404300 7546 404536
rect 7782 404300 7814 404536
rect 7194 368856 7814 404300
rect 7194 368620 7226 368856
rect 7462 368620 7546 368856
rect 7782 368620 7814 368856
rect 7194 368536 7814 368620
rect 7194 368300 7226 368536
rect 7462 368300 7546 368536
rect 7782 368300 7814 368536
rect 7194 332856 7814 368300
rect 7194 332620 7226 332856
rect 7462 332620 7546 332856
rect 7782 332620 7814 332856
rect 7194 332536 7814 332620
rect 7194 332300 7226 332536
rect 7462 332300 7546 332536
rect 7782 332300 7814 332536
rect 7194 296856 7814 332300
rect 7194 296620 7226 296856
rect 7462 296620 7546 296856
rect 7782 296620 7814 296856
rect 7194 296536 7814 296620
rect 7194 296300 7226 296536
rect 7462 296300 7546 296536
rect 7782 296300 7814 296536
rect 7194 260856 7814 296300
rect 7194 260620 7226 260856
rect 7462 260620 7546 260856
rect 7782 260620 7814 260856
rect 7194 260536 7814 260620
rect 7194 260300 7226 260536
rect 7462 260300 7546 260536
rect 7782 260300 7814 260536
rect 7194 224856 7814 260300
rect 7194 224620 7226 224856
rect 7462 224620 7546 224856
rect 7782 224620 7814 224856
rect 7194 224536 7814 224620
rect 7194 224300 7226 224536
rect 7462 224300 7546 224536
rect 7782 224300 7814 224536
rect 7194 188856 7814 224300
rect 7194 188620 7226 188856
rect 7462 188620 7546 188856
rect 7782 188620 7814 188856
rect 7194 188536 7814 188620
rect 7194 188300 7226 188536
rect 7462 188300 7546 188536
rect 7782 188300 7814 188536
rect 7194 152856 7814 188300
rect 7194 152620 7226 152856
rect 7462 152620 7546 152856
rect 7782 152620 7814 152856
rect 7194 152536 7814 152620
rect 7194 152300 7226 152536
rect 7462 152300 7546 152536
rect 7782 152300 7814 152536
rect 7194 116856 7814 152300
rect 7194 116620 7226 116856
rect 7462 116620 7546 116856
rect 7782 116620 7814 116856
rect 7194 116536 7814 116620
rect 7194 116300 7226 116536
rect 7462 116300 7546 116536
rect 7782 116300 7814 116536
rect 7194 80856 7814 116300
rect 7194 80620 7226 80856
rect 7462 80620 7546 80856
rect 7782 80620 7814 80856
rect 7194 80536 7814 80620
rect 7194 80300 7226 80536
rect 7462 80300 7546 80536
rect 7782 80300 7814 80536
rect 7194 44856 7814 80300
rect 7194 44620 7226 44856
rect 7462 44620 7546 44856
rect 7782 44620 7814 44856
rect 7194 44536 7814 44620
rect 7194 44300 7226 44536
rect 7462 44300 7546 44536
rect 7782 44300 7814 44536
rect 7194 8856 7814 44300
rect 7194 8620 7226 8856
rect 7462 8620 7546 8856
rect 7782 8620 7814 8856
rect 7194 8536 7814 8620
rect 7194 8300 7226 8536
rect 7462 8300 7546 8536
rect 7782 8300 7814 8536
rect 7194 -5144 7814 8300
rect 7194 -5380 7226 -5144
rect 7462 -5380 7546 -5144
rect 7782 -5380 7814 -5144
rect 7194 -5464 7814 -5380
rect 7194 -5700 7226 -5464
rect 7462 -5700 7546 -5464
rect 7782 -5700 7814 -5464
rect 7194 -7652 7814 -5700
rect 8434 710600 9054 711592
rect 8434 710364 8466 710600
rect 8702 710364 8786 710600
rect 9022 710364 9054 710600
rect 8434 710280 9054 710364
rect 8434 710044 8466 710280
rect 8702 710044 8786 710280
rect 9022 710044 9054 710280
rect 8434 694096 9054 710044
rect 8434 693860 8466 694096
rect 8702 693860 8786 694096
rect 9022 693860 9054 694096
rect 8434 693776 9054 693860
rect 8434 693540 8466 693776
rect 8702 693540 8786 693776
rect 9022 693540 9054 693776
rect 8434 658096 9054 693540
rect 8434 657860 8466 658096
rect 8702 657860 8786 658096
rect 9022 657860 9054 658096
rect 8434 657776 9054 657860
rect 8434 657540 8466 657776
rect 8702 657540 8786 657776
rect 9022 657540 9054 657776
rect 8434 622096 9054 657540
rect 8434 621860 8466 622096
rect 8702 621860 8786 622096
rect 9022 621860 9054 622096
rect 8434 621776 9054 621860
rect 8434 621540 8466 621776
rect 8702 621540 8786 621776
rect 9022 621540 9054 621776
rect 8434 586096 9054 621540
rect 8434 585860 8466 586096
rect 8702 585860 8786 586096
rect 9022 585860 9054 586096
rect 8434 585776 9054 585860
rect 8434 585540 8466 585776
rect 8702 585540 8786 585776
rect 9022 585540 9054 585776
rect 8434 550096 9054 585540
rect 8434 549860 8466 550096
rect 8702 549860 8786 550096
rect 9022 549860 9054 550096
rect 8434 549776 9054 549860
rect 8434 549540 8466 549776
rect 8702 549540 8786 549776
rect 9022 549540 9054 549776
rect 8434 514096 9054 549540
rect 8434 513860 8466 514096
rect 8702 513860 8786 514096
rect 9022 513860 9054 514096
rect 8434 513776 9054 513860
rect 8434 513540 8466 513776
rect 8702 513540 8786 513776
rect 9022 513540 9054 513776
rect 8434 478096 9054 513540
rect 8434 477860 8466 478096
rect 8702 477860 8786 478096
rect 9022 477860 9054 478096
rect 8434 477776 9054 477860
rect 8434 477540 8466 477776
rect 8702 477540 8786 477776
rect 9022 477540 9054 477776
rect 8434 442096 9054 477540
rect 8434 441860 8466 442096
rect 8702 441860 8786 442096
rect 9022 441860 9054 442096
rect 8434 441776 9054 441860
rect 8434 441540 8466 441776
rect 8702 441540 8786 441776
rect 9022 441540 9054 441776
rect 8434 406096 9054 441540
rect 8434 405860 8466 406096
rect 8702 405860 8786 406096
rect 9022 405860 9054 406096
rect 8434 405776 9054 405860
rect 8434 405540 8466 405776
rect 8702 405540 8786 405776
rect 9022 405540 9054 405776
rect 8434 370096 9054 405540
rect 8434 369860 8466 370096
rect 8702 369860 8786 370096
rect 9022 369860 9054 370096
rect 8434 369776 9054 369860
rect 8434 369540 8466 369776
rect 8702 369540 8786 369776
rect 9022 369540 9054 369776
rect 8434 334096 9054 369540
rect 8434 333860 8466 334096
rect 8702 333860 8786 334096
rect 9022 333860 9054 334096
rect 8434 333776 9054 333860
rect 8434 333540 8466 333776
rect 8702 333540 8786 333776
rect 9022 333540 9054 333776
rect 8434 298096 9054 333540
rect 8434 297860 8466 298096
rect 8702 297860 8786 298096
rect 9022 297860 9054 298096
rect 8434 297776 9054 297860
rect 8434 297540 8466 297776
rect 8702 297540 8786 297776
rect 9022 297540 9054 297776
rect 8434 262096 9054 297540
rect 8434 261860 8466 262096
rect 8702 261860 8786 262096
rect 9022 261860 9054 262096
rect 8434 261776 9054 261860
rect 8434 261540 8466 261776
rect 8702 261540 8786 261776
rect 9022 261540 9054 261776
rect 8434 226096 9054 261540
rect 8434 225860 8466 226096
rect 8702 225860 8786 226096
rect 9022 225860 9054 226096
rect 8434 225776 9054 225860
rect 8434 225540 8466 225776
rect 8702 225540 8786 225776
rect 9022 225540 9054 225776
rect 8434 190096 9054 225540
rect 8434 189860 8466 190096
rect 8702 189860 8786 190096
rect 9022 189860 9054 190096
rect 8434 189776 9054 189860
rect 8434 189540 8466 189776
rect 8702 189540 8786 189776
rect 9022 189540 9054 189776
rect 8434 154096 9054 189540
rect 8434 153860 8466 154096
rect 8702 153860 8786 154096
rect 9022 153860 9054 154096
rect 8434 153776 9054 153860
rect 8434 153540 8466 153776
rect 8702 153540 8786 153776
rect 9022 153540 9054 153776
rect 8434 118096 9054 153540
rect 8434 117860 8466 118096
rect 8702 117860 8786 118096
rect 9022 117860 9054 118096
rect 8434 117776 9054 117860
rect 8434 117540 8466 117776
rect 8702 117540 8786 117776
rect 9022 117540 9054 117776
rect 8434 82096 9054 117540
rect 8434 81860 8466 82096
rect 8702 81860 8786 82096
rect 9022 81860 9054 82096
rect 8434 81776 9054 81860
rect 8434 81540 8466 81776
rect 8702 81540 8786 81776
rect 9022 81540 9054 81776
rect 8434 46096 9054 81540
rect 8434 45860 8466 46096
rect 8702 45860 8786 46096
rect 9022 45860 9054 46096
rect 8434 45776 9054 45860
rect 8434 45540 8466 45776
rect 8702 45540 8786 45776
rect 9022 45540 9054 45776
rect 8434 10096 9054 45540
rect 8434 9860 8466 10096
rect 8702 9860 8786 10096
rect 9022 9860 9054 10096
rect 8434 9776 9054 9860
rect 8434 9540 8466 9776
rect 8702 9540 8786 9776
rect 9022 9540 9054 9776
rect 8434 -6104 9054 9540
rect 8434 -6340 8466 -6104
rect 8702 -6340 8786 -6104
rect 9022 -6340 9054 -6104
rect 8434 -6424 9054 -6340
rect 8434 -6660 8466 -6424
rect 8702 -6660 8786 -6424
rect 9022 -6660 9054 -6424
rect 8434 -7652 9054 -6660
rect 9674 711560 10294 711592
rect 9674 711324 9706 711560
rect 9942 711324 10026 711560
rect 10262 711324 10294 711560
rect 9674 711240 10294 711324
rect 9674 711004 9706 711240
rect 9942 711004 10026 711240
rect 10262 711004 10294 711240
rect 9674 695336 10294 711004
rect 9674 695100 9706 695336
rect 9942 695100 10026 695336
rect 10262 695100 10294 695336
rect 9674 695016 10294 695100
rect 9674 694780 9706 695016
rect 9942 694780 10026 695016
rect 10262 694780 10294 695016
rect 9674 659336 10294 694780
rect 9674 659100 9706 659336
rect 9942 659100 10026 659336
rect 10262 659100 10294 659336
rect 9674 659016 10294 659100
rect 9674 658780 9706 659016
rect 9942 658780 10026 659016
rect 10262 658780 10294 659016
rect 9674 623336 10294 658780
rect 9674 623100 9706 623336
rect 9942 623100 10026 623336
rect 10262 623100 10294 623336
rect 9674 623016 10294 623100
rect 9674 622780 9706 623016
rect 9942 622780 10026 623016
rect 10262 622780 10294 623016
rect 9674 587336 10294 622780
rect 9674 587100 9706 587336
rect 9942 587100 10026 587336
rect 10262 587100 10294 587336
rect 9674 587016 10294 587100
rect 9674 586780 9706 587016
rect 9942 586780 10026 587016
rect 10262 586780 10294 587016
rect 9674 551336 10294 586780
rect 9674 551100 9706 551336
rect 9942 551100 10026 551336
rect 10262 551100 10294 551336
rect 9674 551016 10294 551100
rect 9674 550780 9706 551016
rect 9942 550780 10026 551016
rect 10262 550780 10294 551016
rect 9674 515336 10294 550780
rect 9674 515100 9706 515336
rect 9942 515100 10026 515336
rect 10262 515100 10294 515336
rect 9674 515016 10294 515100
rect 9674 514780 9706 515016
rect 9942 514780 10026 515016
rect 10262 514780 10294 515016
rect 9674 479336 10294 514780
rect 9674 479100 9706 479336
rect 9942 479100 10026 479336
rect 10262 479100 10294 479336
rect 9674 479016 10294 479100
rect 9674 478780 9706 479016
rect 9942 478780 10026 479016
rect 10262 478780 10294 479016
rect 9674 443336 10294 478780
rect 9674 443100 9706 443336
rect 9942 443100 10026 443336
rect 10262 443100 10294 443336
rect 9674 443016 10294 443100
rect 9674 442780 9706 443016
rect 9942 442780 10026 443016
rect 10262 442780 10294 443016
rect 9674 407336 10294 442780
rect 9674 407100 9706 407336
rect 9942 407100 10026 407336
rect 10262 407100 10294 407336
rect 9674 407016 10294 407100
rect 9674 406780 9706 407016
rect 9942 406780 10026 407016
rect 10262 406780 10294 407016
rect 9674 371336 10294 406780
rect 9674 371100 9706 371336
rect 9942 371100 10026 371336
rect 10262 371100 10294 371336
rect 9674 371016 10294 371100
rect 9674 370780 9706 371016
rect 9942 370780 10026 371016
rect 10262 370780 10294 371016
rect 9674 335336 10294 370780
rect 9674 335100 9706 335336
rect 9942 335100 10026 335336
rect 10262 335100 10294 335336
rect 9674 335016 10294 335100
rect 9674 334780 9706 335016
rect 9942 334780 10026 335016
rect 10262 334780 10294 335016
rect 9674 299336 10294 334780
rect 9674 299100 9706 299336
rect 9942 299100 10026 299336
rect 10262 299100 10294 299336
rect 9674 299016 10294 299100
rect 9674 298780 9706 299016
rect 9942 298780 10026 299016
rect 10262 298780 10294 299016
rect 9674 263336 10294 298780
rect 9674 263100 9706 263336
rect 9942 263100 10026 263336
rect 10262 263100 10294 263336
rect 9674 263016 10294 263100
rect 9674 262780 9706 263016
rect 9942 262780 10026 263016
rect 10262 262780 10294 263016
rect 9674 227336 10294 262780
rect 9674 227100 9706 227336
rect 9942 227100 10026 227336
rect 10262 227100 10294 227336
rect 9674 227016 10294 227100
rect 9674 226780 9706 227016
rect 9942 226780 10026 227016
rect 10262 226780 10294 227016
rect 9674 191336 10294 226780
rect 9674 191100 9706 191336
rect 9942 191100 10026 191336
rect 10262 191100 10294 191336
rect 9674 191016 10294 191100
rect 9674 190780 9706 191016
rect 9942 190780 10026 191016
rect 10262 190780 10294 191016
rect 9674 155336 10294 190780
rect 9674 155100 9706 155336
rect 9942 155100 10026 155336
rect 10262 155100 10294 155336
rect 9674 155016 10294 155100
rect 9674 154780 9706 155016
rect 9942 154780 10026 155016
rect 10262 154780 10294 155016
rect 9674 119336 10294 154780
rect 9674 119100 9706 119336
rect 9942 119100 10026 119336
rect 10262 119100 10294 119336
rect 9674 119016 10294 119100
rect 9674 118780 9706 119016
rect 9942 118780 10026 119016
rect 10262 118780 10294 119016
rect 9674 83336 10294 118780
rect 9674 83100 9706 83336
rect 9942 83100 10026 83336
rect 10262 83100 10294 83336
rect 9674 83016 10294 83100
rect 9674 82780 9706 83016
rect 9942 82780 10026 83016
rect 10262 82780 10294 83016
rect 9674 47336 10294 82780
rect 9674 47100 9706 47336
rect 9942 47100 10026 47336
rect 10262 47100 10294 47336
rect 9674 47016 10294 47100
rect 9674 46780 9706 47016
rect 9942 46780 10026 47016
rect 10262 46780 10294 47016
rect 9674 11336 10294 46780
rect 9674 11100 9706 11336
rect 9942 11100 10026 11336
rect 10262 11100 10294 11336
rect 9674 11016 10294 11100
rect 9674 10780 9706 11016
rect 9942 10780 10026 11016
rect 10262 10780 10294 11016
rect 9674 -7064 10294 10780
rect 9674 -7300 9706 -7064
rect 9942 -7300 10026 -7064
rect 10262 -7300 10294 -7064
rect 9674 -7384 10294 -7300
rect 9674 -7620 9706 -7384
rect 9942 -7620 10026 -7384
rect 10262 -7620 10294 -7384
rect 9674 -7652 10294 -7620
rect 36994 704840 37614 711592
rect 36994 704604 37026 704840
rect 37262 704604 37346 704840
rect 37582 704604 37614 704840
rect 36994 704520 37614 704604
rect 36994 704284 37026 704520
rect 37262 704284 37346 704520
rect 37582 704284 37614 704520
rect 36994 686656 37614 704284
rect 36994 686420 37026 686656
rect 37262 686420 37346 686656
rect 37582 686420 37614 686656
rect 36994 686336 37614 686420
rect 36994 686100 37026 686336
rect 37262 686100 37346 686336
rect 37582 686100 37614 686336
rect 36994 650656 37614 686100
rect 36994 650420 37026 650656
rect 37262 650420 37346 650656
rect 37582 650420 37614 650656
rect 36994 650336 37614 650420
rect 36994 650100 37026 650336
rect 37262 650100 37346 650336
rect 37582 650100 37614 650336
rect 36994 614656 37614 650100
rect 36994 614420 37026 614656
rect 37262 614420 37346 614656
rect 37582 614420 37614 614656
rect 36994 614336 37614 614420
rect 36994 614100 37026 614336
rect 37262 614100 37346 614336
rect 37582 614100 37614 614336
rect 36994 578656 37614 614100
rect 36994 578420 37026 578656
rect 37262 578420 37346 578656
rect 37582 578420 37614 578656
rect 36994 578336 37614 578420
rect 36994 578100 37026 578336
rect 37262 578100 37346 578336
rect 37582 578100 37614 578336
rect 36994 542656 37614 578100
rect 36994 542420 37026 542656
rect 37262 542420 37346 542656
rect 37582 542420 37614 542656
rect 36994 542336 37614 542420
rect 36994 542100 37026 542336
rect 37262 542100 37346 542336
rect 37582 542100 37614 542336
rect 36994 506656 37614 542100
rect 36994 506420 37026 506656
rect 37262 506420 37346 506656
rect 37582 506420 37614 506656
rect 36994 506336 37614 506420
rect 36994 506100 37026 506336
rect 37262 506100 37346 506336
rect 37582 506100 37614 506336
rect 36994 470656 37614 506100
rect 36994 470420 37026 470656
rect 37262 470420 37346 470656
rect 37582 470420 37614 470656
rect 36994 470336 37614 470420
rect 36994 470100 37026 470336
rect 37262 470100 37346 470336
rect 37582 470100 37614 470336
rect 36994 434656 37614 470100
rect 36994 434420 37026 434656
rect 37262 434420 37346 434656
rect 37582 434420 37614 434656
rect 36994 434336 37614 434420
rect 36994 434100 37026 434336
rect 37262 434100 37346 434336
rect 37582 434100 37614 434336
rect 36994 398656 37614 434100
rect 36994 398420 37026 398656
rect 37262 398420 37346 398656
rect 37582 398420 37614 398656
rect 36994 398336 37614 398420
rect 36994 398100 37026 398336
rect 37262 398100 37346 398336
rect 37582 398100 37614 398336
rect 36994 362656 37614 398100
rect 36994 362420 37026 362656
rect 37262 362420 37346 362656
rect 37582 362420 37614 362656
rect 36994 362336 37614 362420
rect 36994 362100 37026 362336
rect 37262 362100 37346 362336
rect 37582 362100 37614 362336
rect 36994 326656 37614 362100
rect 36994 326420 37026 326656
rect 37262 326420 37346 326656
rect 37582 326420 37614 326656
rect 36994 326336 37614 326420
rect 36994 326100 37026 326336
rect 37262 326100 37346 326336
rect 37582 326100 37614 326336
rect 36994 290656 37614 326100
rect 36994 290420 37026 290656
rect 37262 290420 37346 290656
rect 37582 290420 37614 290656
rect 36994 290336 37614 290420
rect 36994 290100 37026 290336
rect 37262 290100 37346 290336
rect 37582 290100 37614 290336
rect 36994 254656 37614 290100
rect 36994 254420 37026 254656
rect 37262 254420 37346 254656
rect 37582 254420 37614 254656
rect 36994 254336 37614 254420
rect 36994 254100 37026 254336
rect 37262 254100 37346 254336
rect 37582 254100 37614 254336
rect 36994 218656 37614 254100
rect 36994 218420 37026 218656
rect 37262 218420 37346 218656
rect 37582 218420 37614 218656
rect 36994 218336 37614 218420
rect 36994 218100 37026 218336
rect 37262 218100 37346 218336
rect 37582 218100 37614 218336
rect 36994 182656 37614 218100
rect 36994 182420 37026 182656
rect 37262 182420 37346 182656
rect 37582 182420 37614 182656
rect 36994 182336 37614 182420
rect 36994 182100 37026 182336
rect 37262 182100 37346 182336
rect 37582 182100 37614 182336
rect 36994 146656 37614 182100
rect 36994 146420 37026 146656
rect 37262 146420 37346 146656
rect 37582 146420 37614 146656
rect 36994 146336 37614 146420
rect 36994 146100 37026 146336
rect 37262 146100 37346 146336
rect 37582 146100 37614 146336
rect 36994 110656 37614 146100
rect 36994 110420 37026 110656
rect 37262 110420 37346 110656
rect 37582 110420 37614 110656
rect 36994 110336 37614 110420
rect 36994 110100 37026 110336
rect 37262 110100 37346 110336
rect 37582 110100 37614 110336
rect 36994 74656 37614 110100
rect 36994 74420 37026 74656
rect 37262 74420 37346 74656
rect 37582 74420 37614 74656
rect 36994 74336 37614 74420
rect 36994 74100 37026 74336
rect 37262 74100 37346 74336
rect 37582 74100 37614 74336
rect 36994 38656 37614 74100
rect 36994 38420 37026 38656
rect 37262 38420 37346 38656
rect 37582 38420 37614 38656
rect 36994 38336 37614 38420
rect 36994 38100 37026 38336
rect 37262 38100 37346 38336
rect 37582 38100 37614 38336
rect 36994 2656 37614 38100
rect 36994 2420 37026 2656
rect 37262 2420 37346 2656
rect 37582 2420 37614 2656
rect 36994 2336 37614 2420
rect 36994 2100 37026 2336
rect 37262 2100 37346 2336
rect 37582 2100 37614 2336
rect 36994 -344 37614 2100
rect 36994 -580 37026 -344
rect 37262 -580 37346 -344
rect 37582 -580 37614 -344
rect 36994 -664 37614 -580
rect 36994 -900 37026 -664
rect 37262 -900 37346 -664
rect 37582 -900 37614 -664
rect 36994 -7652 37614 -900
rect 38234 705800 38854 711592
rect 38234 705564 38266 705800
rect 38502 705564 38586 705800
rect 38822 705564 38854 705800
rect 38234 705480 38854 705564
rect 38234 705244 38266 705480
rect 38502 705244 38586 705480
rect 38822 705244 38854 705480
rect 38234 687896 38854 705244
rect 38234 687660 38266 687896
rect 38502 687660 38586 687896
rect 38822 687660 38854 687896
rect 38234 687576 38854 687660
rect 38234 687340 38266 687576
rect 38502 687340 38586 687576
rect 38822 687340 38854 687576
rect 38234 651896 38854 687340
rect 38234 651660 38266 651896
rect 38502 651660 38586 651896
rect 38822 651660 38854 651896
rect 38234 651576 38854 651660
rect 38234 651340 38266 651576
rect 38502 651340 38586 651576
rect 38822 651340 38854 651576
rect 38234 615896 38854 651340
rect 38234 615660 38266 615896
rect 38502 615660 38586 615896
rect 38822 615660 38854 615896
rect 38234 615576 38854 615660
rect 38234 615340 38266 615576
rect 38502 615340 38586 615576
rect 38822 615340 38854 615576
rect 38234 579896 38854 615340
rect 38234 579660 38266 579896
rect 38502 579660 38586 579896
rect 38822 579660 38854 579896
rect 38234 579576 38854 579660
rect 38234 579340 38266 579576
rect 38502 579340 38586 579576
rect 38822 579340 38854 579576
rect 38234 543896 38854 579340
rect 38234 543660 38266 543896
rect 38502 543660 38586 543896
rect 38822 543660 38854 543896
rect 38234 543576 38854 543660
rect 38234 543340 38266 543576
rect 38502 543340 38586 543576
rect 38822 543340 38854 543576
rect 38234 507896 38854 543340
rect 38234 507660 38266 507896
rect 38502 507660 38586 507896
rect 38822 507660 38854 507896
rect 38234 507576 38854 507660
rect 38234 507340 38266 507576
rect 38502 507340 38586 507576
rect 38822 507340 38854 507576
rect 38234 471896 38854 507340
rect 38234 471660 38266 471896
rect 38502 471660 38586 471896
rect 38822 471660 38854 471896
rect 38234 471576 38854 471660
rect 38234 471340 38266 471576
rect 38502 471340 38586 471576
rect 38822 471340 38854 471576
rect 38234 435896 38854 471340
rect 38234 435660 38266 435896
rect 38502 435660 38586 435896
rect 38822 435660 38854 435896
rect 38234 435576 38854 435660
rect 38234 435340 38266 435576
rect 38502 435340 38586 435576
rect 38822 435340 38854 435576
rect 38234 399896 38854 435340
rect 38234 399660 38266 399896
rect 38502 399660 38586 399896
rect 38822 399660 38854 399896
rect 38234 399576 38854 399660
rect 38234 399340 38266 399576
rect 38502 399340 38586 399576
rect 38822 399340 38854 399576
rect 38234 363896 38854 399340
rect 38234 363660 38266 363896
rect 38502 363660 38586 363896
rect 38822 363660 38854 363896
rect 38234 363576 38854 363660
rect 38234 363340 38266 363576
rect 38502 363340 38586 363576
rect 38822 363340 38854 363576
rect 38234 327896 38854 363340
rect 38234 327660 38266 327896
rect 38502 327660 38586 327896
rect 38822 327660 38854 327896
rect 38234 327576 38854 327660
rect 38234 327340 38266 327576
rect 38502 327340 38586 327576
rect 38822 327340 38854 327576
rect 38234 291896 38854 327340
rect 38234 291660 38266 291896
rect 38502 291660 38586 291896
rect 38822 291660 38854 291896
rect 38234 291576 38854 291660
rect 38234 291340 38266 291576
rect 38502 291340 38586 291576
rect 38822 291340 38854 291576
rect 38234 255896 38854 291340
rect 38234 255660 38266 255896
rect 38502 255660 38586 255896
rect 38822 255660 38854 255896
rect 38234 255576 38854 255660
rect 38234 255340 38266 255576
rect 38502 255340 38586 255576
rect 38822 255340 38854 255576
rect 38234 219896 38854 255340
rect 38234 219660 38266 219896
rect 38502 219660 38586 219896
rect 38822 219660 38854 219896
rect 38234 219576 38854 219660
rect 38234 219340 38266 219576
rect 38502 219340 38586 219576
rect 38822 219340 38854 219576
rect 38234 183896 38854 219340
rect 38234 183660 38266 183896
rect 38502 183660 38586 183896
rect 38822 183660 38854 183896
rect 38234 183576 38854 183660
rect 38234 183340 38266 183576
rect 38502 183340 38586 183576
rect 38822 183340 38854 183576
rect 38234 147896 38854 183340
rect 38234 147660 38266 147896
rect 38502 147660 38586 147896
rect 38822 147660 38854 147896
rect 38234 147576 38854 147660
rect 38234 147340 38266 147576
rect 38502 147340 38586 147576
rect 38822 147340 38854 147576
rect 38234 111896 38854 147340
rect 38234 111660 38266 111896
rect 38502 111660 38586 111896
rect 38822 111660 38854 111896
rect 38234 111576 38854 111660
rect 38234 111340 38266 111576
rect 38502 111340 38586 111576
rect 38822 111340 38854 111576
rect 38234 75896 38854 111340
rect 38234 75660 38266 75896
rect 38502 75660 38586 75896
rect 38822 75660 38854 75896
rect 38234 75576 38854 75660
rect 38234 75340 38266 75576
rect 38502 75340 38586 75576
rect 38822 75340 38854 75576
rect 38234 39896 38854 75340
rect 38234 39660 38266 39896
rect 38502 39660 38586 39896
rect 38822 39660 38854 39896
rect 38234 39576 38854 39660
rect 38234 39340 38266 39576
rect 38502 39340 38586 39576
rect 38822 39340 38854 39576
rect 38234 3896 38854 39340
rect 38234 3660 38266 3896
rect 38502 3660 38586 3896
rect 38822 3660 38854 3896
rect 38234 3576 38854 3660
rect 38234 3340 38266 3576
rect 38502 3340 38586 3576
rect 38822 3340 38854 3576
rect 38234 -1304 38854 3340
rect 38234 -1540 38266 -1304
rect 38502 -1540 38586 -1304
rect 38822 -1540 38854 -1304
rect 38234 -1624 38854 -1540
rect 38234 -1860 38266 -1624
rect 38502 -1860 38586 -1624
rect 38822 -1860 38854 -1624
rect 38234 -7652 38854 -1860
rect 39474 706760 40094 711592
rect 39474 706524 39506 706760
rect 39742 706524 39826 706760
rect 40062 706524 40094 706760
rect 39474 706440 40094 706524
rect 39474 706204 39506 706440
rect 39742 706204 39826 706440
rect 40062 706204 40094 706440
rect 39474 689136 40094 706204
rect 39474 688900 39506 689136
rect 39742 688900 39826 689136
rect 40062 688900 40094 689136
rect 39474 688816 40094 688900
rect 39474 688580 39506 688816
rect 39742 688580 39826 688816
rect 40062 688580 40094 688816
rect 39474 653136 40094 688580
rect 39474 652900 39506 653136
rect 39742 652900 39826 653136
rect 40062 652900 40094 653136
rect 39474 652816 40094 652900
rect 39474 652580 39506 652816
rect 39742 652580 39826 652816
rect 40062 652580 40094 652816
rect 39474 617136 40094 652580
rect 39474 616900 39506 617136
rect 39742 616900 39826 617136
rect 40062 616900 40094 617136
rect 39474 616816 40094 616900
rect 39474 616580 39506 616816
rect 39742 616580 39826 616816
rect 40062 616580 40094 616816
rect 39474 581136 40094 616580
rect 39474 580900 39506 581136
rect 39742 580900 39826 581136
rect 40062 580900 40094 581136
rect 39474 580816 40094 580900
rect 39474 580580 39506 580816
rect 39742 580580 39826 580816
rect 40062 580580 40094 580816
rect 39474 545136 40094 580580
rect 39474 544900 39506 545136
rect 39742 544900 39826 545136
rect 40062 544900 40094 545136
rect 39474 544816 40094 544900
rect 39474 544580 39506 544816
rect 39742 544580 39826 544816
rect 40062 544580 40094 544816
rect 39474 509136 40094 544580
rect 39474 508900 39506 509136
rect 39742 508900 39826 509136
rect 40062 508900 40094 509136
rect 39474 508816 40094 508900
rect 39474 508580 39506 508816
rect 39742 508580 39826 508816
rect 40062 508580 40094 508816
rect 39474 473136 40094 508580
rect 39474 472900 39506 473136
rect 39742 472900 39826 473136
rect 40062 472900 40094 473136
rect 39474 472816 40094 472900
rect 39474 472580 39506 472816
rect 39742 472580 39826 472816
rect 40062 472580 40094 472816
rect 39474 437136 40094 472580
rect 39474 436900 39506 437136
rect 39742 436900 39826 437136
rect 40062 436900 40094 437136
rect 39474 436816 40094 436900
rect 39474 436580 39506 436816
rect 39742 436580 39826 436816
rect 40062 436580 40094 436816
rect 39474 401136 40094 436580
rect 39474 400900 39506 401136
rect 39742 400900 39826 401136
rect 40062 400900 40094 401136
rect 39474 400816 40094 400900
rect 39474 400580 39506 400816
rect 39742 400580 39826 400816
rect 40062 400580 40094 400816
rect 39474 365136 40094 400580
rect 39474 364900 39506 365136
rect 39742 364900 39826 365136
rect 40062 364900 40094 365136
rect 39474 364816 40094 364900
rect 39474 364580 39506 364816
rect 39742 364580 39826 364816
rect 40062 364580 40094 364816
rect 39474 329136 40094 364580
rect 39474 328900 39506 329136
rect 39742 328900 39826 329136
rect 40062 328900 40094 329136
rect 39474 328816 40094 328900
rect 39474 328580 39506 328816
rect 39742 328580 39826 328816
rect 40062 328580 40094 328816
rect 39474 293136 40094 328580
rect 39474 292900 39506 293136
rect 39742 292900 39826 293136
rect 40062 292900 40094 293136
rect 39474 292816 40094 292900
rect 39474 292580 39506 292816
rect 39742 292580 39826 292816
rect 40062 292580 40094 292816
rect 39474 257136 40094 292580
rect 39474 256900 39506 257136
rect 39742 256900 39826 257136
rect 40062 256900 40094 257136
rect 39474 256816 40094 256900
rect 39474 256580 39506 256816
rect 39742 256580 39826 256816
rect 40062 256580 40094 256816
rect 39474 221136 40094 256580
rect 39474 220900 39506 221136
rect 39742 220900 39826 221136
rect 40062 220900 40094 221136
rect 39474 220816 40094 220900
rect 39474 220580 39506 220816
rect 39742 220580 39826 220816
rect 40062 220580 40094 220816
rect 39474 185136 40094 220580
rect 39474 184900 39506 185136
rect 39742 184900 39826 185136
rect 40062 184900 40094 185136
rect 39474 184816 40094 184900
rect 39474 184580 39506 184816
rect 39742 184580 39826 184816
rect 40062 184580 40094 184816
rect 39474 149136 40094 184580
rect 39474 148900 39506 149136
rect 39742 148900 39826 149136
rect 40062 148900 40094 149136
rect 39474 148816 40094 148900
rect 39474 148580 39506 148816
rect 39742 148580 39826 148816
rect 40062 148580 40094 148816
rect 39474 113136 40094 148580
rect 39474 112900 39506 113136
rect 39742 112900 39826 113136
rect 40062 112900 40094 113136
rect 39474 112816 40094 112900
rect 39474 112580 39506 112816
rect 39742 112580 39826 112816
rect 40062 112580 40094 112816
rect 39474 77136 40094 112580
rect 39474 76900 39506 77136
rect 39742 76900 39826 77136
rect 40062 76900 40094 77136
rect 39474 76816 40094 76900
rect 39474 76580 39506 76816
rect 39742 76580 39826 76816
rect 40062 76580 40094 76816
rect 39474 41136 40094 76580
rect 39474 40900 39506 41136
rect 39742 40900 39826 41136
rect 40062 40900 40094 41136
rect 39474 40816 40094 40900
rect 39474 40580 39506 40816
rect 39742 40580 39826 40816
rect 40062 40580 40094 40816
rect 39474 5136 40094 40580
rect 39474 4900 39506 5136
rect 39742 4900 39826 5136
rect 40062 4900 40094 5136
rect 39474 4816 40094 4900
rect 39474 4580 39506 4816
rect 39742 4580 39826 4816
rect 40062 4580 40094 4816
rect 39474 -2264 40094 4580
rect 39474 -2500 39506 -2264
rect 39742 -2500 39826 -2264
rect 40062 -2500 40094 -2264
rect 39474 -2584 40094 -2500
rect 39474 -2820 39506 -2584
rect 39742 -2820 39826 -2584
rect 40062 -2820 40094 -2584
rect 39474 -7652 40094 -2820
rect 40714 707720 41334 711592
rect 40714 707484 40746 707720
rect 40982 707484 41066 707720
rect 41302 707484 41334 707720
rect 40714 707400 41334 707484
rect 40714 707164 40746 707400
rect 40982 707164 41066 707400
rect 41302 707164 41334 707400
rect 40714 690376 41334 707164
rect 40714 690140 40746 690376
rect 40982 690140 41066 690376
rect 41302 690140 41334 690376
rect 40714 690056 41334 690140
rect 40714 689820 40746 690056
rect 40982 689820 41066 690056
rect 41302 689820 41334 690056
rect 40714 654376 41334 689820
rect 40714 654140 40746 654376
rect 40982 654140 41066 654376
rect 41302 654140 41334 654376
rect 40714 654056 41334 654140
rect 40714 653820 40746 654056
rect 40982 653820 41066 654056
rect 41302 653820 41334 654056
rect 40714 618376 41334 653820
rect 40714 618140 40746 618376
rect 40982 618140 41066 618376
rect 41302 618140 41334 618376
rect 40714 618056 41334 618140
rect 40714 617820 40746 618056
rect 40982 617820 41066 618056
rect 41302 617820 41334 618056
rect 40714 582376 41334 617820
rect 40714 582140 40746 582376
rect 40982 582140 41066 582376
rect 41302 582140 41334 582376
rect 40714 582056 41334 582140
rect 40714 581820 40746 582056
rect 40982 581820 41066 582056
rect 41302 581820 41334 582056
rect 40714 546376 41334 581820
rect 40714 546140 40746 546376
rect 40982 546140 41066 546376
rect 41302 546140 41334 546376
rect 40714 546056 41334 546140
rect 40714 545820 40746 546056
rect 40982 545820 41066 546056
rect 41302 545820 41334 546056
rect 40714 510376 41334 545820
rect 40714 510140 40746 510376
rect 40982 510140 41066 510376
rect 41302 510140 41334 510376
rect 40714 510056 41334 510140
rect 40714 509820 40746 510056
rect 40982 509820 41066 510056
rect 41302 509820 41334 510056
rect 40714 474376 41334 509820
rect 40714 474140 40746 474376
rect 40982 474140 41066 474376
rect 41302 474140 41334 474376
rect 40714 474056 41334 474140
rect 40714 473820 40746 474056
rect 40982 473820 41066 474056
rect 41302 473820 41334 474056
rect 40714 438376 41334 473820
rect 40714 438140 40746 438376
rect 40982 438140 41066 438376
rect 41302 438140 41334 438376
rect 40714 438056 41334 438140
rect 40714 437820 40746 438056
rect 40982 437820 41066 438056
rect 41302 437820 41334 438056
rect 40714 402376 41334 437820
rect 40714 402140 40746 402376
rect 40982 402140 41066 402376
rect 41302 402140 41334 402376
rect 40714 402056 41334 402140
rect 40714 401820 40746 402056
rect 40982 401820 41066 402056
rect 41302 401820 41334 402056
rect 40714 366376 41334 401820
rect 40714 366140 40746 366376
rect 40982 366140 41066 366376
rect 41302 366140 41334 366376
rect 40714 366056 41334 366140
rect 40714 365820 40746 366056
rect 40982 365820 41066 366056
rect 41302 365820 41334 366056
rect 40714 330376 41334 365820
rect 40714 330140 40746 330376
rect 40982 330140 41066 330376
rect 41302 330140 41334 330376
rect 40714 330056 41334 330140
rect 40714 329820 40746 330056
rect 40982 329820 41066 330056
rect 41302 329820 41334 330056
rect 40714 294376 41334 329820
rect 40714 294140 40746 294376
rect 40982 294140 41066 294376
rect 41302 294140 41334 294376
rect 40714 294056 41334 294140
rect 40714 293820 40746 294056
rect 40982 293820 41066 294056
rect 41302 293820 41334 294056
rect 40714 258376 41334 293820
rect 40714 258140 40746 258376
rect 40982 258140 41066 258376
rect 41302 258140 41334 258376
rect 40714 258056 41334 258140
rect 40714 257820 40746 258056
rect 40982 257820 41066 258056
rect 41302 257820 41334 258056
rect 40714 222376 41334 257820
rect 40714 222140 40746 222376
rect 40982 222140 41066 222376
rect 41302 222140 41334 222376
rect 40714 222056 41334 222140
rect 40714 221820 40746 222056
rect 40982 221820 41066 222056
rect 41302 221820 41334 222056
rect 40714 186376 41334 221820
rect 40714 186140 40746 186376
rect 40982 186140 41066 186376
rect 41302 186140 41334 186376
rect 40714 186056 41334 186140
rect 40714 185820 40746 186056
rect 40982 185820 41066 186056
rect 41302 185820 41334 186056
rect 40714 150376 41334 185820
rect 40714 150140 40746 150376
rect 40982 150140 41066 150376
rect 41302 150140 41334 150376
rect 40714 150056 41334 150140
rect 40714 149820 40746 150056
rect 40982 149820 41066 150056
rect 41302 149820 41334 150056
rect 40714 114376 41334 149820
rect 40714 114140 40746 114376
rect 40982 114140 41066 114376
rect 41302 114140 41334 114376
rect 40714 114056 41334 114140
rect 40714 113820 40746 114056
rect 40982 113820 41066 114056
rect 41302 113820 41334 114056
rect 40714 78376 41334 113820
rect 40714 78140 40746 78376
rect 40982 78140 41066 78376
rect 41302 78140 41334 78376
rect 40714 78056 41334 78140
rect 40714 77820 40746 78056
rect 40982 77820 41066 78056
rect 41302 77820 41334 78056
rect 40714 42376 41334 77820
rect 40714 42140 40746 42376
rect 40982 42140 41066 42376
rect 41302 42140 41334 42376
rect 40714 42056 41334 42140
rect 40714 41820 40746 42056
rect 40982 41820 41066 42056
rect 41302 41820 41334 42056
rect 40714 6376 41334 41820
rect 40714 6140 40746 6376
rect 40982 6140 41066 6376
rect 41302 6140 41334 6376
rect 40714 6056 41334 6140
rect 40714 5820 40746 6056
rect 40982 5820 41066 6056
rect 41302 5820 41334 6056
rect 40714 -3224 41334 5820
rect 40714 -3460 40746 -3224
rect 40982 -3460 41066 -3224
rect 41302 -3460 41334 -3224
rect 40714 -3544 41334 -3460
rect 40714 -3780 40746 -3544
rect 40982 -3780 41066 -3544
rect 41302 -3780 41334 -3544
rect 40714 -7652 41334 -3780
rect 41954 708680 42574 711592
rect 41954 708444 41986 708680
rect 42222 708444 42306 708680
rect 42542 708444 42574 708680
rect 41954 708360 42574 708444
rect 41954 708124 41986 708360
rect 42222 708124 42306 708360
rect 42542 708124 42574 708360
rect 41954 691616 42574 708124
rect 41954 691380 41986 691616
rect 42222 691380 42306 691616
rect 42542 691380 42574 691616
rect 41954 691296 42574 691380
rect 41954 691060 41986 691296
rect 42222 691060 42306 691296
rect 42542 691060 42574 691296
rect 41954 655616 42574 691060
rect 41954 655380 41986 655616
rect 42222 655380 42306 655616
rect 42542 655380 42574 655616
rect 41954 655296 42574 655380
rect 41954 655060 41986 655296
rect 42222 655060 42306 655296
rect 42542 655060 42574 655296
rect 41954 619616 42574 655060
rect 41954 619380 41986 619616
rect 42222 619380 42306 619616
rect 42542 619380 42574 619616
rect 41954 619296 42574 619380
rect 41954 619060 41986 619296
rect 42222 619060 42306 619296
rect 42542 619060 42574 619296
rect 41954 583616 42574 619060
rect 41954 583380 41986 583616
rect 42222 583380 42306 583616
rect 42542 583380 42574 583616
rect 41954 583296 42574 583380
rect 41954 583060 41986 583296
rect 42222 583060 42306 583296
rect 42542 583060 42574 583296
rect 41954 547616 42574 583060
rect 41954 547380 41986 547616
rect 42222 547380 42306 547616
rect 42542 547380 42574 547616
rect 41954 547296 42574 547380
rect 41954 547060 41986 547296
rect 42222 547060 42306 547296
rect 42542 547060 42574 547296
rect 41954 511616 42574 547060
rect 41954 511380 41986 511616
rect 42222 511380 42306 511616
rect 42542 511380 42574 511616
rect 41954 511296 42574 511380
rect 41954 511060 41986 511296
rect 42222 511060 42306 511296
rect 42542 511060 42574 511296
rect 41954 475616 42574 511060
rect 41954 475380 41986 475616
rect 42222 475380 42306 475616
rect 42542 475380 42574 475616
rect 41954 475296 42574 475380
rect 41954 475060 41986 475296
rect 42222 475060 42306 475296
rect 42542 475060 42574 475296
rect 41954 439616 42574 475060
rect 41954 439380 41986 439616
rect 42222 439380 42306 439616
rect 42542 439380 42574 439616
rect 41954 439296 42574 439380
rect 41954 439060 41986 439296
rect 42222 439060 42306 439296
rect 42542 439060 42574 439296
rect 41954 403616 42574 439060
rect 41954 403380 41986 403616
rect 42222 403380 42306 403616
rect 42542 403380 42574 403616
rect 41954 403296 42574 403380
rect 41954 403060 41986 403296
rect 42222 403060 42306 403296
rect 42542 403060 42574 403296
rect 41954 367616 42574 403060
rect 41954 367380 41986 367616
rect 42222 367380 42306 367616
rect 42542 367380 42574 367616
rect 41954 367296 42574 367380
rect 41954 367060 41986 367296
rect 42222 367060 42306 367296
rect 42542 367060 42574 367296
rect 41954 331616 42574 367060
rect 41954 331380 41986 331616
rect 42222 331380 42306 331616
rect 42542 331380 42574 331616
rect 41954 331296 42574 331380
rect 41954 331060 41986 331296
rect 42222 331060 42306 331296
rect 42542 331060 42574 331296
rect 41954 295616 42574 331060
rect 41954 295380 41986 295616
rect 42222 295380 42306 295616
rect 42542 295380 42574 295616
rect 41954 295296 42574 295380
rect 41954 295060 41986 295296
rect 42222 295060 42306 295296
rect 42542 295060 42574 295296
rect 41954 259616 42574 295060
rect 41954 259380 41986 259616
rect 42222 259380 42306 259616
rect 42542 259380 42574 259616
rect 41954 259296 42574 259380
rect 41954 259060 41986 259296
rect 42222 259060 42306 259296
rect 42542 259060 42574 259296
rect 41954 223616 42574 259060
rect 41954 223380 41986 223616
rect 42222 223380 42306 223616
rect 42542 223380 42574 223616
rect 41954 223296 42574 223380
rect 41954 223060 41986 223296
rect 42222 223060 42306 223296
rect 42542 223060 42574 223296
rect 41954 187616 42574 223060
rect 41954 187380 41986 187616
rect 42222 187380 42306 187616
rect 42542 187380 42574 187616
rect 41954 187296 42574 187380
rect 41954 187060 41986 187296
rect 42222 187060 42306 187296
rect 42542 187060 42574 187296
rect 41954 151616 42574 187060
rect 41954 151380 41986 151616
rect 42222 151380 42306 151616
rect 42542 151380 42574 151616
rect 41954 151296 42574 151380
rect 41954 151060 41986 151296
rect 42222 151060 42306 151296
rect 42542 151060 42574 151296
rect 41954 115616 42574 151060
rect 41954 115380 41986 115616
rect 42222 115380 42306 115616
rect 42542 115380 42574 115616
rect 41954 115296 42574 115380
rect 41954 115060 41986 115296
rect 42222 115060 42306 115296
rect 42542 115060 42574 115296
rect 41954 79616 42574 115060
rect 41954 79380 41986 79616
rect 42222 79380 42306 79616
rect 42542 79380 42574 79616
rect 41954 79296 42574 79380
rect 41954 79060 41986 79296
rect 42222 79060 42306 79296
rect 42542 79060 42574 79296
rect 41954 43616 42574 79060
rect 41954 43380 41986 43616
rect 42222 43380 42306 43616
rect 42542 43380 42574 43616
rect 41954 43296 42574 43380
rect 41954 43060 41986 43296
rect 42222 43060 42306 43296
rect 42542 43060 42574 43296
rect 41954 7616 42574 43060
rect 41954 7380 41986 7616
rect 42222 7380 42306 7616
rect 42542 7380 42574 7616
rect 41954 7296 42574 7380
rect 41954 7060 41986 7296
rect 42222 7060 42306 7296
rect 42542 7060 42574 7296
rect 41954 -4184 42574 7060
rect 41954 -4420 41986 -4184
rect 42222 -4420 42306 -4184
rect 42542 -4420 42574 -4184
rect 41954 -4504 42574 -4420
rect 41954 -4740 41986 -4504
rect 42222 -4740 42306 -4504
rect 42542 -4740 42574 -4504
rect 41954 -7652 42574 -4740
rect 43194 709640 43814 711592
rect 43194 709404 43226 709640
rect 43462 709404 43546 709640
rect 43782 709404 43814 709640
rect 43194 709320 43814 709404
rect 43194 709084 43226 709320
rect 43462 709084 43546 709320
rect 43782 709084 43814 709320
rect 43194 692856 43814 709084
rect 43194 692620 43226 692856
rect 43462 692620 43546 692856
rect 43782 692620 43814 692856
rect 43194 692536 43814 692620
rect 43194 692300 43226 692536
rect 43462 692300 43546 692536
rect 43782 692300 43814 692536
rect 43194 656856 43814 692300
rect 43194 656620 43226 656856
rect 43462 656620 43546 656856
rect 43782 656620 43814 656856
rect 43194 656536 43814 656620
rect 43194 656300 43226 656536
rect 43462 656300 43546 656536
rect 43782 656300 43814 656536
rect 43194 620856 43814 656300
rect 43194 620620 43226 620856
rect 43462 620620 43546 620856
rect 43782 620620 43814 620856
rect 43194 620536 43814 620620
rect 43194 620300 43226 620536
rect 43462 620300 43546 620536
rect 43782 620300 43814 620536
rect 43194 584856 43814 620300
rect 43194 584620 43226 584856
rect 43462 584620 43546 584856
rect 43782 584620 43814 584856
rect 43194 584536 43814 584620
rect 43194 584300 43226 584536
rect 43462 584300 43546 584536
rect 43782 584300 43814 584536
rect 43194 548856 43814 584300
rect 43194 548620 43226 548856
rect 43462 548620 43546 548856
rect 43782 548620 43814 548856
rect 43194 548536 43814 548620
rect 43194 548300 43226 548536
rect 43462 548300 43546 548536
rect 43782 548300 43814 548536
rect 43194 512856 43814 548300
rect 43194 512620 43226 512856
rect 43462 512620 43546 512856
rect 43782 512620 43814 512856
rect 43194 512536 43814 512620
rect 43194 512300 43226 512536
rect 43462 512300 43546 512536
rect 43782 512300 43814 512536
rect 43194 476856 43814 512300
rect 43194 476620 43226 476856
rect 43462 476620 43546 476856
rect 43782 476620 43814 476856
rect 43194 476536 43814 476620
rect 43194 476300 43226 476536
rect 43462 476300 43546 476536
rect 43782 476300 43814 476536
rect 43194 440856 43814 476300
rect 43194 440620 43226 440856
rect 43462 440620 43546 440856
rect 43782 440620 43814 440856
rect 43194 440536 43814 440620
rect 43194 440300 43226 440536
rect 43462 440300 43546 440536
rect 43782 440300 43814 440536
rect 43194 404856 43814 440300
rect 43194 404620 43226 404856
rect 43462 404620 43546 404856
rect 43782 404620 43814 404856
rect 43194 404536 43814 404620
rect 43194 404300 43226 404536
rect 43462 404300 43546 404536
rect 43782 404300 43814 404536
rect 43194 368856 43814 404300
rect 43194 368620 43226 368856
rect 43462 368620 43546 368856
rect 43782 368620 43814 368856
rect 43194 368536 43814 368620
rect 43194 368300 43226 368536
rect 43462 368300 43546 368536
rect 43782 368300 43814 368536
rect 43194 332856 43814 368300
rect 43194 332620 43226 332856
rect 43462 332620 43546 332856
rect 43782 332620 43814 332856
rect 43194 332536 43814 332620
rect 43194 332300 43226 332536
rect 43462 332300 43546 332536
rect 43782 332300 43814 332536
rect 43194 296856 43814 332300
rect 43194 296620 43226 296856
rect 43462 296620 43546 296856
rect 43782 296620 43814 296856
rect 43194 296536 43814 296620
rect 43194 296300 43226 296536
rect 43462 296300 43546 296536
rect 43782 296300 43814 296536
rect 43194 260856 43814 296300
rect 43194 260620 43226 260856
rect 43462 260620 43546 260856
rect 43782 260620 43814 260856
rect 43194 260536 43814 260620
rect 43194 260300 43226 260536
rect 43462 260300 43546 260536
rect 43782 260300 43814 260536
rect 43194 224856 43814 260300
rect 43194 224620 43226 224856
rect 43462 224620 43546 224856
rect 43782 224620 43814 224856
rect 43194 224536 43814 224620
rect 43194 224300 43226 224536
rect 43462 224300 43546 224536
rect 43782 224300 43814 224536
rect 43194 188856 43814 224300
rect 43194 188620 43226 188856
rect 43462 188620 43546 188856
rect 43782 188620 43814 188856
rect 43194 188536 43814 188620
rect 43194 188300 43226 188536
rect 43462 188300 43546 188536
rect 43782 188300 43814 188536
rect 43194 152856 43814 188300
rect 43194 152620 43226 152856
rect 43462 152620 43546 152856
rect 43782 152620 43814 152856
rect 43194 152536 43814 152620
rect 43194 152300 43226 152536
rect 43462 152300 43546 152536
rect 43782 152300 43814 152536
rect 43194 116856 43814 152300
rect 43194 116620 43226 116856
rect 43462 116620 43546 116856
rect 43782 116620 43814 116856
rect 43194 116536 43814 116620
rect 43194 116300 43226 116536
rect 43462 116300 43546 116536
rect 43782 116300 43814 116536
rect 43194 80856 43814 116300
rect 43194 80620 43226 80856
rect 43462 80620 43546 80856
rect 43782 80620 43814 80856
rect 43194 80536 43814 80620
rect 43194 80300 43226 80536
rect 43462 80300 43546 80536
rect 43782 80300 43814 80536
rect 43194 44856 43814 80300
rect 43194 44620 43226 44856
rect 43462 44620 43546 44856
rect 43782 44620 43814 44856
rect 43194 44536 43814 44620
rect 43194 44300 43226 44536
rect 43462 44300 43546 44536
rect 43782 44300 43814 44536
rect 43194 8856 43814 44300
rect 43194 8620 43226 8856
rect 43462 8620 43546 8856
rect 43782 8620 43814 8856
rect 43194 8536 43814 8620
rect 43194 8300 43226 8536
rect 43462 8300 43546 8536
rect 43782 8300 43814 8536
rect 43194 -5144 43814 8300
rect 43194 -5380 43226 -5144
rect 43462 -5380 43546 -5144
rect 43782 -5380 43814 -5144
rect 43194 -5464 43814 -5380
rect 43194 -5700 43226 -5464
rect 43462 -5700 43546 -5464
rect 43782 -5700 43814 -5464
rect 43194 -7652 43814 -5700
rect 44434 710600 45054 711592
rect 44434 710364 44466 710600
rect 44702 710364 44786 710600
rect 45022 710364 45054 710600
rect 44434 710280 45054 710364
rect 44434 710044 44466 710280
rect 44702 710044 44786 710280
rect 45022 710044 45054 710280
rect 44434 694096 45054 710044
rect 44434 693860 44466 694096
rect 44702 693860 44786 694096
rect 45022 693860 45054 694096
rect 44434 693776 45054 693860
rect 44434 693540 44466 693776
rect 44702 693540 44786 693776
rect 45022 693540 45054 693776
rect 44434 658096 45054 693540
rect 44434 657860 44466 658096
rect 44702 657860 44786 658096
rect 45022 657860 45054 658096
rect 44434 657776 45054 657860
rect 44434 657540 44466 657776
rect 44702 657540 44786 657776
rect 45022 657540 45054 657776
rect 44434 622096 45054 657540
rect 44434 621860 44466 622096
rect 44702 621860 44786 622096
rect 45022 621860 45054 622096
rect 44434 621776 45054 621860
rect 44434 621540 44466 621776
rect 44702 621540 44786 621776
rect 45022 621540 45054 621776
rect 44434 586096 45054 621540
rect 44434 585860 44466 586096
rect 44702 585860 44786 586096
rect 45022 585860 45054 586096
rect 44434 585776 45054 585860
rect 44434 585540 44466 585776
rect 44702 585540 44786 585776
rect 45022 585540 45054 585776
rect 44434 550096 45054 585540
rect 44434 549860 44466 550096
rect 44702 549860 44786 550096
rect 45022 549860 45054 550096
rect 44434 549776 45054 549860
rect 44434 549540 44466 549776
rect 44702 549540 44786 549776
rect 45022 549540 45054 549776
rect 44434 514096 45054 549540
rect 44434 513860 44466 514096
rect 44702 513860 44786 514096
rect 45022 513860 45054 514096
rect 44434 513776 45054 513860
rect 44434 513540 44466 513776
rect 44702 513540 44786 513776
rect 45022 513540 45054 513776
rect 44434 478096 45054 513540
rect 44434 477860 44466 478096
rect 44702 477860 44786 478096
rect 45022 477860 45054 478096
rect 44434 477776 45054 477860
rect 44434 477540 44466 477776
rect 44702 477540 44786 477776
rect 45022 477540 45054 477776
rect 44434 442096 45054 477540
rect 44434 441860 44466 442096
rect 44702 441860 44786 442096
rect 45022 441860 45054 442096
rect 44434 441776 45054 441860
rect 44434 441540 44466 441776
rect 44702 441540 44786 441776
rect 45022 441540 45054 441776
rect 44434 406096 45054 441540
rect 44434 405860 44466 406096
rect 44702 405860 44786 406096
rect 45022 405860 45054 406096
rect 44434 405776 45054 405860
rect 44434 405540 44466 405776
rect 44702 405540 44786 405776
rect 45022 405540 45054 405776
rect 44434 370096 45054 405540
rect 44434 369860 44466 370096
rect 44702 369860 44786 370096
rect 45022 369860 45054 370096
rect 44434 369776 45054 369860
rect 44434 369540 44466 369776
rect 44702 369540 44786 369776
rect 45022 369540 45054 369776
rect 44434 334096 45054 369540
rect 44434 333860 44466 334096
rect 44702 333860 44786 334096
rect 45022 333860 45054 334096
rect 44434 333776 45054 333860
rect 44434 333540 44466 333776
rect 44702 333540 44786 333776
rect 45022 333540 45054 333776
rect 44434 298096 45054 333540
rect 44434 297860 44466 298096
rect 44702 297860 44786 298096
rect 45022 297860 45054 298096
rect 44434 297776 45054 297860
rect 44434 297540 44466 297776
rect 44702 297540 44786 297776
rect 45022 297540 45054 297776
rect 44434 262096 45054 297540
rect 44434 261860 44466 262096
rect 44702 261860 44786 262096
rect 45022 261860 45054 262096
rect 44434 261776 45054 261860
rect 44434 261540 44466 261776
rect 44702 261540 44786 261776
rect 45022 261540 45054 261776
rect 44434 226096 45054 261540
rect 44434 225860 44466 226096
rect 44702 225860 44786 226096
rect 45022 225860 45054 226096
rect 44434 225776 45054 225860
rect 44434 225540 44466 225776
rect 44702 225540 44786 225776
rect 45022 225540 45054 225776
rect 44434 190096 45054 225540
rect 44434 189860 44466 190096
rect 44702 189860 44786 190096
rect 45022 189860 45054 190096
rect 44434 189776 45054 189860
rect 44434 189540 44466 189776
rect 44702 189540 44786 189776
rect 45022 189540 45054 189776
rect 44434 154096 45054 189540
rect 44434 153860 44466 154096
rect 44702 153860 44786 154096
rect 45022 153860 45054 154096
rect 44434 153776 45054 153860
rect 44434 153540 44466 153776
rect 44702 153540 44786 153776
rect 45022 153540 45054 153776
rect 44434 118096 45054 153540
rect 44434 117860 44466 118096
rect 44702 117860 44786 118096
rect 45022 117860 45054 118096
rect 44434 117776 45054 117860
rect 44434 117540 44466 117776
rect 44702 117540 44786 117776
rect 45022 117540 45054 117776
rect 44434 82096 45054 117540
rect 44434 81860 44466 82096
rect 44702 81860 44786 82096
rect 45022 81860 45054 82096
rect 44434 81776 45054 81860
rect 44434 81540 44466 81776
rect 44702 81540 44786 81776
rect 45022 81540 45054 81776
rect 44434 46096 45054 81540
rect 44434 45860 44466 46096
rect 44702 45860 44786 46096
rect 45022 45860 45054 46096
rect 44434 45776 45054 45860
rect 44434 45540 44466 45776
rect 44702 45540 44786 45776
rect 45022 45540 45054 45776
rect 44434 10096 45054 45540
rect 44434 9860 44466 10096
rect 44702 9860 44786 10096
rect 45022 9860 45054 10096
rect 44434 9776 45054 9860
rect 44434 9540 44466 9776
rect 44702 9540 44786 9776
rect 45022 9540 45054 9776
rect 44434 -6104 45054 9540
rect 44434 -6340 44466 -6104
rect 44702 -6340 44786 -6104
rect 45022 -6340 45054 -6104
rect 44434 -6424 45054 -6340
rect 44434 -6660 44466 -6424
rect 44702 -6660 44786 -6424
rect 45022 -6660 45054 -6424
rect 44434 -7652 45054 -6660
rect 45674 711560 46294 711592
rect 45674 711324 45706 711560
rect 45942 711324 46026 711560
rect 46262 711324 46294 711560
rect 45674 711240 46294 711324
rect 45674 711004 45706 711240
rect 45942 711004 46026 711240
rect 46262 711004 46294 711240
rect 45674 695336 46294 711004
rect 45674 695100 45706 695336
rect 45942 695100 46026 695336
rect 46262 695100 46294 695336
rect 45674 695016 46294 695100
rect 45674 694780 45706 695016
rect 45942 694780 46026 695016
rect 46262 694780 46294 695016
rect 45674 659336 46294 694780
rect 45674 659100 45706 659336
rect 45942 659100 46026 659336
rect 46262 659100 46294 659336
rect 45674 659016 46294 659100
rect 45674 658780 45706 659016
rect 45942 658780 46026 659016
rect 46262 658780 46294 659016
rect 45674 623336 46294 658780
rect 45674 623100 45706 623336
rect 45942 623100 46026 623336
rect 46262 623100 46294 623336
rect 45674 623016 46294 623100
rect 45674 622780 45706 623016
rect 45942 622780 46026 623016
rect 46262 622780 46294 623016
rect 45674 587336 46294 622780
rect 45674 587100 45706 587336
rect 45942 587100 46026 587336
rect 46262 587100 46294 587336
rect 45674 587016 46294 587100
rect 45674 586780 45706 587016
rect 45942 586780 46026 587016
rect 46262 586780 46294 587016
rect 45674 551336 46294 586780
rect 45674 551100 45706 551336
rect 45942 551100 46026 551336
rect 46262 551100 46294 551336
rect 45674 551016 46294 551100
rect 45674 550780 45706 551016
rect 45942 550780 46026 551016
rect 46262 550780 46294 551016
rect 45674 515336 46294 550780
rect 45674 515100 45706 515336
rect 45942 515100 46026 515336
rect 46262 515100 46294 515336
rect 45674 515016 46294 515100
rect 45674 514780 45706 515016
rect 45942 514780 46026 515016
rect 46262 514780 46294 515016
rect 45674 479336 46294 514780
rect 45674 479100 45706 479336
rect 45942 479100 46026 479336
rect 46262 479100 46294 479336
rect 45674 479016 46294 479100
rect 45674 478780 45706 479016
rect 45942 478780 46026 479016
rect 46262 478780 46294 479016
rect 45674 443336 46294 478780
rect 45674 443100 45706 443336
rect 45942 443100 46026 443336
rect 46262 443100 46294 443336
rect 45674 443016 46294 443100
rect 45674 442780 45706 443016
rect 45942 442780 46026 443016
rect 46262 442780 46294 443016
rect 45674 407336 46294 442780
rect 45674 407100 45706 407336
rect 45942 407100 46026 407336
rect 46262 407100 46294 407336
rect 45674 407016 46294 407100
rect 45674 406780 45706 407016
rect 45942 406780 46026 407016
rect 46262 406780 46294 407016
rect 45674 371336 46294 406780
rect 45674 371100 45706 371336
rect 45942 371100 46026 371336
rect 46262 371100 46294 371336
rect 45674 371016 46294 371100
rect 45674 370780 45706 371016
rect 45942 370780 46026 371016
rect 46262 370780 46294 371016
rect 45674 335336 46294 370780
rect 45674 335100 45706 335336
rect 45942 335100 46026 335336
rect 46262 335100 46294 335336
rect 45674 335016 46294 335100
rect 45674 334780 45706 335016
rect 45942 334780 46026 335016
rect 46262 334780 46294 335016
rect 45674 299336 46294 334780
rect 45674 299100 45706 299336
rect 45942 299100 46026 299336
rect 46262 299100 46294 299336
rect 45674 299016 46294 299100
rect 45674 298780 45706 299016
rect 45942 298780 46026 299016
rect 46262 298780 46294 299016
rect 45674 263336 46294 298780
rect 45674 263100 45706 263336
rect 45942 263100 46026 263336
rect 46262 263100 46294 263336
rect 45674 263016 46294 263100
rect 45674 262780 45706 263016
rect 45942 262780 46026 263016
rect 46262 262780 46294 263016
rect 45674 227336 46294 262780
rect 45674 227100 45706 227336
rect 45942 227100 46026 227336
rect 46262 227100 46294 227336
rect 45674 227016 46294 227100
rect 45674 226780 45706 227016
rect 45942 226780 46026 227016
rect 46262 226780 46294 227016
rect 45674 191336 46294 226780
rect 45674 191100 45706 191336
rect 45942 191100 46026 191336
rect 46262 191100 46294 191336
rect 45674 191016 46294 191100
rect 45674 190780 45706 191016
rect 45942 190780 46026 191016
rect 46262 190780 46294 191016
rect 45674 155336 46294 190780
rect 45674 155100 45706 155336
rect 45942 155100 46026 155336
rect 46262 155100 46294 155336
rect 45674 155016 46294 155100
rect 45674 154780 45706 155016
rect 45942 154780 46026 155016
rect 46262 154780 46294 155016
rect 45674 119336 46294 154780
rect 45674 119100 45706 119336
rect 45942 119100 46026 119336
rect 46262 119100 46294 119336
rect 45674 119016 46294 119100
rect 45674 118780 45706 119016
rect 45942 118780 46026 119016
rect 46262 118780 46294 119016
rect 45674 83336 46294 118780
rect 45674 83100 45706 83336
rect 45942 83100 46026 83336
rect 46262 83100 46294 83336
rect 45674 83016 46294 83100
rect 45674 82780 45706 83016
rect 45942 82780 46026 83016
rect 46262 82780 46294 83016
rect 45674 47336 46294 82780
rect 45674 47100 45706 47336
rect 45942 47100 46026 47336
rect 46262 47100 46294 47336
rect 45674 47016 46294 47100
rect 45674 46780 45706 47016
rect 45942 46780 46026 47016
rect 46262 46780 46294 47016
rect 45674 11336 46294 46780
rect 45674 11100 45706 11336
rect 45942 11100 46026 11336
rect 46262 11100 46294 11336
rect 45674 11016 46294 11100
rect 45674 10780 45706 11016
rect 45942 10780 46026 11016
rect 46262 10780 46294 11016
rect 45674 -7064 46294 10780
rect 45674 -7300 45706 -7064
rect 45942 -7300 46026 -7064
rect 46262 -7300 46294 -7064
rect 45674 -7384 46294 -7300
rect 45674 -7620 45706 -7384
rect 45942 -7620 46026 -7384
rect 46262 -7620 46294 -7384
rect 45674 -7652 46294 -7620
rect 72994 704840 73614 711592
rect 72994 704604 73026 704840
rect 73262 704604 73346 704840
rect 73582 704604 73614 704840
rect 72994 704520 73614 704604
rect 72994 704284 73026 704520
rect 73262 704284 73346 704520
rect 73582 704284 73614 704520
rect 72994 686656 73614 704284
rect 72994 686420 73026 686656
rect 73262 686420 73346 686656
rect 73582 686420 73614 686656
rect 72994 686336 73614 686420
rect 72994 686100 73026 686336
rect 73262 686100 73346 686336
rect 73582 686100 73614 686336
rect 72994 650656 73614 686100
rect 72994 650420 73026 650656
rect 73262 650420 73346 650656
rect 73582 650420 73614 650656
rect 72994 650336 73614 650420
rect 72994 650100 73026 650336
rect 73262 650100 73346 650336
rect 73582 650100 73614 650336
rect 72994 614656 73614 650100
rect 72994 614420 73026 614656
rect 73262 614420 73346 614656
rect 73582 614420 73614 614656
rect 72994 614336 73614 614420
rect 72994 614100 73026 614336
rect 73262 614100 73346 614336
rect 73582 614100 73614 614336
rect 72994 578656 73614 614100
rect 72994 578420 73026 578656
rect 73262 578420 73346 578656
rect 73582 578420 73614 578656
rect 72994 578336 73614 578420
rect 72994 578100 73026 578336
rect 73262 578100 73346 578336
rect 73582 578100 73614 578336
rect 72994 542656 73614 578100
rect 72994 542420 73026 542656
rect 73262 542420 73346 542656
rect 73582 542420 73614 542656
rect 72994 542336 73614 542420
rect 72994 542100 73026 542336
rect 73262 542100 73346 542336
rect 73582 542100 73614 542336
rect 72994 506656 73614 542100
rect 72994 506420 73026 506656
rect 73262 506420 73346 506656
rect 73582 506420 73614 506656
rect 72994 506336 73614 506420
rect 72994 506100 73026 506336
rect 73262 506100 73346 506336
rect 73582 506100 73614 506336
rect 72994 470656 73614 506100
rect 72994 470420 73026 470656
rect 73262 470420 73346 470656
rect 73582 470420 73614 470656
rect 72994 470336 73614 470420
rect 72994 470100 73026 470336
rect 73262 470100 73346 470336
rect 73582 470100 73614 470336
rect 72994 434656 73614 470100
rect 72994 434420 73026 434656
rect 73262 434420 73346 434656
rect 73582 434420 73614 434656
rect 72994 434336 73614 434420
rect 72994 434100 73026 434336
rect 73262 434100 73346 434336
rect 73582 434100 73614 434336
rect 72994 398656 73614 434100
rect 72994 398420 73026 398656
rect 73262 398420 73346 398656
rect 73582 398420 73614 398656
rect 72994 398336 73614 398420
rect 72994 398100 73026 398336
rect 73262 398100 73346 398336
rect 73582 398100 73614 398336
rect 72994 362656 73614 398100
rect 72994 362420 73026 362656
rect 73262 362420 73346 362656
rect 73582 362420 73614 362656
rect 72994 362336 73614 362420
rect 72994 362100 73026 362336
rect 73262 362100 73346 362336
rect 73582 362100 73614 362336
rect 72994 326656 73614 362100
rect 72994 326420 73026 326656
rect 73262 326420 73346 326656
rect 73582 326420 73614 326656
rect 72994 326336 73614 326420
rect 72994 326100 73026 326336
rect 73262 326100 73346 326336
rect 73582 326100 73614 326336
rect 72994 290656 73614 326100
rect 72994 290420 73026 290656
rect 73262 290420 73346 290656
rect 73582 290420 73614 290656
rect 72994 290336 73614 290420
rect 72994 290100 73026 290336
rect 73262 290100 73346 290336
rect 73582 290100 73614 290336
rect 72994 254656 73614 290100
rect 72994 254420 73026 254656
rect 73262 254420 73346 254656
rect 73582 254420 73614 254656
rect 72994 254336 73614 254420
rect 72994 254100 73026 254336
rect 73262 254100 73346 254336
rect 73582 254100 73614 254336
rect 72994 218656 73614 254100
rect 72994 218420 73026 218656
rect 73262 218420 73346 218656
rect 73582 218420 73614 218656
rect 72994 218336 73614 218420
rect 72994 218100 73026 218336
rect 73262 218100 73346 218336
rect 73582 218100 73614 218336
rect 72994 182656 73614 218100
rect 72994 182420 73026 182656
rect 73262 182420 73346 182656
rect 73582 182420 73614 182656
rect 72994 182336 73614 182420
rect 72994 182100 73026 182336
rect 73262 182100 73346 182336
rect 73582 182100 73614 182336
rect 72994 146656 73614 182100
rect 72994 146420 73026 146656
rect 73262 146420 73346 146656
rect 73582 146420 73614 146656
rect 72994 146336 73614 146420
rect 72994 146100 73026 146336
rect 73262 146100 73346 146336
rect 73582 146100 73614 146336
rect 72994 110656 73614 146100
rect 72994 110420 73026 110656
rect 73262 110420 73346 110656
rect 73582 110420 73614 110656
rect 72994 110336 73614 110420
rect 72994 110100 73026 110336
rect 73262 110100 73346 110336
rect 73582 110100 73614 110336
rect 72994 74656 73614 110100
rect 72994 74420 73026 74656
rect 73262 74420 73346 74656
rect 73582 74420 73614 74656
rect 72994 74336 73614 74420
rect 72994 74100 73026 74336
rect 73262 74100 73346 74336
rect 73582 74100 73614 74336
rect 72994 38656 73614 74100
rect 72994 38420 73026 38656
rect 73262 38420 73346 38656
rect 73582 38420 73614 38656
rect 72994 38336 73614 38420
rect 72994 38100 73026 38336
rect 73262 38100 73346 38336
rect 73582 38100 73614 38336
rect 72994 2656 73614 38100
rect 72994 2420 73026 2656
rect 73262 2420 73346 2656
rect 73582 2420 73614 2656
rect 72994 2336 73614 2420
rect 72994 2100 73026 2336
rect 73262 2100 73346 2336
rect 73582 2100 73614 2336
rect 72994 -344 73614 2100
rect 72994 -580 73026 -344
rect 73262 -580 73346 -344
rect 73582 -580 73614 -344
rect 72994 -664 73614 -580
rect 72994 -900 73026 -664
rect 73262 -900 73346 -664
rect 73582 -900 73614 -664
rect 72994 -7652 73614 -900
rect 74234 705800 74854 711592
rect 74234 705564 74266 705800
rect 74502 705564 74586 705800
rect 74822 705564 74854 705800
rect 74234 705480 74854 705564
rect 74234 705244 74266 705480
rect 74502 705244 74586 705480
rect 74822 705244 74854 705480
rect 74234 687896 74854 705244
rect 74234 687660 74266 687896
rect 74502 687660 74586 687896
rect 74822 687660 74854 687896
rect 74234 687576 74854 687660
rect 74234 687340 74266 687576
rect 74502 687340 74586 687576
rect 74822 687340 74854 687576
rect 74234 651896 74854 687340
rect 74234 651660 74266 651896
rect 74502 651660 74586 651896
rect 74822 651660 74854 651896
rect 74234 651576 74854 651660
rect 74234 651340 74266 651576
rect 74502 651340 74586 651576
rect 74822 651340 74854 651576
rect 74234 615896 74854 651340
rect 74234 615660 74266 615896
rect 74502 615660 74586 615896
rect 74822 615660 74854 615896
rect 74234 615576 74854 615660
rect 74234 615340 74266 615576
rect 74502 615340 74586 615576
rect 74822 615340 74854 615576
rect 74234 579896 74854 615340
rect 74234 579660 74266 579896
rect 74502 579660 74586 579896
rect 74822 579660 74854 579896
rect 74234 579576 74854 579660
rect 74234 579340 74266 579576
rect 74502 579340 74586 579576
rect 74822 579340 74854 579576
rect 74234 543896 74854 579340
rect 74234 543660 74266 543896
rect 74502 543660 74586 543896
rect 74822 543660 74854 543896
rect 74234 543576 74854 543660
rect 74234 543340 74266 543576
rect 74502 543340 74586 543576
rect 74822 543340 74854 543576
rect 74234 507896 74854 543340
rect 74234 507660 74266 507896
rect 74502 507660 74586 507896
rect 74822 507660 74854 507896
rect 74234 507576 74854 507660
rect 74234 507340 74266 507576
rect 74502 507340 74586 507576
rect 74822 507340 74854 507576
rect 74234 471896 74854 507340
rect 74234 471660 74266 471896
rect 74502 471660 74586 471896
rect 74822 471660 74854 471896
rect 74234 471576 74854 471660
rect 74234 471340 74266 471576
rect 74502 471340 74586 471576
rect 74822 471340 74854 471576
rect 74234 435896 74854 471340
rect 74234 435660 74266 435896
rect 74502 435660 74586 435896
rect 74822 435660 74854 435896
rect 74234 435576 74854 435660
rect 74234 435340 74266 435576
rect 74502 435340 74586 435576
rect 74822 435340 74854 435576
rect 74234 399896 74854 435340
rect 74234 399660 74266 399896
rect 74502 399660 74586 399896
rect 74822 399660 74854 399896
rect 74234 399576 74854 399660
rect 74234 399340 74266 399576
rect 74502 399340 74586 399576
rect 74822 399340 74854 399576
rect 74234 363896 74854 399340
rect 74234 363660 74266 363896
rect 74502 363660 74586 363896
rect 74822 363660 74854 363896
rect 74234 363576 74854 363660
rect 74234 363340 74266 363576
rect 74502 363340 74586 363576
rect 74822 363340 74854 363576
rect 74234 327896 74854 363340
rect 74234 327660 74266 327896
rect 74502 327660 74586 327896
rect 74822 327660 74854 327896
rect 74234 327576 74854 327660
rect 74234 327340 74266 327576
rect 74502 327340 74586 327576
rect 74822 327340 74854 327576
rect 74234 291896 74854 327340
rect 74234 291660 74266 291896
rect 74502 291660 74586 291896
rect 74822 291660 74854 291896
rect 74234 291576 74854 291660
rect 74234 291340 74266 291576
rect 74502 291340 74586 291576
rect 74822 291340 74854 291576
rect 74234 255896 74854 291340
rect 74234 255660 74266 255896
rect 74502 255660 74586 255896
rect 74822 255660 74854 255896
rect 74234 255576 74854 255660
rect 74234 255340 74266 255576
rect 74502 255340 74586 255576
rect 74822 255340 74854 255576
rect 74234 219896 74854 255340
rect 74234 219660 74266 219896
rect 74502 219660 74586 219896
rect 74822 219660 74854 219896
rect 74234 219576 74854 219660
rect 74234 219340 74266 219576
rect 74502 219340 74586 219576
rect 74822 219340 74854 219576
rect 74234 183896 74854 219340
rect 74234 183660 74266 183896
rect 74502 183660 74586 183896
rect 74822 183660 74854 183896
rect 74234 183576 74854 183660
rect 74234 183340 74266 183576
rect 74502 183340 74586 183576
rect 74822 183340 74854 183576
rect 74234 147896 74854 183340
rect 74234 147660 74266 147896
rect 74502 147660 74586 147896
rect 74822 147660 74854 147896
rect 74234 147576 74854 147660
rect 74234 147340 74266 147576
rect 74502 147340 74586 147576
rect 74822 147340 74854 147576
rect 74234 111896 74854 147340
rect 74234 111660 74266 111896
rect 74502 111660 74586 111896
rect 74822 111660 74854 111896
rect 74234 111576 74854 111660
rect 74234 111340 74266 111576
rect 74502 111340 74586 111576
rect 74822 111340 74854 111576
rect 74234 75896 74854 111340
rect 74234 75660 74266 75896
rect 74502 75660 74586 75896
rect 74822 75660 74854 75896
rect 74234 75576 74854 75660
rect 74234 75340 74266 75576
rect 74502 75340 74586 75576
rect 74822 75340 74854 75576
rect 74234 39896 74854 75340
rect 74234 39660 74266 39896
rect 74502 39660 74586 39896
rect 74822 39660 74854 39896
rect 74234 39576 74854 39660
rect 74234 39340 74266 39576
rect 74502 39340 74586 39576
rect 74822 39340 74854 39576
rect 74234 3896 74854 39340
rect 74234 3660 74266 3896
rect 74502 3660 74586 3896
rect 74822 3660 74854 3896
rect 74234 3576 74854 3660
rect 74234 3340 74266 3576
rect 74502 3340 74586 3576
rect 74822 3340 74854 3576
rect 74234 -1304 74854 3340
rect 74234 -1540 74266 -1304
rect 74502 -1540 74586 -1304
rect 74822 -1540 74854 -1304
rect 74234 -1624 74854 -1540
rect 74234 -1860 74266 -1624
rect 74502 -1860 74586 -1624
rect 74822 -1860 74854 -1624
rect 74234 -7652 74854 -1860
rect 75474 706760 76094 711592
rect 75474 706524 75506 706760
rect 75742 706524 75826 706760
rect 76062 706524 76094 706760
rect 75474 706440 76094 706524
rect 75474 706204 75506 706440
rect 75742 706204 75826 706440
rect 76062 706204 76094 706440
rect 75474 689136 76094 706204
rect 75474 688900 75506 689136
rect 75742 688900 75826 689136
rect 76062 688900 76094 689136
rect 75474 688816 76094 688900
rect 75474 688580 75506 688816
rect 75742 688580 75826 688816
rect 76062 688580 76094 688816
rect 75474 653136 76094 688580
rect 75474 652900 75506 653136
rect 75742 652900 75826 653136
rect 76062 652900 76094 653136
rect 75474 652816 76094 652900
rect 75474 652580 75506 652816
rect 75742 652580 75826 652816
rect 76062 652580 76094 652816
rect 75474 617136 76094 652580
rect 75474 616900 75506 617136
rect 75742 616900 75826 617136
rect 76062 616900 76094 617136
rect 75474 616816 76094 616900
rect 75474 616580 75506 616816
rect 75742 616580 75826 616816
rect 76062 616580 76094 616816
rect 75474 581136 76094 616580
rect 75474 580900 75506 581136
rect 75742 580900 75826 581136
rect 76062 580900 76094 581136
rect 75474 580816 76094 580900
rect 75474 580580 75506 580816
rect 75742 580580 75826 580816
rect 76062 580580 76094 580816
rect 75474 545136 76094 580580
rect 75474 544900 75506 545136
rect 75742 544900 75826 545136
rect 76062 544900 76094 545136
rect 75474 544816 76094 544900
rect 75474 544580 75506 544816
rect 75742 544580 75826 544816
rect 76062 544580 76094 544816
rect 75474 509136 76094 544580
rect 75474 508900 75506 509136
rect 75742 508900 75826 509136
rect 76062 508900 76094 509136
rect 75474 508816 76094 508900
rect 75474 508580 75506 508816
rect 75742 508580 75826 508816
rect 76062 508580 76094 508816
rect 75474 473136 76094 508580
rect 75474 472900 75506 473136
rect 75742 472900 75826 473136
rect 76062 472900 76094 473136
rect 75474 472816 76094 472900
rect 75474 472580 75506 472816
rect 75742 472580 75826 472816
rect 76062 472580 76094 472816
rect 75474 437136 76094 472580
rect 75474 436900 75506 437136
rect 75742 436900 75826 437136
rect 76062 436900 76094 437136
rect 75474 436816 76094 436900
rect 75474 436580 75506 436816
rect 75742 436580 75826 436816
rect 76062 436580 76094 436816
rect 75474 401136 76094 436580
rect 75474 400900 75506 401136
rect 75742 400900 75826 401136
rect 76062 400900 76094 401136
rect 75474 400816 76094 400900
rect 75474 400580 75506 400816
rect 75742 400580 75826 400816
rect 76062 400580 76094 400816
rect 75474 365136 76094 400580
rect 75474 364900 75506 365136
rect 75742 364900 75826 365136
rect 76062 364900 76094 365136
rect 75474 364816 76094 364900
rect 75474 364580 75506 364816
rect 75742 364580 75826 364816
rect 76062 364580 76094 364816
rect 75474 329136 76094 364580
rect 75474 328900 75506 329136
rect 75742 328900 75826 329136
rect 76062 328900 76094 329136
rect 75474 328816 76094 328900
rect 75474 328580 75506 328816
rect 75742 328580 75826 328816
rect 76062 328580 76094 328816
rect 75474 293136 76094 328580
rect 75474 292900 75506 293136
rect 75742 292900 75826 293136
rect 76062 292900 76094 293136
rect 75474 292816 76094 292900
rect 75474 292580 75506 292816
rect 75742 292580 75826 292816
rect 76062 292580 76094 292816
rect 75474 257136 76094 292580
rect 75474 256900 75506 257136
rect 75742 256900 75826 257136
rect 76062 256900 76094 257136
rect 75474 256816 76094 256900
rect 75474 256580 75506 256816
rect 75742 256580 75826 256816
rect 76062 256580 76094 256816
rect 75474 221136 76094 256580
rect 75474 220900 75506 221136
rect 75742 220900 75826 221136
rect 76062 220900 76094 221136
rect 75474 220816 76094 220900
rect 75474 220580 75506 220816
rect 75742 220580 75826 220816
rect 76062 220580 76094 220816
rect 75474 185136 76094 220580
rect 75474 184900 75506 185136
rect 75742 184900 75826 185136
rect 76062 184900 76094 185136
rect 75474 184816 76094 184900
rect 75474 184580 75506 184816
rect 75742 184580 75826 184816
rect 76062 184580 76094 184816
rect 75474 149136 76094 184580
rect 75474 148900 75506 149136
rect 75742 148900 75826 149136
rect 76062 148900 76094 149136
rect 75474 148816 76094 148900
rect 75474 148580 75506 148816
rect 75742 148580 75826 148816
rect 76062 148580 76094 148816
rect 75474 113136 76094 148580
rect 75474 112900 75506 113136
rect 75742 112900 75826 113136
rect 76062 112900 76094 113136
rect 75474 112816 76094 112900
rect 75474 112580 75506 112816
rect 75742 112580 75826 112816
rect 76062 112580 76094 112816
rect 75474 77136 76094 112580
rect 75474 76900 75506 77136
rect 75742 76900 75826 77136
rect 76062 76900 76094 77136
rect 75474 76816 76094 76900
rect 75474 76580 75506 76816
rect 75742 76580 75826 76816
rect 76062 76580 76094 76816
rect 75474 41136 76094 76580
rect 75474 40900 75506 41136
rect 75742 40900 75826 41136
rect 76062 40900 76094 41136
rect 75474 40816 76094 40900
rect 75474 40580 75506 40816
rect 75742 40580 75826 40816
rect 76062 40580 76094 40816
rect 75474 5136 76094 40580
rect 75474 4900 75506 5136
rect 75742 4900 75826 5136
rect 76062 4900 76094 5136
rect 75474 4816 76094 4900
rect 75474 4580 75506 4816
rect 75742 4580 75826 4816
rect 76062 4580 76094 4816
rect 75474 -2264 76094 4580
rect 75474 -2500 75506 -2264
rect 75742 -2500 75826 -2264
rect 76062 -2500 76094 -2264
rect 75474 -2584 76094 -2500
rect 75474 -2820 75506 -2584
rect 75742 -2820 75826 -2584
rect 76062 -2820 76094 -2584
rect 75474 -7652 76094 -2820
rect 76714 707720 77334 711592
rect 76714 707484 76746 707720
rect 76982 707484 77066 707720
rect 77302 707484 77334 707720
rect 76714 707400 77334 707484
rect 76714 707164 76746 707400
rect 76982 707164 77066 707400
rect 77302 707164 77334 707400
rect 76714 690376 77334 707164
rect 76714 690140 76746 690376
rect 76982 690140 77066 690376
rect 77302 690140 77334 690376
rect 76714 690056 77334 690140
rect 76714 689820 76746 690056
rect 76982 689820 77066 690056
rect 77302 689820 77334 690056
rect 76714 654376 77334 689820
rect 76714 654140 76746 654376
rect 76982 654140 77066 654376
rect 77302 654140 77334 654376
rect 76714 654056 77334 654140
rect 76714 653820 76746 654056
rect 76982 653820 77066 654056
rect 77302 653820 77334 654056
rect 76714 618376 77334 653820
rect 76714 618140 76746 618376
rect 76982 618140 77066 618376
rect 77302 618140 77334 618376
rect 76714 618056 77334 618140
rect 76714 617820 76746 618056
rect 76982 617820 77066 618056
rect 77302 617820 77334 618056
rect 76714 582376 77334 617820
rect 76714 582140 76746 582376
rect 76982 582140 77066 582376
rect 77302 582140 77334 582376
rect 76714 582056 77334 582140
rect 76714 581820 76746 582056
rect 76982 581820 77066 582056
rect 77302 581820 77334 582056
rect 76714 546376 77334 581820
rect 76714 546140 76746 546376
rect 76982 546140 77066 546376
rect 77302 546140 77334 546376
rect 76714 546056 77334 546140
rect 76714 545820 76746 546056
rect 76982 545820 77066 546056
rect 77302 545820 77334 546056
rect 76714 510376 77334 545820
rect 76714 510140 76746 510376
rect 76982 510140 77066 510376
rect 77302 510140 77334 510376
rect 76714 510056 77334 510140
rect 76714 509820 76746 510056
rect 76982 509820 77066 510056
rect 77302 509820 77334 510056
rect 76714 474376 77334 509820
rect 76714 474140 76746 474376
rect 76982 474140 77066 474376
rect 77302 474140 77334 474376
rect 76714 474056 77334 474140
rect 76714 473820 76746 474056
rect 76982 473820 77066 474056
rect 77302 473820 77334 474056
rect 76714 438376 77334 473820
rect 76714 438140 76746 438376
rect 76982 438140 77066 438376
rect 77302 438140 77334 438376
rect 76714 438056 77334 438140
rect 76714 437820 76746 438056
rect 76982 437820 77066 438056
rect 77302 437820 77334 438056
rect 76714 402376 77334 437820
rect 76714 402140 76746 402376
rect 76982 402140 77066 402376
rect 77302 402140 77334 402376
rect 76714 402056 77334 402140
rect 76714 401820 76746 402056
rect 76982 401820 77066 402056
rect 77302 401820 77334 402056
rect 76714 366376 77334 401820
rect 76714 366140 76746 366376
rect 76982 366140 77066 366376
rect 77302 366140 77334 366376
rect 76714 366056 77334 366140
rect 76714 365820 76746 366056
rect 76982 365820 77066 366056
rect 77302 365820 77334 366056
rect 76714 330376 77334 365820
rect 76714 330140 76746 330376
rect 76982 330140 77066 330376
rect 77302 330140 77334 330376
rect 76714 330056 77334 330140
rect 76714 329820 76746 330056
rect 76982 329820 77066 330056
rect 77302 329820 77334 330056
rect 76714 294376 77334 329820
rect 76714 294140 76746 294376
rect 76982 294140 77066 294376
rect 77302 294140 77334 294376
rect 76714 294056 77334 294140
rect 76714 293820 76746 294056
rect 76982 293820 77066 294056
rect 77302 293820 77334 294056
rect 76714 258376 77334 293820
rect 76714 258140 76746 258376
rect 76982 258140 77066 258376
rect 77302 258140 77334 258376
rect 76714 258056 77334 258140
rect 76714 257820 76746 258056
rect 76982 257820 77066 258056
rect 77302 257820 77334 258056
rect 76714 222376 77334 257820
rect 76714 222140 76746 222376
rect 76982 222140 77066 222376
rect 77302 222140 77334 222376
rect 76714 222056 77334 222140
rect 76714 221820 76746 222056
rect 76982 221820 77066 222056
rect 77302 221820 77334 222056
rect 76714 186376 77334 221820
rect 76714 186140 76746 186376
rect 76982 186140 77066 186376
rect 77302 186140 77334 186376
rect 76714 186056 77334 186140
rect 76714 185820 76746 186056
rect 76982 185820 77066 186056
rect 77302 185820 77334 186056
rect 76714 150376 77334 185820
rect 76714 150140 76746 150376
rect 76982 150140 77066 150376
rect 77302 150140 77334 150376
rect 76714 150056 77334 150140
rect 76714 149820 76746 150056
rect 76982 149820 77066 150056
rect 77302 149820 77334 150056
rect 76714 114376 77334 149820
rect 76714 114140 76746 114376
rect 76982 114140 77066 114376
rect 77302 114140 77334 114376
rect 76714 114056 77334 114140
rect 76714 113820 76746 114056
rect 76982 113820 77066 114056
rect 77302 113820 77334 114056
rect 76714 78376 77334 113820
rect 76714 78140 76746 78376
rect 76982 78140 77066 78376
rect 77302 78140 77334 78376
rect 76714 78056 77334 78140
rect 76714 77820 76746 78056
rect 76982 77820 77066 78056
rect 77302 77820 77334 78056
rect 76714 42376 77334 77820
rect 76714 42140 76746 42376
rect 76982 42140 77066 42376
rect 77302 42140 77334 42376
rect 76714 42056 77334 42140
rect 76714 41820 76746 42056
rect 76982 41820 77066 42056
rect 77302 41820 77334 42056
rect 76714 6376 77334 41820
rect 76714 6140 76746 6376
rect 76982 6140 77066 6376
rect 77302 6140 77334 6376
rect 76714 6056 77334 6140
rect 76714 5820 76746 6056
rect 76982 5820 77066 6056
rect 77302 5820 77334 6056
rect 76714 -3224 77334 5820
rect 76714 -3460 76746 -3224
rect 76982 -3460 77066 -3224
rect 77302 -3460 77334 -3224
rect 76714 -3544 77334 -3460
rect 76714 -3780 76746 -3544
rect 76982 -3780 77066 -3544
rect 77302 -3780 77334 -3544
rect 76714 -7652 77334 -3780
rect 77954 708680 78574 711592
rect 77954 708444 77986 708680
rect 78222 708444 78306 708680
rect 78542 708444 78574 708680
rect 77954 708360 78574 708444
rect 77954 708124 77986 708360
rect 78222 708124 78306 708360
rect 78542 708124 78574 708360
rect 77954 691616 78574 708124
rect 77954 691380 77986 691616
rect 78222 691380 78306 691616
rect 78542 691380 78574 691616
rect 77954 691296 78574 691380
rect 77954 691060 77986 691296
rect 78222 691060 78306 691296
rect 78542 691060 78574 691296
rect 77954 655616 78574 691060
rect 77954 655380 77986 655616
rect 78222 655380 78306 655616
rect 78542 655380 78574 655616
rect 77954 655296 78574 655380
rect 77954 655060 77986 655296
rect 78222 655060 78306 655296
rect 78542 655060 78574 655296
rect 77954 619616 78574 655060
rect 77954 619380 77986 619616
rect 78222 619380 78306 619616
rect 78542 619380 78574 619616
rect 77954 619296 78574 619380
rect 77954 619060 77986 619296
rect 78222 619060 78306 619296
rect 78542 619060 78574 619296
rect 77954 583616 78574 619060
rect 77954 583380 77986 583616
rect 78222 583380 78306 583616
rect 78542 583380 78574 583616
rect 77954 583296 78574 583380
rect 77954 583060 77986 583296
rect 78222 583060 78306 583296
rect 78542 583060 78574 583296
rect 77954 547616 78574 583060
rect 77954 547380 77986 547616
rect 78222 547380 78306 547616
rect 78542 547380 78574 547616
rect 77954 547296 78574 547380
rect 77954 547060 77986 547296
rect 78222 547060 78306 547296
rect 78542 547060 78574 547296
rect 77954 511616 78574 547060
rect 77954 511380 77986 511616
rect 78222 511380 78306 511616
rect 78542 511380 78574 511616
rect 77954 511296 78574 511380
rect 77954 511060 77986 511296
rect 78222 511060 78306 511296
rect 78542 511060 78574 511296
rect 77954 475616 78574 511060
rect 77954 475380 77986 475616
rect 78222 475380 78306 475616
rect 78542 475380 78574 475616
rect 77954 475296 78574 475380
rect 77954 475060 77986 475296
rect 78222 475060 78306 475296
rect 78542 475060 78574 475296
rect 77954 439616 78574 475060
rect 77954 439380 77986 439616
rect 78222 439380 78306 439616
rect 78542 439380 78574 439616
rect 77954 439296 78574 439380
rect 77954 439060 77986 439296
rect 78222 439060 78306 439296
rect 78542 439060 78574 439296
rect 77954 403616 78574 439060
rect 77954 403380 77986 403616
rect 78222 403380 78306 403616
rect 78542 403380 78574 403616
rect 77954 403296 78574 403380
rect 77954 403060 77986 403296
rect 78222 403060 78306 403296
rect 78542 403060 78574 403296
rect 77954 367616 78574 403060
rect 77954 367380 77986 367616
rect 78222 367380 78306 367616
rect 78542 367380 78574 367616
rect 77954 367296 78574 367380
rect 77954 367060 77986 367296
rect 78222 367060 78306 367296
rect 78542 367060 78574 367296
rect 77954 331616 78574 367060
rect 77954 331380 77986 331616
rect 78222 331380 78306 331616
rect 78542 331380 78574 331616
rect 77954 331296 78574 331380
rect 77954 331060 77986 331296
rect 78222 331060 78306 331296
rect 78542 331060 78574 331296
rect 77954 295616 78574 331060
rect 77954 295380 77986 295616
rect 78222 295380 78306 295616
rect 78542 295380 78574 295616
rect 77954 295296 78574 295380
rect 77954 295060 77986 295296
rect 78222 295060 78306 295296
rect 78542 295060 78574 295296
rect 77954 259616 78574 295060
rect 77954 259380 77986 259616
rect 78222 259380 78306 259616
rect 78542 259380 78574 259616
rect 77954 259296 78574 259380
rect 77954 259060 77986 259296
rect 78222 259060 78306 259296
rect 78542 259060 78574 259296
rect 77954 223616 78574 259060
rect 77954 223380 77986 223616
rect 78222 223380 78306 223616
rect 78542 223380 78574 223616
rect 77954 223296 78574 223380
rect 77954 223060 77986 223296
rect 78222 223060 78306 223296
rect 78542 223060 78574 223296
rect 77954 187616 78574 223060
rect 77954 187380 77986 187616
rect 78222 187380 78306 187616
rect 78542 187380 78574 187616
rect 77954 187296 78574 187380
rect 77954 187060 77986 187296
rect 78222 187060 78306 187296
rect 78542 187060 78574 187296
rect 77954 151616 78574 187060
rect 77954 151380 77986 151616
rect 78222 151380 78306 151616
rect 78542 151380 78574 151616
rect 77954 151296 78574 151380
rect 77954 151060 77986 151296
rect 78222 151060 78306 151296
rect 78542 151060 78574 151296
rect 77954 115616 78574 151060
rect 77954 115380 77986 115616
rect 78222 115380 78306 115616
rect 78542 115380 78574 115616
rect 77954 115296 78574 115380
rect 77954 115060 77986 115296
rect 78222 115060 78306 115296
rect 78542 115060 78574 115296
rect 77954 79616 78574 115060
rect 77954 79380 77986 79616
rect 78222 79380 78306 79616
rect 78542 79380 78574 79616
rect 77954 79296 78574 79380
rect 77954 79060 77986 79296
rect 78222 79060 78306 79296
rect 78542 79060 78574 79296
rect 77954 43616 78574 79060
rect 77954 43380 77986 43616
rect 78222 43380 78306 43616
rect 78542 43380 78574 43616
rect 77954 43296 78574 43380
rect 77954 43060 77986 43296
rect 78222 43060 78306 43296
rect 78542 43060 78574 43296
rect 77954 7616 78574 43060
rect 77954 7380 77986 7616
rect 78222 7380 78306 7616
rect 78542 7380 78574 7616
rect 77954 7296 78574 7380
rect 77954 7060 77986 7296
rect 78222 7060 78306 7296
rect 78542 7060 78574 7296
rect 77954 -4184 78574 7060
rect 77954 -4420 77986 -4184
rect 78222 -4420 78306 -4184
rect 78542 -4420 78574 -4184
rect 77954 -4504 78574 -4420
rect 77954 -4740 77986 -4504
rect 78222 -4740 78306 -4504
rect 78542 -4740 78574 -4504
rect 77954 -7652 78574 -4740
rect 79194 709640 79814 711592
rect 79194 709404 79226 709640
rect 79462 709404 79546 709640
rect 79782 709404 79814 709640
rect 79194 709320 79814 709404
rect 79194 709084 79226 709320
rect 79462 709084 79546 709320
rect 79782 709084 79814 709320
rect 79194 692856 79814 709084
rect 79194 692620 79226 692856
rect 79462 692620 79546 692856
rect 79782 692620 79814 692856
rect 79194 692536 79814 692620
rect 79194 692300 79226 692536
rect 79462 692300 79546 692536
rect 79782 692300 79814 692536
rect 79194 656856 79814 692300
rect 79194 656620 79226 656856
rect 79462 656620 79546 656856
rect 79782 656620 79814 656856
rect 79194 656536 79814 656620
rect 79194 656300 79226 656536
rect 79462 656300 79546 656536
rect 79782 656300 79814 656536
rect 79194 620856 79814 656300
rect 79194 620620 79226 620856
rect 79462 620620 79546 620856
rect 79782 620620 79814 620856
rect 79194 620536 79814 620620
rect 79194 620300 79226 620536
rect 79462 620300 79546 620536
rect 79782 620300 79814 620536
rect 79194 584856 79814 620300
rect 79194 584620 79226 584856
rect 79462 584620 79546 584856
rect 79782 584620 79814 584856
rect 79194 584536 79814 584620
rect 79194 584300 79226 584536
rect 79462 584300 79546 584536
rect 79782 584300 79814 584536
rect 79194 548856 79814 584300
rect 79194 548620 79226 548856
rect 79462 548620 79546 548856
rect 79782 548620 79814 548856
rect 79194 548536 79814 548620
rect 79194 548300 79226 548536
rect 79462 548300 79546 548536
rect 79782 548300 79814 548536
rect 79194 512856 79814 548300
rect 79194 512620 79226 512856
rect 79462 512620 79546 512856
rect 79782 512620 79814 512856
rect 79194 512536 79814 512620
rect 79194 512300 79226 512536
rect 79462 512300 79546 512536
rect 79782 512300 79814 512536
rect 79194 476856 79814 512300
rect 79194 476620 79226 476856
rect 79462 476620 79546 476856
rect 79782 476620 79814 476856
rect 79194 476536 79814 476620
rect 79194 476300 79226 476536
rect 79462 476300 79546 476536
rect 79782 476300 79814 476536
rect 79194 440856 79814 476300
rect 79194 440620 79226 440856
rect 79462 440620 79546 440856
rect 79782 440620 79814 440856
rect 79194 440536 79814 440620
rect 79194 440300 79226 440536
rect 79462 440300 79546 440536
rect 79782 440300 79814 440536
rect 79194 404856 79814 440300
rect 79194 404620 79226 404856
rect 79462 404620 79546 404856
rect 79782 404620 79814 404856
rect 79194 404536 79814 404620
rect 79194 404300 79226 404536
rect 79462 404300 79546 404536
rect 79782 404300 79814 404536
rect 79194 368856 79814 404300
rect 79194 368620 79226 368856
rect 79462 368620 79546 368856
rect 79782 368620 79814 368856
rect 79194 368536 79814 368620
rect 79194 368300 79226 368536
rect 79462 368300 79546 368536
rect 79782 368300 79814 368536
rect 79194 332856 79814 368300
rect 79194 332620 79226 332856
rect 79462 332620 79546 332856
rect 79782 332620 79814 332856
rect 79194 332536 79814 332620
rect 79194 332300 79226 332536
rect 79462 332300 79546 332536
rect 79782 332300 79814 332536
rect 79194 296856 79814 332300
rect 79194 296620 79226 296856
rect 79462 296620 79546 296856
rect 79782 296620 79814 296856
rect 79194 296536 79814 296620
rect 79194 296300 79226 296536
rect 79462 296300 79546 296536
rect 79782 296300 79814 296536
rect 79194 260856 79814 296300
rect 79194 260620 79226 260856
rect 79462 260620 79546 260856
rect 79782 260620 79814 260856
rect 79194 260536 79814 260620
rect 79194 260300 79226 260536
rect 79462 260300 79546 260536
rect 79782 260300 79814 260536
rect 79194 224856 79814 260300
rect 79194 224620 79226 224856
rect 79462 224620 79546 224856
rect 79782 224620 79814 224856
rect 79194 224536 79814 224620
rect 79194 224300 79226 224536
rect 79462 224300 79546 224536
rect 79782 224300 79814 224536
rect 79194 188856 79814 224300
rect 79194 188620 79226 188856
rect 79462 188620 79546 188856
rect 79782 188620 79814 188856
rect 79194 188536 79814 188620
rect 79194 188300 79226 188536
rect 79462 188300 79546 188536
rect 79782 188300 79814 188536
rect 79194 152856 79814 188300
rect 79194 152620 79226 152856
rect 79462 152620 79546 152856
rect 79782 152620 79814 152856
rect 79194 152536 79814 152620
rect 79194 152300 79226 152536
rect 79462 152300 79546 152536
rect 79782 152300 79814 152536
rect 79194 116856 79814 152300
rect 79194 116620 79226 116856
rect 79462 116620 79546 116856
rect 79782 116620 79814 116856
rect 79194 116536 79814 116620
rect 79194 116300 79226 116536
rect 79462 116300 79546 116536
rect 79782 116300 79814 116536
rect 79194 80856 79814 116300
rect 79194 80620 79226 80856
rect 79462 80620 79546 80856
rect 79782 80620 79814 80856
rect 79194 80536 79814 80620
rect 79194 80300 79226 80536
rect 79462 80300 79546 80536
rect 79782 80300 79814 80536
rect 79194 44856 79814 80300
rect 79194 44620 79226 44856
rect 79462 44620 79546 44856
rect 79782 44620 79814 44856
rect 79194 44536 79814 44620
rect 79194 44300 79226 44536
rect 79462 44300 79546 44536
rect 79782 44300 79814 44536
rect 79194 8856 79814 44300
rect 79194 8620 79226 8856
rect 79462 8620 79546 8856
rect 79782 8620 79814 8856
rect 79194 8536 79814 8620
rect 79194 8300 79226 8536
rect 79462 8300 79546 8536
rect 79782 8300 79814 8536
rect 79194 -5144 79814 8300
rect 79194 -5380 79226 -5144
rect 79462 -5380 79546 -5144
rect 79782 -5380 79814 -5144
rect 79194 -5464 79814 -5380
rect 79194 -5700 79226 -5464
rect 79462 -5700 79546 -5464
rect 79782 -5700 79814 -5464
rect 79194 -7652 79814 -5700
rect 80434 710600 81054 711592
rect 80434 710364 80466 710600
rect 80702 710364 80786 710600
rect 81022 710364 81054 710600
rect 80434 710280 81054 710364
rect 80434 710044 80466 710280
rect 80702 710044 80786 710280
rect 81022 710044 81054 710280
rect 80434 694096 81054 710044
rect 80434 693860 80466 694096
rect 80702 693860 80786 694096
rect 81022 693860 81054 694096
rect 80434 693776 81054 693860
rect 80434 693540 80466 693776
rect 80702 693540 80786 693776
rect 81022 693540 81054 693776
rect 80434 658096 81054 693540
rect 80434 657860 80466 658096
rect 80702 657860 80786 658096
rect 81022 657860 81054 658096
rect 80434 657776 81054 657860
rect 80434 657540 80466 657776
rect 80702 657540 80786 657776
rect 81022 657540 81054 657776
rect 80434 622096 81054 657540
rect 80434 621860 80466 622096
rect 80702 621860 80786 622096
rect 81022 621860 81054 622096
rect 80434 621776 81054 621860
rect 80434 621540 80466 621776
rect 80702 621540 80786 621776
rect 81022 621540 81054 621776
rect 80434 586096 81054 621540
rect 80434 585860 80466 586096
rect 80702 585860 80786 586096
rect 81022 585860 81054 586096
rect 80434 585776 81054 585860
rect 80434 585540 80466 585776
rect 80702 585540 80786 585776
rect 81022 585540 81054 585776
rect 80434 550096 81054 585540
rect 80434 549860 80466 550096
rect 80702 549860 80786 550096
rect 81022 549860 81054 550096
rect 80434 549776 81054 549860
rect 80434 549540 80466 549776
rect 80702 549540 80786 549776
rect 81022 549540 81054 549776
rect 80434 514096 81054 549540
rect 80434 513860 80466 514096
rect 80702 513860 80786 514096
rect 81022 513860 81054 514096
rect 80434 513776 81054 513860
rect 80434 513540 80466 513776
rect 80702 513540 80786 513776
rect 81022 513540 81054 513776
rect 80434 478096 81054 513540
rect 80434 477860 80466 478096
rect 80702 477860 80786 478096
rect 81022 477860 81054 478096
rect 80434 477776 81054 477860
rect 80434 477540 80466 477776
rect 80702 477540 80786 477776
rect 81022 477540 81054 477776
rect 80434 442096 81054 477540
rect 80434 441860 80466 442096
rect 80702 441860 80786 442096
rect 81022 441860 81054 442096
rect 80434 441776 81054 441860
rect 80434 441540 80466 441776
rect 80702 441540 80786 441776
rect 81022 441540 81054 441776
rect 80434 406096 81054 441540
rect 80434 405860 80466 406096
rect 80702 405860 80786 406096
rect 81022 405860 81054 406096
rect 80434 405776 81054 405860
rect 80434 405540 80466 405776
rect 80702 405540 80786 405776
rect 81022 405540 81054 405776
rect 80434 370096 81054 405540
rect 80434 369860 80466 370096
rect 80702 369860 80786 370096
rect 81022 369860 81054 370096
rect 80434 369776 81054 369860
rect 80434 369540 80466 369776
rect 80702 369540 80786 369776
rect 81022 369540 81054 369776
rect 80434 334096 81054 369540
rect 80434 333860 80466 334096
rect 80702 333860 80786 334096
rect 81022 333860 81054 334096
rect 80434 333776 81054 333860
rect 80434 333540 80466 333776
rect 80702 333540 80786 333776
rect 81022 333540 81054 333776
rect 80434 298096 81054 333540
rect 80434 297860 80466 298096
rect 80702 297860 80786 298096
rect 81022 297860 81054 298096
rect 80434 297776 81054 297860
rect 80434 297540 80466 297776
rect 80702 297540 80786 297776
rect 81022 297540 81054 297776
rect 80434 262096 81054 297540
rect 80434 261860 80466 262096
rect 80702 261860 80786 262096
rect 81022 261860 81054 262096
rect 80434 261776 81054 261860
rect 80434 261540 80466 261776
rect 80702 261540 80786 261776
rect 81022 261540 81054 261776
rect 80434 226096 81054 261540
rect 80434 225860 80466 226096
rect 80702 225860 80786 226096
rect 81022 225860 81054 226096
rect 80434 225776 81054 225860
rect 80434 225540 80466 225776
rect 80702 225540 80786 225776
rect 81022 225540 81054 225776
rect 80434 190096 81054 225540
rect 80434 189860 80466 190096
rect 80702 189860 80786 190096
rect 81022 189860 81054 190096
rect 80434 189776 81054 189860
rect 80434 189540 80466 189776
rect 80702 189540 80786 189776
rect 81022 189540 81054 189776
rect 80434 154096 81054 189540
rect 80434 153860 80466 154096
rect 80702 153860 80786 154096
rect 81022 153860 81054 154096
rect 80434 153776 81054 153860
rect 80434 153540 80466 153776
rect 80702 153540 80786 153776
rect 81022 153540 81054 153776
rect 80434 118096 81054 153540
rect 80434 117860 80466 118096
rect 80702 117860 80786 118096
rect 81022 117860 81054 118096
rect 80434 117776 81054 117860
rect 80434 117540 80466 117776
rect 80702 117540 80786 117776
rect 81022 117540 81054 117776
rect 80434 82096 81054 117540
rect 80434 81860 80466 82096
rect 80702 81860 80786 82096
rect 81022 81860 81054 82096
rect 80434 81776 81054 81860
rect 80434 81540 80466 81776
rect 80702 81540 80786 81776
rect 81022 81540 81054 81776
rect 80434 46096 81054 81540
rect 80434 45860 80466 46096
rect 80702 45860 80786 46096
rect 81022 45860 81054 46096
rect 80434 45776 81054 45860
rect 80434 45540 80466 45776
rect 80702 45540 80786 45776
rect 81022 45540 81054 45776
rect 80434 10096 81054 45540
rect 80434 9860 80466 10096
rect 80702 9860 80786 10096
rect 81022 9860 81054 10096
rect 80434 9776 81054 9860
rect 80434 9540 80466 9776
rect 80702 9540 80786 9776
rect 81022 9540 81054 9776
rect 80434 -6104 81054 9540
rect 80434 -6340 80466 -6104
rect 80702 -6340 80786 -6104
rect 81022 -6340 81054 -6104
rect 80434 -6424 81054 -6340
rect 80434 -6660 80466 -6424
rect 80702 -6660 80786 -6424
rect 81022 -6660 81054 -6424
rect 80434 -7652 81054 -6660
rect 81674 711560 82294 711592
rect 81674 711324 81706 711560
rect 81942 711324 82026 711560
rect 82262 711324 82294 711560
rect 81674 711240 82294 711324
rect 81674 711004 81706 711240
rect 81942 711004 82026 711240
rect 82262 711004 82294 711240
rect 81674 695336 82294 711004
rect 81674 695100 81706 695336
rect 81942 695100 82026 695336
rect 82262 695100 82294 695336
rect 81674 695016 82294 695100
rect 81674 694780 81706 695016
rect 81942 694780 82026 695016
rect 82262 694780 82294 695016
rect 81674 659336 82294 694780
rect 81674 659100 81706 659336
rect 81942 659100 82026 659336
rect 82262 659100 82294 659336
rect 81674 659016 82294 659100
rect 81674 658780 81706 659016
rect 81942 658780 82026 659016
rect 82262 658780 82294 659016
rect 81674 623336 82294 658780
rect 81674 623100 81706 623336
rect 81942 623100 82026 623336
rect 82262 623100 82294 623336
rect 81674 623016 82294 623100
rect 81674 622780 81706 623016
rect 81942 622780 82026 623016
rect 82262 622780 82294 623016
rect 81674 587336 82294 622780
rect 81674 587100 81706 587336
rect 81942 587100 82026 587336
rect 82262 587100 82294 587336
rect 81674 587016 82294 587100
rect 81674 586780 81706 587016
rect 81942 586780 82026 587016
rect 82262 586780 82294 587016
rect 81674 551336 82294 586780
rect 81674 551100 81706 551336
rect 81942 551100 82026 551336
rect 82262 551100 82294 551336
rect 81674 551016 82294 551100
rect 81674 550780 81706 551016
rect 81942 550780 82026 551016
rect 82262 550780 82294 551016
rect 81674 515336 82294 550780
rect 81674 515100 81706 515336
rect 81942 515100 82026 515336
rect 82262 515100 82294 515336
rect 81674 515016 82294 515100
rect 81674 514780 81706 515016
rect 81942 514780 82026 515016
rect 82262 514780 82294 515016
rect 81674 479336 82294 514780
rect 81674 479100 81706 479336
rect 81942 479100 82026 479336
rect 82262 479100 82294 479336
rect 81674 479016 82294 479100
rect 81674 478780 81706 479016
rect 81942 478780 82026 479016
rect 82262 478780 82294 479016
rect 81674 443336 82294 478780
rect 81674 443100 81706 443336
rect 81942 443100 82026 443336
rect 82262 443100 82294 443336
rect 81674 443016 82294 443100
rect 81674 442780 81706 443016
rect 81942 442780 82026 443016
rect 82262 442780 82294 443016
rect 81674 407336 82294 442780
rect 81674 407100 81706 407336
rect 81942 407100 82026 407336
rect 82262 407100 82294 407336
rect 81674 407016 82294 407100
rect 81674 406780 81706 407016
rect 81942 406780 82026 407016
rect 82262 406780 82294 407016
rect 81674 371336 82294 406780
rect 81674 371100 81706 371336
rect 81942 371100 82026 371336
rect 82262 371100 82294 371336
rect 81674 371016 82294 371100
rect 81674 370780 81706 371016
rect 81942 370780 82026 371016
rect 82262 370780 82294 371016
rect 81674 335336 82294 370780
rect 81674 335100 81706 335336
rect 81942 335100 82026 335336
rect 82262 335100 82294 335336
rect 81674 335016 82294 335100
rect 81674 334780 81706 335016
rect 81942 334780 82026 335016
rect 82262 334780 82294 335016
rect 81674 299336 82294 334780
rect 81674 299100 81706 299336
rect 81942 299100 82026 299336
rect 82262 299100 82294 299336
rect 81674 299016 82294 299100
rect 81674 298780 81706 299016
rect 81942 298780 82026 299016
rect 82262 298780 82294 299016
rect 81674 263336 82294 298780
rect 81674 263100 81706 263336
rect 81942 263100 82026 263336
rect 82262 263100 82294 263336
rect 81674 263016 82294 263100
rect 81674 262780 81706 263016
rect 81942 262780 82026 263016
rect 82262 262780 82294 263016
rect 81674 227336 82294 262780
rect 81674 227100 81706 227336
rect 81942 227100 82026 227336
rect 82262 227100 82294 227336
rect 81674 227016 82294 227100
rect 81674 226780 81706 227016
rect 81942 226780 82026 227016
rect 82262 226780 82294 227016
rect 81674 191336 82294 226780
rect 81674 191100 81706 191336
rect 81942 191100 82026 191336
rect 82262 191100 82294 191336
rect 81674 191016 82294 191100
rect 81674 190780 81706 191016
rect 81942 190780 82026 191016
rect 82262 190780 82294 191016
rect 81674 155336 82294 190780
rect 81674 155100 81706 155336
rect 81942 155100 82026 155336
rect 82262 155100 82294 155336
rect 81674 155016 82294 155100
rect 81674 154780 81706 155016
rect 81942 154780 82026 155016
rect 82262 154780 82294 155016
rect 81674 119336 82294 154780
rect 81674 119100 81706 119336
rect 81942 119100 82026 119336
rect 82262 119100 82294 119336
rect 81674 119016 82294 119100
rect 81674 118780 81706 119016
rect 81942 118780 82026 119016
rect 82262 118780 82294 119016
rect 81674 83336 82294 118780
rect 81674 83100 81706 83336
rect 81942 83100 82026 83336
rect 82262 83100 82294 83336
rect 81674 83016 82294 83100
rect 81674 82780 81706 83016
rect 81942 82780 82026 83016
rect 82262 82780 82294 83016
rect 81674 47336 82294 82780
rect 81674 47100 81706 47336
rect 81942 47100 82026 47336
rect 82262 47100 82294 47336
rect 81674 47016 82294 47100
rect 81674 46780 81706 47016
rect 81942 46780 82026 47016
rect 82262 46780 82294 47016
rect 81674 11336 82294 46780
rect 81674 11100 81706 11336
rect 81942 11100 82026 11336
rect 82262 11100 82294 11336
rect 81674 11016 82294 11100
rect 81674 10780 81706 11016
rect 81942 10780 82026 11016
rect 82262 10780 82294 11016
rect 81674 -7064 82294 10780
rect 81674 -7300 81706 -7064
rect 81942 -7300 82026 -7064
rect 82262 -7300 82294 -7064
rect 81674 -7384 82294 -7300
rect 81674 -7620 81706 -7384
rect 81942 -7620 82026 -7384
rect 82262 -7620 82294 -7384
rect 81674 -7652 82294 -7620
rect 108994 704840 109614 711592
rect 108994 704604 109026 704840
rect 109262 704604 109346 704840
rect 109582 704604 109614 704840
rect 108994 704520 109614 704604
rect 108994 704284 109026 704520
rect 109262 704284 109346 704520
rect 109582 704284 109614 704520
rect 108994 686656 109614 704284
rect 108994 686420 109026 686656
rect 109262 686420 109346 686656
rect 109582 686420 109614 686656
rect 108994 686336 109614 686420
rect 108994 686100 109026 686336
rect 109262 686100 109346 686336
rect 109582 686100 109614 686336
rect 108994 650656 109614 686100
rect 108994 650420 109026 650656
rect 109262 650420 109346 650656
rect 109582 650420 109614 650656
rect 108994 650336 109614 650420
rect 108994 650100 109026 650336
rect 109262 650100 109346 650336
rect 109582 650100 109614 650336
rect 108994 614656 109614 650100
rect 108994 614420 109026 614656
rect 109262 614420 109346 614656
rect 109582 614420 109614 614656
rect 108994 614336 109614 614420
rect 108994 614100 109026 614336
rect 109262 614100 109346 614336
rect 109582 614100 109614 614336
rect 108994 578656 109614 614100
rect 108994 578420 109026 578656
rect 109262 578420 109346 578656
rect 109582 578420 109614 578656
rect 108994 578336 109614 578420
rect 108994 578100 109026 578336
rect 109262 578100 109346 578336
rect 109582 578100 109614 578336
rect 108994 542656 109614 578100
rect 108994 542420 109026 542656
rect 109262 542420 109346 542656
rect 109582 542420 109614 542656
rect 108994 542336 109614 542420
rect 108994 542100 109026 542336
rect 109262 542100 109346 542336
rect 109582 542100 109614 542336
rect 108994 506656 109614 542100
rect 108994 506420 109026 506656
rect 109262 506420 109346 506656
rect 109582 506420 109614 506656
rect 108994 506336 109614 506420
rect 108994 506100 109026 506336
rect 109262 506100 109346 506336
rect 109582 506100 109614 506336
rect 108994 470656 109614 506100
rect 108994 470420 109026 470656
rect 109262 470420 109346 470656
rect 109582 470420 109614 470656
rect 108994 470336 109614 470420
rect 108994 470100 109026 470336
rect 109262 470100 109346 470336
rect 109582 470100 109614 470336
rect 108994 434656 109614 470100
rect 108994 434420 109026 434656
rect 109262 434420 109346 434656
rect 109582 434420 109614 434656
rect 108994 434336 109614 434420
rect 108994 434100 109026 434336
rect 109262 434100 109346 434336
rect 109582 434100 109614 434336
rect 108994 398656 109614 434100
rect 108994 398420 109026 398656
rect 109262 398420 109346 398656
rect 109582 398420 109614 398656
rect 108994 398336 109614 398420
rect 108994 398100 109026 398336
rect 109262 398100 109346 398336
rect 109582 398100 109614 398336
rect 108994 362656 109614 398100
rect 108994 362420 109026 362656
rect 109262 362420 109346 362656
rect 109582 362420 109614 362656
rect 108994 362336 109614 362420
rect 108994 362100 109026 362336
rect 109262 362100 109346 362336
rect 109582 362100 109614 362336
rect 108994 326656 109614 362100
rect 108994 326420 109026 326656
rect 109262 326420 109346 326656
rect 109582 326420 109614 326656
rect 108994 326336 109614 326420
rect 108994 326100 109026 326336
rect 109262 326100 109346 326336
rect 109582 326100 109614 326336
rect 108994 290656 109614 326100
rect 108994 290420 109026 290656
rect 109262 290420 109346 290656
rect 109582 290420 109614 290656
rect 108994 290336 109614 290420
rect 108994 290100 109026 290336
rect 109262 290100 109346 290336
rect 109582 290100 109614 290336
rect 108994 254656 109614 290100
rect 108994 254420 109026 254656
rect 109262 254420 109346 254656
rect 109582 254420 109614 254656
rect 108994 254336 109614 254420
rect 108994 254100 109026 254336
rect 109262 254100 109346 254336
rect 109582 254100 109614 254336
rect 108994 218656 109614 254100
rect 108994 218420 109026 218656
rect 109262 218420 109346 218656
rect 109582 218420 109614 218656
rect 108994 218336 109614 218420
rect 108994 218100 109026 218336
rect 109262 218100 109346 218336
rect 109582 218100 109614 218336
rect 108994 182656 109614 218100
rect 108994 182420 109026 182656
rect 109262 182420 109346 182656
rect 109582 182420 109614 182656
rect 108994 182336 109614 182420
rect 108994 182100 109026 182336
rect 109262 182100 109346 182336
rect 109582 182100 109614 182336
rect 108994 146656 109614 182100
rect 108994 146420 109026 146656
rect 109262 146420 109346 146656
rect 109582 146420 109614 146656
rect 108994 146336 109614 146420
rect 108994 146100 109026 146336
rect 109262 146100 109346 146336
rect 109582 146100 109614 146336
rect 108994 110656 109614 146100
rect 108994 110420 109026 110656
rect 109262 110420 109346 110656
rect 109582 110420 109614 110656
rect 108994 110336 109614 110420
rect 108994 110100 109026 110336
rect 109262 110100 109346 110336
rect 109582 110100 109614 110336
rect 108994 74656 109614 110100
rect 108994 74420 109026 74656
rect 109262 74420 109346 74656
rect 109582 74420 109614 74656
rect 108994 74336 109614 74420
rect 108994 74100 109026 74336
rect 109262 74100 109346 74336
rect 109582 74100 109614 74336
rect 108994 38656 109614 74100
rect 108994 38420 109026 38656
rect 109262 38420 109346 38656
rect 109582 38420 109614 38656
rect 108994 38336 109614 38420
rect 108994 38100 109026 38336
rect 109262 38100 109346 38336
rect 109582 38100 109614 38336
rect 108994 2656 109614 38100
rect 108994 2420 109026 2656
rect 109262 2420 109346 2656
rect 109582 2420 109614 2656
rect 108994 2336 109614 2420
rect 108994 2100 109026 2336
rect 109262 2100 109346 2336
rect 109582 2100 109614 2336
rect 108994 -344 109614 2100
rect 108994 -580 109026 -344
rect 109262 -580 109346 -344
rect 109582 -580 109614 -344
rect 108994 -664 109614 -580
rect 108994 -900 109026 -664
rect 109262 -900 109346 -664
rect 109582 -900 109614 -664
rect 108994 -7652 109614 -900
rect 110234 705800 110854 711592
rect 110234 705564 110266 705800
rect 110502 705564 110586 705800
rect 110822 705564 110854 705800
rect 110234 705480 110854 705564
rect 110234 705244 110266 705480
rect 110502 705244 110586 705480
rect 110822 705244 110854 705480
rect 110234 687896 110854 705244
rect 110234 687660 110266 687896
rect 110502 687660 110586 687896
rect 110822 687660 110854 687896
rect 110234 687576 110854 687660
rect 110234 687340 110266 687576
rect 110502 687340 110586 687576
rect 110822 687340 110854 687576
rect 110234 651896 110854 687340
rect 110234 651660 110266 651896
rect 110502 651660 110586 651896
rect 110822 651660 110854 651896
rect 110234 651576 110854 651660
rect 110234 651340 110266 651576
rect 110502 651340 110586 651576
rect 110822 651340 110854 651576
rect 110234 615896 110854 651340
rect 110234 615660 110266 615896
rect 110502 615660 110586 615896
rect 110822 615660 110854 615896
rect 110234 615576 110854 615660
rect 110234 615340 110266 615576
rect 110502 615340 110586 615576
rect 110822 615340 110854 615576
rect 110234 579896 110854 615340
rect 110234 579660 110266 579896
rect 110502 579660 110586 579896
rect 110822 579660 110854 579896
rect 110234 579576 110854 579660
rect 110234 579340 110266 579576
rect 110502 579340 110586 579576
rect 110822 579340 110854 579576
rect 110234 543896 110854 579340
rect 110234 543660 110266 543896
rect 110502 543660 110586 543896
rect 110822 543660 110854 543896
rect 110234 543576 110854 543660
rect 110234 543340 110266 543576
rect 110502 543340 110586 543576
rect 110822 543340 110854 543576
rect 110234 507896 110854 543340
rect 110234 507660 110266 507896
rect 110502 507660 110586 507896
rect 110822 507660 110854 507896
rect 110234 507576 110854 507660
rect 110234 507340 110266 507576
rect 110502 507340 110586 507576
rect 110822 507340 110854 507576
rect 110234 471896 110854 507340
rect 110234 471660 110266 471896
rect 110502 471660 110586 471896
rect 110822 471660 110854 471896
rect 110234 471576 110854 471660
rect 110234 471340 110266 471576
rect 110502 471340 110586 471576
rect 110822 471340 110854 471576
rect 110234 435896 110854 471340
rect 110234 435660 110266 435896
rect 110502 435660 110586 435896
rect 110822 435660 110854 435896
rect 110234 435576 110854 435660
rect 110234 435340 110266 435576
rect 110502 435340 110586 435576
rect 110822 435340 110854 435576
rect 110234 399896 110854 435340
rect 110234 399660 110266 399896
rect 110502 399660 110586 399896
rect 110822 399660 110854 399896
rect 110234 399576 110854 399660
rect 110234 399340 110266 399576
rect 110502 399340 110586 399576
rect 110822 399340 110854 399576
rect 110234 363896 110854 399340
rect 110234 363660 110266 363896
rect 110502 363660 110586 363896
rect 110822 363660 110854 363896
rect 110234 363576 110854 363660
rect 110234 363340 110266 363576
rect 110502 363340 110586 363576
rect 110822 363340 110854 363576
rect 110234 327896 110854 363340
rect 110234 327660 110266 327896
rect 110502 327660 110586 327896
rect 110822 327660 110854 327896
rect 110234 327576 110854 327660
rect 110234 327340 110266 327576
rect 110502 327340 110586 327576
rect 110822 327340 110854 327576
rect 110234 291896 110854 327340
rect 110234 291660 110266 291896
rect 110502 291660 110586 291896
rect 110822 291660 110854 291896
rect 110234 291576 110854 291660
rect 110234 291340 110266 291576
rect 110502 291340 110586 291576
rect 110822 291340 110854 291576
rect 110234 255896 110854 291340
rect 110234 255660 110266 255896
rect 110502 255660 110586 255896
rect 110822 255660 110854 255896
rect 110234 255576 110854 255660
rect 110234 255340 110266 255576
rect 110502 255340 110586 255576
rect 110822 255340 110854 255576
rect 110234 219896 110854 255340
rect 110234 219660 110266 219896
rect 110502 219660 110586 219896
rect 110822 219660 110854 219896
rect 110234 219576 110854 219660
rect 110234 219340 110266 219576
rect 110502 219340 110586 219576
rect 110822 219340 110854 219576
rect 110234 183896 110854 219340
rect 110234 183660 110266 183896
rect 110502 183660 110586 183896
rect 110822 183660 110854 183896
rect 110234 183576 110854 183660
rect 110234 183340 110266 183576
rect 110502 183340 110586 183576
rect 110822 183340 110854 183576
rect 110234 147896 110854 183340
rect 110234 147660 110266 147896
rect 110502 147660 110586 147896
rect 110822 147660 110854 147896
rect 110234 147576 110854 147660
rect 110234 147340 110266 147576
rect 110502 147340 110586 147576
rect 110822 147340 110854 147576
rect 110234 111896 110854 147340
rect 110234 111660 110266 111896
rect 110502 111660 110586 111896
rect 110822 111660 110854 111896
rect 110234 111576 110854 111660
rect 110234 111340 110266 111576
rect 110502 111340 110586 111576
rect 110822 111340 110854 111576
rect 110234 75896 110854 111340
rect 110234 75660 110266 75896
rect 110502 75660 110586 75896
rect 110822 75660 110854 75896
rect 110234 75576 110854 75660
rect 110234 75340 110266 75576
rect 110502 75340 110586 75576
rect 110822 75340 110854 75576
rect 110234 39896 110854 75340
rect 110234 39660 110266 39896
rect 110502 39660 110586 39896
rect 110822 39660 110854 39896
rect 110234 39576 110854 39660
rect 110234 39340 110266 39576
rect 110502 39340 110586 39576
rect 110822 39340 110854 39576
rect 110234 3896 110854 39340
rect 110234 3660 110266 3896
rect 110502 3660 110586 3896
rect 110822 3660 110854 3896
rect 110234 3576 110854 3660
rect 110234 3340 110266 3576
rect 110502 3340 110586 3576
rect 110822 3340 110854 3576
rect 110234 -1304 110854 3340
rect 110234 -1540 110266 -1304
rect 110502 -1540 110586 -1304
rect 110822 -1540 110854 -1304
rect 110234 -1624 110854 -1540
rect 110234 -1860 110266 -1624
rect 110502 -1860 110586 -1624
rect 110822 -1860 110854 -1624
rect 110234 -7652 110854 -1860
rect 111474 706760 112094 711592
rect 111474 706524 111506 706760
rect 111742 706524 111826 706760
rect 112062 706524 112094 706760
rect 111474 706440 112094 706524
rect 111474 706204 111506 706440
rect 111742 706204 111826 706440
rect 112062 706204 112094 706440
rect 111474 689136 112094 706204
rect 111474 688900 111506 689136
rect 111742 688900 111826 689136
rect 112062 688900 112094 689136
rect 111474 688816 112094 688900
rect 111474 688580 111506 688816
rect 111742 688580 111826 688816
rect 112062 688580 112094 688816
rect 111474 653136 112094 688580
rect 111474 652900 111506 653136
rect 111742 652900 111826 653136
rect 112062 652900 112094 653136
rect 111474 652816 112094 652900
rect 111474 652580 111506 652816
rect 111742 652580 111826 652816
rect 112062 652580 112094 652816
rect 111474 617136 112094 652580
rect 111474 616900 111506 617136
rect 111742 616900 111826 617136
rect 112062 616900 112094 617136
rect 111474 616816 112094 616900
rect 111474 616580 111506 616816
rect 111742 616580 111826 616816
rect 112062 616580 112094 616816
rect 111474 581136 112094 616580
rect 111474 580900 111506 581136
rect 111742 580900 111826 581136
rect 112062 580900 112094 581136
rect 111474 580816 112094 580900
rect 111474 580580 111506 580816
rect 111742 580580 111826 580816
rect 112062 580580 112094 580816
rect 111474 545136 112094 580580
rect 111474 544900 111506 545136
rect 111742 544900 111826 545136
rect 112062 544900 112094 545136
rect 111474 544816 112094 544900
rect 111474 544580 111506 544816
rect 111742 544580 111826 544816
rect 112062 544580 112094 544816
rect 111474 509136 112094 544580
rect 111474 508900 111506 509136
rect 111742 508900 111826 509136
rect 112062 508900 112094 509136
rect 111474 508816 112094 508900
rect 111474 508580 111506 508816
rect 111742 508580 111826 508816
rect 112062 508580 112094 508816
rect 111474 473136 112094 508580
rect 111474 472900 111506 473136
rect 111742 472900 111826 473136
rect 112062 472900 112094 473136
rect 111474 472816 112094 472900
rect 111474 472580 111506 472816
rect 111742 472580 111826 472816
rect 112062 472580 112094 472816
rect 111474 437136 112094 472580
rect 111474 436900 111506 437136
rect 111742 436900 111826 437136
rect 112062 436900 112094 437136
rect 111474 436816 112094 436900
rect 111474 436580 111506 436816
rect 111742 436580 111826 436816
rect 112062 436580 112094 436816
rect 111474 401136 112094 436580
rect 111474 400900 111506 401136
rect 111742 400900 111826 401136
rect 112062 400900 112094 401136
rect 111474 400816 112094 400900
rect 111474 400580 111506 400816
rect 111742 400580 111826 400816
rect 112062 400580 112094 400816
rect 111474 365136 112094 400580
rect 111474 364900 111506 365136
rect 111742 364900 111826 365136
rect 112062 364900 112094 365136
rect 111474 364816 112094 364900
rect 111474 364580 111506 364816
rect 111742 364580 111826 364816
rect 112062 364580 112094 364816
rect 111474 329136 112094 364580
rect 111474 328900 111506 329136
rect 111742 328900 111826 329136
rect 112062 328900 112094 329136
rect 111474 328816 112094 328900
rect 111474 328580 111506 328816
rect 111742 328580 111826 328816
rect 112062 328580 112094 328816
rect 111474 293136 112094 328580
rect 111474 292900 111506 293136
rect 111742 292900 111826 293136
rect 112062 292900 112094 293136
rect 111474 292816 112094 292900
rect 111474 292580 111506 292816
rect 111742 292580 111826 292816
rect 112062 292580 112094 292816
rect 111474 257136 112094 292580
rect 111474 256900 111506 257136
rect 111742 256900 111826 257136
rect 112062 256900 112094 257136
rect 111474 256816 112094 256900
rect 111474 256580 111506 256816
rect 111742 256580 111826 256816
rect 112062 256580 112094 256816
rect 111474 221136 112094 256580
rect 111474 220900 111506 221136
rect 111742 220900 111826 221136
rect 112062 220900 112094 221136
rect 111474 220816 112094 220900
rect 111474 220580 111506 220816
rect 111742 220580 111826 220816
rect 112062 220580 112094 220816
rect 111474 185136 112094 220580
rect 111474 184900 111506 185136
rect 111742 184900 111826 185136
rect 112062 184900 112094 185136
rect 111474 184816 112094 184900
rect 111474 184580 111506 184816
rect 111742 184580 111826 184816
rect 112062 184580 112094 184816
rect 111474 149136 112094 184580
rect 111474 148900 111506 149136
rect 111742 148900 111826 149136
rect 112062 148900 112094 149136
rect 111474 148816 112094 148900
rect 111474 148580 111506 148816
rect 111742 148580 111826 148816
rect 112062 148580 112094 148816
rect 111474 113136 112094 148580
rect 111474 112900 111506 113136
rect 111742 112900 111826 113136
rect 112062 112900 112094 113136
rect 111474 112816 112094 112900
rect 111474 112580 111506 112816
rect 111742 112580 111826 112816
rect 112062 112580 112094 112816
rect 111474 77136 112094 112580
rect 111474 76900 111506 77136
rect 111742 76900 111826 77136
rect 112062 76900 112094 77136
rect 111474 76816 112094 76900
rect 111474 76580 111506 76816
rect 111742 76580 111826 76816
rect 112062 76580 112094 76816
rect 111474 41136 112094 76580
rect 111474 40900 111506 41136
rect 111742 40900 111826 41136
rect 112062 40900 112094 41136
rect 111474 40816 112094 40900
rect 111474 40580 111506 40816
rect 111742 40580 111826 40816
rect 112062 40580 112094 40816
rect 111474 5136 112094 40580
rect 111474 4900 111506 5136
rect 111742 4900 111826 5136
rect 112062 4900 112094 5136
rect 111474 4816 112094 4900
rect 111474 4580 111506 4816
rect 111742 4580 111826 4816
rect 112062 4580 112094 4816
rect 111474 -2264 112094 4580
rect 111474 -2500 111506 -2264
rect 111742 -2500 111826 -2264
rect 112062 -2500 112094 -2264
rect 111474 -2584 112094 -2500
rect 111474 -2820 111506 -2584
rect 111742 -2820 111826 -2584
rect 112062 -2820 112094 -2584
rect 111474 -7652 112094 -2820
rect 112714 707720 113334 711592
rect 112714 707484 112746 707720
rect 112982 707484 113066 707720
rect 113302 707484 113334 707720
rect 112714 707400 113334 707484
rect 112714 707164 112746 707400
rect 112982 707164 113066 707400
rect 113302 707164 113334 707400
rect 112714 690376 113334 707164
rect 112714 690140 112746 690376
rect 112982 690140 113066 690376
rect 113302 690140 113334 690376
rect 112714 690056 113334 690140
rect 112714 689820 112746 690056
rect 112982 689820 113066 690056
rect 113302 689820 113334 690056
rect 112714 654376 113334 689820
rect 112714 654140 112746 654376
rect 112982 654140 113066 654376
rect 113302 654140 113334 654376
rect 112714 654056 113334 654140
rect 112714 653820 112746 654056
rect 112982 653820 113066 654056
rect 113302 653820 113334 654056
rect 112714 618376 113334 653820
rect 112714 618140 112746 618376
rect 112982 618140 113066 618376
rect 113302 618140 113334 618376
rect 112714 618056 113334 618140
rect 112714 617820 112746 618056
rect 112982 617820 113066 618056
rect 113302 617820 113334 618056
rect 112714 582376 113334 617820
rect 112714 582140 112746 582376
rect 112982 582140 113066 582376
rect 113302 582140 113334 582376
rect 112714 582056 113334 582140
rect 112714 581820 112746 582056
rect 112982 581820 113066 582056
rect 113302 581820 113334 582056
rect 112714 546376 113334 581820
rect 112714 546140 112746 546376
rect 112982 546140 113066 546376
rect 113302 546140 113334 546376
rect 112714 546056 113334 546140
rect 112714 545820 112746 546056
rect 112982 545820 113066 546056
rect 113302 545820 113334 546056
rect 112714 510376 113334 545820
rect 112714 510140 112746 510376
rect 112982 510140 113066 510376
rect 113302 510140 113334 510376
rect 112714 510056 113334 510140
rect 112714 509820 112746 510056
rect 112982 509820 113066 510056
rect 113302 509820 113334 510056
rect 112714 474376 113334 509820
rect 112714 474140 112746 474376
rect 112982 474140 113066 474376
rect 113302 474140 113334 474376
rect 112714 474056 113334 474140
rect 112714 473820 112746 474056
rect 112982 473820 113066 474056
rect 113302 473820 113334 474056
rect 112714 438376 113334 473820
rect 112714 438140 112746 438376
rect 112982 438140 113066 438376
rect 113302 438140 113334 438376
rect 112714 438056 113334 438140
rect 112714 437820 112746 438056
rect 112982 437820 113066 438056
rect 113302 437820 113334 438056
rect 112714 402376 113334 437820
rect 112714 402140 112746 402376
rect 112982 402140 113066 402376
rect 113302 402140 113334 402376
rect 112714 402056 113334 402140
rect 112714 401820 112746 402056
rect 112982 401820 113066 402056
rect 113302 401820 113334 402056
rect 112714 366376 113334 401820
rect 112714 366140 112746 366376
rect 112982 366140 113066 366376
rect 113302 366140 113334 366376
rect 112714 366056 113334 366140
rect 112714 365820 112746 366056
rect 112982 365820 113066 366056
rect 113302 365820 113334 366056
rect 112714 330376 113334 365820
rect 112714 330140 112746 330376
rect 112982 330140 113066 330376
rect 113302 330140 113334 330376
rect 112714 330056 113334 330140
rect 112714 329820 112746 330056
rect 112982 329820 113066 330056
rect 113302 329820 113334 330056
rect 112714 294376 113334 329820
rect 112714 294140 112746 294376
rect 112982 294140 113066 294376
rect 113302 294140 113334 294376
rect 112714 294056 113334 294140
rect 112714 293820 112746 294056
rect 112982 293820 113066 294056
rect 113302 293820 113334 294056
rect 112714 258376 113334 293820
rect 112714 258140 112746 258376
rect 112982 258140 113066 258376
rect 113302 258140 113334 258376
rect 112714 258056 113334 258140
rect 112714 257820 112746 258056
rect 112982 257820 113066 258056
rect 113302 257820 113334 258056
rect 112714 222376 113334 257820
rect 112714 222140 112746 222376
rect 112982 222140 113066 222376
rect 113302 222140 113334 222376
rect 112714 222056 113334 222140
rect 112714 221820 112746 222056
rect 112982 221820 113066 222056
rect 113302 221820 113334 222056
rect 112714 186376 113334 221820
rect 112714 186140 112746 186376
rect 112982 186140 113066 186376
rect 113302 186140 113334 186376
rect 112714 186056 113334 186140
rect 112714 185820 112746 186056
rect 112982 185820 113066 186056
rect 113302 185820 113334 186056
rect 112714 150376 113334 185820
rect 112714 150140 112746 150376
rect 112982 150140 113066 150376
rect 113302 150140 113334 150376
rect 112714 150056 113334 150140
rect 112714 149820 112746 150056
rect 112982 149820 113066 150056
rect 113302 149820 113334 150056
rect 112714 114376 113334 149820
rect 112714 114140 112746 114376
rect 112982 114140 113066 114376
rect 113302 114140 113334 114376
rect 112714 114056 113334 114140
rect 112714 113820 112746 114056
rect 112982 113820 113066 114056
rect 113302 113820 113334 114056
rect 112714 78376 113334 113820
rect 112714 78140 112746 78376
rect 112982 78140 113066 78376
rect 113302 78140 113334 78376
rect 112714 78056 113334 78140
rect 112714 77820 112746 78056
rect 112982 77820 113066 78056
rect 113302 77820 113334 78056
rect 112714 42376 113334 77820
rect 112714 42140 112746 42376
rect 112982 42140 113066 42376
rect 113302 42140 113334 42376
rect 112714 42056 113334 42140
rect 112714 41820 112746 42056
rect 112982 41820 113066 42056
rect 113302 41820 113334 42056
rect 112714 6376 113334 41820
rect 112714 6140 112746 6376
rect 112982 6140 113066 6376
rect 113302 6140 113334 6376
rect 112714 6056 113334 6140
rect 112714 5820 112746 6056
rect 112982 5820 113066 6056
rect 113302 5820 113334 6056
rect 112714 -3224 113334 5820
rect 112714 -3460 112746 -3224
rect 112982 -3460 113066 -3224
rect 113302 -3460 113334 -3224
rect 112714 -3544 113334 -3460
rect 112714 -3780 112746 -3544
rect 112982 -3780 113066 -3544
rect 113302 -3780 113334 -3544
rect 112714 -7652 113334 -3780
rect 113954 708680 114574 711592
rect 113954 708444 113986 708680
rect 114222 708444 114306 708680
rect 114542 708444 114574 708680
rect 113954 708360 114574 708444
rect 113954 708124 113986 708360
rect 114222 708124 114306 708360
rect 114542 708124 114574 708360
rect 113954 691616 114574 708124
rect 113954 691380 113986 691616
rect 114222 691380 114306 691616
rect 114542 691380 114574 691616
rect 113954 691296 114574 691380
rect 113954 691060 113986 691296
rect 114222 691060 114306 691296
rect 114542 691060 114574 691296
rect 113954 655616 114574 691060
rect 113954 655380 113986 655616
rect 114222 655380 114306 655616
rect 114542 655380 114574 655616
rect 113954 655296 114574 655380
rect 113954 655060 113986 655296
rect 114222 655060 114306 655296
rect 114542 655060 114574 655296
rect 113954 619616 114574 655060
rect 113954 619380 113986 619616
rect 114222 619380 114306 619616
rect 114542 619380 114574 619616
rect 113954 619296 114574 619380
rect 113954 619060 113986 619296
rect 114222 619060 114306 619296
rect 114542 619060 114574 619296
rect 113954 583616 114574 619060
rect 113954 583380 113986 583616
rect 114222 583380 114306 583616
rect 114542 583380 114574 583616
rect 113954 583296 114574 583380
rect 113954 583060 113986 583296
rect 114222 583060 114306 583296
rect 114542 583060 114574 583296
rect 113954 547616 114574 583060
rect 113954 547380 113986 547616
rect 114222 547380 114306 547616
rect 114542 547380 114574 547616
rect 113954 547296 114574 547380
rect 113954 547060 113986 547296
rect 114222 547060 114306 547296
rect 114542 547060 114574 547296
rect 113954 511616 114574 547060
rect 113954 511380 113986 511616
rect 114222 511380 114306 511616
rect 114542 511380 114574 511616
rect 113954 511296 114574 511380
rect 113954 511060 113986 511296
rect 114222 511060 114306 511296
rect 114542 511060 114574 511296
rect 113954 475616 114574 511060
rect 113954 475380 113986 475616
rect 114222 475380 114306 475616
rect 114542 475380 114574 475616
rect 113954 475296 114574 475380
rect 113954 475060 113986 475296
rect 114222 475060 114306 475296
rect 114542 475060 114574 475296
rect 113954 439616 114574 475060
rect 113954 439380 113986 439616
rect 114222 439380 114306 439616
rect 114542 439380 114574 439616
rect 113954 439296 114574 439380
rect 113954 439060 113986 439296
rect 114222 439060 114306 439296
rect 114542 439060 114574 439296
rect 113954 403616 114574 439060
rect 113954 403380 113986 403616
rect 114222 403380 114306 403616
rect 114542 403380 114574 403616
rect 113954 403296 114574 403380
rect 113954 403060 113986 403296
rect 114222 403060 114306 403296
rect 114542 403060 114574 403296
rect 113954 367616 114574 403060
rect 113954 367380 113986 367616
rect 114222 367380 114306 367616
rect 114542 367380 114574 367616
rect 113954 367296 114574 367380
rect 113954 367060 113986 367296
rect 114222 367060 114306 367296
rect 114542 367060 114574 367296
rect 113954 331616 114574 367060
rect 113954 331380 113986 331616
rect 114222 331380 114306 331616
rect 114542 331380 114574 331616
rect 113954 331296 114574 331380
rect 113954 331060 113986 331296
rect 114222 331060 114306 331296
rect 114542 331060 114574 331296
rect 113954 295616 114574 331060
rect 113954 295380 113986 295616
rect 114222 295380 114306 295616
rect 114542 295380 114574 295616
rect 113954 295296 114574 295380
rect 113954 295060 113986 295296
rect 114222 295060 114306 295296
rect 114542 295060 114574 295296
rect 113954 259616 114574 295060
rect 113954 259380 113986 259616
rect 114222 259380 114306 259616
rect 114542 259380 114574 259616
rect 113954 259296 114574 259380
rect 113954 259060 113986 259296
rect 114222 259060 114306 259296
rect 114542 259060 114574 259296
rect 113954 223616 114574 259060
rect 113954 223380 113986 223616
rect 114222 223380 114306 223616
rect 114542 223380 114574 223616
rect 113954 223296 114574 223380
rect 113954 223060 113986 223296
rect 114222 223060 114306 223296
rect 114542 223060 114574 223296
rect 113954 187616 114574 223060
rect 113954 187380 113986 187616
rect 114222 187380 114306 187616
rect 114542 187380 114574 187616
rect 113954 187296 114574 187380
rect 113954 187060 113986 187296
rect 114222 187060 114306 187296
rect 114542 187060 114574 187296
rect 113954 151616 114574 187060
rect 113954 151380 113986 151616
rect 114222 151380 114306 151616
rect 114542 151380 114574 151616
rect 113954 151296 114574 151380
rect 113954 151060 113986 151296
rect 114222 151060 114306 151296
rect 114542 151060 114574 151296
rect 113954 115616 114574 151060
rect 113954 115380 113986 115616
rect 114222 115380 114306 115616
rect 114542 115380 114574 115616
rect 113954 115296 114574 115380
rect 113954 115060 113986 115296
rect 114222 115060 114306 115296
rect 114542 115060 114574 115296
rect 113954 79616 114574 115060
rect 113954 79380 113986 79616
rect 114222 79380 114306 79616
rect 114542 79380 114574 79616
rect 113954 79296 114574 79380
rect 113954 79060 113986 79296
rect 114222 79060 114306 79296
rect 114542 79060 114574 79296
rect 113954 43616 114574 79060
rect 113954 43380 113986 43616
rect 114222 43380 114306 43616
rect 114542 43380 114574 43616
rect 113954 43296 114574 43380
rect 113954 43060 113986 43296
rect 114222 43060 114306 43296
rect 114542 43060 114574 43296
rect 113954 7616 114574 43060
rect 113954 7380 113986 7616
rect 114222 7380 114306 7616
rect 114542 7380 114574 7616
rect 113954 7296 114574 7380
rect 113954 7060 113986 7296
rect 114222 7060 114306 7296
rect 114542 7060 114574 7296
rect 113954 -4184 114574 7060
rect 113954 -4420 113986 -4184
rect 114222 -4420 114306 -4184
rect 114542 -4420 114574 -4184
rect 113954 -4504 114574 -4420
rect 113954 -4740 113986 -4504
rect 114222 -4740 114306 -4504
rect 114542 -4740 114574 -4504
rect 113954 -7652 114574 -4740
rect 115194 709640 115814 711592
rect 115194 709404 115226 709640
rect 115462 709404 115546 709640
rect 115782 709404 115814 709640
rect 115194 709320 115814 709404
rect 115194 709084 115226 709320
rect 115462 709084 115546 709320
rect 115782 709084 115814 709320
rect 115194 692856 115814 709084
rect 115194 692620 115226 692856
rect 115462 692620 115546 692856
rect 115782 692620 115814 692856
rect 115194 692536 115814 692620
rect 115194 692300 115226 692536
rect 115462 692300 115546 692536
rect 115782 692300 115814 692536
rect 115194 656856 115814 692300
rect 115194 656620 115226 656856
rect 115462 656620 115546 656856
rect 115782 656620 115814 656856
rect 115194 656536 115814 656620
rect 115194 656300 115226 656536
rect 115462 656300 115546 656536
rect 115782 656300 115814 656536
rect 115194 620856 115814 656300
rect 115194 620620 115226 620856
rect 115462 620620 115546 620856
rect 115782 620620 115814 620856
rect 115194 620536 115814 620620
rect 115194 620300 115226 620536
rect 115462 620300 115546 620536
rect 115782 620300 115814 620536
rect 115194 584856 115814 620300
rect 115194 584620 115226 584856
rect 115462 584620 115546 584856
rect 115782 584620 115814 584856
rect 115194 584536 115814 584620
rect 115194 584300 115226 584536
rect 115462 584300 115546 584536
rect 115782 584300 115814 584536
rect 115194 548856 115814 584300
rect 115194 548620 115226 548856
rect 115462 548620 115546 548856
rect 115782 548620 115814 548856
rect 115194 548536 115814 548620
rect 115194 548300 115226 548536
rect 115462 548300 115546 548536
rect 115782 548300 115814 548536
rect 115194 512856 115814 548300
rect 115194 512620 115226 512856
rect 115462 512620 115546 512856
rect 115782 512620 115814 512856
rect 115194 512536 115814 512620
rect 115194 512300 115226 512536
rect 115462 512300 115546 512536
rect 115782 512300 115814 512536
rect 115194 476856 115814 512300
rect 115194 476620 115226 476856
rect 115462 476620 115546 476856
rect 115782 476620 115814 476856
rect 115194 476536 115814 476620
rect 115194 476300 115226 476536
rect 115462 476300 115546 476536
rect 115782 476300 115814 476536
rect 115194 440856 115814 476300
rect 115194 440620 115226 440856
rect 115462 440620 115546 440856
rect 115782 440620 115814 440856
rect 115194 440536 115814 440620
rect 115194 440300 115226 440536
rect 115462 440300 115546 440536
rect 115782 440300 115814 440536
rect 115194 404856 115814 440300
rect 115194 404620 115226 404856
rect 115462 404620 115546 404856
rect 115782 404620 115814 404856
rect 115194 404536 115814 404620
rect 115194 404300 115226 404536
rect 115462 404300 115546 404536
rect 115782 404300 115814 404536
rect 115194 368856 115814 404300
rect 115194 368620 115226 368856
rect 115462 368620 115546 368856
rect 115782 368620 115814 368856
rect 115194 368536 115814 368620
rect 115194 368300 115226 368536
rect 115462 368300 115546 368536
rect 115782 368300 115814 368536
rect 115194 332856 115814 368300
rect 115194 332620 115226 332856
rect 115462 332620 115546 332856
rect 115782 332620 115814 332856
rect 115194 332536 115814 332620
rect 115194 332300 115226 332536
rect 115462 332300 115546 332536
rect 115782 332300 115814 332536
rect 115194 296856 115814 332300
rect 115194 296620 115226 296856
rect 115462 296620 115546 296856
rect 115782 296620 115814 296856
rect 115194 296536 115814 296620
rect 115194 296300 115226 296536
rect 115462 296300 115546 296536
rect 115782 296300 115814 296536
rect 115194 260856 115814 296300
rect 115194 260620 115226 260856
rect 115462 260620 115546 260856
rect 115782 260620 115814 260856
rect 115194 260536 115814 260620
rect 115194 260300 115226 260536
rect 115462 260300 115546 260536
rect 115782 260300 115814 260536
rect 115194 224856 115814 260300
rect 115194 224620 115226 224856
rect 115462 224620 115546 224856
rect 115782 224620 115814 224856
rect 115194 224536 115814 224620
rect 115194 224300 115226 224536
rect 115462 224300 115546 224536
rect 115782 224300 115814 224536
rect 115194 188856 115814 224300
rect 115194 188620 115226 188856
rect 115462 188620 115546 188856
rect 115782 188620 115814 188856
rect 115194 188536 115814 188620
rect 115194 188300 115226 188536
rect 115462 188300 115546 188536
rect 115782 188300 115814 188536
rect 115194 152856 115814 188300
rect 115194 152620 115226 152856
rect 115462 152620 115546 152856
rect 115782 152620 115814 152856
rect 115194 152536 115814 152620
rect 115194 152300 115226 152536
rect 115462 152300 115546 152536
rect 115782 152300 115814 152536
rect 115194 116856 115814 152300
rect 115194 116620 115226 116856
rect 115462 116620 115546 116856
rect 115782 116620 115814 116856
rect 115194 116536 115814 116620
rect 115194 116300 115226 116536
rect 115462 116300 115546 116536
rect 115782 116300 115814 116536
rect 115194 80856 115814 116300
rect 115194 80620 115226 80856
rect 115462 80620 115546 80856
rect 115782 80620 115814 80856
rect 115194 80536 115814 80620
rect 115194 80300 115226 80536
rect 115462 80300 115546 80536
rect 115782 80300 115814 80536
rect 115194 44856 115814 80300
rect 115194 44620 115226 44856
rect 115462 44620 115546 44856
rect 115782 44620 115814 44856
rect 115194 44536 115814 44620
rect 115194 44300 115226 44536
rect 115462 44300 115546 44536
rect 115782 44300 115814 44536
rect 115194 8856 115814 44300
rect 115194 8620 115226 8856
rect 115462 8620 115546 8856
rect 115782 8620 115814 8856
rect 115194 8536 115814 8620
rect 115194 8300 115226 8536
rect 115462 8300 115546 8536
rect 115782 8300 115814 8536
rect 115194 -5144 115814 8300
rect 115194 -5380 115226 -5144
rect 115462 -5380 115546 -5144
rect 115782 -5380 115814 -5144
rect 115194 -5464 115814 -5380
rect 115194 -5700 115226 -5464
rect 115462 -5700 115546 -5464
rect 115782 -5700 115814 -5464
rect 115194 -7652 115814 -5700
rect 116434 710600 117054 711592
rect 116434 710364 116466 710600
rect 116702 710364 116786 710600
rect 117022 710364 117054 710600
rect 116434 710280 117054 710364
rect 116434 710044 116466 710280
rect 116702 710044 116786 710280
rect 117022 710044 117054 710280
rect 116434 694096 117054 710044
rect 116434 693860 116466 694096
rect 116702 693860 116786 694096
rect 117022 693860 117054 694096
rect 116434 693776 117054 693860
rect 116434 693540 116466 693776
rect 116702 693540 116786 693776
rect 117022 693540 117054 693776
rect 116434 658096 117054 693540
rect 116434 657860 116466 658096
rect 116702 657860 116786 658096
rect 117022 657860 117054 658096
rect 116434 657776 117054 657860
rect 116434 657540 116466 657776
rect 116702 657540 116786 657776
rect 117022 657540 117054 657776
rect 116434 622096 117054 657540
rect 116434 621860 116466 622096
rect 116702 621860 116786 622096
rect 117022 621860 117054 622096
rect 116434 621776 117054 621860
rect 116434 621540 116466 621776
rect 116702 621540 116786 621776
rect 117022 621540 117054 621776
rect 116434 586096 117054 621540
rect 116434 585860 116466 586096
rect 116702 585860 116786 586096
rect 117022 585860 117054 586096
rect 116434 585776 117054 585860
rect 116434 585540 116466 585776
rect 116702 585540 116786 585776
rect 117022 585540 117054 585776
rect 116434 550096 117054 585540
rect 116434 549860 116466 550096
rect 116702 549860 116786 550096
rect 117022 549860 117054 550096
rect 116434 549776 117054 549860
rect 116434 549540 116466 549776
rect 116702 549540 116786 549776
rect 117022 549540 117054 549776
rect 116434 514096 117054 549540
rect 116434 513860 116466 514096
rect 116702 513860 116786 514096
rect 117022 513860 117054 514096
rect 116434 513776 117054 513860
rect 116434 513540 116466 513776
rect 116702 513540 116786 513776
rect 117022 513540 117054 513776
rect 116434 478096 117054 513540
rect 116434 477860 116466 478096
rect 116702 477860 116786 478096
rect 117022 477860 117054 478096
rect 116434 477776 117054 477860
rect 116434 477540 116466 477776
rect 116702 477540 116786 477776
rect 117022 477540 117054 477776
rect 116434 442096 117054 477540
rect 116434 441860 116466 442096
rect 116702 441860 116786 442096
rect 117022 441860 117054 442096
rect 116434 441776 117054 441860
rect 116434 441540 116466 441776
rect 116702 441540 116786 441776
rect 117022 441540 117054 441776
rect 116434 406096 117054 441540
rect 116434 405860 116466 406096
rect 116702 405860 116786 406096
rect 117022 405860 117054 406096
rect 116434 405776 117054 405860
rect 116434 405540 116466 405776
rect 116702 405540 116786 405776
rect 117022 405540 117054 405776
rect 116434 370096 117054 405540
rect 116434 369860 116466 370096
rect 116702 369860 116786 370096
rect 117022 369860 117054 370096
rect 116434 369776 117054 369860
rect 116434 369540 116466 369776
rect 116702 369540 116786 369776
rect 117022 369540 117054 369776
rect 116434 334096 117054 369540
rect 116434 333860 116466 334096
rect 116702 333860 116786 334096
rect 117022 333860 117054 334096
rect 116434 333776 117054 333860
rect 116434 333540 116466 333776
rect 116702 333540 116786 333776
rect 117022 333540 117054 333776
rect 116434 298096 117054 333540
rect 116434 297860 116466 298096
rect 116702 297860 116786 298096
rect 117022 297860 117054 298096
rect 116434 297776 117054 297860
rect 116434 297540 116466 297776
rect 116702 297540 116786 297776
rect 117022 297540 117054 297776
rect 116434 262096 117054 297540
rect 116434 261860 116466 262096
rect 116702 261860 116786 262096
rect 117022 261860 117054 262096
rect 116434 261776 117054 261860
rect 116434 261540 116466 261776
rect 116702 261540 116786 261776
rect 117022 261540 117054 261776
rect 116434 226096 117054 261540
rect 116434 225860 116466 226096
rect 116702 225860 116786 226096
rect 117022 225860 117054 226096
rect 116434 225776 117054 225860
rect 116434 225540 116466 225776
rect 116702 225540 116786 225776
rect 117022 225540 117054 225776
rect 116434 190096 117054 225540
rect 116434 189860 116466 190096
rect 116702 189860 116786 190096
rect 117022 189860 117054 190096
rect 116434 189776 117054 189860
rect 116434 189540 116466 189776
rect 116702 189540 116786 189776
rect 117022 189540 117054 189776
rect 116434 154096 117054 189540
rect 116434 153860 116466 154096
rect 116702 153860 116786 154096
rect 117022 153860 117054 154096
rect 116434 153776 117054 153860
rect 116434 153540 116466 153776
rect 116702 153540 116786 153776
rect 117022 153540 117054 153776
rect 116434 118096 117054 153540
rect 116434 117860 116466 118096
rect 116702 117860 116786 118096
rect 117022 117860 117054 118096
rect 116434 117776 117054 117860
rect 116434 117540 116466 117776
rect 116702 117540 116786 117776
rect 117022 117540 117054 117776
rect 116434 82096 117054 117540
rect 116434 81860 116466 82096
rect 116702 81860 116786 82096
rect 117022 81860 117054 82096
rect 116434 81776 117054 81860
rect 116434 81540 116466 81776
rect 116702 81540 116786 81776
rect 117022 81540 117054 81776
rect 116434 46096 117054 81540
rect 116434 45860 116466 46096
rect 116702 45860 116786 46096
rect 117022 45860 117054 46096
rect 116434 45776 117054 45860
rect 116434 45540 116466 45776
rect 116702 45540 116786 45776
rect 117022 45540 117054 45776
rect 116434 10096 117054 45540
rect 116434 9860 116466 10096
rect 116702 9860 116786 10096
rect 117022 9860 117054 10096
rect 116434 9776 117054 9860
rect 116434 9540 116466 9776
rect 116702 9540 116786 9776
rect 117022 9540 117054 9776
rect 116434 -6104 117054 9540
rect 116434 -6340 116466 -6104
rect 116702 -6340 116786 -6104
rect 117022 -6340 117054 -6104
rect 116434 -6424 117054 -6340
rect 116434 -6660 116466 -6424
rect 116702 -6660 116786 -6424
rect 117022 -6660 117054 -6424
rect 116434 -7652 117054 -6660
rect 117674 711560 118294 711592
rect 117674 711324 117706 711560
rect 117942 711324 118026 711560
rect 118262 711324 118294 711560
rect 117674 711240 118294 711324
rect 117674 711004 117706 711240
rect 117942 711004 118026 711240
rect 118262 711004 118294 711240
rect 117674 695336 118294 711004
rect 117674 695100 117706 695336
rect 117942 695100 118026 695336
rect 118262 695100 118294 695336
rect 117674 695016 118294 695100
rect 117674 694780 117706 695016
rect 117942 694780 118026 695016
rect 118262 694780 118294 695016
rect 117674 659336 118294 694780
rect 117674 659100 117706 659336
rect 117942 659100 118026 659336
rect 118262 659100 118294 659336
rect 117674 659016 118294 659100
rect 117674 658780 117706 659016
rect 117942 658780 118026 659016
rect 118262 658780 118294 659016
rect 117674 623336 118294 658780
rect 117674 623100 117706 623336
rect 117942 623100 118026 623336
rect 118262 623100 118294 623336
rect 117674 623016 118294 623100
rect 117674 622780 117706 623016
rect 117942 622780 118026 623016
rect 118262 622780 118294 623016
rect 117674 587336 118294 622780
rect 117674 587100 117706 587336
rect 117942 587100 118026 587336
rect 118262 587100 118294 587336
rect 117674 587016 118294 587100
rect 117674 586780 117706 587016
rect 117942 586780 118026 587016
rect 118262 586780 118294 587016
rect 117674 551336 118294 586780
rect 117674 551100 117706 551336
rect 117942 551100 118026 551336
rect 118262 551100 118294 551336
rect 117674 551016 118294 551100
rect 117674 550780 117706 551016
rect 117942 550780 118026 551016
rect 118262 550780 118294 551016
rect 117674 515336 118294 550780
rect 117674 515100 117706 515336
rect 117942 515100 118026 515336
rect 118262 515100 118294 515336
rect 117674 515016 118294 515100
rect 117674 514780 117706 515016
rect 117942 514780 118026 515016
rect 118262 514780 118294 515016
rect 117674 479336 118294 514780
rect 117674 479100 117706 479336
rect 117942 479100 118026 479336
rect 118262 479100 118294 479336
rect 117674 479016 118294 479100
rect 117674 478780 117706 479016
rect 117942 478780 118026 479016
rect 118262 478780 118294 479016
rect 117674 443336 118294 478780
rect 117674 443100 117706 443336
rect 117942 443100 118026 443336
rect 118262 443100 118294 443336
rect 117674 443016 118294 443100
rect 117674 442780 117706 443016
rect 117942 442780 118026 443016
rect 118262 442780 118294 443016
rect 117674 407336 118294 442780
rect 117674 407100 117706 407336
rect 117942 407100 118026 407336
rect 118262 407100 118294 407336
rect 117674 407016 118294 407100
rect 117674 406780 117706 407016
rect 117942 406780 118026 407016
rect 118262 406780 118294 407016
rect 117674 371336 118294 406780
rect 117674 371100 117706 371336
rect 117942 371100 118026 371336
rect 118262 371100 118294 371336
rect 117674 371016 118294 371100
rect 117674 370780 117706 371016
rect 117942 370780 118026 371016
rect 118262 370780 118294 371016
rect 117674 335336 118294 370780
rect 117674 335100 117706 335336
rect 117942 335100 118026 335336
rect 118262 335100 118294 335336
rect 117674 335016 118294 335100
rect 117674 334780 117706 335016
rect 117942 334780 118026 335016
rect 118262 334780 118294 335016
rect 117674 299336 118294 334780
rect 117674 299100 117706 299336
rect 117942 299100 118026 299336
rect 118262 299100 118294 299336
rect 117674 299016 118294 299100
rect 117674 298780 117706 299016
rect 117942 298780 118026 299016
rect 118262 298780 118294 299016
rect 117674 263336 118294 298780
rect 117674 263100 117706 263336
rect 117942 263100 118026 263336
rect 118262 263100 118294 263336
rect 117674 263016 118294 263100
rect 117674 262780 117706 263016
rect 117942 262780 118026 263016
rect 118262 262780 118294 263016
rect 117674 227336 118294 262780
rect 117674 227100 117706 227336
rect 117942 227100 118026 227336
rect 118262 227100 118294 227336
rect 117674 227016 118294 227100
rect 117674 226780 117706 227016
rect 117942 226780 118026 227016
rect 118262 226780 118294 227016
rect 117674 191336 118294 226780
rect 117674 191100 117706 191336
rect 117942 191100 118026 191336
rect 118262 191100 118294 191336
rect 117674 191016 118294 191100
rect 117674 190780 117706 191016
rect 117942 190780 118026 191016
rect 118262 190780 118294 191016
rect 117674 155336 118294 190780
rect 117674 155100 117706 155336
rect 117942 155100 118026 155336
rect 118262 155100 118294 155336
rect 117674 155016 118294 155100
rect 117674 154780 117706 155016
rect 117942 154780 118026 155016
rect 118262 154780 118294 155016
rect 117674 119336 118294 154780
rect 117674 119100 117706 119336
rect 117942 119100 118026 119336
rect 118262 119100 118294 119336
rect 117674 119016 118294 119100
rect 117674 118780 117706 119016
rect 117942 118780 118026 119016
rect 118262 118780 118294 119016
rect 117674 83336 118294 118780
rect 117674 83100 117706 83336
rect 117942 83100 118026 83336
rect 118262 83100 118294 83336
rect 117674 83016 118294 83100
rect 117674 82780 117706 83016
rect 117942 82780 118026 83016
rect 118262 82780 118294 83016
rect 117674 47336 118294 82780
rect 117674 47100 117706 47336
rect 117942 47100 118026 47336
rect 118262 47100 118294 47336
rect 117674 47016 118294 47100
rect 117674 46780 117706 47016
rect 117942 46780 118026 47016
rect 118262 46780 118294 47016
rect 117674 11336 118294 46780
rect 117674 11100 117706 11336
rect 117942 11100 118026 11336
rect 118262 11100 118294 11336
rect 117674 11016 118294 11100
rect 117674 10780 117706 11016
rect 117942 10780 118026 11016
rect 118262 10780 118294 11016
rect 117674 -7064 118294 10780
rect 117674 -7300 117706 -7064
rect 117942 -7300 118026 -7064
rect 118262 -7300 118294 -7064
rect 117674 -7384 118294 -7300
rect 117674 -7620 117706 -7384
rect 117942 -7620 118026 -7384
rect 118262 -7620 118294 -7384
rect 117674 -7652 118294 -7620
rect 144994 704840 145614 711592
rect 144994 704604 145026 704840
rect 145262 704604 145346 704840
rect 145582 704604 145614 704840
rect 144994 704520 145614 704604
rect 144994 704284 145026 704520
rect 145262 704284 145346 704520
rect 145582 704284 145614 704520
rect 144994 686656 145614 704284
rect 144994 686420 145026 686656
rect 145262 686420 145346 686656
rect 145582 686420 145614 686656
rect 144994 686336 145614 686420
rect 144994 686100 145026 686336
rect 145262 686100 145346 686336
rect 145582 686100 145614 686336
rect 144994 650656 145614 686100
rect 144994 650420 145026 650656
rect 145262 650420 145346 650656
rect 145582 650420 145614 650656
rect 144994 650336 145614 650420
rect 144994 650100 145026 650336
rect 145262 650100 145346 650336
rect 145582 650100 145614 650336
rect 144994 614656 145614 650100
rect 144994 614420 145026 614656
rect 145262 614420 145346 614656
rect 145582 614420 145614 614656
rect 144994 614336 145614 614420
rect 144994 614100 145026 614336
rect 145262 614100 145346 614336
rect 145582 614100 145614 614336
rect 144994 578656 145614 614100
rect 144994 578420 145026 578656
rect 145262 578420 145346 578656
rect 145582 578420 145614 578656
rect 144994 578336 145614 578420
rect 144994 578100 145026 578336
rect 145262 578100 145346 578336
rect 145582 578100 145614 578336
rect 144994 542656 145614 578100
rect 144994 542420 145026 542656
rect 145262 542420 145346 542656
rect 145582 542420 145614 542656
rect 144994 542336 145614 542420
rect 144994 542100 145026 542336
rect 145262 542100 145346 542336
rect 145582 542100 145614 542336
rect 144994 506656 145614 542100
rect 144994 506420 145026 506656
rect 145262 506420 145346 506656
rect 145582 506420 145614 506656
rect 144994 506336 145614 506420
rect 144994 506100 145026 506336
rect 145262 506100 145346 506336
rect 145582 506100 145614 506336
rect 144994 470656 145614 506100
rect 144994 470420 145026 470656
rect 145262 470420 145346 470656
rect 145582 470420 145614 470656
rect 144994 470336 145614 470420
rect 144994 470100 145026 470336
rect 145262 470100 145346 470336
rect 145582 470100 145614 470336
rect 144994 434656 145614 470100
rect 144994 434420 145026 434656
rect 145262 434420 145346 434656
rect 145582 434420 145614 434656
rect 144994 434336 145614 434420
rect 144994 434100 145026 434336
rect 145262 434100 145346 434336
rect 145582 434100 145614 434336
rect 144994 398656 145614 434100
rect 144994 398420 145026 398656
rect 145262 398420 145346 398656
rect 145582 398420 145614 398656
rect 144994 398336 145614 398420
rect 144994 398100 145026 398336
rect 145262 398100 145346 398336
rect 145582 398100 145614 398336
rect 144994 362656 145614 398100
rect 144994 362420 145026 362656
rect 145262 362420 145346 362656
rect 145582 362420 145614 362656
rect 144994 362336 145614 362420
rect 144994 362100 145026 362336
rect 145262 362100 145346 362336
rect 145582 362100 145614 362336
rect 144994 326656 145614 362100
rect 144994 326420 145026 326656
rect 145262 326420 145346 326656
rect 145582 326420 145614 326656
rect 144994 326336 145614 326420
rect 144994 326100 145026 326336
rect 145262 326100 145346 326336
rect 145582 326100 145614 326336
rect 144994 290656 145614 326100
rect 144994 290420 145026 290656
rect 145262 290420 145346 290656
rect 145582 290420 145614 290656
rect 144994 290336 145614 290420
rect 144994 290100 145026 290336
rect 145262 290100 145346 290336
rect 145582 290100 145614 290336
rect 144994 254656 145614 290100
rect 144994 254420 145026 254656
rect 145262 254420 145346 254656
rect 145582 254420 145614 254656
rect 144994 254336 145614 254420
rect 144994 254100 145026 254336
rect 145262 254100 145346 254336
rect 145582 254100 145614 254336
rect 144994 218656 145614 254100
rect 144994 218420 145026 218656
rect 145262 218420 145346 218656
rect 145582 218420 145614 218656
rect 144994 218336 145614 218420
rect 144994 218100 145026 218336
rect 145262 218100 145346 218336
rect 145582 218100 145614 218336
rect 144994 182656 145614 218100
rect 144994 182420 145026 182656
rect 145262 182420 145346 182656
rect 145582 182420 145614 182656
rect 144994 182336 145614 182420
rect 144994 182100 145026 182336
rect 145262 182100 145346 182336
rect 145582 182100 145614 182336
rect 144994 146656 145614 182100
rect 144994 146420 145026 146656
rect 145262 146420 145346 146656
rect 145582 146420 145614 146656
rect 144994 146336 145614 146420
rect 144994 146100 145026 146336
rect 145262 146100 145346 146336
rect 145582 146100 145614 146336
rect 144994 110656 145614 146100
rect 144994 110420 145026 110656
rect 145262 110420 145346 110656
rect 145582 110420 145614 110656
rect 144994 110336 145614 110420
rect 144994 110100 145026 110336
rect 145262 110100 145346 110336
rect 145582 110100 145614 110336
rect 144994 74656 145614 110100
rect 144994 74420 145026 74656
rect 145262 74420 145346 74656
rect 145582 74420 145614 74656
rect 144994 74336 145614 74420
rect 144994 74100 145026 74336
rect 145262 74100 145346 74336
rect 145582 74100 145614 74336
rect 144994 38656 145614 74100
rect 144994 38420 145026 38656
rect 145262 38420 145346 38656
rect 145582 38420 145614 38656
rect 144994 38336 145614 38420
rect 144994 38100 145026 38336
rect 145262 38100 145346 38336
rect 145582 38100 145614 38336
rect 144994 2656 145614 38100
rect 144994 2420 145026 2656
rect 145262 2420 145346 2656
rect 145582 2420 145614 2656
rect 144994 2336 145614 2420
rect 144994 2100 145026 2336
rect 145262 2100 145346 2336
rect 145582 2100 145614 2336
rect 144994 -344 145614 2100
rect 144994 -580 145026 -344
rect 145262 -580 145346 -344
rect 145582 -580 145614 -344
rect 144994 -664 145614 -580
rect 144994 -900 145026 -664
rect 145262 -900 145346 -664
rect 145582 -900 145614 -664
rect 144994 -7652 145614 -900
rect 146234 705800 146854 711592
rect 146234 705564 146266 705800
rect 146502 705564 146586 705800
rect 146822 705564 146854 705800
rect 146234 705480 146854 705564
rect 146234 705244 146266 705480
rect 146502 705244 146586 705480
rect 146822 705244 146854 705480
rect 146234 687896 146854 705244
rect 146234 687660 146266 687896
rect 146502 687660 146586 687896
rect 146822 687660 146854 687896
rect 146234 687576 146854 687660
rect 146234 687340 146266 687576
rect 146502 687340 146586 687576
rect 146822 687340 146854 687576
rect 146234 651896 146854 687340
rect 146234 651660 146266 651896
rect 146502 651660 146586 651896
rect 146822 651660 146854 651896
rect 146234 651576 146854 651660
rect 146234 651340 146266 651576
rect 146502 651340 146586 651576
rect 146822 651340 146854 651576
rect 146234 615896 146854 651340
rect 146234 615660 146266 615896
rect 146502 615660 146586 615896
rect 146822 615660 146854 615896
rect 146234 615576 146854 615660
rect 146234 615340 146266 615576
rect 146502 615340 146586 615576
rect 146822 615340 146854 615576
rect 146234 579896 146854 615340
rect 146234 579660 146266 579896
rect 146502 579660 146586 579896
rect 146822 579660 146854 579896
rect 146234 579576 146854 579660
rect 146234 579340 146266 579576
rect 146502 579340 146586 579576
rect 146822 579340 146854 579576
rect 146234 543896 146854 579340
rect 146234 543660 146266 543896
rect 146502 543660 146586 543896
rect 146822 543660 146854 543896
rect 146234 543576 146854 543660
rect 146234 543340 146266 543576
rect 146502 543340 146586 543576
rect 146822 543340 146854 543576
rect 146234 507896 146854 543340
rect 146234 507660 146266 507896
rect 146502 507660 146586 507896
rect 146822 507660 146854 507896
rect 146234 507576 146854 507660
rect 146234 507340 146266 507576
rect 146502 507340 146586 507576
rect 146822 507340 146854 507576
rect 146234 471896 146854 507340
rect 146234 471660 146266 471896
rect 146502 471660 146586 471896
rect 146822 471660 146854 471896
rect 146234 471576 146854 471660
rect 146234 471340 146266 471576
rect 146502 471340 146586 471576
rect 146822 471340 146854 471576
rect 146234 435896 146854 471340
rect 146234 435660 146266 435896
rect 146502 435660 146586 435896
rect 146822 435660 146854 435896
rect 146234 435576 146854 435660
rect 146234 435340 146266 435576
rect 146502 435340 146586 435576
rect 146822 435340 146854 435576
rect 146234 399896 146854 435340
rect 146234 399660 146266 399896
rect 146502 399660 146586 399896
rect 146822 399660 146854 399896
rect 146234 399576 146854 399660
rect 146234 399340 146266 399576
rect 146502 399340 146586 399576
rect 146822 399340 146854 399576
rect 146234 363896 146854 399340
rect 146234 363660 146266 363896
rect 146502 363660 146586 363896
rect 146822 363660 146854 363896
rect 146234 363576 146854 363660
rect 146234 363340 146266 363576
rect 146502 363340 146586 363576
rect 146822 363340 146854 363576
rect 146234 327896 146854 363340
rect 146234 327660 146266 327896
rect 146502 327660 146586 327896
rect 146822 327660 146854 327896
rect 146234 327576 146854 327660
rect 146234 327340 146266 327576
rect 146502 327340 146586 327576
rect 146822 327340 146854 327576
rect 146234 291896 146854 327340
rect 146234 291660 146266 291896
rect 146502 291660 146586 291896
rect 146822 291660 146854 291896
rect 146234 291576 146854 291660
rect 146234 291340 146266 291576
rect 146502 291340 146586 291576
rect 146822 291340 146854 291576
rect 146234 255896 146854 291340
rect 146234 255660 146266 255896
rect 146502 255660 146586 255896
rect 146822 255660 146854 255896
rect 146234 255576 146854 255660
rect 146234 255340 146266 255576
rect 146502 255340 146586 255576
rect 146822 255340 146854 255576
rect 146234 219896 146854 255340
rect 146234 219660 146266 219896
rect 146502 219660 146586 219896
rect 146822 219660 146854 219896
rect 146234 219576 146854 219660
rect 146234 219340 146266 219576
rect 146502 219340 146586 219576
rect 146822 219340 146854 219576
rect 146234 183896 146854 219340
rect 146234 183660 146266 183896
rect 146502 183660 146586 183896
rect 146822 183660 146854 183896
rect 146234 183576 146854 183660
rect 146234 183340 146266 183576
rect 146502 183340 146586 183576
rect 146822 183340 146854 183576
rect 146234 147896 146854 183340
rect 146234 147660 146266 147896
rect 146502 147660 146586 147896
rect 146822 147660 146854 147896
rect 146234 147576 146854 147660
rect 146234 147340 146266 147576
rect 146502 147340 146586 147576
rect 146822 147340 146854 147576
rect 146234 111896 146854 147340
rect 146234 111660 146266 111896
rect 146502 111660 146586 111896
rect 146822 111660 146854 111896
rect 146234 111576 146854 111660
rect 146234 111340 146266 111576
rect 146502 111340 146586 111576
rect 146822 111340 146854 111576
rect 146234 75896 146854 111340
rect 146234 75660 146266 75896
rect 146502 75660 146586 75896
rect 146822 75660 146854 75896
rect 146234 75576 146854 75660
rect 146234 75340 146266 75576
rect 146502 75340 146586 75576
rect 146822 75340 146854 75576
rect 146234 39896 146854 75340
rect 146234 39660 146266 39896
rect 146502 39660 146586 39896
rect 146822 39660 146854 39896
rect 146234 39576 146854 39660
rect 146234 39340 146266 39576
rect 146502 39340 146586 39576
rect 146822 39340 146854 39576
rect 146234 3896 146854 39340
rect 146234 3660 146266 3896
rect 146502 3660 146586 3896
rect 146822 3660 146854 3896
rect 146234 3576 146854 3660
rect 146234 3340 146266 3576
rect 146502 3340 146586 3576
rect 146822 3340 146854 3576
rect 146234 -1304 146854 3340
rect 146234 -1540 146266 -1304
rect 146502 -1540 146586 -1304
rect 146822 -1540 146854 -1304
rect 146234 -1624 146854 -1540
rect 146234 -1860 146266 -1624
rect 146502 -1860 146586 -1624
rect 146822 -1860 146854 -1624
rect 146234 -7652 146854 -1860
rect 147474 706760 148094 711592
rect 147474 706524 147506 706760
rect 147742 706524 147826 706760
rect 148062 706524 148094 706760
rect 147474 706440 148094 706524
rect 147474 706204 147506 706440
rect 147742 706204 147826 706440
rect 148062 706204 148094 706440
rect 147474 689136 148094 706204
rect 147474 688900 147506 689136
rect 147742 688900 147826 689136
rect 148062 688900 148094 689136
rect 147474 688816 148094 688900
rect 147474 688580 147506 688816
rect 147742 688580 147826 688816
rect 148062 688580 148094 688816
rect 147474 653136 148094 688580
rect 147474 652900 147506 653136
rect 147742 652900 147826 653136
rect 148062 652900 148094 653136
rect 147474 652816 148094 652900
rect 147474 652580 147506 652816
rect 147742 652580 147826 652816
rect 148062 652580 148094 652816
rect 147474 617136 148094 652580
rect 147474 616900 147506 617136
rect 147742 616900 147826 617136
rect 148062 616900 148094 617136
rect 147474 616816 148094 616900
rect 147474 616580 147506 616816
rect 147742 616580 147826 616816
rect 148062 616580 148094 616816
rect 147474 581136 148094 616580
rect 147474 580900 147506 581136
rect 147742 580900 147826 581136
rect 148062 580900 148094 581136
rect 147474 580816 148094 580900
rect 147474 580580 147506 580816
rect 147742 580580 147826 580816
rect 148062 580580 148094 580816
rect 147474 545136 148094 580580
rect 147474 544900 147506 545136
rect 147742 544900 147826 545136
rect 148062 544900 148094 545136
rect 147474 544816 148094 544900
rect 147474 544580 147506 544816
rect 147742 544580 147826 544816
rect 148062 544580 148094 544816
rect 147474 509136 148094 544580
rect 147474 508900 147506 509136
rect 147742 508900 147826 509136
rect 148062 508900 148094 509136
rect 147474 508816 148094 508900
rect 147474 508580 147506 508816
rect 147742 508580 147826 508816
rect 148062 508580 148094 508816
rect 147474 473136 148094 508580
rect 147474 472900 147506 473136
rect 147742 472900 147826 473136
rect 148062 472900 148094 473136
rect 147474 472816 148094 472900
rect 147474 472580 147506 472816
rect 147742 472580 147826 472816
rect 148062 472580 148094 472816
rect 147474 437136 148094 472580
rect 147474 436900 147506 437136
rect 147742 436900 147826 437136
rect 148062 436900 148094 437136
rect 147474 436816 148094 436900
rect 147474 436580 147506 436816
rect 147742 436580 147826 436816
rect 148062 436580 148094 436816
rect 147474 401136 148094 436580
rect 147474 400900 147506 401136
rect 147742 400900 147826 401136
rect 148062 400900 148094 401136
rect 147474 400816 148094 400900
rect 147474 400580 147506 400816
rect 147742 400580 147826 400816
rect 148062 400580 148094 400816
rect 147474 365136 148094 400580
rect 147474 364900 147506 365136
rect 147742 364900 147826 365136
rect 148062 364900 148094 365136
rect 147474 364816 148094 364900
rect 147474 364580 147506 364816
rect 147742 364580 147826 364816
rect 148062 364580 148094 364816
rect 147474 329136 148094 364580
rect 147474 328900 147506 329136
rect 147742 328900 147826 329136
rect 148062 328900 148094 329136
rect 147474 328816 148094 328900
rect 147474 328580 147506 328816
rect 147742 328580 147826 328816
rect 148062 328580 148094 328816
rect 147474 293136 148094 328580
rect 147474 292900 147506 293136
rect 147742 292900 147826 293136
rect 148062 292900 148094 293136
rect 147474 292816 148094 292900
rect 147474 292580 147506 292816
rect 147742 292580 147826 292816
rect 148062 292580 148094 292816
rect 147474 257136 148094 292580
rect 147474 256900 147506 257136
rect 147742 256900 147826 257136
rect 148062 256900 148094 257136
rect 147474 256816 148094 256900
rect 147474 256580 147506 256816
rect 147742 256580 147826 256816
rect 148062 256580 148094 256816
rect 147474 221136 148094 256580
rect 147474 220900 147506 221136
rect 147742 220900 147826 221136
rect 148062 220900 148094 221136
rect 147474 220816 148094 220900
rect 147474 220580 147506 220816
rect 147742 220580 147826 220816
rect 148062 220580 148094 220816
rect 147474 185136 148094 220580
rect 147474 184900 147506 185136
rect 147742 184900 147826 185136
rect 148062 184900 148094 185136
rect 147474 184816 148094 184900
rect 147474 184580 147506 184816
rect 147742 184580 147826 184816
rect 148062 184580 148094 184816
rect 147474 149136 148094 184580
rect 147474 148900 147506 149136
rect 147742 148900 147826 149136
rect 148062 148900 148094 149136
rect 147474 148816 148094 148900
rect 147474 148580 147506 148816
rect 147742 148580 147826 148816
rect 148062 148580 148094 148816
rect 147474 113136 148094 148580
rect 147474 112900 147506 113136
rect 147742 112900 147826 113136
rect 148062 112900 148094 113136
rect 147474 112816 148094 112900
rect 147474 112580 147506 112816
rect 147742 112580 147826 112816
rect 148062 112580 148094 112816
rect 147474 77136 148094 112580
rect 147474 76900 147506 77136
rect 147742 76900 147826 77136
rect 148062 76900 148094 77136
rect 147474 76816 148094 76900
rect 147474 76580 147506 76816
rect 147742 76580 147826 76816
rect 148062 76580 148094 76816
rect 147474 41136 148094 76580
rect 147474 40900 147506 41136
rect 147742 40900 147826 41136
rect 148062 40900 148094 41136
rect 147474 40816 148094 40900
rect 147474 40580 147506 40816
rect 147742 40580 147826 40816
rect 148062 40580 148094 40816
rect 147474 5136 148094 40580
rect 147474 4900 147506 5136
rect 147742 4900 147826 5136
rect 148062 4900 148094 5136
rect 147474 4816 148094 4900
rect 147474 4580 147506 4816
rect 147742 4580 147826 4816
rect 148062 4580 148094 4816
rect 147474 -2264 148094 4580
rect 147474 -2500 147506 -2264
rect 147742 -2500 147826 -2264
rect 148062 -2500 148094 -2264
rect 147474 -2584 148094 -2500
rect 147474 -2820 147506 -2584
rect 147742 -2820 147826 -2584
rect 148062 -2820 148094 -2584
rect 147474 -7652 148094 -2820
rect 148714 707720 149334 711592
rect 148714 707484 148746 707720
rect 148982 707484 149066 707720
rect 149302 707484 149334 707720
rect 148714 707400 149334 707484
rect 148714 707164 148746 707400
rect 148982 707164 149066 707400
rect 149302 707164 149334 707400
rect 148714 690376 149334 707164
rect 148714 690140 148746 690376
rect 148982 690140 149066 690376
rect 149302 690140 149334 690376
rect 148714 690056 149334 690140
rect 148714 689820 148746 690056
rect 148982 689820 149066 690056
rect 149302 689820 149334 690056
rect 148714 654376 149334 689820
rect 148714 654140 148746 654376
rect 148982 654140 149066 654376
rect 149302 654140 149334 654376
rect 148714 654056 149334 654140
rect 148714 653820 148746 654056
rect 148982 653820 149066 654056
rect 149302 653820 149334 654056
rect 148714 618376 149334 653820
rect 148714 618140 148746 618376
rect 148982 618140 149066 618376
rect 149302 618140 149334 618376
rect 148714 618056 149334 618140
rect 148714 617820 148746 618056
rect 148982 617820 149066 618056
rect 149302 617820 149334 618056
rect 148714 582376 149334 617820
rect 148714 582140 148746 582376
rect 148982 582140 149066 582376
rect 149302 582140 149334 582376
rect 148714 582056 149334 582140
rect 148714 581820 148746 582056
rect 148982 581820 149066 582056
rect 149302 581820 149334 582056
rect 148714 546376 149334 581820
rect 148714 546140 148746 546376
rect 148982 546140 149066 546376
rect 149302 546140 149334 546376
rect 148714 546056 149334 546140
rect 148714 545820 148746 546056
rect 148982 545820 149066 546056
rect 149302 545820 149334 546056
rect 148714 510376 149334 545820
rect 148714 510140 148746 510376
rect 148982 510140 149066 510376
rect 149302 510140 149334 510376
rect 148714 510056 149334 510140
rect 148714 509820 148746 510056
rect 148982 509820 149066 510056
rect 149302 509820 149334 510056
rect 148714 474376 149334 509820
rect 148714 474140 148746 474376
rect 148982 474140 149066 474376
rect 149302 474140 149334 474376
rect 148714 474056 149334 474140
rect 148714 473820 148746 474056
rect 148982 473820 149066 474056
rect 149302 473820 149334 474056
rect 148714 438376 149334 473820
rect 148714 438140 148746 438376
rect 148982 438140 149066 438376
rect 149302 438140 149334 438376
rect 148714 438056 149334 438140
rect 148714 437820 148746 438056
rect 148982 437820 149066 438056
rect 149302 437820 149334 438056
rect 148714 402376 149334 437820
rect 148714 402140 148746 402376
rect 148982 402140 149066 402376
rect 149302 402140 149334 402376
rect 148714 402056 149334 402140
rect 148714 401820 148746 402056
rect 148982 401820 149066 402056
rect 149302 401820 149334 402056
rect 148714 366376 149334 401820
rect 148714 366140 148746 366376
rect 148982 366140 149066 366376
rect 149302 366140 149334 366376
rect 148714 366056 149334 366140
rect 148714 365820 148746 366056
rect 148982 365820 149066 366056
rect 149302 365820 149334 366056
rect 148714 330376 149334 365820
rect 148714 330140 148746 330376
rect 148982 330140 149066 330376
rect 149302 330140 149334 330376
rect 148714 330056 149334 330140
rect 148714 329820 148746 330056
rect 148982 329820 149066 330056
rect 149302 329820 149334 330056
rect 148714 294376 149334 329820
rect 148714 294140 148746 294376
rect 148982 294140 149066 294376
rect 149302 294140 149334 294376
rect 148714 294056 149334 294140
rect 148714 293820 148746 294056
rect 148982 293820 149066 294056
rect 149302 293820 149334 294056
rect 148714 258376 149334 293820
rect 148714 258140 148746 258376
rect 148982 258140 149066 258376
rect 149302 258140 149334 258376
rect 148714 258056 149334 258140
rect 148714 257820 148746 258056
rect 148982 257820 149066 258056
rect 149302 257820 149334 258056
rect 148714 222376 149334 257820
rect 148714 222140 148746 222376
rect 148982 222140 149066 222376
rect 149302 222140 149334 222376
rect 148714 222056 149334 222140
rect 148714 221820 148746 222056
rect 148982 221820 149066 222056
rect 149302 221820 149334 222056
rect 148714 186376 149334 221820
rect 148714 186140 148746 186376
rect 148982 186140 149066 186376
rect 149302 186140 149334 186376
rect 148714 186056 149334 186140
rect 148714 185820 148746 186056
rect 148982 185820 149066 186056
rect 149302 185820 149334 186056
rect 148714 150376 149334 185820
rect 148714 150140 148746 150376
rect 148982 150140 149066 150376
rect 149302 150140 149334 150376
rect 148714 150056 149334 150140
rect 148714 149820 148746 150056
rect 148982 149820 149066 150056
rect 149302 149820 149334 150056
rect 148714 114376 149334 149820
rect 148714 114140 148746 114376
rect 148982 114140 149066 114376
rect 149302 114140 149334 114376
rect 148714 114056 149334 114140
rect 148714 113820 148746 114056
rect 148982 113820 149066 114056
rect 149302 113820 149334 114056
rect 148714 78376 149334 113820
rect 148714 78140 148746 78376
rect 148982 78140 149066 78376
rect 149302 78140 149334 78376
rect 148714 78056 149334 78140
rect 148714 77820 148746 78056
rect 148982 77820 149066 78056
rect 149302 77820 149334 78056
rect 148714 42376 149334 77820
rect 148714 42140 148746 42376
rect 148982 42140 149066 42376
rect 149302 42140 149334 42376
rect 148714 42056 149334 42140
rect 148714 41820 148746 42056
rect 148982 41820 149066 42056
rect 149302 41820 149334 42056
rect 148714 6376 149334 41820
rect 148714 6140 148746 6376
rect 148982 6140 149066 6376
rect 149302 6140 149334 6376
rect 148714 6056 149334 6140
rect 148714 5820 148746 6056
rect 148982 5820 149066 6056
rect 149302 5820 149334 6056
rect 148714 -3224 149334 5820
rect 148714 -3460 148746 -3224
rect 148982 -3460 149066 -3224
rect 149302 -3460 149334 -3224
rect 148714 -3544 149334 -3460
rect 148714 -3780 148746 -3544
rect 148982 -3780 149066 -3544
rect 149302 -3780 149334 -3544
rect 148714 -7652 149334 -3780
rect 149954 708680 150574 711592
rect 149954 708444 149986 708680
rect 150222 708444 150306 708680
rect 150542 708444 150574 708680
rect 149954 708360 150574 708444
rect 149954 708124 149986 708360
rect 150222 708124 150306 708360
rect 150542 708124 150574 708360
rect 149954 691616 150574 708124
rect 149954 691380 149986 691616
rect 150222 691380 150306 691616
rect 150542 691380 150574 691616
rect 149954 691296 150574 691380
rect 149954 691060 149986 691296
rect 150222 691060 150306 691296
rect 150542 691060 150574 691296
rect 149954 655616 150574 691060
rect 149954 655380 149986 655616
rect 150222 655380 150306 655616
rect 150542 655380 150574 655616
rect 149954 655296 150574 655380
rect 149954 655060 149986 655296
rect 150222 655060 150306 655296
rect 150542 655060 150574 655296
rect 149954 619616 150574 655060
rect 149954 619380 149986 619616
rect 150222 619380 150306 619616
rect 150542 619380 150574 619616
rect 149954 619296 150574 619380
rect 149954 619060 149986 619296
rect 150222 619060 150306 619296
rect 150542 619060 150574 619296
rect 149954 583616 150574 619060
rect 149954 583380 149986 583616
rect 150222 583380 150306 583616
rect 150542 583380 150574 583616
rect 149954 583296 150574 583380
rect 149954 583060 149986 583296
rect 150222 583060 150306 583296
rect 150542 583060 150574 583296
rect 149954 547616 150574 583060
rect 149954 547380 149986 547616
rect 150222 547380 150306 547616
rect 150542 547380 150574 547616
rect 149954 547296 150574 547380
rect 149954 547060 149986 547296
rect 150222 547060 150306 547296
rect 150542 547060 150574 547296
rect 149954 511616 150574 547060
rect 149954 511380 149986 511616
rect 150222 511380 150306 511616
rect 150542 511380 150574 511616
rect 149954 511296 150574 511380
rect 149954 511060 149986 511296
rect 150222 511060 150306 511296
rect 150542 511060 150574 511296
rect 149954 475616 150574 511060
rect 149954 475380 149986 475616
rect 150222 475380 150306 475616
rect 150542 475380 150574 475616
rect 149954 475296 150574 475380
rect 149954 475060 149986 475296
rect 150222 475060 150306 475296
rect 150542 475060 150574 475296
rect 149954 439616 150574 475060
rect 149954 439380 149986 439616
rect 150222 439380 150306 439616
rect 150542 439380 150574 439616
rect 149954 439296 150574 439380
rect 149954 439060 149986 439296
rect 150222 439060 150306 439296
rect 150542 439060 150574 439296
rect 149954 403616 150574 439060
rect 149954 403380 149986 403616
rect 150222 403380 150306 403616
rect 150542 403380 150574 403616
rect 149954 403296 150574 403380
rect 149954 403060 149986 403296
rect 150222 403060 150306 403296
rect 150542 403060 150574 403296
rect 149954 367616 150574 403060
rect 149954 367380 149986 367616
rect 150222 367380 150306 367616
rect 150542 367380 150574 367616
rect 149954 367296 150574 367380
rect 149954 367060 149986 367296
rect 150222 367060 150306 367296
rect 150542 367060 150574 367296
rect 149954 331616 150574 367060
rect 149954 331380 149986 331616
rect 150222 331380 150306 331616
rect 150542 331380 150574 331616
rect 149954 331296 150574 331380
rect 149954 331060 149986 331296
rect 150222 331060 150306 331296
rect 150542 331060 150574 331296
rect 149954 295616 150574 331060
rect 149954 295380 149986 295616
rect 150222 295380 150306 295616
rect 150542 295380 150574 295616
rect 149954 295296 150574 295380
rect 149954 295060 149986 295296
rect 150222 295060 150306 295296
rect 150542 295060 150574 295296
rect 149954 259616 150574 295060
rect 149954 259380 149986 259616
rect 150222 259380 150306 259616
rect 150542 259380 150574 259616
rect 149954 259296 150574 259380
rect 149954 259060 149986 259296
rect 150222 259060 150306 259296
rect 150542 259060 150574 259296
rect 149954 223616 150574 259060
rect 149954 223380 149986 223616
rect 150222 223380 150306 223616
rect 150542 223380 150574 223616
rect 149954 223296 150574 223380
rect 149954 223060 149986 223296
rect 150222 223060 150306 223296
rect 150542 223060 150574 223296
rect 149954 187616 150574 223060
rect 149954 187380 149986 187616
rect 150222 187380 150306 187616
rect 150542 187380 150574 187616
rect 149954 187296 150574 187380
rect 149954 187060 149986 187296
rect 150222 187060 150306 187296
rect 150542 187060 150574 187296
rect 149954 151616 150574 187060
rect 149954 151380 149986 151616
rect 150222 151380 150306 151616
rect 150542 151380 150574 151616
rect 149954 151296 150574 151380
rect 149954 151060 149986 151296
rect 150222 151060 150306 151296
rect 150542 151060 150574 151296
rect 149954 115616 150574 151060
rect 149954 115380 149986 115616
rect 150222 115380 150306 115616
rect 150542 115380 150574 115616
rect 149954 115296 150574 115380
rect 149954 115060 149986 115296
rect 150222 115060 150306 115296
rect 150542 115060 150574 115296
rect 149954 79616 150574 115060
rect 149954 79380 149986 79616
rect 150222 79380 150306 79616
rect 150542 79380 150574 79616
rect 149954 79296 150574 79380
rect 149954 79060 149986 79296
rect 150222 79060 150306 79296
rect 150542 79060 150574 79296
rect 149954 43616 150574 79060
rect 149954 43380 149986 43616
rect 150222 43380 150306 43616
rect 150542 43380 150574 43616
rect 149954 43296 150574 43380
rect 149954 43060 149986 43296
rect 150222 43060 150306 43296
rect 150542 43060 150574 43296
rect 149954 7616 150574 43060
rect 149954 7380 149986 7616
rect 150222 7380 150306 7616
rect 150542 7380 150574 7616
rect 149954 7296 150574 7380
rect 149954 7060 149986 7296
rect 150222 7060 150306 7296
rect 150542 7060 150574 7296
rect 149954 -4184 150574 7060
rect 149954 -4420 149986 -4184
rect 150222 -4420 150306 -4184
rect 150542 -4420 150574 -4184
rect 149954 -4504 150574 -4420
rect 149954 -4740 149986 -4504
rect 150222 -4740 150306 -4504
rect 150542 -4740 150574 -4504
rect 149954 -7652 150574 -4740
rect 151194 709640 151814 711592
rect 151194 709404 151226 709640
rect 151462 709404 151546 709640
rect 151782 709404 151814 709640
rect 151194 709320 151814 709404
rect 151194 709084 151226 709320
rect 151462 709084 151546 709320
rect 151782 709084 151814 709320
rect 151194 692856 151814 709084
rect 151194 692620 151226 692856
rect 151462 692620 151546 692856
rect 151782 692620 151814 692856
rect 151194 692536 151814 692620
rect 151194 692300 151226 692536
rect 151462 692300 151546 692536
rect 151782 692300 151814 692536
rect 151194 656856 151814 692300
rect 151194 656620 151226 656856
rect 151462 656620 151546 656856
rect 151782 656620 151814 656856
rect 151194 656536 151814 656620
rect 151194 656300 151226 656536
rect 151462 656300 151546 656536
rect 151782 656300 151814 656536
rect 151194 620856 151814 656300
rect 151194 620620 151226 620856
rect 151462 620620 151546 620856
rect 151782 620620 151814 620856
rect 151194 620536 151814 620620
rect 151194 620300 151226 620536
rect 151462 620300 151546 620536
rect 151782 620300 151814 620536
rect 151194 584856 151814 620300
rect 151194 584620 151226 584856
rect 151462 584620 151546 584856
rect 151782 584620 151814 584856
rect 151194 584536 151814 584620
rect 151194 584300 151226 584536
rect 151462 584300 151546 584536
rect 151782 584300 151814 584536
rect 151194 548856 151814 584300
rect 151194 548620 151226 548856
rect 151462 548620 151546 548856
rect 151782 548620 151814 548856
rect 151194 548536 151814 548620
rect 151194 548300 151226 548536
rect 151462 548300 151546 548536
rect 151782 548300 151814 548536
rect 151194 512856 151814 548300
rect 151194 512620 151226 512856
rect 151462 512620 151546 512856
rect 151782 512620 151814 512856
rect 151194 512536 151814 512620
rect 151194 512300 151226 512536
rect 151462 512300 151546 512536
rect 151782 512300 151814 512536
rect 151194 476856 151814 512300
rect 151194 476620 151226 476856
rect 151462 476620 151546 476856
rect 151782 476620 151814 476856
rect 151194 476536 151814 476620
rect 151194 476300 151226 476536
rect 151462 476300 151546 476536
rect 151782 476300 151814 476536
rect 151194 440856 151814 476300
rect 151194 440620 151226 440856
rect 151462 440620 151546 440856
rect 151782 440620 151814 440856
rect 151194 440536 151814 440620
rect 151194 440300 151226 440536
rect 151462 440300 151546 440536
rect 151782 440300 151814 440536
rect 151194 404856 151814 440300
rect 151194 404620 151226 404856
rect 151462 404620 151546 404856
rect 151782 404620 151814 404856
rect 151194 404536 151814 404620
rect 151194 404300 151226 404536
rect 151462 404300 151546 404536
rect 151782 404300 151814 404536
rect 151194 368856 151814 404300
rect 151194 368620 151226 368856
rect 151462 368620 151546 368856
rect 151782 368620 151814 368856
rect 151194 368536 151814 368620
rect 151194 368300 151226 368536
rect 151462 368300 151546 368536
rect 151782 368300 151814 368536
rect 151194 332856 151814 368300
rect 151194 332620 151226 332856
rect 151462 332620 151546 332856
rect 151782 332620 151814 332856
rect 151194 332536 151814 332620
rect 151194 332300 151226 332536
rect 151462 332300 151546 332536
rect 151782 332300 151814 332536
rect 151194 296856 151814 332300
rect 151194 296620 151226 296856
rect 151462 296620 151546 296856
rect 151782 296620 151814 296856
rect 151194 296536 151814 296620
rect 151194 296300 151226 296536
rect 151462 296300 151546 296536
rect 151782 296300 151814 296536
rect 151194 260856 151814 296300
rect 151194 260620 151226 260856
rect 151462 260620 151546 260856
rect 151782 260620 151814 260856
rect 151194 260536 151814 260620
rect 151194 260300 151226 260536
rect 151462 260300 151546 260536
rect 151782 260300 151814 260536
rect 151194 224856 151814 260300
rect 151194 224620 151226 224856
rect 151462 224620 151546 224856
rect 151782 224620 151814 224856
rect 151194 224536 151814 224620
rect 151194 224300 151226 224536
rect 151462 224300 151546 224536
rect 151782 224300 151814 224536
rect 151194 188856 151814 224300
rect 151194 188620 151226 188856
rect 151462 188620 151546 188856
rect 151782 188620 151814 188856
rect 151194 188536 151814 188620
rect 151194 188300 151226 188536
rect 151462 188300 151546 188536
rect 151782 188300 151814 188536
rect 151194 152856 151814 188300
rect 151194 152620 151226 152856
rect 151462 152620 151546 152856
rect 151782 152620 151814 152856
rect 151194 152536 151814 152620
rect 151194 152300 151226 152536
rect 151462 152300 151546 152536
rect 151782 152300 151814 152536
rect 151194 116856 151814 152300
rect 151194 116620 151226 116856
rect 151462 116620 151546 116856
rect 151782 116620 151814 116856
rect 151194 116536 151814 116620
rect 151194 116300 151226 116536
rect 151462 116300 151546 116536
rect 151782 116300 151814 116536
rect 151194 80856 151814 116300
rect 151194 80620 151226 80856
rect 151462 80620 151546 80856
rect 151782 80620 151814 80856
rect 151194 80536 151814 80620
rect 151194 80300 151226 80536
rect 151462 80300 151546 80536
rect 151782 80300 151814 80536
rect 151194 44856 151814 80300
rect 151194 44620 151226 44856
rect 151462 44620 151546 44856
rect 151782 44620 151814 44856
rect 151194 44536 151814 44620
rect 151194 44300 151226 44536
rect 151462 44300 151546 44536
rect 151782 44300 151814 44536
rect 151194 8856 151814 44300
rect 151194 8620 151226 8856
rect 151462 8620 151546 8856
rect 151782 8620 151814 8856
rect 151194 8536 151814 8620
rect 151194 8300 151226 8536
rect 151462 8300 151546 8536
rect 151782 8300 151814 8536
rect 151194 -5144 151814 8300
rect 151194 -5380 151226 -5144
rect 151462 -5380 151546 -5144
rect 151782 -5380 151814 -5144
rect 151194 -5464 151814 -5380
rect 151194 -5700 151226 -5464
rect 151462 -5700 151546 -5464
rect 151782 -5700 151814 -5464
rect 151194 -7652 151814 -5700
rect 152434 710600 153054 711592
rect 152434 710364 152466 710600
rect 152702 710364 152786 710600
rect 153022 710364 153054 710600
rect 152434 710280 153054 710364
rect 152434 710044 152466 710280
rect 152702 710044 152786 710280
rect 153022 710044 153054 710280
rect 152434 694096 153054 710044
rect 152434 693860 152466 694096
rect 152702 693860 152786 694096
rect 153022 693860 153054 694096
rect 152434 693776 153054 693860
rect 152434 693540 152466 693776
rect 152702 693540 152786 693776
rect 153022 693540 153054 693776
rect 152434 658096 153054 693540
rect 152434 657860 152466 658096
rect 152702 657860 152786 658096
rect 153022 657860 153054 658096
rect 152434 657776 153054 657860
rect 152434 657540 152466 657776
rect 152702 657540 152786 657776
rect 153022 657540 153054 657776
rect 152434 622096 153054 657540
rect 152434 621860 152466 622096
rect 152702 621860 152786 622096
rect 153022 621860 153054 622096
rect 152434 621776 153054 621860
rect 152434 621540 152466 621776
rect 152702 621540 152786 621776
rect 153022 621540 153054 621776
rect 152434 586096 153054 621540
rect 152434 585860 152466 586096
rect 152702 585860 152786 586096
rect 153022 585860 153054 586096
rect 152434 585776 153054 585860
rect 152434 585540 152466 585776
rect 152702 585540 152786 585776
rect 153022 585540 153054 585776
rect 152434 550096 153054 585540
rect 152434 549860 152466 550096
rect 152702 549860 152786 550096
rect 153022 549860 153054 550096
rect 152434 549776 153054 549860
rect 152434 549540 152466 549776
rect 152702 549540 152786 549776
rect 153022 549540 153054 549776
rect 152434 514096 153054 549540
rect 152434 513860 152466 514096
rect 152702 513860 152786 514096
rect 153022 513860 153054 514096
rect 152434 513776 153054 513860
rect 152434 513540 152466 513776
rect 152702 513540 152786 513776
rect 153022 513540 153054 513776
rect 152434 478096 153054 513540
rect 152434 477860 152466 478096
rect 152702 477860 152786 478096
rect 153022 477860 153054 478096
rect 152434 477776 153054 477860
rect 152434 477540 152466 477776
rect 152702 477540 152786 477776
rect 153022 477540 153054 477776
rect 152434 442096 153054 477540
rect 152434 441860 152466 442096
rect 152702 441860 152786 442096
rect 153022 441860 153054 442096
rect 152434 441776 153054 441860
rect 152434 441540 152466 441776
rect 152702 441540 152786 441776
rect 153022 441540 153054 441776
rect 152434 406096 153054 441540
rect 152434 405860 152466 406096
rect 152702 405860 152786 406096
rect 153022 405860 153054 406096
rect 152434 405776 153054 405860
rect 152434 405540 152466 405776
rect 152702 405540 152786 405776
rect 153022 405540 153054 405776
rect 152434 370096 153054 405540
rect 152434 369860 152466 370096
rect 152702 369860 152786 370096
rect 153022 369860 153054 370096
rect 152434 369776 153054 369860
rect 152434 369540 152466 369776
rect 152702 369540 152786 369776
rect 153022 369540 153054 369776
rect 152434 334096 153054 369540
rect 152434 333860 152466 334096
rect 152702 333860 152786 334096
rect 153022 333860 153054 334096
rect 152434 333776 153054 333860
rect 152434 333540 152466 333776
rect 152702 333540 152786 333776
rect 153022 333540 153054 333776
rect 152434 298096 153054 333540
rect 152434 297860 152466 298096
rect 152702 297860 152786 298096
rect 153022 297860 153054 298096
rect 152434 297776 153054 297860
rect 152434 297540 152466 297776
rect 152702 297540 152786 297776
rect 153022 297540 153054 297776
rect 152434 262096 153054 297540
rect 152434 261860 152466 262096
rect 152702 261860 152786 262096
rect 153022 261860 153054 262096
rect 152434 261776 153054 261860
rect 152434 261540 152466 261776
rect 152702 261540 152786 261776
rect 153022 261540 153054 261776
rect 152434 226096 153054 261540
rect 152434 225860 152466 226096
rect 152702 225860 152786 226096
rect 153022 225860 153054 226096
rect 152434 225776 153054 225860
rect 152434 225540 152466 225776
rect 152702 225540 152786 225776
rect 153022 225540 153054 225776
rect 152434 190096 153054 225540
rect 152434 189860 152466 190096
rect 152702 189860 152786 190096
rect 153022 189860 153054 190096
rect 152434 189776 153054 189860
rect 152434 189540 152466 189776
rect 152702 189540 152786 189776
rect 153022 189540 153054 189776
rect 152434 154096 153054 189540
rect 152434 153860 152466 154096
rect 152702 153860 152786 154096
rect 153022 153860 153054 154096
rect 152434 153776 153054 153860
rect 152434 153540 152466 153776
rect 152702 153540 152786 153776
rect 153022 153540 153054 153776
rect 152434 118096 153054 153540
rect 152434 117860 152466 118096
rect 152702 117860 152786 118096
rect 153022 117860 153054 118096
rect 152434 117776 153054 117860
rect 152434 117540 152466 117776
rect 152702 117540 152786 117776
rect 153022 117540 153054 117776
rect 152434 82096 153054 117540
rect 152434 81860 152466 82096
rect 152702 81860 152786 82096
rect 153022 81860 153054 82096
rect 152434 81776 153054 81860
rect 152434 81540 152466 81776
rect 152702 81540 152786 81776
rect 153022 81540 153054 81776
rect 152434 46096 153054 81540
rect 152434 45860 152466 46096
rect 152702 45860 152786 46096
rect 153022 45860 153054 46096
rect 152434 45776 153054 45860
rect 152434 45540 152466 45776
rect 152702 45540 152786 45776
rect 153022 45540 153054 45776
rect 152434 10096 153054 45540
rect 152434 9860 152466 10096
rect 152702 9860 152786 10096
rect 153022 9860 153054 10096
rect 152434 9776 153054 9860
rect 152434 9540 152466 9776
rect 152702 9540 152786 9776
rect 153022 9540 153054 9776
rect 152434 -6104 153054 9540
rect 152434 -6340 152466 -6104
rect 152702 -6340 152786 -6104
rect 153022 -6340 153054 -6104
rect 152434 -6424 153054 -6340
rect 152434 -6660 152466 -6424
rect 152702 -6660 152786 -6424
rect 153022 -6660 153054 -6424
rect 152434 -7652 153054 -6660
rect 153674 711560 154294 711592
rect 153674 711324 153706 711560
rect 153942 711324 154026 711560
rect 154262 711324 154294 711560
rect 153674 711240 154294 711324
rect 153674 711004 153706 711240
rect 153942 711004 154026 711240
rect 154262 711004 154294 711240
rect 153674 695336 154294 711004
rect 153674 695100 153706 695336
rect 153942 695100 154026 695336
rect 154262 695100 154294 695336
rect 153674 695016 154294 695100
rect 153674 694780 153706 695016
rect 153942 694780 154026 695016
rect 154262 694780 154294 695016
rect 153674 659336 154294 694780
rect 153674 659100 153706 659336
rect 153942 659100 154026 659336
rect 154262 659100 154294 659336
rect 153674 659016 154294 659100
rect 153674 658780 153706 659016
rect 153942 658780 154026 659016
rect 154262 658780 154294 659016
rect 153674 623336 154294 658780
rect 153674 623100 153706 623336
rect 153942 623100 154026 623336
rect 154262 623100 154294 623336
rect 153674 623016 154294 623100
rect 153674 622780 153706 623016
rect 153942 622780 154026 623016
rect 154262 622780 154294 623016
rect 153674 587336 154294 622780
rect 153674 587100 153706 587336
rect 153942 587100 154026 587336
rect 154262 587100 154294 587336
rect 153674 587016 154294 587100
rect 153674 586780 153706 587016
rect 153942 586780 154026 587016
rect 154262 586780 154294 587016
rect 153674 551336 154294 586780
rect 153674 551100 153706 551336
rect 153942 551100 154026 551336
rect 154262 551100 154294 551336
rect 153674 551016 154294 551100
rect 153674 550780 153706 551016
rect 153942 550780 154026 551016
rect 154262 550780 154294 551016
rect 153674 515336 154294 550780
rect 153674 515100 153706 515336
rect 153942 515100 154026 515336
rect 154262 515100 154294 515336
rect 153674 515016 154294 515100
rect 153674 514780 153706 515016
rect 153942 514780 154026 515016
rect 154262 514780 154294 515016
rect 153674 479336 154294 514780
rect 153674 479100 153706 479336
rect 153942 479100 154026 479336
rect 154262 479100 154294 479336
rect 153674 479016 154294 479100
rect 153674 478780 153706 479016
rect 153942 478780 154026 479016
rect 154262 478780 154294 479016
rect 153674 443336 154294 478780
rect 153674 443100 153706 443336
rect 153942 443100 154026 443336
rect 154262 443100 154294 443336
rect 153674 443016 154294 443100
rect 153674 442780 153706 443016
rect 153942 442780 154026 443016
rect 154262 442780 154294 443016
rect 153674 407336 154294 442780
rect 153674 407100 153706 407336
rect 153942 407100 154026 407336
rect 154262 407100 154294 407336
rect 153674 407016 154294 407100
rect 153674 406780 153706 407016
rect 153942 406780 154026 407016
rect 154262 406780 154294 407016
rect 153674 371336 154294 406780
rect 153674 371100 153706 371336
rect 153942 371100 154026 371336
rect 154262 371100 154294 371336
rect 153674 371016 154294 371100
rect 153674 370780 153706 371016
rect 153942 370780 154026 371016
rect 154262 370780 154294 371016
rect 153674 335336 154294 370780
rect 153674 335100 153706 335336
rect 153942 335100 154026 335336
rect 154262 335100 154294 335336
rect 153674 335016 154294 335100
rect 153674 334780 153706 335016
rect 153942 334780 154026 335016
rect 154262 334780 154294 335016
rect 153674 299336 154294 334780
rect 153674 299100 153706 299336
rect 153942 299100 154026 299336
rect 154262 299100 154294 299336
rect 153674 299016 154294 299100
rect 153674 298780 153706 299016
rect 153942 298780 154026 299016
rect 154262 298780 154294 299016
rect 153674 263336 154294 298780
rect 153674 263100 153706 263336
rect 153942 263100 154026 263336
rect 154262 263100 154294 263336
rect 153674 263016 154294 263100
rect 153674 262780 153706 263016
rect 153942 262780 154026 263016
rect 154262 262780 154294 263016
rect 153674 227336 154294 262780
rect 153674 227100 153706 227336
rect 153942 227100 154026 227336
rect 154262 227100 154294 227336
rect 153674 227016 154294 227100
rect 153674 226780 153706 227016
rect 153942 226780 154026 227016
rect 154262 226780 154294 227016
rect 153674 191336 154294 226780
rect 153674 191100 153706 191336
rect 153942 191100 154026 191336
rect 154262 191100 154294 191336
rect 153674 191016 154294 191100
rect 153674 190780 153706 191016
rect 153942 190780 154026 191016
rect 154262 190780 154294 191016
rect 153674 155336 154294 190780
rect 153674 155100 153706 155336
rect 153942 155100 154026 155336
rect 154262 155100 154294 155336
rect 153674 155016 154294 155100
rect 153674 154780 153706 155016
rect 153942 154780 154026 155016
rect 154262 154780 154294 155016
rect 153674 119336 154294 154780
rect 153674 119100 153706 119336
rect 153942 119100 154026 119336
rect 154262 119100 154294 119336
rect 153674 119016 154294 119100
rect 153674 118780 153706 119016
rect 153942 118780 154026 119016
rect 154262 118780 154294 119016
rect 153674 83336 154294 118780
rect 153674 83100 153706 83336
rect 153942 83100 154026 83336
rect 154262 83100 154294 83336
rect 153674 83016 154294 83100
rect 153674 82780 153706 83016
rect 153942 82780 154026 83016
rect 154262 82780 154294 83016
rect 153674 47336 154294 82780
rect 153674 47100 153706 47336
rect 153942 47100 154026 47336
rect 154262 47100 154294 47336
rect 153674 47016 154294 47100
rect 153674 46780 153706 47016
rect 153942 46780 154026 47016
rect 154262 46780 154294 47016
rect 153674 11336 154294 46780
rect 153674 11100 153706 11336
rect 153942 11100 154026 11336
rect 154262 11100 154294 11336
rect 153674 11016 154294 11100
rect 153674 10780 153706 11016
rect 153942 10780 154026 11016
rect 154262 10780 154294 11016
rect 153674 -7064 154294 10780
rect 153674 -7300 153706 -7064
rect 153942 -7300 154026 -7064
rect 154262 -7300 154294 -7064
rect 153674 -7384 154294 -7300
rect 153674 -7620 153706 -7384
rect 153942 -7620 154026 -7384
rect 154262 -7620 154294 -7384
rect 153674 -7652 154294 -7620
rect 180994 704840 181614 711592
rect 180994 704604 181026 704840
rect 181262 704604 181346 704840
rect 181582 704604 181614 704840
rect 180994 704520 181614 704604
rect 180994 704284 181026 704520
rect 181262 704284 181346 704520
rect 181582 704284 181614 704520
rect 180994 686656 181614 704284
rect 180994 686420 181026 686656
rect 181262 686420 181346 686656
rect 181582 686420 181614 686656
rect 180994 686336 181614 686420
rect 180994 686100 181026 686336
rect 181262 686100 181346 686336
rect 181582 686100 181614 686336
rect 180994 650656 181614 686100
rect 180994 650420 181026 650656
rect 181262 650420 181346 650656
rect 181582 650420 181614 650656
rect 180994 650336 181614 650420
rect 180994 650100 181026 650336
rect 181262 650100 181346 650336
rect 181582 650100 181614 650336
rect 180994 614656 181614 650100
rect 180994 614420 181026 614656
rect 181262 614420 181346 614656
rect 181582 614420 181614 614656
rect 180994 614336 181614 614420
rect 180994 614100 181026 614336
rect 181262 614100 181346 614336
rect 181582 614100 181614 614336
rect 180994 578656 181614 614100
rect 180994 578420 181026 578656
rect 181262 578420 181346 578656
rect 181582 578420 181614 578656
rect 180994 578336 181614 578420
rect 180994 578100 181026 578336
rect 181262 578100 181346 578336
rect 181582 578100 181614 578336
rect 180994 542656 181614 578100
rect 180994 542420 181026 542656
rect 181262 542420 181346 542656
rect 181582 542420 181614 542656
rect 180994 542336 181614 542420
rect 180994 542100 181026 542336
rect 181262 542100 181346 542336
rect 181582 542100 181614 542336
rect 180994 506656 181614 542100
rect 180994 506420 181026 506656
rect 181262 506420 181346 506656
rect 181582 506420 181614 506656
rect 180994 506336 181614 506420
rect 180994 506100 181026 506336
rect 181262 506100 181346 506336
rect 181582 506100 181614 506336
rect 180994 470656 181614 506100
rect 180994 470420 181026 470656
rect 181262 470420 181346 470656
rect 181582 470420 181614 470656
rect 180994 470336 181614 470420
rect 180994 470100 181026 470336
rect 181262 470100 181346 470336
rect 181582 470100 181614 470336
rect 180994 434656 181614 470100
rect 180994 434420 181026 434656
rect 181262 434420 181346 434656
rect 181582 434420 181614 434656
rect 180994 434336 181614 434420
rect 180994 434100 181026 434336
rect 181262 434100 181346 434336
rect 181582 434100 181614 434336
rect 180994 398656 181614 434100
rect 180994 398420 181026 398656
rect 181262 398420 181346 398656
rect 181582 398420 181614 398656
rect 180994 398336 181614 398420
rect 180994 398100 181026 398336
rect 181262 398100 181346 398336
rect 181582 398100 181614 398336
rect 180994 362656 181614 398100
rect 180994 362420 181026 362656
rect 181262 362420 181346 362656
rect 181582 362420 181614 362656
rect 180994 362336 181614 362420
rect 180994 362100 181026 362336
rect 181262 362100 181346 362336
rect 181582 362100 181614 362336
rect 180994 326656 181614 362100
rect 180994 326420 181026 326656
rect 181262 326420 181346 326656
rect 181582 326420 181614 326656
rect 180994 326336 181614 326420
rect 180994 326100 181026 326336
rect 181262 326100 181346 326336
rect 181582 326100 181614 326336
rect 180994 290656 181614 326100
rect 180994 290420 181026 290656
rect 181262 290420 181346 290656
rect 181582 290420 181614 290656
rect 180994 290336 181614 290420
rect 180994 290100 181026 290336
rect 181262 290100 181346 290336
rect 181582 290100 181614 290336
rect 180994 254656 181614 290100
rect 180994 254420 181026 254656
rect 181262 254420 181346 254656
rect 181582 254420 181614 254656
rect 180994 254336 181614 254420
rect 180994 254100 181026 254336
rect 181262 254100 181346 254336
rect 181582 254100 181614 254336
rect 180994 218656 181614 254100
rect 180994 218420 181026 218656
rect 181262 218420 181346 218656
rect 181582 218420 181614 218656
rect 180994 218336 181614 218420
rect 180994 218100 181026 218336
rect 181262 218100 181346 218336
rect 181582 218100 181614 218336
rect 180994 182656 181614 218100
rect 180994 182420 181026 182656
rect 181262 182420 181346 182656
rect 181582 182420 181614 182656
rect 180994 182336 181614 182420
rect 180994 182100 181026 182336
rect 181262 182100 181346 182336
rect 181582 182100 181614 182336
rect 180994 146656 181614 182100
rect 180994 146420 181026 146656
rect 181262 146420 181346 146656
rect 181582 146420 181614 146656
rect 180994 146336 181614 146420
rect 180994 146100 181026 146336
rect 181262 146100 181346 146336
rect 181582 146100 181614 146336
rect 180994 110656 181614 146100
rect 180994 110420 181026 110656
rect 181262 110420 181346 110656
rect 181582 110420 181614 110656
rect 180994 110336 181614 110420
rect 180994 110100 181026 110336
rect 181262 110100 181346 110336
rect 181582 110100 181614 110336
rect 180994 74656 181614 110100
rect 180994 74420 181026 74656
rect 181262 74420 181346 74656
rect 181582 74420 181614 74656
rect 180994 74336 181614 74420
rect 180994 74100 181026 74336
rect 181262 74100 181346 74336
rect 181582 74100 181614 74336
rect 180994 38656 181614 74100
rect 180994 38420 181026 38656
rect 181262 38420 181346 38656
rect 181582 38420 181614 38656
rect 180994 38336 181614 38420
rect 180994 38100 181026 38336
rect 181262 38100 181346 38336
rect 181582 38100 181614 38336
rect 180994 2656 181614 38100
rect 180994 2420 181026 2656
rect 181262 2420 181346 2656
rect 181582 2420 181614 2656
rect 180994 2336 181614 2420
rect 180994 2100 181026 2336
rect 181262 2100 181346 2336
rect 181582 2100 181614 2336
rect 180994 -344 181614 2100
rect 180994 -580 181026 -344
rect 181262 -580 181346 -344
rect 181582 -580 181614 -344
rect 180994 -664 181614 -580
rect 180994 -900 181026 -664
rect 181262 -900 181346 -664
rect 181582 -900 181614 -664
rect 180994 -7652 181614 -900
rect 182234 705800 182854 711592
rect 182234 705564 182266 705800
rect 182502 705564 182586 705800
rect 182822 705564 182854 705800
rect 182234 705480 182854 705564
rect 182234 705244 182266 705480
rect 182502 705244 182586 705480
rect 182822 705244 182854 705480
rect 182234 687896 182854 705244
rect 182234 687660 182266 687896
rect 182502 687660 182586 687896
rect 182822 687660 182854 687896
rect 182234 687576 182854 687660
rect 182234 687340 182266 687576
rect 182502 687340 182586 687576
rect 182822 687340 182854 687576
rect 182234 651896 182854 687340
rect 182234 651660 182266 651896
rect 182502 651660 182586 651896
rect 182822 651660 182854 651896
rect 182234 651576 182854 651660
rect 182234 651340 182266 651576
rect 182502 651340 182586 651576
rect 182822 651340 182854 651576
rect 182234 615896 182854 651340
rect 182234 615660 182266 615896
rect 182502 615660 182586 615896
rect 182822 615660 182854 615896
rect 182234 615576 182854 615660
rect 182234 615340 182266 615576
rect 182502 615340 182586 615576
rect 182822 615340 182854 615576
rect 182234 579896 182854 615340
rect 182234 579660 182266 579896
rect 182502 579660 182586 579896
rect 182822 579660 182854 579896
rect 182234 579576 182854 579660
rect 182234 579340 182266 579576
rect 182502 579340 182586 579576
rect 182822 579340 182854 579576
rect 182234 543896 182854 579340
rect 182234 543660 182266 543896
rect 182502 543660 182586 543896
rect 182822 543660 182854 543896
rect 182234 543576 182854 543660
rect 182234 543340 182266 543576
rect 182502 543340 182586 543576
rect 182822 543340 182854 543576
rect 182234 507896 182854 543340
rect 182234 507660 182266 507896
rect 182502 507660 182586 507896
rect 182822 507660 182854 507896
rect 182234 507576 182854 507660
rect 182234 507340 182266 507576
rect 182502 507340 182586 507576
rect 182822 507340 182854 507576
rect 182234 471896 182854 507340
rect 182234 471660 182266 471896
rect 182502 471660 182586 471896
rect 182822 471660 182854 471896
rect 182234 471576 182854 471660
rect 182234 471340 182266 471576
rect 182502 471340 182586 471576
rect 182822 471340 182854 471576
rect 182234 435896 182854 471340
rect 182234 435660 182266 435896
rect 182502 435660 182586 435896
rect 182822 435660 182854 435896
rect 182234 435576 182854 435660
rect 182234 435340 182266 435576
rect 182502 435340 182586 435576
rect 182822 435340 182854 435576
rect 182234 399896 182854 435340
rect 182234 399660 182266 399896
rect 182502 399660 182586 399896
rect 182822 399660 182854 399896
rect 182234 399576 182854 399660
rect 182234 399340 182266 399576
rect 182502 399340 182586 399576
rect 182822 399340 182854 399576
rect 182234 363896 182854 399340
rect 182234 363660 182266 363896
rect 182502 363660 182586 363896
rect 182822 363660 182854 363896
rect 182234 363576 182854 363660
rect 182234 363340 182266 363576
rect 182502 363340 182586 363576
rect 182822 363340 182854 363576
rect 182234 327896 182854 363340
rect 182234 327660 182266 327896
rect 182502 327660 182586 327896
rect 182822 327660 182854 327896
rect 182234 327576 182854 327660
rect 182234 327340 182266 327576
rect 182502 327340 182586 327576
rect 182822 327340 182854 327576
rect 182234 291896 182854 327340
rect 182234 291660 182266 291896
rect 182502 291660 182586 291896
rect 182822 291660 182854 291896
rect 182234 291576 182854 291660
rect 182234 291340 182266 291576
rect 182502 291340 182586 291576
rect 182822 291340 182854 291576
rect 182234 255896 182854 291340
rect 182234 255660 182266 255896
rect 182502 255660 182586 255896
rect 182822 255660 182854 255896
rect 182234 255576 182854 255660
rect 182234 255340 182266 255576
rect 182502 255340 182586 255576
rect 182822 255340 182854 255576
rect 182234 219896 182854 255340
rect 182234 219660 182266 219896
rect 182502 219660 182586 219896
rect 182822 219660 182854 219896
rect 182234 219576 182854 219660
rect 182234 219340 182266 219576
rect 182502 219340 182586 219576
rect 182822 219340 182854 219576
rect 182234 183896 182854 219340
rect 182234 183660 182266 183896
rect 182502 183660 182586 183896
rect 182822 183660 182854 183896
rect 182234 183576 182854 183660
rect 182234 183340 182266 183576
rect 182502 183340 182586 183576
rect 182822 183340 182854 183576
rect 182234 147896 182854 183340
rect 182234 147660 182266 147896
rect 182502 147660 182586 147896
rect 182822 147660 182854 147896
rect 182234 147576 182854 147660
rect 182234 147340 182266 147576
rect 182502 147340 182586 147576
rect 182822 147340 182854 147576
rect 182234 111896 182854 147340
rect 182234 111660 182266 111896
rect 182502 111660 182586 111896
rect 182822 111660 182854 111896
rect 182234 111576 182854 111660
rect 182234 111340 182266 111576
rect 182502 111340 182586 111576
rect 182822 111340 182854 111576
rect 182234 75896 182854 111340
rect 182234 75660 182266 75896
rect 182502 75660 182586 75896
rect 182822 75660 182854 75896
rect 182234 75576 182854 75660
rect 182234 75340 182266 75576
rect 182502 75340 182586 75576
rect 182822 75340 182854 75576
rect 182234 39896 182854 75340
rect 182234 39660 182266 39896
rect 182502 39660 182586 39896
rect 182822 39660 182854 39896
rect 182234 39576 182854 39660
rect 182234 39340 182266 39576
rect 182502 39340 182586 39576
rect 182822 39340 182854 39576
rect 182234 3896 182854 39340
rect 182234 3660 182266 3896
rect 182502 3660 182586 3896
rect 182822 3660 182854 3896
rect 182234 3576 182854 3660
rect 182234 3340 182266 3576
rect 182502 3340 182586 3576
rect 182822 3340 182854 3576
rect 182234 -1304 182854 3340
rect 182234 -1540 182266 -1304
rect 182502 -1540 182586 -1304
rect 182822 -1540 182854 -1304
rect 182234 -1624 182854 -1540
rect 182234 -1860 182266 -1624
rect 182502 -1860 182586 -1624
rect 182822 -1860 182854 -1624
rect 182234 -7652 182854 -1860
rect 183474 706760 184094 711592
rect 183474 706524 183506 706760
rect 183742 706524 183826 706760
rect 184062 706524 184094 706760
rect 183474 706440 184094 706524
rect 183474 706204 183506 706440
rect 183742 706204 183826 706440
rect 184062 706204 184094 706440
rect 183474 689136 184094 706204
rect 183474 688900 183506 689136
rect 183742 688900 183826 689136
rect 184062 688900 184094 689136
rect 183474 688816 184094 688900
rect 183474 688580 183506 688816
rect 183742 688580 183826 688816
rect 184062 688580 184094 688816
rect 183474 653136 184094 688580
rect 183474 652900 183506 653136
rect 183742 652900 183826 653136
rect 184062 652900 184094 653136
rect 183474 652816 184094 652900
rect 183474 652580 183506 652816
rect 183742 652580 183826 652816
rect 184062 652580 184094 652816
rect 183474 617136 184094 652580
rect 183474 616900 183506 617136
rect 183742 616900 183826 617136
rect 184062 616900 184094 617136
rect 183474 616816 184094 616900
rect 183474 616580 183506 616816
rect 183742 616580 183826 616816
rect 184062 616580 184094 616816
rect 183474 581136 184094 616580
rect 183474 580900 183506 581136
rect 183742 580900 183826 581136
rect 184062 580900 184094 581136
rect 183474 580816 184094 580900
rect 183474 580580 183506 580816
rect 183742 580580 183826 580816
rect 184062 580580 184094 580816
rect 183474 545136 184094 580580
rect 183474 544900 183506 545136
rect 183742 544900 183826 545136
rect 184062 544900 184094 545136
rect 183474 544816 184094 544900
rect 183474 544580 183506 544816
rect 183742 544580 183826 544816
rect 184062 544580 184094 544816
rect 183474 509136 184094 544580
rect 183474 508900 183506 509136
rect 183742 508900 183826 509136
rect 184062 508900 184094 509136
rect 183474 508816 184094 508900
rect 183474 508580 183506 508816
rect 183742 508580 183826 508816
rect 184062 508580 184094 508816
rect 183474 473136 184094 508580
rect 183474 472900 183506 473136
rect 183742 472900 183826 473136
rect 184062 472900 184094 473136
rect 183474 472816 184094 472900
rect 183474 472580 183506 472816
rect 183742 472580 183826 472816
rect 184062 472580 184094 472816
rect 183474 437136 184094 472580
rect 183474 436900 183506 437136
rect 183742 436900 183826 437136
rect 184062 436900 184094 437136
rect 183474 436816 184094 436900
rect 183474 436580 183506 436816
rect 183742 436580 183826 436816
rect 184062 436580 184094 436816
rect 183474 401136 184094 436580
rect 183474 400900 183506 401136
rect 183742 400900 183826 401136
rect 184062 400900 184094 401136
rect 183474 400816 184094 400900
rect 183474 400580 183506 400816
rect 183742 400580 183826 400816
rect 184062 400580 184094 400816
rect 183474 365136 184094 400580
rect 183474 364900 183506 365136
rect 183742 364900 183826 365136
rect 184062 364900 184094 365136
rect 183474 364816 184094 364900
rect 183474 364580 183506 364816
rect 183742 364580 183826 364816
rect 184062 364580 184094 364816
rect 183474 329136 184094 364580
rect 183474 328900 183506 329136
rect 183742 328900 183826 329136
rect 184062 328900 184094 329136
rect 183474 328816 184094 328900
rect 183474 328580 183506 328816
rect 183742 328580 183826 328816
rect 184062 328580 184094 328816
rect 183474 293136 184094 328580
rect 183474 292900 183506 293136
rect 183742 292900 183826 293136
rect 184062 292900 184094 293136
rect 183474 292816 184094 292900
rect 183474 292580 183506 292816
rect 183742 292580 183826 292816
rect 184062 292580 184094 292816
rect 183474 257136 184094 292580
rect 183474 256900 183506 257136
rect 183742 256900 183826 257136
rect 184062 256900 184094 257136
rect 183474 256816 184094 256900
rect 183474 256580 183506 256816
rect 183742 256580 183826 256816
rect 184062 256580 184094 256816
rect 183474 221136 184094 256580
rect 183474 220900 183506 221136
rect 183742 220900 183826 221136
rect 184062 220900 184094 221136
rect 183474 220816 184094 220900
rect 183474 220580 183506 220816
rect 183742 220580 183826 220816
rect 184062 220580 184094 220816
rect 183474 185136 184094 220580
rect 183474 184900 183506 185136
rect 183742 184900 183826 185136
rect 184062 184900 184094 185136
rect 183474 184816 184094 184900
rect 183474 184580 183506 184816
rect 183742 184580 183826 184816
rect 184062 184580 184094 184816
rect 183474 149136 184094 184580
rect 183474 148900 183506 149136
rect 183742 148900 183826 149136
rect 184062 148900 184094 149136
rect 183474 148816 184094 148900
rect 183474 148580 183506 148816
rect 183742 148580 183826 148816
rect 184062 148580 184094 148816
rect 183474 113136 184094 148580
rect 183474 112900 183506 113136
rect 183742 112900 183826 113136
rect 184062 112900 184094 113136
rect 183474 112816 184094 112900
rect 183474 112580 183506 112816
rect 183742 112580 183826 112816
rect 184062 112580 184094 112816
rect 183474 77136 184094 112580
rect 183474 76900 183506 77136
rect 183742 76900 183826 77136
rect 184062 76900 184094 77136
rect 183474 76816 184094 76900
rect 183474 76580 183506 76816
rect 183742 76580 183826 76816
rect 184062 76580 184094 76816
rect 183474 41136 184094 76580
rect 183474 40900 183506 41136
rect 183742 40900 183826 41136
rect 184062 40900 184094 41136
rect 183474 40816 184094 40900
rect 183474 40580 183506 40816
rect 183742 40580 183826 40816
rect 184062 40580 184094 40816
rect 183474 5136 184094 40580
rect 183474 4900 183506 5136
rect 183742 4900 183826 5136
rect 184062 4900 184094 5136
rect 183474 4816 184094 4900
rect 183474 4580 183506 4816
rect 183742 4580 183826 4816
rect 184062 4580 184094 4816
rect 183474 -2264 184094 4580
rect 183474 -2500 183506 -2264
rect 183742 -2500 183826 -2264
rect 184062 -2500 184094 -2264
rect 183474 -2584 184094 -2500
rect 183474 -2820 183506 -2584
rect 183742 -2820 183826 -2584
rect 184062 -2820 184094 -2584
rect 183474 -7652 184094 -2820
rect 184714 707720 185334 711592
rect 184714 707484 184746 707720
rect 184982 707484 185066 707720
rect 185302 707484 185334 707720
rect 184714 707400 185334 707484
rect 184714 707164 184746 707400
rect 184982 707164 185066 707400
rect 185302 707164 185334 707400
rect 184714 690376 185334 707164
rect 184714 690140 184746 690376
rect 184982 690140 185066 690376
rect 185302 690140 185334 690376
rect 184714 690056 185334 690140
rect 184714 689820 184746 690056
rect 184982 689820 185066 690056
rect 185302 689820 185334 690056
rect 184714 654376 185334 689820
rect 184714 654140 184746 654376
rect 184982 654140 185066 654376
rect 185302 654140 185334 654376
rect 184714 654056 185334 654140
rect 184714 653820 184746 654056
rect 184982 653820 185066 654056
rect 185302 653820 185334 654056
rect 184714 618376 185334 653820
rect 184714 618140 184746 618376
rect 184982 618140 185066 618376
rect 185302 618140 185334 618376
rect 184714 618056 185334 618140
rect 184714 617820 184746 618056
rect 184982 617820 185066 618056
rect 185302 617820 185334 618056
rect 184714 582376 185334 617820
rect 184714 582140 184746 582376
rect 184982 582140 185066 582376
rect 185302 582140 185334 582376
rect 184714 582056 185334 582140
rect 184714 581820 184746 582056
rect 184982 581820 185066 582056
rect 185302 581820 185334 582056
rect 184714 546376 185334 581820
rect 184714 546140 184746 546376
rect 184982 546140 185066 546376
rect 185302 546140 185334 546376
rect 184714 546056 185334 546140
rect 184714 545820 184746 546056
rect 184982 545820 185066 546056
rect 185302 545820 185334 546056
rect 184714 510376 185334 545820
rect 184714 510140 184746 510376
rect 184982 510140 185066 510376
rect 185302 510140 185334 510376
rect 184714 510056 185334 510140
rect 184714 509820 184746 510056
rect 184982 509820 185066 510056
rect 185302 509820 185334 510056
rect 184714 474376 185334 509820
rect 184714 474140 184746 474376
rect 184982 474140 185066 474376
rect 185302 474140 185334 474376
rect 184714 474056 185334 474140
rect 184714 473820 184746 474056
rect 184982 473820 185066 474056
rect 185302 473820 185334 474056
rect 184714 438376 185334 473820
rect 184714 438140 184746 438376
rect 184982 438140 185066 438376
rect 185302 438140 185334 438376
rect 184714 438056 185334 438140
rect 184714 437820 184746 438056
rect 184982 437820 185066 438056
rect 185302 437820 185334 438056
rect 184714 402376 185334 437820
rect 184714 402140 184746 402376
rect 184982 402140 185066 402376
rect 185302 402140 185334 402376
rect 184714 402056 185334 402140
rect 184714 401820 184746 402056
rect 184982 401820 185066 402056
rect 185302 401820 185334 402056
rect 184714 366376 185334 401820
rect 184714 366140 184746 366376
rect 184982 366140 185066 366376
rect 185302 366140 185334 366376
rect 184714 366056 185334 366140
rect 184714 365820 184746 366056
rect 184982 365820 185066 366056
rect 185302 365820 185334 366056
rect 184714 330376 185334 365820
rect 184714 330140 184746 330376
rect 184982 330140 185066 330376
rect 185302 330140 185334 330376
rect 184714 330056 185334 330140
rect 184714 329820 184746 330056
rect 184982 329820 185066 330056
rect 185302 329820 185334 330056
rect 184714 294376 185334 329820
rect 184714 294140 184746 294376
rect 184982 294140 185066 294376
rect 185302 294140 185334 294376
rect 184714 294056 185334 294140
rect 184714 293820 184746 294056
rect 184982 293820 185066 294056
rect 185302 293820 185334 294056
rect 184714 258376 185334 293820
rect 184714 258140 184746 258376
rect 184982 258140 185066 258376
rect 185302 258140 185334 258376
rect 184714 258056 185334 258140
rect 184714 257820 184746 258056
rect 184982 257820 185066 258056
rect 185302 257820 185334 258056
rect 184714 222376 185334 257820
rect 184714 222140 184746 222376
rect 184982 222140 185066 222376
rect 185302 222140 185334 222376
rect 184714 222056 185334 222140
rect 184714 221820 184746 222056
rect 184982 221820 185066 222056
rect 185302 221820 185334 222056
rect 184714 186376 185334 221820
rect 184714 186140 184746 186376
rect 184982 186140 185066 186376
rect 185302 186140 185334 186376
rect 184714 186056 185334 186140
rect 184714 185820 184746 186056
rect 184982 185820 185066 186056
rect 185302 185820 185334 186056
rect 184714 150376 185334 185820
rect 184714 150140 184746 150376
rect 184982 150140 185066 150376
rect 185302 150140 185334 150376
rect 184714 150056 185334 150140
rect 184714 149820 184746 150056
rect 184982 149820 185066 150056
rect 185302 149820 185334 150056
rect 184714 114376 185334 149820
rect 184714 114140 184746 114376
rect 184982 114140 185066 114376
rect 185302 114140 185334 114376
rect 184714 114056 185334 114140
rect 184714 113820 184746 114056
rect 184982 113820 185066 114056
rect 185302 113820 185334 114056
rect 184714 78376 185334 113820
rect 184714 78140 184746 78376
rect 184982 78140 185066 78376
rect 185302 78140 185334 78376
rect 184714 78056 185334 78140
rect 184714 77820 184746 78056
rect 184982 77820 185066 78056
rect 185302 77820 185334 78056
rect 184714 42376 185334 77820
rect 184714 42140 184746 42376
rect 184982 42140 185066 42376
rect 185302 42140 185334 42376
rect 184714 42056 185334 42140
rect 184714 41820 184746 42056
rect 184982 41820 185066 42056
rect 185302 41820 185334 42056
rect 184714 6376 185334 41820
rect 184714 6140 184746 6376
rect 184982 6140 185066 6376
rect 185302 6140 185334 6376
rect 184714 6056 185334 6140
rect 184714 5820 184746 6056
rect 184982 5820 185066 6056
rect 185302 5820 185334 6056
rect 184714 -3224 185334 5820
rect 184714 -3460 184746 -3224
rect 184982 -3460 185066 -3224
rect 185302 -3460 185334 -3224
rect 184714 -3544 185334 -3460
rect 184714 -3780 184746 -3544
rect 184982 -3780 185066 -3544
rect 185302 -3780 185334 -3544
rect 184714 -7652 185334 -3780
rect 185954 708680 186574 711592
rect 185954 708444 185986 708680
rect 186222 708444 186306 708680
rect 186542 708444 186574 708680
rect 185954 708360 186574 708444
rect 185954 708124 185986 708360
rect 186222 708124 186306 708360
rect 186542 708124 186574 708360
rect 185954 691616 186574 708124
rect 185954 691380 185986 691616
rect 186222 691380 186306 691616
rect 186542 691380 186574 691616
rect 185954 691296 186574 691380
rect 185954 691060 185986 691296
rect 186222 691060 186306 691296
rect 186542 691060 186574 691296
rect 185954 655616 186574 691060
rect 185954 655380 185986 655616
rect 186222 655380 186306 655616
rect 186542 655380 186574 655616
rect 185954 655296 186574 655380
rect 185954 655060 185986 655296
rect 186222 655060 186306 655296
rect 186542 655060 186574 655296
rect 185954 619616 186574 655060
rect 185954 619380 185986 619616
rect 186222 619380 186306 619616
rect 186542 619380 186574 619616
rect 185954 619296 186574 619380
rect 185954 619060 185986 619296
rect 186222 619060 186306 619296
rect 186542 619060 186574 619296
rect 185954 583616 186574 619060
rect 185954 583380 185986 583616
rect 186222 583380 186306 583616
rect 186542 583380 186574 583616
rect 185954 583296 186574 583380
rect 185954 583060 185986 583296
rect 186222 583060 186306 583296
rect 186542 583060 186574 583296
rect 185954 547616 186574 583060
rect 185954 547380 185986 547616
rect 186222 547380 186306 547616
rect 186542 547380 186574 547616
rect 185954 547296 186574 547380
rect 185954 547060 185986 547296
rect 186222 547060 186306 547296
rect 186542 547060 186574 547296
rect 185954 511616 186574 547060
rect 185954 511380 185986 511616
rect 186222 511380 186306 511616
rect 186542 511380 186574 511616
rect 185954 511296 186574 511380
rect 185954 511060 185986 511296
rect 186222 511060 186306 511296
rect 186542 511060 186574 511296
rect 185954 475616 186574 511060
rect 185954 475380 185986 475616
rect 186222 475380 186306 475616
rect 186542 475380 186574 475616
rect 185954 475296 186574 475380
rect 185954 475060 185986 475296
rect 186222 475060 186306 475296
rect 186542 475060 186574 475296
rect 185954 439616 186574 475060
rect 185954 439380 185986 439616
rect 186222 439380 186306 439616
rect 186542 439380 186574 439616
rect 185954 439296 186574 439380
rect 185954 439060 185986 439296
rect 186222 439060 186306 439296
rect 186542 439060 186574 439296
rect 185954 403616 186574 439060
rect 185954 403380 185986 403616
rect 186222 403380 186306 403616
rect 186542 403380 186574 403616
rect 185954 403296 186574 403380
rect 185954 403060 185986 403296
rect 186222 403060 186306 403296
rect 186542 403060 186574 403296
rect 185954 367616 186574 403060
rect 185954 367380 185986 367616
rect 186222 367380 186306 367616
rect 186542 367380 186574 367616
rect 185954 367296 186574 367380
rect 185954 367060 185986 367296
rect 186222 367060 186306 367296
rect 186542 367060 186574 367296
rect 185954 331616 186574 367060
rect 185954 331380 185986 331616
rect 186222 331380 186306 331616
rect 186542 331380 186574 331616
rect 185954 331296 186574 331380
rect 185954 331060 185986 331296
rect 186222 331060 186306 331296
rect 186542 331060 186574 331296
rect 185954 295616 186574 331060
rect 185954 295380 185986 295616
rect 186222 295380 186306 295616
rect 186542 295380 186574 295616
rect 185954 295296 186574 295380
rect 185954 295060 185986 295296
rect 186222 295060 186306 295296
rect 186542 295060 186574 295296
rect 185954 259616 186574 295060
rect 185954 259380 185986 259616
rect 186222 259380 186306 259616
rect 186542 259380 186574 259616
rect 185954 259296 186574 259380
rect 185954 259060 185986 259296
rect 186222 259060 186306 259296
rect 186542 259060 186574 259296
rect 185954 223616 186574 259060
rect 185954 223380 185986 223616
rect 186222 223380 186306 223616
rect 186542 223380 186574 223616
rect 185954 223296 186574 223380
rect 185954 223060 185986 223296
rect 186222 223060 186306 223296
rect 186542 223060 186574 223296
rect 185954 187616 186574 223060
rect 185954 187380 185986 187616
rect 186222 187380 186306 187616
rect 186542 187380 186574 187616
rect 185954 187296 186574 187380
rect 185954 187060 185986 187296
rect 186222 187060 186306 187296
rect 186542 187060 186574 187296
rect 185954 151616 186574 187060
rect 185954 151380 185986 151616
rect 186222 151380 186306 151616
rect 186542 151380 186574 151616
rect 185954 151296 186574 151380
rect 185954 151060 185986 151296
rect 186222 151060 186306 151296
rect 186542 151060 186574 151296
rect 185954 115616 186574 151060
rect 185954 115380 185986 115616
rect 186222 115380 186306 115616
rect 186542 115380 186574 115616
rect 185954 115296 186574 115380
rect 185954 115060 185986 115296
rect 186222 115060 186306 115296
rect 186542 115060 186574 115296
rect 185954 79616 186574 115060
rect 185954 79380 185986 79616
rect 186222 79380 186306 79616
rect 186542 79380 186574 79616
rect 185954 79296 186574 79380
rect 185954 79060 185986 79296
rect 186222 79060 186306 79296
rect 186542 79060 186574 79296
rect 185954 43616 186574 79060
rect 185954 43380 185986 43616
rect 186222 43380 186306 43616
rect 186542 43380 186574 43616
rect 185954 43296 186574 43380
rect 185954 43060 185986 43296
rect 186222 43060 186306 43296
rect 186542 43060 186574 43296
rect 185954 7616 186574 43060
rect 185954 7380 185986 7616
rect 186222 7380 186306 7616
rect 186542 7380 186574 7616
rect 185954 7296 186574 7380
rect 185954 7060 185986 7296
rect 186222 7060 186306 7296
rect 186542 7060 186574 7296
rect 185954 -4184 186574 7060
rect 185954 -4420 185986 -4184
rect 186222 -4420 186306 -4184
rect 186542 -4420 186574 -4184
rect 185954 -4504 186574 -4420
rect 185954 -4740 185986 -4504
rect 186222 -4740 186306 -4504
rect 186542 -4740 186574 -4504
rect 185954 -7652 186574 -4740
rect 187194 709640 187814 711592
rect 187194 709404 187226 709640
rect 187462 709404 187546 709640
rect 187782 709404 187814 709640
rect 187194 709320 187814 709404
rect 187194 709084 187226 709320
rect 187462 709084 187546 709320
rect 187782 709084 187814 709320
rect 187194 692856 187814 709084
rect 187194 692620 187226 692856
rect 187462 692620 187546 692856
rect 187782 692620 187814 692856
rect 187194 692536 187814 692620
rect 187194 692300 187226 692536
rect 187462 692300 187546 692536
rect 187782 692300 187814 692536
rect 187194 656856 187814 692300
rect 187194 656620 187226 656856
rect 187462 656620 187546 656856
rect 187782 656620 187814 656856
rect 187194 656536 187814 656620
rect 187194 656300 187226 656536
rect 187462 656300 187546 656536
rect 187782 656300 187814 656536
rect 187194 620856 187814 656300
rect 187194 620620 187226 620856
rect 187462 620620 187546 620856
rect 187782 620620 187814 620856
rect 187194 620536 187814 620620
rect 187194 620300 187226 620536
rect 187462 620300 187546 620536
rect 187782 620300 187814 620536
rect 187194 584856 187814 620300
rect 187194 584620 187226 584856
rect 187462 584620 187546 584856
rect 187782 584620 187814 584856
rect 187194 584536 187814 584620
rect 187194 584300 187226 584536
rect 187462 584300 187546 584536
rect 187782 584300 187814 584536
rect 187194 548856 187814 584300
rect 187194 548620 187226 548856
rect 187462 548620 187546 548856
rect 187782 548620 187814 548856
rect 187194 548536 187814 548620
rect 187194 548300 187226 548536
rect 187462 548300 187546 548536
rect 187782 548300 187814 548536
rect 187194 512856 187814 548300
rect 187194 512620 187226 512856
rect 187462 512620 187546 512856
rect 187782 512620 187814 512856
rect 187194 512536 187814 512620
rect 187194 512300 187226 512536
rect 187462 512300 187546 512536
rect 187782 512300 187814 512536
rect 187194 476856 187814 512300
rect 187194 476620 187226 476856
rect 187462 476620 187546 476856
rect 187782 476620 187814 476856
rect 187194 476536 187814 476620
rect 187194 476300 187226 476536
rect 187462 476300 187546 476536
rect 187782 476300 187814 476536
rect 187194 440856 187814 476300
rect 187194 440620 187226 440856
rect 187462 440620 187546 440856
rect 187782 440620 187814 440856
rect 187194 440536 187814 440620
rect 187194 440300 187226 440536
rect 187462 440300 187546 440536
rect 187782 440300 187814 440536
rect 187194 404856 187814 440300
rect 187194 404620 187226 404856
rect 187462 404620 187546 404856
rect 187782 404620 187814 404856
rect 187194 404536 187814 404620
rect 187194 404300 187226 404536
rect 187462 404300 187546 404536
rect 187782 404300 187814 404536
rect 187194 368856 187814 404300
rect 187194 368620 187226 368856
rect 187462 368620 187546 368856
rect 187782 368620 187814 368856
rect 187194 368536 187814 368620
rect 187194 368300 187226 368536
rect 187462 368300 187546 368536
rect 187782 368300 187814 368536
rect 187194 332856 187814 368300
rect 187194 332620 187226 332856
rect 187462 332620 187546 332856
rect 187782 332620 187814 332856
rect 187194 332536 187814 332620
rect 187194 332300 187226 332536
rect 187462 332300 187546 332536
rect 187782 332300 187814 332536
rect 187194 296856 187814 332300
rect 187194 296620 187226 296856
rect 187462 296620 187546 296856
rect 187782 296620 187814 296856
rect 187194 296536 187814 296620
rect 187194 296300 187226 296536
rect 187462 296300 187546 296536
rect 187782 296300 187814 296536
rect 187194 260856 187814 296300
rect 187194 260620 187226 260856
rect 187462 260620 187546 260856
rect 187782 260620 187814 260856
rect 187194 260536 187814 260620
rect 187194 260300 187226 260536
rect 187462 260300 187546 260536
rect 187782 260300 187814 260536
rect 187194 224856 187814 260300
rect 187194 224620 187226 224856
rect 187462 224620 187546 224856
rect 187782 224620 187814 224856
rect 187194 224536 187814 224620
rect 187194 224300 187226 224536
rect 187462 224300 187546 224536
rect 187782 224300 187814 224536
rect 187194 188856 187814 224300
rect 187194 188620 187226 188856
rect 187462 188620 187546 188856
rect 187782 188620 187814 188856
rect 187194 188536 187814 188620
rect 187194 188300 187226 188536
rect 187462 188300 187546 188536
rect 187782 188300 187814 188536
rect 187194 152856 187814 188300
rect 187194 152620 187226 152856
rect 187462 152620 187546 152856
rect 187782 152620 187814 152856
rect 187194 152536 187814 152620
rect 187194 152300 187226 152536
rect 187462 152300 187546 152536
rect 187782 152300 187814 152536
rect 187194 116856 187814 152300
rect 187194 116620 187226 116856
rect 187462 116620 187546 116856
rect 187782 116620 187814 116856
rect 187194 116536 187814 116620
rect 187194 116300 187226 116536
rect 187462 116300 187546 116536
rect 187782 116300 187814 116536
rect 187194 80856 187814 116300
rect 187194 80620 187226 80856
rect 187462 80620 187546 80856
rect 187782 80620 187814 80856
rect 187194 80536 187814 80620
rect 187194 80300 187226 80536
rect 187462 80300 187546 80536
rect 187782 80300 187814 80536
rect 187194 44856 187814 80300
rect 187194 44620 187226 44856
rect 187462 44620 187546 44856
rect 187782 44620 187814 44856
rect 187194 44536 187814 44620
rect 187194 44300 187226 44536
rect 187462 44300 187546 44536
rect 187782 44300 187814 44536
rect 187194 8856 187814 44300
rect 187194 8620 187226 8856
rect 187462 8620 187546 8856
rect 187782 8620 187814 8856
rect 187194 8536 187814 8620
rect 187194 8300 187226 8536
rect 187462 8300 187546 8536
rect 187782 8300 187814 8536
rect 187194 -5144 187814 8300
rect 187194 -5380 187226 -5144
rect 187462 -5380 187546 -5144
rect 187782 -5380 187814 -5144
rect 187194 -5464 187814 -5380
rect 187194 -5700 187226 -5464
rect 187462 -5700 187546 -5464
rect 187782 -5700 187814 -5464
rect 187194 -7652 187814 -5700
rect 188434 710600 189054 711592
rect 188434 710364 188466 710600
rect 188702 710364 188786 710600
rect 189022 710364 189054 710600
rect 188434 710280 189054 710364
rect 188434 710044 188466 710280
rect 188702 710044 188786 710280
rect 189022 710044 189054 710280
rect 188434 694096 189054 710044
rect 188434 693860 188466 694096
rect 188702 693860 188786 694096
rect 189022 693860 189054 694096
rect 188434 693776 189054 693860
rect 188434 693540 188466 693776
rect 188702 693540 188786 693776
rect 189022 693540 189054 693776
rect 188434 658096 189054 693540
rect 188434 657860 188466 658096
rect 188702 657860 188786 658096
rect 189022 657860 189054 658096
rect 188434 657776 189054 657860
rect 188434 657540 188466 657776
rect 188702 657540 188786 657776
rect 189022 657540 189054 657776
rect 188434 622096 189054 657540
rect 188434 621860 188466 622096
rect 188702 621860 188786 622096
rect 189022 621860 189054 622096
rect 188434 621776 189054 621860
rect 188434 621540 188466 621776
rect 188702 621540 188786 621776
rect 189022 621540 189054 621776
rect 188434 586096 189054 621540
rect 188434 585860 188466 586096
rect 188702 585860 188786 586096
rect 189022 585860 189054 586096
rect 188434 585776 189054 585860
rect 188434 585540 188466 585776
rect 188702 585540 188786 585776
rect 189022 585540 189054 585776
rect 188434 550096 189054 585540
rect 188434 549860 188466 550096
rect 188702 549860 188786 550096
rect 189022 549860 189054 550096
rect 188434 549776 189054 549860
rect 188434 549540 188466 549776
rect 188702 549540 188786 549776
rect 189022 549540 189054 549776
rect 188434 514096 189054 549540
rect 188434 513860 188466 514096
rect 188702 513860 188786 514096
rect 189022 513860 189054 514096
rect 188434 513776 189054 513860
rect 188434 513540 188466 513776
rect 188702 513540 188786 513776
rect 189022 513540 189054 513776
rect 188434 478096 189054 513540
rect 188434 477860 188466 478096
rect 188702 477860 188786 478096
rect 189022 477860 189054 478096
rect 188434 477776 189054 477860
rect 188434 477540 188466 477776
rect 188702 477540 188786 477776
rect 189022 477540 189054 477776
rect 188434 442096 189054 477540
rect 188434 441860 188466 442096
rect 188702 441860 188786 442096
rect 189022 441860 189054 442096
rect 188434 441776 189054 441860
rect 188434 441540 188466 441776
rect 188702 441540 188786 441776
rect 189022 441540 189054 441776
rect 188434 406096 189054 441540
rect 188434 405860 188466 406096
rect 188702 405860 188786 406096
rect 189022 405860 189054 406096
rect 188434 405776 189054 405860
rect 188434 405540 188466 405776
rect 188702 405540 188786 405776
rect 189022 405540 189054 405776
rect 188434 370096 189054 405540
rect 188434 369860 188466 370096
rect 188702 369860 188786 370096
rect 189022 369860 189054 370096
rect 188434 369776 189054 369860
rect 188434 369540 188466 369776
rect 188702 369540 188786 369776
rect 189022 369540 189054 369776
rect 188434 334096 189054 369540
rect 188434 333860 188466 334096
rect 188702 333860 188786 334096
rect 189022 333860 189054 334096
rect 188434 333776 189054 333860
rect 188434 333540 188466 333776
rect 188702 333540 188786 333776
rect 189022 333540 189054 333776
rect 188434 298096 189054 333540
rect 188434 297860 188466 298096
rect 188702 297860 188786 298096
rect 189022 297860 189054 298096
rect 188434 297776 189054 297860
rect 188434 297540 188466 297776
rect 188702 297540 188786 297776
rect 189022 297540 189054 297776
rect 188434 262096 189054 297540
rect 188434 261860 188466 262096
rect 188702 261860 188786 262096
rect 189022 261860 189054 262096
rect 188434 261776 189054 261860
rect 188434 261540 188466 261776
rect 188702 261540 188786 261776
rect 189022 261540 189054 261776
rect 188434 226096 189054 261540
rect 188434 225860 188466 226096
rect 188702 225860 188786 226096
rect 189022 225860 189054 226096
rect 188434 225776 189054 225860
rect 188434 225540 188466 225776
rect 188702 225540 188786 225776
rect 189022 225540 189054 225776
rect 188434 190096 189054 225540
rect 188434 189860 188466 190096
rect 188702 189860 188786 190096
rect 189022 189860 189054 190096
rect 188434 189776 189054 189860
rect 188434 189540 188466 189776
rect 188702 189540 188786 189776
rect 189022 189540 189054 189776
rect 188434 154096 189054 189540
rect 188434 153860 188466 154096
rect 188702 153860 188786 154096
rect 189022 153860 189054 154096
rect 188434 153776 189054 153860
rect 188434 153540 188466 153776
rect 188702 153540 188786 153776
rect 189022 153540 189054 153776
rect 188434 118096 189054 153540
rect 188434 117860 188466 118096
rect 188702 117860 188786 118096
rect 189022 117860 189054 118096
rect 188434 117776 189054 117860
rect 188434 117540 188466 117776
rect 188702 117540 188786 117776
rect 189022 117540 189054 117776
rect 188434 82096 189054 117540
rect 188434 81860 188466 82096
rect 188702 81860 188786 82096
rect 189022 81860 189054 82096
rect 188434 81776 189054 81860
rect 188434 81540 188466 81776
rect 188702 81540 188786 81776
rect 189022 81540 189054 81776
rect 188434 46096 189054 81540
rect 188434 45860 188466 46096
rect 188702 45860 188786 46096
rect 189022 45860 189054 46096
rect 188434 45776 189054 45860
rect 188434 45540 188466 45776
rect 188702 45540 188786 45776
rect 189022 45540 189054 45776
rect 188434 10096 189054 45540
rect 188434 9860 188466 10096
rect 188702 9860 188786 10096
rect 189022 9860 189054 10096
rect 188434 9776 189054 9860
rect 188434 9540 188466 9776
rect 188702 9540 188786 9776
rect 189022 9540 189054 9776
rect 188434 -6104 189054 9540
rect 188434 -6340 188466 -6104
rect 188702 -6340 188786 -6104
rect 189022 -6340 189054 -6104
rect 188434 -6424 189054 -6340
rect 188434 -6660 188466 -6424
rect 188702 -6660 188786 -6424
rect 189022 -6660 189054 -6424
rect 188434 -7652 189054 -6660
rect 189674 711560 190294 711592
rect 189674 711324 189706 711560
rect 189942 711324 190026 711560
rect 190262 711324 190294 711560
rect 189674 711240 190294 711324
rect 189674 711004 189706 711240
rect 189942 711004 190026 711240
rect 190262 711004 190294 711240
rect 189674 695336 190294 711004
rect 189674 695100 189706 695336
rect 189942 695100 190026 695336
rect 190262 695100 190294 695336
rect 189674 695016 190294 695100
rect 189674 694780 189706 695016
rect 189942 694780 190026 695016
rect 190262 694780 190294 695016
rect 189674 659336 190294 694780
rect 189674 659100 189706 659336
rect 189942 659100 190026 659336
rect 190262 659100 190294 659336
rect 189674 659016 190294 659100
rect 189674 658780 189706 659016
rect 189942 658780 190026 659016
rect 190262 658780 190294 659016
rect 189674 623336 190294 658780
rect 189674 623100 189706 623336
rect 189942 623100 190026 623336
rect 190262 623100 190294 623336
rect 189674 623016 190294 623100
rect 189674 622780 189706 623016
rect 189942 622780 190026 623016
rect 190262 622780 190294 623016
rect 189674 587336 190294 622780
rect 189674 587100 189706 587336
rect 189942 587100 190026 587336
rect 190262 587100 190294 587336
rect 189674 587016 190294 587100
rect 189674 586780 189706 587016
rect 189942 586780 190026 587016
rect 190262 586780 190294 587016
rect 189674 551336 190294 586780
rect 189674 551100 189706 551336
rect 189942 551100 190026 551336
rect 190262 551100 190294 551336
rect 189674 551016 190294 551100
rect 189674 550780 189706 551016
rect 189942 550780 190026 551016
rect 190262 550780 190294 551016
rect 189674 515336 190294 550780
rect 189674 515100 189706 515336
rect 189942 515100 190026 515336
rect 190262 515100 190294 515336
rect 189674 515016 190294 515100
rect 189674 514780 189706 515016
rect 189942 514780 190026 515016
rect 190262 514780 190294 515016
rect 189674 479336 190294 514780
rect 189674 479100 189706 479336
rect 189942 479100 190026 479336
rect 190262 479100 190294 479336
rect 189674 479016 190294 479100
rect 189674 478780 189706 479016
rect 189942 478780 190026 479016
rect 190262 478780 190294 479016
rect 189674 443336 190294 478780
rect 189674 443100 189706 443336
rect 189942 443100 190026 443336
rect 190262 443100 190294 443336
rect 189674 443016 190294 443100
rect 189674 442780 189706 443016
rect 189942 442780 190026 443016
rect 190262 442780 190294 443016
rect 189674 407336 190294 442780
rect 189674 407100 189706 407336
rect 189942 407100 190026 407336
rect 190262 407100 190294 407336
rect 189674 407016 190294 407100
rect 189674 406780 189706 407016
rect 189942 406780 190026 407016
rect 190262 406780 190294 407016
rect 189674 371336 190294 406780
rect 189674 371100 189706 371336
rect 189942 371100 190026 371336
rect 190262 371100 190294 371336
rect 189674 371016 190294 371100
rect 189674 370780 189706 371016
rect 189942 370780 190026 371016
rect 190262 370780 190294 371016
rect 189674 335336 190294 370780
rect 189674 335100 189706 335336
rect 189942 335100 190026 335336
rect 190262 335100 190294 335336
rect 189674 335016 190294 335100
rect 189674 334780 189706 335016
rect 189942 334780 190026 335016
rect 190262 334780 190294 335016
rect 189674 299336 190294 334780
rect 189674 299100 189706 299336
rect 189942 299100 190026 299336
rect 190262 299100 190294 299336
rect 189674 299016 190294 299100
rect 189674 298780 189706 299016
rect 189942 298780 190026 299016
rect 190262 298780 190294 299016
rect 189674 263336 190294 298780
rect 189674 263100 189706 263336
rect 189942 263100 190026 263336
rect 190262 263100 190294 263336
rect 189674 263016 190294 263100
rect 189674 262780 189706 263016
rect 189942 262780 190026 263016
rect 190262 262780 190294 263016
rect 189674 227336 190294 262780
rect 189674 227100 189706 227336
rect 189942 227100 190026 227336
rect 190262 227100 190294 227336
rect 189674 227016 190294 227100
rect 189674 226780 189706 227016
rect 189942 226780 190026 227016
rect 190262 226780 190294 227016
rect 189674 191336 190294 226780
rect 189674 191100 189706 191336
rect 189942 191100 190026 191336
rect 190262 191100 190294 191336
rect 189674 191016 190294 191100
rect 189674 190780 189706 191016
rect 189942 190780 190026 191016
rect 190262 190780 190294 191016
rect 189674 155336 190294 190780
rect 189674 155100 189706 155336
rect 189942 155100 190026 155336
rect 190262 155100 190294 155336
rect 189674 155016 190294 155100
rect 189674 154780 189706 155016
rect 189942 154780 190026 155016
rect 190262 154780 190294 155016
rect 189674 119336 190294 154780
rect 189674 119100 189706 119336
rect 189942 119100 190026 119336
rect 190262 119100 190294 119336
rect 189674 119016 190294 119100
rect 189674 118780 189706 119016
rect 189942 118780 190026 119016
rect 190262 118780 190294 119016
rect 189674 83336 190294 118780
rect 189674 83100 189706 83336
rect 189942 83100 190026 83336
rect 190262 83100 190294 83336
rect 189674 83016 190294 83100
rect 189674 82780 189706 83016
rect 189942 82780 190026 83016
rect 190262 82780 190294 83016
rect 189674 47336 190294 82780
rect 189674 47100 189706 47336
rect 189942 47100 190026 47336
rect 190262 47100 190294 47336
rect 189674 47016 190294 47100
rect 189674 46780 189706 47016
rect 189942 46780 190026 47016
rect 190262 46780 190294 47016
rect 189674 11336 190294 46780
rect 189674 11100 189706 11336
rect 189942 11100 190026 11336
rect 190262 11100 190294 11336
rect 189674 11016 190294 11100
rect 189674 10780 189706 11016
rect 189942 10780 190026 11016
rect 190262 10780 190294 11016
rect 189674 -7064 190294 10780
rect 189674 -7300 189706 -7064
rect 189942 -7300 190026 -7064
rect 190262 -7300 190294 -7064
rect 189674 -7384 190294 -7300
rect 189674 -7620 189706 -7384
rect 189942 -7620 190026 -7384
rect 190262 -7620 190294 -7384
rect 189674 -7652 190294 -7620
rect 216994 704840 217614 711592
rect 216994 704604 217026 704840
rect 217262 704604 217346 704840
rect 217582 704604 217614 704840
rect 216994 704520 217614 704604
rect 216994 704284 217026 704520
rect 217262 704284 217346 704520
rect 217582 704284 217614 704520
rect 216994 686656 217614 704284
rect 216994 686420 217026 686656
rect 217262 686420 217346 686656
rect 217582 686420 217614 686656
rect 216994 686336 217614 686420
rect 216994 686100 217026 686336
rect 217262 686100 217346 686336
rect 217582 686100 217614 686336
rect 216994 650656 217614 686100
rect 216994 650420 217026 650656
rect 217262 650420 217346 650656
rect 217582 650420 217614 650656
rect 216994 650336 217614 650420
rect 216994 650100 217026 650336
rect 217262 650100 217346 650336
rect 217582 650100 217614 650336
rect 216994 614656 217614 650100
rect 216994 614420 217026 614656
rect 217262 614420 217346 614656
rect 217582 614420 217614 614656
rect 216994 614336 217614 614420
rect 216994 614100 217026 614336
rect 217262 614100 217346 614336
rect 217582 614100 217614 614336
rect 216994 578656 217614 614100
rect 216994 578420 217026 578656
rect 217262 578420 217346 578656
rect 217582 578420 217614 578656
rect 216994 578336 217614 578420
rect 216994 578100 217026 578336
rect 217262 578100 217346 578336
rect 217582 578100 217614 578336
rect 216994 542656 217614 578100
rect 216994 542420 217026 542656
rect 217262 542420 217346 542656
rect 217582 542420 217614 542656
rect 216994 542336 217614 542420
rect 216994 542100 217026 542336
rect 217262 542100 217346 542336
rect 217582 542100 217614 542336
rect 216994 506656 217614 542100
rect 216994 506420 217026 506656
rect 217262 506420 217346 506656
rect 217582 506420 217614 506656
rect 216994 506336 217614 506420
rect 216994 506100 217026 506336
rect 217262 506100 217346 506336
rect 217582 506100 217614 506336
rect 216994 470656 217614 506100
rect 216994 470420 217026 470656
rect 217262 470420 217346 470656
rect 217582 470420 217614 470656
rect 216994 470336 217614 470420
rect 216994 470100 217026 470336
rect 217262 470100 217346 470336
rect 217582 470100 217614 470336
rect 216994 434656 217614 470100
rect 216994 434420 217026 434656
rect 217262 434420 217346 434656
rect 217582 434420 217614 434656
rect 216994 434336 217614 434420
rect 216994 434100 217026 434336
rect 217262 434100 217346 434336
rect 217582 434100 217614 434336
rect 216994 398656 217614 434100
rect 216994 398420 217026 398656
rect 217262 398420 217346 398656
rect 217582 398420 217614 398656
rect 216994 398336 217614 398420
rect 216994 398100 217026 398336
rect 217262 398100 217346 398336
rect 217582 398100 217614 398336
rect 216994 362656 217614 398100
rect 216994 362420 217026 362656
rect 217262 362420 217346 362656
rect 217582 362420 217614 362656
rect 216994 362336 217614 362420
rect 216994 362100 217026 362336
rect 217262 362100 217346 362336
rect 217582 362100 217614 362336
rect 216994 326656 217614 362100
rect 216994 326420 217026 326656
rect 217262 326420 217346 326656
rect 217582 326420 217614 326656
rect 216994 326336 217614 326420
rect 216994 326100 217026 326336
rect 217262 326100 217346 326336
rect 217582 326100 217614 326336
rect 216994 290656 217614 326100
rect 216994 290420 217026 290656
rect 217262 290420 217346 290656
rect 217582 290420 217614 290656
rect 216994 290336 217614 290420
rect 216994 290100 217026 290336
rect 217262 290100 217346 290336
rect 217582 290100 217614 290336
rect 216994 254656 217614 290100
rect 216994 254420 217026 254656
rect 217262 254420 217346 254656
rect 217582 254420 217614 254656
rect 216994 254336 217614 254420
rect 216994 254100 217026 254336
rect 217262 254100 217346 254336
rect 217582 254100 217614 254336
rect 216994 218656 217614 254100
rect 216994 218420 217026 218656
rect 217262 218420 217346 218656
rect 217582 218420 217614 218656
rect 216994 218336 217614 218420
rect 216994 218100 217026 218336
rect 217262 218100 217346 218336
rect 217582 218100 217614 218336
rect 216994 182656 217614 218100
rect 216994 182420 217026 182656
rect 217262 182420 217346 182656
rect 217582 182420 217614 182656
rect 216994 182336 217614 182420
rect 216994 182100 217026 182336
rect 217262 182100 217346 182336
rect 217582 182100 217614 182336
rect 216994 146656 217614 182100
rect 216994 146420 217026 146656
rect 217262 146420 217346 146656
rect 217582 146420 217614 146656
rect 216994 146336 217614 146420
rect 216994 146100 217026 146336
rect 217262 146100 217346 146336
rect 217582 146100 217614 146336
rect 216994 110656 217614 146100
rect 216994 110420 217026 110656
rect 217262 110420 217346 110656
rect 217582 110420 217614 110656
rect 216994 110336 217614 110420
rect 216994 110100 217026 110336
rect 217262 110100 217346 110336
rect 217582 110100 217614 110336
rect 216994 74656 217614 110100
rect 216994 74420 217026 74656
rect 217262 74420 217346 74656
rect 217582 74420 217614 74656
rect 216994 74336 217614 74420
rect 216994 74100 217026 74336
rect 217262 74100 217346 74336
rect 217582 74100 217614 74336
rect 216994 38656 217614 74100
rect 216994 38420 217026 38656
rect 217262 38420 217346 38656
rect 217582 38420 217614 38656
rect 216994 38336 217614 38420
rect 216994 38100 217026 38336
rect 217262 38100 217346 38336
rect 217582 38100 217614 38336
rect 216994 2656 217614 38100
rect 216994 2420 217026 2656
rect 217262 2420 217346 2656
rect 217582 2420 217614 2656
rect 216994 2336 217614 2420
rect 216994 2100 217026 2336
rect 217262 2100 217346 2336
rect 217582 2100 217614 2336
rect 216994 -344 217614 2100
rect 216994 -580 217026 -344
rect 217262 -580 217346 -344
rect 217582 -580 217614 -344
rect 216994 -664 217614 -580
rect 216994 -900 217026 -664
rect 217262 -900 217346 -664
rect 217582 -900 217614 -664
rect 216994 -7652 217614 -900
rect 218234 705800 218854 711592
rect 218234 705564 218266 705800
rect 218502 705564 218586 705800
rect 218822 705564 218854 705800
rect 218234 705480 218854 705564
rect 218234 705244 218266 705480
rect 218502 705244 218586 705480
rect 218822 705244 218854 705480
rect 218234 687896 218854 705244
rect 218234 687660 218266 687896
rect 218502 687660 218586 687896
rect 218822 687660 218854 687896
rect 218234 687576 218854 687660
rect 218234 687340 218266 687576
rect 218502 687340 218586 687576
rect 218822 687340 218854 687576
rect 218234 651896 218854 687340
rect 218234 651660 218266 651896
rect 218502 651660 218586 651896
rect 218822 651660 218854 651896
rect 218234 651576 218854 651660
rect 218234 651340 218266 651576
rect 218502 651340 218586 651576
rect 218822 651340 218854 651576
rect 218234 615896 218854 651340
rect 218234 615660 218266 615896
rect 218502 615660 218586 615896
rect 218822 615660 218854 615896
rect 218234 615576 218854 615660
rect 218234 615340 218266 615576
rect 218502 615340 218586 615576
rect 218822 615340 218854 615576
rect 218234 579896 218854 615340
rect 218234 579660 218266 579896
rect 218502 579660 218586 579896
rect 218822 579660 218854 579896
rect 218234 579576 218854 579660
rect 218234 579340 218266 579576
rect 218502 579340 218586 579576
rect 218822 579340 218854 579576
rect 218234 543896 218854 579340
rect 218234 543660 218266 543896
rect 218502 543660 218586 543896
rect 218822 543660 218854 543896
rect 218234 543576 218854 543660
rect 218234 543340 218266 543576
rect 218502 543340 218586 543576
rect 218822 543340 218854 543576
rect 218234 507896 218854 543340
rect 218234 507660 218266 507896
rect 218502 507660 218586 507896
rect 218822 507660 218854 507896
rect 218234 507576 218854 507660
rect 218234 507340 218266 507576
rect 218502 507340 218586 507576
rect 218822 507340 218854 507576
rect 218234 471896 218854 507340
rect 218234 471660 218266 471896
rect 218502 471660 218586 471896
rect 218822 471660 218854 471896
rect 218234 471576 218854 471660
rect 218234 471340 218266 471576
rect 218502 471340 218586 471576
rect 218822 471340 218854 471576
rect 218234 435896 218854 471340
rect 218234 435660 218266 435896
rect 218502 435660 218586 435896
rect 218822 435660 218854 435896
rect 218234 435576 218854 435660
rect 218234 435340 218266 435576
rect 218502 435340 218586 435576
rect 218822 435340 218854 435576
rect 218234 399896 218854 435340
rect 218234 399660 218266 399896
rect 218502 399660 218586 399896
rect 218822 399660 218854 399896
rect 218234 399576 218854 399660
rect 218234 399340 218266 399576
rect 218502 399340 218586 399576
rect 218822 399340 218854 399576
rect 218234 363896 218854 399340
rect 218234 363660 218266 363896
rect 218502 363660 218586 363896
rect 218822 363660 218854 363896
rect 218234 363576 218854 363660
rect 218234 363340 218266 363576
rect 218502 363340 218586 363576
rect 218822 363340 218854 363576
rect 218234 327896 218854 363340
rect 218234 327660 218266 327896
rect 218502 327660 218586 327896
rect 218822 327660 218854 327896
rect 218234 327576 218854 327660
rect 218234 327340 218266 327576
rect 218502 327340 218586 327576
rect 218822 327340 218854 327576
rect 218234 291896 218854 327340
rect 218234 291660 218266 291896
rect 218502 291660 218586 291896
rect 218822 291660 218854 291896
rect 218234 291576 218854 291660
rect 218234 291340 218266 291576
rect 218502 291340 218586 291576
rect 218822 291340 218854 291576
rect 218234 255896 218854 291340
rect 218234 255660 218266 255896
rect 218502 255660 218586 255896
rect 218822 255660 218854 255896
rect 218234 255576 218854 255660
rect 218234 255340 218266 255576
rect 218502 255340 218586 255576
rect 218822 255340 218854 255576
rect 218234 219896 218854 255340
rect 218234 219660 218266 219896
rect 218502 219660 218586 219896
rect 218822 219660 218854 219896
rect 218234 219576 218854 219660
rect 218234 219340 218266 219576
rect 218502 219340 218586 219576
rect 218822 219340 218854 219576
rect 218234 183896 218854 219340
rect 218234 183660 218266 183896
rect 218502 183660 218586 183896
rect 218822 183660 218854 183896
rect 218234 183576 218854 183660
rect 218234 183340 218266 183576
rect 218502 183340 218586 183576
rect 218822 183340 218854 183576
rect 218234 147896 218854 183340
rect 218234 147660 218266 147896
rect 218502 147660 218586 147896
rect 218822 147660 218854 147896
rect 218234 147576 218854 147660
rect 218234 147340 218266 147576
rect 218502 147340 218586 147576
rect 218822 147340 218854 147576
rect 218234 111896 218854 147340
rect 218234 111660 218266 111896
rect 218502 111660 218586 111896
rect 218822 111660 218854 111896
rect 218234 111576 218854 111660
rect 218234 111340 218266 111576
rect 218502 111340 218586 111576
rect 218822 111340 218854 111576
rect 218234 75896 218854 111340
rect 218234 75660 218266 75896
rect 218502 75660 218586 75896
rect 218822 75660 218854 75896
rect 218234 75576 218854 75660
rect 218234 75340 218266 75576
rect 218502 75340 218586 75576
rect 218822 75340 218854 75576
rect 218234 39896 218854 75340
rect 218234 39660 218266 39896
rect 218502 39660 218586 39896
rect 218822 39660 218854 39896
rect 218234 39576 218854 39660
rect 218234 39340 218266 39576
rect 218502 39340 218586 39576
rect 218822 39340 218854 39576
rect 218234 3896 218854 39340
rect 218234 3660 218266 3896
rect 218502 3660 218586 3896
rect 218822 3660 218854 3896
rect 218234 3576 218854 3660
rect 218234 3340 218266 3576
rect 218502 3340 218586 3576
rect 218822 3340 218854 3576
rect 218234 -1304 218854 3340
rect 218234 -1540 218266 -1304
rect 218502 -1540 218586 -1304
rect 218822 -1540 218854 -1304
rect 218234 -1624 218854 -1540
rect 218234 -1860 218266 -1624
rect 218502 -1860 218586 -1624
rect 218822 -1860 218854 -1624
rect 218234 -7652 218854 -1860
rect 219474 706760 220094 711592
rect 219474 706524 219506 706760
rect 219742 706524 219826 706760
rect 220062 706524 220094 706760
rect 219474 706440 220094 706524
rect 219474 706204 219506 706440
rect 219742 706204 219826 706440
rect 220062 706204 220094 706440
rect 219474 689136 220094 706204
rect 219474 688900 219506 689136
rect 219742 688900 219826 689136
rect 220062 688900 220094 689136
rect 219474 688816 220094 688900
rect 219474 688580 219506 688816
rect 219742 688580 219826 688816
rect 220062 688580 220094 688816
rect 219474 653136 220094 688580
rect 219474 652900 219506 653136
rect 219742 652900 219826 653136
rect 220062 652900 220094 653136
rect 219474 652816 220094 652900
rect 219474 652580 219506 652816
rect 219742 652580 219826 652816
rect 220062 652580 220094 652816
rect 219474 617136 220094 652580
rect 219474 616900 219506 617136
rect 219742 616900 219826 617136
rect 220062 616900 220094 617136
rect 219474 616816 220094 616900
rect 219474 616580 219506 616816
rect 219742 616580 219826 616816
rect 220062 616580 220094 616816
rect 219474 581136 220094 616580
rect 219474 580900 219506 581136
rect 219742 580900 219826 581136
rect 220062 580900 220094 581136
rect 219474 580816 220094 580900
rect 219474 580580 219506 580816
rect 219742 580580 219826 580816
rect 220062 580580 220094 580816
rect 219474 545136 220094 580580
rect 219474 544900 219506 545136
rect 219742 544900 219826 545136
rect 220062 544900 220094 545136
rect 219474 544816 220094 544900
rect 219474 544580 219506 544816
rect 219742 544580 219826 544816
rect 220062 544580 220094 544816
rect 219474 509136 220094 544580
rect 219474 508900 219506 509136
rect 219742 508900 219826 509136
rect 220062 508900 220094 509136
rect 219474 508816 220094 508900
rect 219474 508580 219506 508816
rect 219742 508580 219826 508816
rect 220062 508580 220094 508816
rect 219474 473136 220094 508580
rect 219474 472900 219506 473136
rect 219742 472900 219826 473136
rect 220062 472900 220094 473136
rect 219474 472816 220094 472900
rect 219474 472580 219506 472816
rect 219742 472580 219826 472816
rect 220062 472580 220094 472816
rect 219474 437136 220094 472580
rect 219474 436900 219506 437136
rect 219742 436900 219826 437136
rect 220062 436900 220094 437136
rect 219474 436816 220094 436900
rect 219474 436580 219506 436816
rect 219742 436580 219826 436816
rect 220062 436580 220094 436816
rect 219474 401136 220094 436580
rect 219474 400900 219506 401136
rect 219742 400900 219826 401136
rect 220062 400900 220094 401136
rect 219474 400816 220094 400900
rect 219474 400580 219506 400816
rect 219742 400580 219826 400816
rect 220062 400580 220094 400816
rect 219474 365136 220094 400580
rect 219474 364900 219506 365136
rect 219742 364900 219826 365136
rect 220062 364900 220094 365136
rect 219474 364816 220094 364900
rect 219474 364580 219506 364816
rect 219742 364580 219826 364816
rect 220062 364580 220094 364816
rect 219474 329136 220094 364580
rect 219474 328900 219506 329136
rect 219742 328900 219826 329136
rect 220062 328900 220094 329136
rect 219474 328816 220094 328900
rect 219474 328580 219506 328816
rect 219742 328580 219826 328816
rect 220062 328580 220094 328816
rect 219474 293136 220094 328580
rect 219474 292900 219506 293136
rect 219742 292900 219826 293136
rect 220062 292900 220094 293136
rect 219474 292816 220094 292900
rect 219474 292580 219506 292816
rect 219742 292580 219826 292816
rect 220062 292580 220094 292816
rect 219474 257136 220094 292580
rect 219474 256900 219506 257136
rect 219742 256900 219826 257136
rect 220062 256900 220094 257136
rect 219474 256816 220094 256900
rect 219474 256580 219506 256816
rect 219742 256580 219826 256816
rect 220062 256580 220094 256816
rect 219474 221136 220094 256580
rect 219474 220900 219506 221136
rect 219742 220900 219826 221136
rect 220062 220900 220094 221136
rect 219474 220816 220094 220900
rect 219474 220580 219506 220816
rect 219742 220580 219826 220816
rect 220062 220580 220094 220816
rect 219474 185136 220094 220580
rect 219474 184900 219506 185136
rect 219742 184900 219826 185136
rect 220062 184900 220094 185136
rect 219474 184816 220094 184900
rect 219474 184580 219506 184816
rect 219742 184580 219826 184816
rect 220062 184580 220094 184816
rect 219474 149136 220094 184580
rect 219474 148900 219506 149136
rect 219742 148900 219826 149136
rect 220062 148900 220094 149136
rect 219474 148816 220094 148900
rect 219474 148580 219506 148816
rect 219742 148580 219826 148816
rect 220062 148580 220094 148816
rect 219474 113136 220094 148580
rect 219474 112900 219506 113136
rect 219742 112900 219826 113136
rect 220062 112900 220094 113136
rect 219474 112816 220094 112900
rect 219474 112580 219506 112816
rect 219742 112580 219826 112816
rect 220062 112580 220094 112816
rect 219474 77136 220094 112580
rect 219474 76900 219506 77136
rect 219742 76900 219826 77136
rect 220062 76900 220094 77136
rect 219474 76816 220094 76900
rect 219474 76580 219506 76816
rect 219742 76580 219826 76816
rect 220062 76580 220094 76816
rect 219474 41136 220094 76580
rect 219474 40900 219506 41136
rect 219742 40900 219826 41136
rect 220062 40900 220094 41136
rect 219474 40816 220094 40900
rect 219474 40580 219506 40816
rect 219742 40580 219826 40816
rect 220062 40580 220094 40816
rect 219474 5136 220094 40580
rect 219474 4900 219506 5136
rect 219742 4900 219826 5136
rect 220062 4900 220094 5136
rect 219474 4816 220094 4900
rect 219474 4580 219506 4816
rect 219742 4580 219826 4816
rect 220062 4580 220094 4816
rect 219474 -2264 220094 4580
rect 219474 -2500 219506 -2264
rect 219742 -2500 219826 -2264
rect 220062 -2500 220094 -2264
rect 219474 -2584 220094 -2500
rect 219474 -2820 219506 -2584
rect 219742 -2820 219826 -2584
rect 220062 -2820 220094 -2584
rect 219474 -7652 220094 -2820
rect 220714 707720 221334 711592
rect 220714 707484 220746 707720
rect 220982 707484 221066 707720
rect 221302 707484 221334 707720
rect 220714 707400 221334 707484
rect 220714 707164 220746 707400
rect 220982 707164 221066 707400
rect 221302 707164 221334 707400
rect 220714 690376 221334 707164
rect 220714 690140 220746 690376
rect 220982 690140 221066 690376
rect 221302 690140 221334 690376
rect 220714 690056 221334 690140
rect 220714 689820 220746 690056
rect 220982 689820 221066 690056
rect 221302 689820 221334 690056
rect 220714 654376 221334 689820
rect 220714 654140 220746 654376
rect 220982 654140 221066 654376
rect 221302 654140 221334 654376
rect 220714 654056 221334 654140
rect 220714 653820 220746 654056
rect 220982 653820 221066 654056
rect 221302 653820 221334 654056
rect 220714 618376 221334 653820
rect 220714 618140 220746 618376
rect 220982 618140 221066 618376
rect 221302 618140 221334 618376
rect 220714 618056 221334 618140
rect 220714 617820 220746 618056
rect 220982 617820 221066 618056
rect 221302 617820 221334 618056
rect 220714 582376 221334 617820
rect 220714 582140 220746 582376
rect 220982 582140 221066 582376
rect 221302 582140 221334 582376
rect 220714 582056 221334 582140
rect 220714 581820 220746 582056
rect 220982 581820 221066 582056
rect 221302 581820 221334 582056
rect 220714 546376 221334 581820
rect 220714 546140 220746 546376
rect 220982 546140 221066 546376
rect 221302 546140 221334 546376
rect 220714 546056 221334 546140
rect 220714 545820 220746 546056
rect 220982 545820 221066 546056
rect 221302 545820 221334 546056
rect 220714 510376 221334 545820
rect 220714 510140 220746 510376
rect 220982 510140 221066 510376
rect 221302 510140 221334 510376
rect 220714 510056 221334 510140
rect 220714 509820 220746 510056
rect 220982 509820 221066 510056
rect 221302 509820 221334 510056
rect 220714 474376 221334 509820
rect 220714 474140 220746 474376
rect 220982 474140 221066 474376
rect 221302 474140 221334 474376
rect 220714 474056 221334 474140
rect 220714 473820 220746 474056
rect 220982 473820 221066 474056
rect 221302 473820 221334 474056
rect 220714 438376 221334 473820
rect 220714 438140 220746 438376
rect 220982 438140 221066 438376
rect 221302 438140 221334 438376
rect 220714 438056 221334 438140
rect 220714 437820 220746 438056
rect 220982 437820 221066 438056
rect 221302 437820 221334 438056
rect 220714 402376 221334 437820
rect 220714 402140 220746 402376
rect 220982 402140 221066 402376
rect 221302 402140 221334 402376
rect 220714 402056 221334 402140
rect 220714 401820 220746 402056
rect 220982 401820 221066 402056
rect 221302 401820 221334 402056
rect 220714 366376 221334 401820
rect 220714 366140 220746 366376
rect 220982 366140 221066 366376
rect 221302 366140 221334 366376
rect 220714 366056 221334 366140
rect 220714 365820 220746 366056
rect 220982 365820 221066 366056
rect 221302 365820 221334 366056
rect 220714 330376 221334 365820
rect 220714 330140 220746 330376
rect 220982 330140 221066 330376
rect 221302 330140 221334 330376
rect 220714 330056 221334 330140
rect 220714 329820 220746 330056
rect 220982 329820 221066 330056
rect 221302 329820 221334 330056
rect 220714 294376 221334 329820
rect 220714 294140 220746 294376
rect 220982 294140 221066 294376
rect 221302 294140 221334 294376
rect 220714 294056 221334 294140
rect 220714 293820 220746 294056
rect 220982 293820 221066 294056
rect 221302 293820 221334 294056
rect 220714 258376 221334 293820
rect 220714 258140 220746 258376
rect 220982 258140 221066 258376
rect 221302 258140 221334 258376
rect 220714 258056 221334 258140
rect 220714 257820 220746 258056
rect 220982 257820 221066 258056
rect 221302 257820 221334 258056
rect 220714 222376 221334 257820
rect 220714 222140 220746 222376
rect 220982 222140 221066 222376
rect 221302 222140 221334 222376
rect 220714 222056 221334 222140
rect 220714 221820 220746 222056
rect 220982 221820 221066 222056
rect 221302 221820 221334 222056
rect 220714 186376 221334 221820
rect 220714 186140 220746 186376
rect 220982 186140 221066 186376
rect 221302 186140 221334 186376
rect 220714 186056 221334 186140
rect 220714 185820 220746 186056
rect 220982 185820 221066 186056
rect 221302 185820 221334 186056
rect 220714 150376 221334 185820
rect 220714 150140 220746 150376
rect 220982 150140 221066 150376
rect 221302 150140 221334 150376
rect 220714 150056 221334 150140
rect 220714 149820 220746 150056
rect 220982 149820 221066 150056
rect 221302 149820 221334 150056
rect 220714 114376 221334 149820
rect 220714 114140 220746 114376
rect 220982 114140 221066 114376
rect 221302 114140 221334 114376
rect 220714 114056 221334 114140
rect 220714 113820 220746 114056
rect 220982 113820 221066 114056
rect 221302 113820 221334 114056
rect 220714 78376 221334 113820
rect 220714 78140 220746 78376
rect 220982 78140 221066 78376
rect 221302 78140 221334 78376
rect 220714 78056 221334 78140
rect 220714 77820 220746 78056
rect 220982 77820 221066 78056
rect 221302 77820 221334 78056
rect 220714 42376 221334 77820
rect 220714 42140 220746 42376
rect 220982 42140 221066 42376
rect 221302 42140 221334 42376
rect 220714 42056 221334 42140
rect 220714 41820 220746 42056
rect 220982 41820 221066 42056
rect 221302 41820 221334 42056
rect 220714 6376 221334 41820
rect 220714 6140 220746 6376
rect 220982 6140 221066 6376
rect 221302 6140 221334 6376
rect 220714 6056 221334 6140
rect 220714 5820 220746 6056
rect 220982 5820 221066 6056
rect 221302 5820 221334 6056
rect 220714 -3224 221334 5820
rect 220714 -3460 220746 -3224
rect 220982 -3460 221066 -3224
rect 221302 -3460 221334 -3224
rect 220714 -3544 221334 -3460
rect 220714 -3780 220746 -3544
rect 220982 -3780 221066 -3544
rect 221302 -3780 221334 -3544
rect 220714 -7652 221334 -3780
rect 221954 708680 222574 711592
rect 221954 708444 221986 708680
rect 222222 708444 222306 708680
rect 222542 708444 222574 708680
rect 221954 708360 222574 708444
rect 221954 708124 221986 708360
rect 222222 708124 222306 708360
rect 222542 708124 222574 708360
rect 221954 691616 222574 708124
rect 221954 691380 221986 691616
rect 222222 691380 222306 691616
rect 222542 691380 222574 691616
rect 221954 691296 222574 691380
rect 221954 691060 221986 691296
rect 222222 691060 222306 691296
rect 222542 691060 222574 691296
rect 221954 655616 222574 691060
rect 221954 655380 221986 655616
rect 222222 655380 222306 655616
rect 222542 655380 222574 655616
rect 221954 655296 222574 655380
rect 221954 655060 221986 655296
rect 222222 655060 222306 655296
rect 222542 655060 222574 655296
rect 221954 619616 222574 655060
rect 221954 619380 221986 619616
rect 222222 619380 222306 619616
rect 222542 619380 222574 619616
rect 221954 619296 222574 619380
rect 221954 619060 221986 619296
rect 222222 619060 222306 619296
rect 222542 619060 222574 619296
rect 221954 583616 222574 619060
rect 221954 583380 221986 583616
rect 222222 583380 222306 583616
rect 222542 583380 222574 583616
rect 221954 583296 222574 583380
rect 221954 583060 221986 583296
rect 222222 583060 222306 583296
rect 222542 583060 222574 583296
rect 221954 547616 222574 583060
rect 221954 547380 221986 547616
rect 222222 547380 222306 547616
rect 222542 547380 222574 547616
rect 221954 547296 222574 547380
rect 221954 547060 221986 547296
rect 222222 547060 222306 547296
rect 222542 547060 222574 547296
rect 221954 511616 222574 547060
rect 221954 511380 221986 511616
rect 222222 511380 222306 511616
rect 222542 511380 222574 511616
rect 221954 511296 222574 511380
rect 221954 511060 221986 511296
rect 222222 511060 222306 511296
rect 222542 511060 222574 511296
rect 221954 475616 222574 511060
rect 221954 475380 221986 475616
rect 222222 475380 222306 475616
rect 222542 475380 222574 475616
rect 221954 475296 222574 475380
rect 221954 475060 221986 475296
rect 222222 475060 222306 475296
rect 222542 475060 222574 475296
rect 221954 439616 222574 475060
rect 221954 439380 221986 439616
rect 222222 439380 222306 439616
rect 222542 439380 222574 439616
rect 221954 439296 222574 439380
rect 221954 439060 221986 439296
rect 222222 439060 222306 439296
rect 222542 439060 222574 439296
rect 221954 403616 222574 439060
rect 221954 403380 221986 403616
rect 222222 403380 222306 403616
rect 222542 403380 222574 403616
rect 221954 403296 222574 403380
rect 221954 403060 221986 403296
rect 222222 403060 222306 403296
rect 222542 403060 222574 403296
rect 221954 367616 222574 403060
rect 221954 367380 221986 367616
rect 222222 367380 222306 367616
rect 222542 367380 222574 367616
rect 221954 367296 222574 367380
rect 221954 367060 221986 367296
rect 222222 367060 222306 367296
rect 222542 367060 222574 367296
rect 221954 331616 222574 367060
rect 221954 331380 221986 331616
rect 222222 331380 222306 331616
rect 222542 331380 222574 331616
rect 221954 331296 222574 331380
rect 221954 331060 221986 331296
rect 222222 331060 222306 331296
rect 222542 331060 222574 331296
rect 221954 295616 222574 331060
rect 221954 295380 221986 295616
rect 222222 295380 222306 295616
rect 222542 295380 222574 295616
rect 221954 295296 222574 295380
rect 221954 295060 221986 295296
rect 222222 295060 222306 295296
rect 222542 295060 222574 295296
rect 221954 259616 222574 295060
rect 221954 259380 221986 259616
rect 222222 259380 222306 259616
rect 222542 259380 222574 259616
rect 221954 259296 222574 259380
rect 221954 259060 221986 259296
rect 222222 259060 222306 259296
rect 222542 259060 222574 259296
rect 221954 223616 222574 259060
rect 221954 223380 221986 223616
rect 222222 223380 222306 223616
rect 222542 223380 222574 223616
rect 221954 223296 222574 223380
rect 221954 223060 221986 223296
rect 222222 223060 222306 223296
rect 222542 223060 222574 223296
rect 221954 187616 222574 223060
rect 221954 187380 221986 187616
rect 222222 187380 222306 187616
rect 222542 187380 222574 187616
rect 221954 187296 222574 187380
rect 221954 187060 221986 187296
rect 222222 187060 222306 187296
rect 222542 187060 222574 187296
rect 221954 151616 222574 187060
rect 221954 151380 221986 151616
rect 222222 151380 222306 151616
rect 222542 151380 222574 151616
rect 221954 151296 222574 151380
rect 221954 151060 221986 151296
rect 222222 151060 222306 151296
rect 222542 151060 222574 151296
rect 221954 115616 222574 151060
rect 221954 115380 221986 115616
rect 222222 115380 222306 115616
rect 222542 115380 222574 115616
rect 221954 115296 222574 115380
rect 221954 115060 221986 115296
rect 222222 115060 222306 115296
rect 222542 115060 222574 115296
rect 221954 79616 222574 115060
rect 221954 79380 221986 79616
rect 222222 79380 222306 79616
rect 222542 79380 222574 79616
rect 221954 79296 222574 79380
rect 221954 79060 221986 79296
rect 222222 79060 222306 79296
rect 222542 79060 222574 79296
rect 221954 43616 222574 79060
rect 221954 43380 221986 43616
rect 222222 43380 222306 43616
rect 222542 43380 222574 43616
rect 221954 43296 222574 43380
rect 221954 43060 221986 43296
rect 222222 43060 222306 43296
rect 222542 43060 222574 43296
rect 221954 7616 222574 43060
rect 221954 7380 221986 7616
rect 222222 7380 222306 7616
rect 222542 7380 222574 7616
rect 221954 7296 222574 7380
rect 221954 7060 221986 7296
rect 222222 7060 222306 7296
rect 222542 7060 222574 7296
rect 221954 -4184 222574 7060
rect 221954 -4420 221986 -4184
rect 222222 -4420 222306 -4184
rect 222542 -4420 222574 -4184
rect 221954 -4504 222574 -4420
rect 221954 -4740 221986 -4504
rect 222222 -4740 222306 -4504
rect 222542 -4740 222574 -4504
rect 221954 -7652 222574 -4740
rect 223194 709640 223814 711592
rect 223194 709404 223226 709640
rect 223462 709404 223546 709640
rect 223782 709404 223814 709640
rect 223194 709320 223814 709404
rect 223194 709084 223226 709320
rect 223462 709084 223546 709320
rect 223782 709084 223814 709320
rect 223194 692856 223814 709084
rect 223194 692620 223226 692856
rect 223462 692620 223546 692856
rect 223782 692620 223814 692856
rect 223194 692536 223814 692620
rect 223194 692300 223226 692536
rect 223462 692300 223546 692536
rect 223782 692300 223814 692536
rect 223194 656856 223814 692300
rect 223194 656620 223226 656856
rect 223462 656620 223546 656856
rect 223782 656620 223814 656856
rect 223194 656536 223814 656620
rect 223194 656300 223226 656536
rect 223462 656300 223546 656536
rect 223782 656300 223814 656536
rect 223194 620856 223814 656300
rect 223194 620620 223226 620856
rect 223462 620620 223546 620856
rect 223782 620620 223814 620856
rect 223194 620536 223814 620620
rect 223194 620300 223226 620536
rect 223462 620300 223546 620536
rect 223782 620300 223814 620536
rect 223194 584856 223814 620300
rect 223194 584620 223226 584856
rect 223462 584620 223546 584856
rect 223782 584620 223814 584856
rect 223194 584536 223814 584620
rect 223194 584300 223226 584536
rect 223462 584300 223546 584536
rect 223782 584300 223814 584536
rect 223194 548856 223814 584300
rect 223194 548620 223226 548856
rect 223462 548620 223546 548856
rect 223782 548620 223814 548856
rect 223194 548536 223814 548620
rect 223194 548300 223226 548536
rect 223462 548300 223546 548536
rect 223782 548300 223814 548536
rect 223194 512856 223814 548300
rect 223194 512620 223226 512856
rect 223462 512620 223546 512856
rect 223782 512620 223814 512856
rect 223194 512536 223814 512620
rect 223194 512300 223226 512536
rect 223462 512300 223546 512536
rect 223782 512300 223814 512536
rect 223194 476856 223814 512300
rect 223194 476620 223226 476856
rect 223462 476620 223546 476856
rect 223782 476620 223814 476856
rect 223194 476536 223814 476620
rect 223194 476300 223226 476536
rect 223462 476300 223546 476536
rect 223782 476300 223814 476536
rect 223194 440856 223814 476300
rect 223194 440620 223226 440856
rect 223462 440620 223546 440856
rect 223782 440620 223814 440856
rect 223194 440536 223814 440620
rect 223194 440300 223226 440536
rect 223462 440300 223546 440536
rect 223782 440300 223814 440536
rect 223194 404856 223814 440300
rect 223194 404620 223226 404856
rect 223462 404620 223546 404856
rect 223782 404620 223814 404856
rect 223194 404536 223814 404620
rect 223194 404300 223226 404536
rect 223462 404300 223546 404536
rect 223782 404300 223814 404536
rect 223194 368856 223814 404300
rect 223194 368620 223226 368856
rect 223462 368620 223546 368856
rect 223782 368620 223814 368856
rect 223194 368536 223814 368620
rect 223194 368300 223226 368536
rect 223462 368300 223546 368536
rect 223782 368300 223814 368536
rect 223194 332856 223814 368300
rect 223194 332620 223226 332856
rect 223462 332620 223546 332856
rect 223782 332620 223814 332856
rect 223194 332536 223814 332620
rect 223194 332300 223226 332536
rect 223462 332300 223546 332536
rect 223782 332300 223814 332536
rect 223194 296856 223814 332300
rect 223194 296620 223226 296856
rect 223462 296620 223546 296856
rect 223782 296620 223814 296856
rect 223194 296536 223814 296620
rect 223194 296300 223226 296536
rect 223462 296300 223546 296536
rect 223782 296300 223814 296536
rect 223194 260856 223814 296300
rect 223194 260620 223226 260856
rect 223462 260620 223546 260856
rect 223782 260620 223814 260856
rect 223194 260536 223814 260620
rect 223194 260300 223226 260536
rect 223462 260300 223546 260536
rect 223782 260300 223814 260536
rect 223194 224856 223814 260300
rect 223194 224620 223226 224856
rect 223462 224620 223546 224856
rect 223782 224620 223814 224856
rect 223194 224536 223814 224620
rect 223194 224300 223226 224536
rect 223462 224300 223546 224536
rect 223782 224300 223814 224536
rect 223194 188856 223814 224300
rect 223194 188620 223226 188856
rect 223462 188620 223546 188856
rect 223782 188620 223814 188856
rect 223194 188536 223814 188620
rect 223194 188300 223226 188536
rect 223462 188300 223546 188536
rect 223782 188300 223814 188536
rect 223194 152856 223814 188300
rect 223194 152620 223226 152856
rect 223462 152620 223546 152856
rect 223782 152620 223814 152856
rect 223194 152536 223814 152620
rect 223194 152300 223226 152536
rect 223462 152300 223546 152536
rect 223782 152300 223814 152536
rect 223194 116856 223814 152300
rect 223194 116620 223226 116856
rect 223462 116620 223546 116856
rect 223782 116620 223814 116856
rect 223194 116536 223814 116620
rect 223194 116300 223226 116536
rect 223462 116300 223546 116536
rect 223782 116300 223814 116536
rect 223194 80856 223814 116300
rect 223194 80620 223226 80856
rect 223462 80620 223546 80856
rect 223782 80620 223814 80856
rect 223194 80536 223814 80620
rect 223194 80300 223226 80536
rect 223462 80300 223546 80536
rect 223782 80300 223814 80536
rect 223194 44856 223814 80300
rect 223194 44620 223226 44856
rect 223462 44620 223546 44856
rect 223782 44620 223814 44856
rect 223194 44536 223814 44620
rect 223194 44300 223226 44536
rect 223462 44300 223546 44536
rect 223782 44300 223814 44536
rect 223194 8856 223814 44300
rect 223194 8620 223226 8856
rect 223462 8620 223546 8856
rect 223782 8620 223814 8856
rect 223194 8536 223814 8620
rect 223194 8300 223226 8536
rect 223462 8300 223546 8536
rect 223782 8300 223814 8536
rect 223194 -5144 223814 8300
rect 223194 -5380 223226 -5144
rect 223462 -5380 223546 -5144
rect 223782 -5380 223814 -5144
rect 223194 -5464 223814 -5380
rect 223194 -5700 223226 -5464
rect 223462 -5700 223546 -5464
rect 223782 -5700 223814 -5464
rect 223194 -7652 223814 -5700
rect 224434 710600 225054 711592
rect 224434 710364 224466 710600
rect 224702 710364 224786 710600
rect 225022 710364 225054 710600
rect 224434 710280 225054 710364
rect 224434 710044 224466 710280
rect 224702 710044 224786 710280
rect 225022 710044 225054 710280
rect 224434 694096 225054 710044
rect 224434 693860 224466 694096
rect 224702 693860 224786 694096
rect 225022 693860 225054 694096
rect 224434 693776 225054 693860
rect 224434 693540 224466 693776
rect 224702 693540 224786 693776
rect 225022 693540 225054 693776
rect 224434 658096 225054 693540
rect 224434 657860 224466 658096
rect 224702 657860 224786 658096
rect 225022 657860 225054 658096
rect 224434 657776 225054 657860
rect 224434 657540 224466 657776
rect 224702 657540 224786 657776
rect 225022 657540 225054 657776
rect 224434 622096 225054 657540
rect 224434 621860 224466 622096
rect 224702 621860 224786 622096
rect 225022 621860 225054 622096
rect 224434 621776 225054 621860
rect 224434 621540 224466 621776
rect 224702 621540 224786 621776
rect 225022 621540 225054 621776
rect 224434 586096 225054 621540
rect 224434 585860 224466 586096
rect 224702 585860 224786 586096
rect 225022 585860 225054 586096
rect 224434 585776 225054 585860
rect 224434 585540 224466 585776
rect 224702 585540 224786 585776
rect 225022 585540 225054 585776
rect 224434 550096 225054 585540
rect 224434 549860 224466 550096
rect 224702 549860 224786 550096
rect 225022 549860 225054 550096
rect 224434 549776 225054 549860
rect 224434 549540 224466 549776
rect 224702 549540 224786 549776
rect 225022 549540 225054 549776
rect 224434 514096 225054 549540
rect 224434 513860 224466 514096
rect 224702 513860 224786 514096
rect 225022 513860 225054 514096
rect 224434 513776 225054 513860
rect 224434 513540 224466 513776
rect 224702 513540 224786 513776
rect 225022 513540 225054 513776
rect 224434 478096 225054 513540
rect 224434 477860 224466 478096
rect 224702 477860 224786 478096
rect 225022 477860 225054 478096
rect 224434 477776 225054 477860
rect 224434 477540 224466 477776
rect 224702 477540 224786 477776
rect 225022 477540 225054 477776
rect 224434 442096 225054 477540
rect 224434 441860 224466 442096
rect 224702 441860 224786 442096
rect 225022 441860 225054 442096
rect 224434 441776 225054 441860
rect 224434 441540 224466 441776
rect 224702 441540 224786 441776
rect 225022 441540 225054 441776
rect 224434 406096 225054 441540
rect 224434 405860 224466 406096
rect 224702 405860 224786 406096
rect 225022 405860 225054 406096
rect 224434 405776 225054 405860
rect 224434 405540 224466 405776
rect 224702 405540 224786 405776
rect 225022 405540 225054 405776
rect 224434 370096 225054 405540
rect 224434 369860 224466 370096
rect 224702 369860 224786 370096
rect 225022 369860 225054 370096
rect 224434 369776 225054 369860
rect 224434 369540 224466 369776
rect 224702 369540 224786 369776
rect 225022 369540 225054 369776
rect 224434 334096 225054 369540
rect 224434 333860 224466 334096
rect 224702 333860 224786 334096
rect 225022 333860 225054 334096
rect 224434 333776 225054 333860
rect 224434 333540 224466 333776
rect 224702 333540 224786 333776
rect 225022 333540 225054 333776
rect 224434 298096 225054 333540
rect 224434 297860 224466 298096
rect 224702 297860 224786 298096
rect 225022 297860 225054 298096
rect 224434 297776 225054 297860
rect 224434 297540 224466 297776
rect 224702 297540 224786 297776
rect 225022 297540 225054 297776
rect 224434 262096 225054 297540
rect 224434 261860 224466 262096
rect 224702 261860 224786 262096
rect 225022 261860 225054 262096
rect 224434 261776 225054 261860
rect 224434 261540 224466 261776
rect 224702 261540 224786 261776
rect 225022 261540 225054 261776
rect 224434 226096 225054 261540
rect 224434 225860 224466 226096
rect 224702 225860 224786 226096
rect 225022 225860 225054 226096
rect 224434 225776 225054 225860
rect 224434 225540 224466 225776
rect 224702 225540 224786 225776
rect 225022 225540 225054 225776
rect 224434 190096 225054 225540
rect 224434 189860 224466 190096
rect 224702 189860 224786 190096
rect 225022 189860 225054 190096
rect 224434 189776 225054 189860
rect 224434 189540 224466 189776
rect 224702 189540 224786 189776
rect 225022 189540 225054 189776
rect 224434 154096 225054 189540
rect 224434 153860 224466 154096
rect 224702 153860 224786 154096
rect 225022 153860 225054 154096
rect 224434 153776 225054 153860
rect 224434 153540 224466 153776
rect 224702 153540 224786 153776
rect 225022 153540 225054 153776
rect 224434 118096 225054 153540
rect 224434 117860 224466 118096
rect 224702 117860 224786 118096
rect 225022 117860 225054 118096
rect 224434 117776 225054 117860
rect 224434 117540 224466 117776
rect 224702 117540 224786 117776
rect 225022 117540 225054 117776
rect 224434 82096 225054 117540
rect 224434 81860 224466 82096
rect 224702 81860 224786 82096
rect 225022 81860 225054 82096
rect 224434 81776 225054 81860
rect 224434 81540 224466 81776
rect 224702 81540 224786 81776
rect 225022 81540 225054 81776
rect 224434 46096 225054 81540
rect 224434 45860 224466 46096
rect 224702 45860 224786 46096
rect 225022 45860 225054 46096
rect 224434 45776 225054 45860
rect 224434 45540 224466 45776
rect 224702 45540 224786 45776
rect 225022 45540 225054 45776
rect 224434 10096 225054 45540
rect 224434 9860 224466 10096
rect 224702 9860 224786 10096
rect 225022 9860 225054 10096
rect 224434 9776 225054 9860
rect 224434 9540 224466 9776
rect 224702 9540 224786 9776
rect 225022 9540 225054 9776
rect 224434 -6104 225054 9540
rect 224434 -6340 224466 -6104
rect 224702 -6340 224786 -6104
rect 225022 -6340 225054 -6104
rect 224434 -6424 225054 -6340
rect 224434 -6660 224466 -6424
rect 224702 -6660 224786 -6424
rect 225022 -6660 225054 -6424
rect 224434 -7652 225054 -6660
rect 225674 711560 226294 711592
rect 225674 711324 225706 711560
rect 225942 711324 226026 711560
rect 226262 711324 226294 711560
rect 225674 711240 226294 711324
rect 225674 711004 225706 711240
rect 225942 711004 226026 711240
rect 226262 711004 226294 711240
rect 225674 695336 226294 711004
rect 225674 695100 225706 695336
rect 225942 695100 226026 695336
rect 226262 695100 226294 695336
rect 225674 695016 226294 695100
rect 225674 694780 225706 695016
rect 225942 694780 226026 695016
rect 226262 694780 226294 695016
rect 225674 659336 226294 694780
rect 225674 659100 225706 659336
rect 225942 659100 226026 659336
rect 226262 659100 226294 659336
rect 225674 659016 226294 659100
rect 225674 658780 225706 659016
rect 225942 658780 226026 659016
rect 226262 658780 226294 659016
rect 225674 623336 226294 658780
rect 225674 623100 225706 623336
rect 225942 623100 226026 623336
rect 226262 623100 226294 623336
rect 225674 623016 226294 623100
rect 225674 622780 225706 623016
rect 225942 622780 226026 623016
rect 226262 622780 226294 623016
rect 225674 587336 226294 622780
rect 225674 587100 225706 587336
rect 225942 587100 226026 587336
rect 226262 587100 226294 587336
rect 225674 587016 226294 587100
rect 225674 586780 225706 587016
rect 225942 586780 226026 587016
rect 226262 586780 226294 587016
rect 225674 551336 226294 586780
rect 225674 551100 225706 551336
rect 225942 551100 226026 551336
rect 226262 551100 226294 551336
rect 225674 551016 226294 551100
rect 225674 550780 225706 551016
rect 225942 550780 226026 551016
rect 226262 550780 226294 551016
rect 225674 515336 226294 550780
rect 225674 515100 225706 515336
rect 225942 515100 226026 515336
rect 226262 515100 226294 515336
rect 225674 515016 226294 515100
rect 225674 514780 225706 515016
rect 225942 514780 226026 515016
rect 226262 514780 226294 515016
rect 225674 479336 226294 514780
rect 225674 479100 225706 479336
rect 225942 479100 226026 479336
rect 226262 479100 226294 479336
rect 225674 479016 226294 479100
rect 225674 478780 225706 479016
rect 225942 478780 226026 479016
rect 226262 478780 226294 479016
rect 225674 443336 226294 478780
rect 225674 443100 225706 443336
rect 225942 443100 226026 443336
rect 226262 443100 226294 443336
rect 225674 443016 226294 443100
rect 225674 442780 225706 443016
rect 225942 442780 226026 443016
rect 226262 442780 226294 443016
rect 225674 407336 226294 442780
rect 225674 407100 225706 407336
rect 225942 407100 226026 407336
rect 226262 407100 226294 407336
rect 225674 407016 226294 407100
rect 225674 406780 225706 407016
rect 225942 406780 226026 407016
rect 226262 406780 226294 407016
rect 225674 371336 226294 406780
rect 225674 371100 225706 371336
rect 225942 371100 226026 371336
rect 226262 371100 226294 371336
rect 225674 371016 226294 371100
rect 225674 370780 225706 371016
rect 225942 370780 226026 371016
rect 226262 370780 226294 371016
rect 225674 335336 226294 370780
rect 225674 335100 225706 335336
rect 225942 335100 226026 335336
rect 226262 335100 226294 335336
rect 225674 335016 226294 335100
rect 225674 334780 225706 335016
rect 225942 334780 226026 335016
rect 226262 334780 226294 335016
rect 225674 299336 226294 334780
rect 225674 299100 225706 299336
rect 225942 299100 226026 299336
rect 226262 299100 226294 299336
rect 225674 299016 226294 299100
rect 225674 298780 225706 299016
rect 225942 298780 226026 299016
rect 226262 298780 226294 299016
rect 225674 263336 226294 298780
rect 225674 263100 225706 263336
rect 225942 263100 226026 263336
rect 226262 263100 226294 263336
rect 225674 263016 226294 263100
rect 225674 262780 225706 263016
rect 225942 262780 226026 263016
rect 226262 262780 226294 263016
rect 225674 227336 226294 262780
rect 225674 227100 225706 227336
rect 225942 227100 226026 227336
rect 226262 227100 226294 227336
rect 225674 227016 226294 227100
rect 225674 226780 225706 227016
rect 225942 226780 226026 227016
rect 226262 226780 226294 227016
rect 225674 191336 226294 226780
rect 225674 191100 225706 191336
rect 225942 191100 226026 191336
rect 226262 191100 226294 191336
rect 225674 191016 226294 191100
rect 225674 190780 225706 191016
rect 225942 190780 226026 191016
rect 226262 190780 226294 191016
rect 225674 155336 226294 190780
rect 225674 155100 225706 155336
rect 225942 155100 226026 155336
rect 226262 155100 226294 155336
rect 225674 155016 226294 155100
rect 225674 154780 225706 155016
rect 225942 154780 226026 155016
rect 226262 154780 226294 155016
rect 225674 119336 226294 154780
rect 225674 119100 225706 119336
rect 225942 119100 226026 119336
rect 226262 119100 226294 119336
rect 225674 119016 226294 119100
rect 225674 118780 225706 119016
rect 225942 118780 226026 119016
rect 226262 118780 226294 119016
rect 225674 83336 226294 118780
rect 225674 83100 225706 83336
rect 225942 83100 226026 83336
rect 226262 83100 226294 83336
rect 225674 83016 226294 83100
rect 225674 82780 225706 83016
rect 225942 82780 226026 83016
rect 226262 82780 226294 83016
rect 225674 47336 226294 82780
rect 225674 47100 225706 47336
rect 225942 47100 226026 47336
rect 226262 47100 226294 47336
rect 225674 47016 226294 47100
rect 225674 46780 225706 47016
rect 225942 46780 226026 47016
rect 226262 46780 226294 47016
rect 225674 11336 226294 46780
rect 225674 11100 225706 11336
rect 225942 11100 226026 11336
rect 226262 11100 226294 11336
rect 225674 11016 226294 11100
rect 225674 10780 225706 11016
rect 225942 10780 226026 11016
rect 226262 10780 226294 11016
rect 225674 -7064 226294 10780
rect 225674 -7300 225706 -7064
rect 225942 -7300 226026 -7064
rect 226262 -7300 226294 -7064
rect 225674 -7384 226294 -7300
rect 225674 -7620 225706 -7384
rect 225942 -7620 226026 -7384
rect 226262 -7620 226294 -7384
rect 225674 -7652 226294 -7620
rect 252994 704840 253614 711592
rect 252994 704604 253026 704840
rect 253262 704604 253346 704840
rect 253582 704604 253614 704840
rect 252994 704520 253614 704604
rect 252994 704284 253026 704520
rect 253262 704284 253346 704520
rect 253582 704284 253614 704520
rect 252994 702568 253614 704284
rect 252994 702504 253032 702568
rect 253096 702504 253112 702568
rect 253176 702504 253192 702568
rect 253256 702504 253272 702568
rect 253336 702504 253352 702568
rect 253416 702504 253432 702568
rect 253496 702504 253512 702568
rect 253576 702504 253614 702568
rect 252994 702488 253614 702504
rect 252994 702424 253032 702488
rect 253096 702424 253112 702488
rect 253176 702424 253192 702488
rect 253256 702424 253272 702488
rect 253336 702424 253352 702488
rect 253416 702424 253432 702488
rect 253496 702424 253512 702488
rect 253576 702424 253614 702488
rect 252994 702408 253614 702424
rect 252994 702344 253032 702408
rect 253096 702344 253112 702408
rect 253176 702344 253192 702408
rect 253256 702344 253272 702408
rect 253336 702344 253352 702408
rect 253416 702344 253432 702408
rect 253496 702344 253512 702408
rect 253576 702344 253614 702408
rect 252994 702328 253614 702344
rect 252994 702264 253032 702328
rect 253096 702264 253112 702328
rect 253176 702264 253192 702328
rect 253256 702264 253272 702328
rect 253336 702264 253352 702328
rect 253416 702264 253432 702328
rect 253496 702264 253512 702328
rect 253576 702264 253614 702328
rect 252994 686656 253614 702264
rect 252994 686420 253026 686656
rect 253262 686420 253346 686656
rect 253582 686420 253614 686656
rect 252994 686336 253614 686420
rect 252994 686100 253026 686336
rect 253262 686100 253346 686336
rect 253582 686100 253614 686336
rect 252994 650656 253614 686100
rect 252994 650420 253026 650656
rect 253262 650420 253346 650656
rect 253582 650420 253614 650656
rect 252994 650336 253614 650420
rect 252994 650100 253026 650336
rect 253262 650100 253346 650336
rect 253582 650100 253614 650336
rect 252994 614656 253614 650100
rect 252994 614420 253026 614656
rect 253262 614420 253346 614656
rect 253582 614420 253614 614656
rect 252994 614336 253614 614420
rect 252994 614100 253026 614336
rect 253262 614100 253346 614336
rect 253582 614100 253614 614336
rect 252994 578656 253614 614100
rect 252994 578420 253026 578656
rect 253262 578420 253346 578656
rect 253582 578420 253614 578656
rect 252994 578336 253614 578420
rect 252994 578100 253026 578336
rect 253262 578100 253346 578336
rect 253582 578100 253614 578336
rect 252994 542656 253614 578100
rect 252994 542420 253026 542656
rect 253262 542420 253346 542656
rect 253582 542420 253614 542656
rect 252994 542336 253614 542420
rect 252994 542100 253026 542336
rect 253262 542100 253346 542336
rect 253582 542100 253614 542336
rect 252994 506656 253614 542100
rect 252994 506420 253026 506656
rect 253262 506420 253346 506656
rect 253582 506420 253614 506656
rect 252994 506336 253614 506420
rect 252994 506100 253026 506336
rect 253262 506100 253346 506336
rect 253582 506100 253614 506336
rect 252994 470656 253614 506100
rect 252994 470420 253026 470656
rect 253262 470420 253346 470656
rect 253582 470420 253614 470656
rect 252994 470336 253614 470420
rect 252994 470100 253026 470336
rect 253262 470100 253346 470336
rect 253582 470100 253614 470336
rect 252994 434656 253614 470100
rect 252994 434420 253026 434656
rect 253262 434420 253346 434656
rect 253582 434420 253614 434656
rect 252994 434336 253614 434420
rect 252994 434100 253026 434336
rect 253262 434100 253346 434336
rect 253582 434100 253614 434336
rect 252994 398656 253614 434100
rect 252994 398420 253026 398656
rect 253262 398420 253346 398656
rect 253582 398420 253614 398656
rect 252994 398336 253614 398420
rect 252994 398100 253026 398336
rect 253262 398100 253346 398336
rect 253582 398100 253614 398336
rect 252994 362656 253614 398100
rect 252994 362420 253026 362656
rect 253262 362420 253346 362656
rect 253582 362420 253614 362656
rect 252994 362336 253614 362420
rect 252994 362100 253026 362336
rect 253262 362100 253346 362336
rect 253582 362100 253614 362336
rect 252994 326656 253614 362100
rect 252994 326420 253026 326656
rect 253262 326420 253346 326656
rect 253582 326420 253614 326656
rect 252994 326336 253614 326420
rect 252994 326100 253026 326336
rect 253262 326100 253346 326336
rect 253582 326100 253614 326336
rect 252994 290656 253614 326100
rect 252994 290420 253026 290656
rect 253262 290420 253346 290656
rect 253582 290420 253614 290656
rect 252994 290336 253614 290420
rect 252994 290100 253026 290336
rect 253262 290100 253346 290336
rect 253582 290100 253614 290336
rect 252994 254656 253614 290100
rect 252994 254420 253026 254656
rect 253262 254420 253346 254656
rect 253582 254420 253614 254656
rect 252994 254336 253614 254420
rect 252994 254100 253026 254336
rect 253262 254100 253346 254336
rect 253582 254100 253614 254336
rect 252994 218656 253614 254100
rect 252994 218420 253026 218656
rect 253262 218420 253346 218656
rect 253582 218420 253614 218656
rect 252994 218336 253614 218420
rect 252994 218100 253026 218336
rect 253262 218100 253346 218336
rect 253582 218100 253614 218336
rect 252994 182656 253614 218100
rect 252994 182420 253026 182656
rect 253262 182420 253346 182656
rect 253582 182420 253614 182656
rect 252994 182336 253614 182420
rect 252994 182100 253026 182336
rect 253262 182100 253346 182336
rect 253582 182100 253614 182336
rect 252994 146656 253614 182100
rect 252994 146420 253026 146656
rect 253262 146420 253346 146656
rect 253582 146420 253614 146656
rect 252994 146336 253614 146420
rect 252994 146100 253026 146336
rect 253262 146100 253346 146336
rect 253582 146100 253614 146336
rect 252994 110656 253614 146100
rect 252994 110420 253026 110656
rect 253262 110420 253346 110656
rect 253582 110420 253614 110656
rect 252994 110336 253614 110420
rect 252994 110100 253026 110336
rect 253262 110100 253346 110336
rect 253582 110100 253614 110336
rect 252994 74656 253614 110100
rect 252994 74420 253026 74656
rect 253262 74420 253346 74656
rect 253582 74420 253614 74656
rect 252994 74336 253614 74420
rect 252994 74100 253026 74336
rect 253262 74100 253346 74336
rect 253582 74100 253614 74336
rect 252994 38656 253614 74100
rect 252994 38420 253026 38656
rect 253262 38420 253346 38656
rect 253582 38420 253614 38656
rect 252994 38336 253614 38420
rect 252994 38100 253026 38336
rect 253262 38100 253346 38336
rect 253582 38100 253614 38336
rect 252994 2656 253614 38100
rect 252994 2420 253026 2656
rect 253262 2420 253346 2656
rect 253582 2420 253614 2656
rect 252994 2336 253614 2420
rect 252994 2100 253026 2336
rect 253262 2100 253346 2336
rect 253582 2100 253614 2336
rect 252994 -344 253614 2100
rect 252994 -580 253026 -344
rect 253262 -580 253346 -344
rect 253582 -580 253614 -344
rect 252994 -664 253614 -580
rect 252994 -900 253026 -664
rect 253262 -900 253346 -664
rect 253582 -900 253614 -664
rect 252994 -7652 253614 -900
rect 254234 705800 254854 711592
rect 254234 705564 254266 705800
rect 254502 705564 254586 705800
rect 254822 705564 254854 705800
rect 254234 705480 254854 705564
rect 254234 705244 254266 705480
rect 254502 705244 254586 705480
rect 254822 705244 254854 705480
rect 254234 703336 254854 705244
rect 254234 703272 254272 703336
rect 254336 703272 254352 703336
rect 254416 703272 254432 703336
rect 254496 703272 254512 703336
rect 254576 703272 254592 703336
rect 254656 703272 254672 703336
rect 254736 703272 254752 703336
rect 254816 703272 254854 703336
rect 254234 703256 254854 703272
rect 254234 703192 254272 703256
rect 254336 703192 254352 703256
rect 254416 703192 254432 703256
rect 254496 703192 254512 703256
rect 254576 703192 254592 703256
rect 254656 703192 254672 703256
rect 254736 703192 254752 703256
rect 254816 703192 254854 703256
rect 254234 703176 254854 703192
rect 254234 703112 254272 703176
rect 254336 703112 254352 703176
rect 254416 703112 254432 703176
rect 254496 703112 254512 703176
rect 254576 703112 254592 703176
rect 254656 703112 254672 703176
rect 254736 703112 254752 703176
rect 254816 703112 254854 703176
rect 254234 703096 254854 703112
rect 254234 703032 254272 703096
rect 254336 703032 254352 703096
rect 254416 703032 254432 703096
rect 254496 703032 254512 703096
rect 254576 703032 254592 703096
rect 254656 703032 254672 703096
rect 254736 703032 254752 703096
rect 254816 703032 254854 703096
rect 254234 687896 254854 703032
rect 254234 687660 254266 687896
rect 254502 687660 254586 687896
rect 254822 687660 254854 687896
rect 254234 687576 254854 687660
rect 254234 687340 254266 687576
rect 254502 687340 254586 687576
rect 254822 687340 254854 687576
rect 254234 651896 254854 687340
rect 254234 651660 254266 651896
rect 254502 651660 254586 651896
rect 254822 651660 254854 651896
rect 254234 651576 254854 651660
rect 254234 651340 254266 651576
rect 254502 651340 254586 651576
rect 254822 651340 254854 651576
rect 254234 615896 254854 651340
rect 254234 615660 254266 615896
rect 254502 615660 254586 615896
rect 254822 615660 254854 615896
rect 254234 615576 254854 615660
rect 254234 615340 254266 615576
rect 254502 615340 254586 615576
rect 254822 615340 254854 615576
rect 254234 579896 254854 615340
rect 254234 579660 254266 579896
rect 254502 579660 254586 579896
rect 254822 579660 254854 579896
rect 254234 579576 254854 579660
rect 254234 579340 254266 579576
rect 254502 579340 254586 579576
rect 254822 579340 254854 579576
rect 254234 543896 254854 579340
rect 254234 543660 254266 543896
rect 254502 543660 254586 543896
rect 254822 543660 254854 543896
rect 254234 543576 254854 543660
rect 254234 543340 254266 543576
rect 254502 543340 254586 543576
rect 254822 543340 254854 543576
rect 254234 507896 254854 543340
rect 254234 507660 254266 507896
rect 254502 507660 254586 507896
rect 254822 507660 254854 507896
rect 254234 507576 254854 507660
rect 254234 507340 254266 507576
rect 254502 507340 254586 507576
rect 254822 507340 254854 507576
rect 254234 471896 254854 507340
rect 254234 471660 254266 471896
rect 254502 471660 254586 471896
rect 254822 471660 254854 471896
rect 254234 471576 254854 471660
rect 254234 471340 254266 471576
rect 254502 471340 254586 471576
rect 254822 471340 254854 471576
rect 254234 435896 254854 471340
rect 254234 435660 254266 435896
rect 254502 435660 254586 435896
rect 254822 435660 254854 435896
rect 254234 435576 254854 435660
rect 254234 435340 254266 435576
rect 254502 435340 254586 435576
rect 254822 435340 254854 435576
rect 254234 399896 254854 435340
rect 254234 399660 254266 399896
rect 254502 399660 254586 399896
rect 254822 399660 254854 399896
rect 254234 399576 254854 399660
rect 254234 399340 254266 399576
rect 254502 399340 254586 399576
rect 254822 399340 254854 399576
rect 254234 363896 254854 399340
rect 254234 363660 254266 363896
rect 254502 363660 254586 363896
rect 254822 363660 254854 363896
rect 254234 363576 254854 363660
rect 254234 363340 254266 363576
rect 254502 363340 254586 363576
rect 254822 363340 254854 363576
rect 254234 327896 254854 363340
rect 254234 327660 254266 327896
rect 254502 327660 254586 327896
rect 254822 327660 254854 327896
rect 254234 327576 254854 327660
rect 254234 327340 254266 327576
rect 254502 327340 254586 327576
rect 254822 327340 254854 327576
rect 254234 291896 254854 327340
rect 254234 291660 254266 291896
rect 254502 291660 254586 291896
rect 254822 291660 254854 291896
rect 254234 291576 254854 291660
rect 254234 291340 254266 291576
rect 254502 291340 254586 291576
rect 254822 291340 254854 291576
rect 254234 255896 254854 291340
rect 254234 255660 254266 255896
rect 254502 255660 254586 255896
rect 254822 255660 254854 255896
rect 254234 255576 254854 255660
rect 254234 255340 254266 255576
rect 254502 255340 254586 255576
rect 254822 255340 254854 255576
rect 254234 219896 254854 255340
rect 254234 219660 254266 219896
rect 254502 219660 254586 219896
rect 254822 219660 254854 219896
rect 254234 219576 254854 219660
rect 254234 219340 254266 219576
rect 254502 219340 254586 219576
rect 254822 219340 254854 219576
rect 254234 183896 254854 219340
rect 254234 183660 254266 183896
rect 254502 183660 254586 183896
rect 254822 183660 254854 183896
rect 254234 183576 254854 183660
rect 254234 183340 254266 183576
rect 254502 183340 254586 183576
rect 254822 183340 254854 183576
rect 254234 147896 254854 183340
rect 254234 147660 254266 147896
rect 254502 147660 254586 147896
rect 254822 147660 254854 147896
rect 254234 147576 254854 147660
rect 254234 147340 254266 147576
rect 254502 147340 254586 147576
rect 254822 147340 254854 147576
rect 254234 111896 254854 147340
rect 254234 111660 254266 111896
rect 254502 111660 254586 111896
rect 254822 111660 254854 111896
rect 254234 111576 254854 111660
rect 254234 111340 254266 111576
rect 254502 111340 254586 111576
rect 254822 111340 254854 111576
rect 254234 75896 254854 111340
rect 254234 75660 254266 75896
rect 254502 75660 254586 75896
rect 254822 75660 254854 75896
rect 254234 75576 254854 75660
rect 254234 75340 254266 75576
rect 254502 75340 254586 75576
rect 254822 75340 254854 75576
rect 254234 39896 254854 75340
rect 254234 39660 254266 39896
rect 254502 39660 254586 39896
rect 254822 39660 254854 39896
rect 254234 39576 254854 39660
rect 254234 39340 254266 39576
rect 254502 39340 254586 39576
rect 254822 39340 254854 39576
rect 254234 3896 254854 39340
rect 254234 3660 254266 3896
rect 254502 3660 254586 3896
rect 254822 3660 254854 3896
rect 254234 3576 254854 3660
rect 254234 3340 254266 3576
rect 254502 3340 254586 3576
rect 254822 3340 254854 3576
rect 254234 -1304 254854 3340
rect 254234 -1540 254266 -1304
rect 254502 -1540 254586 -1304
rect 254822 -1540 254854 -1304
rect 254234 -1624 254854 -1540
rect 254234 -1860 254266 -1624
rect 254502 -1860 254586 -1624
rect 254822 -1860 254854 -1624
rect 254234 -7652 254854 -1860
rect 255474 706760 256094 711592
rect 255474 706524 255506 706760
rect 255742 706524 255826 706760
rect 256062 706524 256094 706760
rect 255474 706440 256094 706524
rect 255474 706204 255506 706440
rect 255742 706204 255826 706440
rect 256062 706204 256094 706440
rect 255474 689136 256094 706204
rect 255474 688900 255506 689136
rect 255742 688900 255826 689136
rect 256062 688900 256094 689136
rect 255474 688816 256094 688900
rect 255474 688580 255506 688816
rect 255742 688580 255826 688816
rect 256062 688580 256094 688816
rect 255474 653136 256094 688580
rect 255474 652900 255506 653136
rect 255742 652900 255826 653136
rect 256062 652900 256094 653136
rect 255474 652816 256094 652900
rect 255474 652580 255506 652816
rect 255742 652580 255826 652816
rect 256062 652580 256094 652816
rect 255474 617136 256094 652580
rect 255474 616900 255506 617136
rect 255742 616900 255826 617136
rect 256062 616900 256094 617136
rect 255474 616816 256094 616900
rect 255474 616580 255506 616816
rect 255742 616580 255826 616816
rect 256062 616580 256094 616816
rect 255474 581136 256094 616580
rect 255474 580900 255506 581136
rect 255742 580900 255826 581136
rect 256062 580900 256094 581136
rect 255474 580816 256094 580900
rect 255474 580580 255506 580816
rect 255742 580580 255826 580816
rect 256062 580580 256094 580816
rect 255474 545136 256094 580580
rect 255474 544900 255506 545136
rect 255742 544900 255826 545136
rect 256062 544900 256094 545136
rect 255474 544816 256094 544900
rect 255474 544580 255506 544816
rect 255742 544580 255826 544816
rect 256062 544580 256094 544816
rect 255474 509136 256094 544580
rect 255474 508900 255506 509136
rect 255742 508900 255826 509136
rect 256062 508900 256094 509136
rect 255474 508816 256094 508900
rect 255474 508580 255506 508816
rect 255742 508580 255826 508816
rect 256062 508580 256094 508816
rect 255474 473136 256094 508580
rect 255474 472900 255506 473136
rect 255742 472900 255826 473136
rect 256062 472900 256094 473136
rect 255474 472816 256094 472900
rect 255474 472580 255506 472816
rect 255742 472580 255826 472816
rect 256062 472580 256094 472816
rect 255474 437136 256094 472580
rect 255474 436900 255506 437136
rect 255742 436900 255826 437136
rect 256062 436900 256094 437136
rect 255474 436816 256094 436900
rect 255474 436580 255506 436816
rect 255742 436580 255826 436816
rect 256062 436580 256094 436816
rect 255474 401136 256094 436580
rect 255474 400900 255506 401136
rect 255742 400900 255826 401136
rect 256062 400900 256094 401136
rect 255474 400816 256094 400900
rect 255474 400580 255506 400816
rect 255742 400580 255826 400816
rect 256062 400580 256094 400816
rect 255474 365136 256094 400580
rect 255474 364900 255506 365136
rect 255742 364900 255826 365136
rect 256062 364900 256094 365136
rect 255474 364816 256094 364900
rect 255474 364580 255506 364816
rect 255742 364580 255826 364816
rect 256062 364580 256094 364816
rect 255474 329136 256094 364580
rect 255474 328900 255506 329136
rect 255742 328900 255826 329136
rect 256062 328900 256094 329136
rect 255474 328816 256094 328900
rect 255474 328580 255506 328816
rect 255742 328580 255826 328816
rect 256062 328580 256094 328816
rect 255474 293136 256094 328580
rect 255474 292900 255506 293136
rect 255742 292900 255826 293136
rect 256062 292900 256094 293136
rect 255474 292816 256094 292900
rect 255474 292580 255506 292816
rect 255742 292580 255826 292816
rect 256062 292580 256094 292816
rect 255474 257136 256094 292580
rect 255474 256900 255506 257136
rect 255742 256900 255826 257136
rect 256062 256900 256094 257136
rect 255474 256816 256094 256900
rect 255474 256580 255506 256816
rect 255742 256580 255826 256816
rect 256062 256580 256094 256816
rect 255474 221136 256094 256580
rect 255474 220900 255506 221136
rect 255742 220900 255826 221136
rect 256062 220900 256094 221136
rect 255474 220816 256094 220900
rect 255474 220580 255506 220816
rect 255742 220580 255826 220816
rect 256062 220580 256094 220816
rect 255474 185136 256094 220580
rect 255474 184900 255506 185136
rect 255742 184900 255826 185136
rect 256062 184900 256094 185136
rect 255474 184816 256094 184900
rect 255474 184580 255506 184816
rect 255742 184580 255826 184816
rect 256062 184580 256094 184816
rect 255474 149136 256094 184580
rect 255474 148900 255506 149136
rect 255742 148900 255826 149136
rect 256062 148900 256094 149136
rect 255474 148816 256094 148900
rect 255474 148580 255506 148816
rect 255742 148580 255826 148816
rect 256062 148580 256094 148816
rect 255474 113136 256094 148580
rect 255474 112900 255506 113136
rect 255742 112900 255826 113136
rect 256062 112900 256094 113136
rect 255474 112816 256094 112900
rect 255474 112580 255506 112816
rect 255742 112580 255826 112816
rect 256062 112580 256094 112816
rect 255474 77136 256094 112580
rect 255474 76900 255506 77136
rect 255742 76900 255826 77136
rect 256062 76900 256094 77136
rect 255474 76816 256094 76900
rect 255474 76580 255506 76816
rect 255742 76580 255826 76816
rect 256062 76580 256094 76816
rect 255474 41136 256094 76580
rect 255474 40900 255506 41136
rect 255742 40900 255826 41136
rect 256062 40900 256094 41136
rect 255474 40816 256094 40900
rect 255474 40580 255506 40816
rect 255742 40580 255826 40816
rect 256062 40580 256094 40816
rect 255474 5136 256094 40580
rect 255474 4900 255506 5136
rect 255742 4900 255826 5136
rect 256062 4900 256094 5136
rect 255474 4816 256094 4900
rect 255474 4580 255506 4816
rect 255742 4580 255826 4816
rect 256062 4580 256094 4816
rect 255474 -2264 256094 4580
rect 255474 -2500 255506 -2264
rect 255742 -2500 255826 -2264
rect 256062 -2500 256094 -2264
rect 255474 -2584 256094 -2500
rect 255474 -2820 255506 -2584
rect 255742 -2820 255826 -2584
rect 256062 -2820 256094 -2584
rect 255474 -7652 256094 -2820
rect 256714 707720 257334 711592
rect 256714 707484 256746 707720
rect 256982 707484 257066 707720
rect 257302 707484 257334 707720
rect 256714 707400 257334 707484
rect 256714 707164 256746 707400
rect 256982 707164 257066 707400
rect 257302 707164 257334 707400
rect 256714 690376 257334 707164
rect 256714 690140 256746 690376
rect 256982 690140 257066 690376
rect 257302 690140 257334 690376
rect 256714 690056 257334 690140
rect 256714 689820 256746 690056
rect 256982 689820 257066 690056
rect 257302 689820 257334 690056
rect 256714 654376 257334 689820
rect 256714 654140 256746 654376
rect 256982 654140 257066 654376
rect 257302 654140 257334 654376
rect 256714 654056 257334 654140
rect 256714 653820 256746 654056
rect 256982 653820 257066 654056
rect 257302 653820 257334 654056
rect 256714 618376 257334 653820
rect 256714 618140 256746 618376
rect 256982 618140 257066 618376
rect 257302 618140 257334 618376
rect 256714 618056 257334 618140
rect 256714 617820 256746 618056
rect 256982 617820 257066 618056
rect 257302 617820 257334 618056
rect 256714 582376 257334 617820
rect 256714 582140 256746 582376
rect 256982 582140 257066 582376
rect 257302 582140 257334 582376
rect 256714 582056 257334 582140
rect 256714 581820 256746 582056
rect 256982 581820 257066 582056
rect 257302 581820 257334 582056
rect 256714 546376 257334 581820
rect 256714 546140 256746 546376
rect 256982 546140 257066 546376
rect 257302 546140 257334 546376
rect 256714 546056 257334 546140
rect 256714 545820 256746 546056
rect 256982 545820 257066 546056
rect 257302 545820 257334 546056
rect 256714 510376 257334 545820
rect 256714 510140 256746 510376
rect 256982 510140 257066 510376
rect 257302 510140 257334 510376
rect 256714 510056 257334 510140
rect 256714 509820 256746 510056
rect 256982 509820 257066 510056
rect 257302 509820 257334 510056
rect 256714 474376 257334 509820
rect 256714 474140 256746 474376
rect 256982 474140 257066 474376
rect 257302 474140 257334 474376
rect 256714 474056 257334 474140
rect 256714 473820 256746 474056
rect 256982 473820 257066 474056
rect 257302 473820 257334 474056
rect 256714 438376 257334 473820
rect 256714 438140 256746 438376
rect 256982 438140 257066 438376
rect 257302 438140 257334 438376
rect 256714 438056 257334 438140
rect 256714 437820 256746 438056
rect 256982 437820 257066 438056
rect 257302 437820 257334 438056
rect 256714 402376 257334 437820
rect 256714 402140 256746 402376
rect 256982 402140 257066 402376
rect 257302 402140 257334 402376
rect 256714 402056 257334 402140
rect 256714 401820 256746 402056
rect 256982 401820 257066 402056
rect 257302 401820 257334 402056
rect 256714 366376 257334 401820
rect 256714 366140 256746 366376
rect 256982 366140 257066 366376
rect 257302 366140 257334 366376
rect 256714 366056 257334 366140
rect 256714 365820 256746 366056
rect 256982 365820 257066 366056
rect 257302 365820 257334 366056
rect 256714 330376 257334 365820
rect 256714 330140 256746 330376
rect 256982 330140 257066 330376
rect 257302 330140 257334 330376
rect 256714 330056 257334 330140
rect 256714 329820 256746 330056
rect 256982 329820 257066 330056
rect 257302 329820 257334 330056
rect 256714 294376 257334 329820
rect 256714 294140 256746 294376
rect 256982 294140 257066 294376
rect 257302 294140 257334 294376
rect 256714 294056 257334 294140
rect 256714 293820 256746 294056
rect 256982 293820 257066 294056
rect 257302 293820 257334 294056
rect 256714 258376 257334 293820
rect 256714 258140 256746 258376
rect 256982 258140 257066 258376
rect 257302 258140 257334 258376
rect 256714 258056 257334 258140
rect 256714 257820 256746 258056
rect 256982 257820 257066 258056
rect 257302 257820 257334 258056
rect 256714 222376 257334 257820
rect 256714 222140 256746 222376
rect 256982 222140 257066 222376
rect 257302 222140 257334 222376
rect 256714 222056 257334 222140
rect 256714 221820 256746 222056
rect 256982 221820 257066 222056
rect 257302 221820 257334 222056
rect 256714 186376 257334 221820
rect 256714 186140 256746 186376
rect 256982 186140 257066 186376
rect 257302 186140 257334 186376
rect 256714 186056 257334 186140
rect 256714 185820 256746 186056
rect 256982 185820 257066 186056
rect 257302 185820 257334 186056
rect 256714 150376 257334 185820
rect 256714 150140 256746 150376
rect 256982 150140 257066 150376
rect 257302 150140 257334 150376
rect 256714 150056 257334 150140
rect 256714 149820 256746 150056
rect 256982 149820 257066 150056
rect 257302 149820 257334 150056
rect 256714 114376 257334 149820
rect 256714 114140 256746 114376
rect 256982 114140 257066 114376
rect 257302 114140 257334 114376
rect 256714 114056 257334 114140
rect 256714 113820 256746 114056
rect 256982 113820 257066 114056
rect 257302 113820 257334 114056
rect 256714 78376 257334 113820
rect 256714 78140 256746 78376
rect 256982 78140 257066 78376
rect 257302 78140 257334 78376
rect 256714 78056 257334 78140
rect 256714 77820 256746 78056
rect 256982 77820 257066 78056
rect 257302 77820 257334 78056
rect 256714 42376 257334 77820
rect 256714 42140 256746 42376
rect 256982 42140 257066 42376
rect 257302 42140 257334 42376
rect 256714 42056 257334 42140
rect 256714 41820 256746 42056
rect 256982 41820 257066 42056
rect 257302 41820 257334 42056
rect 256714 6376 257334 41820
rect 256714 6140 256746 6376
rect 256982 6140 257066 6376
rect 257302 6140 257334 6376
rect 256714 6056 257334 6140
rect 256714 5820 256746 6056
rect 256982 5820 257066 6056
rect 257302 5820 257334 6056
rect 256714 -3224 257334 5820
rect 256714 -3460 256746 -3224
rect 256982 -3460 257066 -3224
rect 257302 -3460 257334 -3224
rect 256714 -3544 257334 -3460
rect 256714 -3780 256746 -3544
rect 256982 -3780 257066 -3544
rect 257302 -3780 257334 -3544
rect 256714 -7652 257334 -3780
rect 257954 708680 258574 711592
rect 257954 708444 257986 708680
rect 258222 708444 258306 708680
rect 258542 708444 258574 708680
rect 257954 708360 258574 708444
rect 257954 708124 257986 708360
rect 258222 708124 258306 708360
rect 258542 708124 258574 708360
rect 257954 691616 258574 708124
rect 257954 691380 257986 691616
rect 258222 691380 258306 691616
rect 258542 691380 258574 691616
rect 257954 691296 258574 691380
rect 257954 691060 257986 691296
rect 258222 691060 258306 691296
rect 258542 691060 258574 691296
rect 257954 655616 258574 691060
rect 257954 655380 257986 655616
rect 258222 655380 258306 655616
rect 258542 655380 258574 655616
rect 257954 655296 258574 655380
rect 257954 655060 257986 655296
rect 258222 655060 258306 655296
rect 258542 655060 258574 655296
rect 257954 619616 258574 655060
rect 257954 619380 257986 619616
rect 258222 619380 258306 619616
rect 258542 619380 258574 619616
rect 257954 619296 258574 619380
rect 257954 619060 257986 619296
rect 258222 619060 258306 619296
rect 258542 619060 258574 619296
rect 257954 583616 258574 619060
rect 257954 583380 257986 583616
rect 258222 583380 258306 583616
rect 258542 583380 258574 583616
rect 257954 583296 258574 583380
rect 257954 583060 257986 583296
rect 258222 583060 258306 583296
rect 258542 583060 258574 583296
rect 257954 547616 258574 583060
rect 257954 547380 257986 547616
rect 258222 547380 258306 547616
rect 258542 547380 258574 547616
rect 257954 547296 258574 547380
rect 257954 547060 257986 547296
rect 258222 547060 258306 547296
rect 258542 547060 258574 547296
rect 257954 511616 258574 547060
rect 257954 511380 257986 511616
rect 258222 511380 258306 511616
rect 258542 511380 258574 511616
rect 257954 511296 258574 511380
rect 257954 511060 257986 511296
rect 258222 511060 258306 511296
rect 258542 511060 258574 511296
rect 257954 475616 258574 511060
rect 257954 475380 257986 475616
rect 258222 475380 258306 475616
rect 258542 475380 258574 475616
rect 257954 475296 258574 475380
rect 257954 475060 257986 475296
rect 258222 475060 258306 475296
rect 258542 475060 258574 475296
rect 257954 439616 258574 475060
rect 257954 439380 257986 439616
rect 258222 439380 258306 439616
rect 258542 439380 258574 439616
rect 257954 439296 258574 439380
rect 257954 439060 257986 439296
rect 258222 439060 258306 439296
rect 258542 439060 258574 439296
rect 257954 403616 258574 439060
rect 257954 403380 257986 403616
rect 258222 403380 258306 403616
rect 258542 403380 258574 403616
rect 257954 403296 258574 403380
rect 257954 403060 257986 403296
rect 258222 403060 258306 403296
rect 258542 403060 258574 403296
rect 257954 367616 258574 403060
rect 257954 367380 257986 367616
rect 258222 367380 258306 367616
rect 258542 367380 258574 367616
rect 257954 367296 258574 367380
rect 257954 367060 257986 367296
rect 258222 367060 258306 367296
rect 258542 367060 258574 367296
rect 257954 331616 258574 367060
rect 257954 331380 257986 331616
rect 258222 331380 258306 331616
rect 258542 331380 258574 331616
rect 257954 331296 258574 331380
rect 257954 331060 257986 331296
rect 258222 331060 258306 331296
rect 258542 331060 258574 331296
rect 257954 295616 258574 331060
rect 257954 295380 257986 295616
rect 258222 295380 258306 295616
rect 258542 295380 258574 295616
rect 257954 295296 258574 295380
rect 257954 295060 257986 295296
rect 258222 295060 258306 295296
rect 258542 295060 258574 295296
rect 257954 259616 258574 295060
rect 257954 259380 257986 259616
rect 258222 259380 258306 259616
rect 258542 259380 258574 259616
rect 257954 259296 258574 259380
rect 257954 259060 257986 259296
rect 258222 259060 258306 259296
rect 258542 259060 258574 259296
rect 257954 223616 258574 259060
rect 257954 223380 257986 223616
rect 258222 223380 258306 223616
rect 258542 223380 258574 223616
rect 257954 223296 258574 223380
rect 257954 223060 257986 223296
rect 258222 223060 258306 223296
rect 258542 223060 258574 223296
rect 257954 187616 258574 223060
rect 257954 187380 257986 187616
rect 258222 187380 258306 187616
rect 258542 187380 258574 187616
rect 257954 187296 258574 187380
rect 257954 187060 257986 187296
rect 258222 187060 258306 187296
rect 258542 187060 258574 187296
rect 257954 151616 258574 187060
rect 257954 151380 257986 151616
rect 258222 151380 258306 151616
rect 258542 151380 258574 151616
rect 257954 151296 258574 151380
rect 257954 151060 257986 151296
rect 258222 151060 258306 151296
rect 258542 151060 258574 151296
rect 257954 115616 258574 151060
rect 257954 115380 257986 115616
rect 258222 115380 258306 115616
rect 258542 115380 258574 115616
rect 257954 115296 258574 115380
rect 257954 115060 257986 115296
rect 258222 115060 258306 115296
rect 258542 115060 258574 115296
rect 257954 79616 258574 115060
rect 257954 79380 257986 79616
rect 258222 79380 258306 79616
rect 258542 79380 258574 79616
rect 257954 79296 258574 79380
rect 257954 79060 257986 79296
rect 258222 79060 258306 79296
rect 258542 79060 258574 79296
rect 257954 43616 258574 79060
rect 257954 43380 257986 43616
rect 258222 43380 258306 43616
rect 258542 43380 258574 43616
rect 257954 43296 258574 43380
rect 257954 43060 257986 43296
rect 258222 43060 258306 43296
rect 258542 43060 258574 43296
rect 257954 7616 258574 43060
rect 257954 7380 257986 7616
rect 258222 7380 258306 7616
rect 258542 7380 258574 7616
rect 257954 7296 258574 7380
rect 257954 7060 257986 7296
rect 258222 7060 258306 7296
rect 258542 7060 258574 7296
rect 257954 -4184 258574 7060
rect 257954 -4420 257986 -4184
rect 258222 -4420 258306 -4184
rect 258542 -4420 258574 -4184
rect 257954 -4504 258574 -4420
rect 257954 -4740 257986 -4504
rect 258222 -4740 258306 -4504
rect 258542 -4740 258574 -4504
rect 257954 -7652 258574 -4740
rect 259194 709640 259814 711592
rect 259194 709404 259226 709640
rect 259462 709404 259546 709640
rect 259782 709404 259814 709640
rect 259194 709320 259814 709404
rect 259194 709084 259226 709320
rect 259462 709084 259546 709320
rect 259782 709084 259814 709320
rect 259194 692856 259814 709084
rect 259194 692620 259226 692856
rect 259462 692620 259546 692856
rect 259782 692620 259814 692856
rect 259194 692536 259814 692620
rect 259194 692300 259226 692536
rect 259462 692300 259546 692536
rect 259782 692300 259814 692536
rect 259194 656856 259814 692300
rect 259194 656620 259226 656856
rect 259462 656620 259546 656856
rect 259782 656620 259814 656856
rect 259194 656536 259814 656620
rect 259194 656300 259226 656536
rect 259462 656300 259546 656536
rect 259782 656300 259814 656536
rect 259194 620856 259814 656300
rect 259194 620620 259226 620856
rect 259462 620620 259546 620856
rect 259782 620620 259814 620856
rect 259194 620536 259814 620620
rect 259194 620300 259226 620536
rect 259462 620300 259546 620536
rect 259782 620300 259814 620536
rect 259194 584856 259814 620300
rect 259194 584620 259226 584856
rect 259462 584620 259546 584856
rect 259782 584620 259814 584856
rect 259194 584536 259814 584620
rect 259194 584300 259226 584536
rect 259462 584300 259546 584536
rect 259782 584300 259814 584536
rect 259194 548856 259814 584300
rect 259194 548620 259226 548856
rect 259462 548620 259546 548856
rect 259782 548620 259814 548856
rect 259194 548536 259814 548620
rect 259194 548300 259226 548536
rect 259462 548300 259546 548536
rect 259782 548300 259814 548536
rect 259194 512856 259814 548300
rect 259194 512620 259226 512856
rect 259462 512620 259546 512856
rect 259782 512620 259814 512856
rect 259194 512536 259814 512620
rect 259194 512300 259226 512536
rect 259462 512300 259546 512536
rect 259782 512300 259814 512536
rect 259194 476856 259814 512300
rect 259194 476620 259226 476856
rect 259462 476620 259546 476856
rect 259782 476620 259814 476856
rect 259194 476536 259814 476620
rect 259194 476300 259226 476536
rect 259462 476300 259546 476536
rect 259782 476300 259814 476536
rect 259194 440856 259814 476300
rect 259194 440620 259226 440856
rect 259462 440620 259546 440856
rect 259782 440620 259814 440856
rect 259194 440536 259814 440620
rect 259194 440300 259226 440536
rect 259462 440300 259546 440536
rect 259782 440300 259814 440536
rect 259194 404856 259814 440300
rect 259194 404620 259226 404856
rect 259462 404620 259546 404856
rect 259782 404620 259814 404856
rect 259194 404536 259814 404620
rect 259194 404300 259226 404536
rect 259462 404300 259546 404536
rect 259782 404300 259814 404536
rect 259194 368856 259814 404300
rect 259194 368620 259226 368856
rect 259462 368620 259546 368856
rect 259782 368620 259814 368856
rect 259194 368536 259814 368620
rect 259194 368300 259226 368536
rect 259462 368300 259546 368536
rect 259782 368300 259814 368536
rect 259194 332856 259814 368300
rect 259194 332620 259226 332856
rect 259462 332620 259546 332856
rect 259782 332620 259814 332856
rect 259194 332536 259814 332620
rect 259194 332300 259226 332536
rect 259462 332300 259546 332536
rect 259782 332300 259814 332536
rect 259194 296856 259814 332300
rect 259194 296620 259226 296856
rect 259462 296620 259546 296856
rect 259782 296620 259814 296856
rect 259194 296536 259814 296620
rect 259194 296300 259226 296536
rect 259462 296300 259546 296536
rect 259782 296300 259814 296536
rect 259194 260856 259814 296300
rect 259194 260620 259226 260856
rect 259462 260620 259546 260856
rect 259782 260620 259814 260856
rect 259194 260536 259814 260620
rect 259194 260300 259226 260536
rect 259462 260300 259546 260536
rect 259782 260300 259814 260536
rect 259194 224856 259814 260300
rect 259194 224620 259226 224856
rect 259462 224620 259546 224856
rect 259782 224620 259814 224856
rect 259194 224536 259814 224620
rect 259194 224300 259226 224536
rect 259462 224300 259546 224536
rect 259782 224300 259814 224536
rect 259194 188856 259814 224300
rect 259194 188620 259226 188856
rect 259462 188620 259546 188856
rect 259782 188620 259814 188856
rect 259194 188536 259814 188620
rect 259194 188300 259226 188536
rect 259462 188300 259546 188536
rect 259782 188300 259814 188536
rect 259194 152856 259814 188300
rect 259194 152620 259226 152856
rect 259462 152620 259546 152856
rect 259782 152620 259814 152856
rect 259194 152536 259814 152620
rect 259194 152300 259226 152536
rect 259462 152300 259546 152536
rect 259782 152300 259814 152536
rect 259194 116856 259814 152300
rect 259194 116620 259226 116856
rect 259462 116620 259546 116856
rect 259782 116620 259814 116856
rect 259194 116536 259814 116620
rect 259194 116300 259226 116536
rect 259462 116300 259546 116536
rect 259782 116300 259814 116536
rect 259194 80856 259814 116300
rect 259194 80620 259226 80856
rect 259462 80620 259546 80856
rect 259782 80620 259814 80856
rect 259194 80536 259814 80620
rect 259194 80300 259226 80536
rect 259462 80300 259546 80536
rect 259782 80300 259814 80536
rect 259194 44856 259814 80300
rect 259194 44620 259226 44856
rect 259462 44620 259546 44856
rect 259782 44620 259814 44856
rect 259194 44536 259814 44620
rect 259194 44300 259226 44536
rect 259462 44300 259546 44536
rect 259782 44300 259814 44536
rect 259194 8856 259814 44300
rect 259194 8620 259226 8856
rect 259462 8620 259546 8856
rect 259782 8620 259814 8856
rect 259194 8536 259814 8620
rect 259194 8300 259226 8536
rect 259462 8300 259546 8536
rect 259782 8300 259814 8536
rect 259194 -5144 259814 8300
rect 259194 -5380 259226 -5144
rect 259462 -5380 259546 -5144
rect 259782 -5380 259814 -5144
rect 259194 -5464 259814 -5380
rect 259194 -5700 259226 -5464
rect 259462 -5700 259546 -5464
rect 259782 -5700 259814 -5464
rect 259194 -7652 259814 -5700
rect 260434 710600 261054 711592
rect 260434 710364 260466 710600
rect 260702 710364 260786 710600
rect 261022 710364 261054 710600
rect 260434 710280 261054 710364
rect 260434 710044 260466 710280
rect 260702 710044 260786 710280
rect 261022 710044 261054 710280
rect 260434 694096 261054 710044
rect 260434 693860 260466 694096
rect 260702 693860 260786 694096
rect 261022 693860 261054 694096
rect 260434 693776 261054 693860
rect 260434 693540 260466 693776
rect 260702 693540 260786 693776
rect 261022 693540 261054 693776
rect 260434 658096 261054 693540
rect 260434 657860 260466 658096
rect 260702 657860 260786 658096
rect 261022 657860 261054 658096
rect 260434 657776 261054 657860
rect 260434 657540 260466 657776
rect 260702 657540 260786 657776
rect 261022 657540 261054 657776
rect 260434 622096 261054 657540
rect 260434 621860 260466 622096
rect 260702 621860 260786 622096
rect 261022 621860 261054 622096
rect 260434 621776 261054 621860
rect 260434 621540 260466 621776
rect 260702 621540 260786 621776
rect 261022 621540 261054 621776
rect 260434 586096 261054 621540
rect 260434 585860 260466 586096
rect 260702 585860 260786 586096
rect 261022 585860 261054 586096
rect 260434 585776 261054 585860
rect 260434 585540 260466 585776
rect 260702 585540 260786 585776
rect 261022 585540 261054 585776
rect 260434 550096 261054 585540
rect 260434 549860 260466 550096
rect 260702 549860 260786 550096
rect 261022 549860 261054 550096
rect 260434 549776 261054 549860
rect 260434 549540 260466 549776
rect 260702 549540 260786 549776
rect 261022 549540 261054 549776
rect 260434 514096 261054 549540
rect 260434 513860 260466 514096
rect 260702 513860 260786 514096
rect 261022 513860 261054 514096
rect 260434 513776 261054 513860
rect 260434 513540 260466 513776
rect 260702 513540 260786 513776
rect 261022 513540 261054 513776
rect 260434 478096 261054 513540
rect 260434 477860 260466 478096
rect 260702 477860 260786 478096
rect 261022 477860 261054 478096
rect 260434 477776 261054 477860
rect 260434 477540 260466 477776
rect 260702 477540 260786 477776
rect 261022 477540 261054 477776
rect 260434 442096 261054 477540
rect 260434 441860 260466 442096
rect 260702 441860 260786 442096
rect 261022 441860 261054 442096
rect 260434 441776 261054 441860
rect 260434 441540 260466 441776
rect 260702 441540 260786 441776
rect 261022 441540 261054 441776
rect 260434 406096 261054 441540
rect 260434 405860 260466 406096
rect 260702 405860 260786 406096
rect 261022 405860 261054 406096
rect 260434 405776 261054 405860
rect 260434 405540 260466 405776
rect 260702 405540 260786 405776
rect 261022 405540 261054 405776
rect 260434 370096 261054 405540
rect 260434 369860 260466 370096
rect 260702 369860 260786 370096
rect 261022 369860 261054 370096
rect 260434 369776 261054 369860
rect 260434 369540 260466 369776
rect 260702 369540 260786 369776
rect 261022 369540 261054 369776
rect 260434 334096 261054 369540
rect 260434 333860 260466 334096
rect 260702 333860 260786 334096
rect 261022 333860 261054 334096
rect 260434 333776 261054 333860
rect 260434 333540 260466 333776
rect 260702 333540 260786 333776
rect 261022 333540 261054 333776
rect 260434 298096 261054 333540
rect 260434 297860 260466 298096
rect 260702 297860 260786 298096
rect 261022 297860 261054 298096
rect 260434 297776 261054 297860
rect 260434 297540 260466 297776
rect 260702 297540 260786 297776
rect 261022 297540 261054 297776
rect 260434 262096 261054 297540
rect 260434 261860 260466 262096
rect 260702 261860 260786 262096
rect 261022 261860 261054 262096
rect 260434 261776 261054 261860
rect 260434 261540 260466 261776
rect 260702 261540 260786 261776
rect 261022 261540 261054 261776
rect 260434 226096 261054 261540
rect 260434 225860 260466 226096
rect 260702 225860 260786 226096
rect 261022 225860 261054 226096
rect 260434 225776 261054 225860
rect 260434 225540 260466 225776
rect 260702 225540 260786 225776
rect 261022 225540 261054 225776
rect 260434 190096 261054 225540
rect 260434 189860 260466 190096
rect 260702 189860 260786 190096
rect 261022 189860 261054 190096
rect 260434 189776 261054 189860
rect 260434 189540 260466 189776
rect 260702 189540 260786 189776
rect 261022 189540 261054 189776
rect 260434 154096 261054 189540
rect 260434 153860 260466 154096
rect 260702 153860 260786 154096
rect 261022 153860 261054 154096
rect 260434 153776 261054 153860
rect 260434 153540 260466 153776
rect 260702 153540 260786 153776
rect 261022 153540 261054 153776
rect 260434 118096 261054 153540
rect 260434 117860 260466 118096
rect 260702 117860 260786 118096
rect 261022 117860 261054 118096
rect 260434 117776 261054 117860
rect 260434 117540 260466 117776
rect 260702 117540 260786 117776
rect 261022 117540 261054 117776
rect 260434 82096 261054 117540
rect 260434 81860 260466 82096
rect 260702 81860 260786 82096
rect 261022 81860 261054 82096
rect 260434 81776 261054 81860
rect 260434 81540 260466 81776
rect 260702 81540 260786 81776
rect 261022 81540 261054 81776
rect 260434 46096 261054 81540
rect 260434 45860 260466 46096
rect 260702 45860 260786 46096
rect 261022 45860 261054 46096
rect 260434 45776 261054 45860
rect 260434 45540 260466 45776
rect 260702 45540 260786 45776
rect 261022 45540 261054 45776
rect 260434 10096 261054 45540
rect 260434 9860 260466 10096
rect 260702 9860 260786 10096
rect 261022 9860 261054 10096
rect 260434 9776 261054 9860
rect 260434 9540 260466 9776
rect 260702 9540 260786 9776
rect 261022 9540 261054 9776
rect 260434 -6104 261054 9540
rect 260434 -6340 260466 -6104
rect 260702 -6340 260786 -6104
rect 261022 -6340 261054 -6104
rect 260434 -6424 261054 -6340
rect 260434 -6660 260466 -6424
rect 260702 -6660 260786 -6424
rect 261022 -6660 261054 -6424
rect 260434 -7652 261054 -6660
rect 261674 711560 262294 711592
rect 261674 711324 261706 711560
rect 261942 711324 262026 711560
rect 262262 711324 262294 711560
rect 261674 711240 262294 711324
rect 261674 711004 261706 711240
rect 261942 711004 262026 711240
rect 262262 711004 262294 711240
rect 261674 695336 262294 711004
rect 261674 695100 261706 695336
rect 261942 695100 262026 695336
rect 262262 695100 262294 695336
rect 261674 695016 262294 695100
rect 261674 694780 261706 695016
rect 261942 694780 262026 695016
rect 262262 694780 262294 695016
rect 261674 659336 262294 694780
rect 261674 659100 261706 659336
rect 261942 659100 262026 659336
rect 262262 659100 262294 659336
rect 261674 659016 262294 659100
rect 261674 658780 261706 659016
rect 261942 658780 262026 659016
rect 262262 658780 262294 659016
rect 261674 623336 262294 658780
rect 261674 623100 261706 623336
rect 261942 623100 262026 623336
rect 262262 623100 262294 623336
rect 261674 623016 262294 623100
rect 261674 622780 261706 623016
rect 261942 622780 262026 623016
rect 262262 622780 262294 623016
rect 261674 587336 262294 622780
rect 261674 587100 261706 587336
rect 261942 587100 262026 587336
rect 262262 587100 262294 587336
rect 261674 587016 262294 587100
rect 261674 586780 261706 587016
rect 261942 586780 262026 587016
rect 262262 586780 262294 587016
rect 261674 551336 262294 586780
rect 261674 551100 261706 551336
rect 261942 551100 262026 551336
rect 262262 551100 262294 551336
rect 261674 551016 262294 551100
rect 261674 550780 261706 551016
rect 261942 550780 262026 551016
rect 262262 550780 262294 551016
rect 261674 515336 262294 550780
rect 261674 515100 261706 515336
rect 261942 515100 262026 515336
rect 262262 515100 262294 515336
rect 261674 515016 262294 515100
rect 261674 514780 261706 515016
rect 261942 514780 262026 515016
rect 262262 514780 262294 515016
rect 261674 479336 262294 514780
rect 261674 479100 261706 479336
rect 261942 479100 262026 479336
rect 262262 479100 262294 479336
rect 261674 479016 262294 479100
rect 261674 478780 261706 479016
rect 261942 478780 262026 479016
rect 262262 478780 262294 479016
rect 261674 443336 262294 478780
rect 261674 443100 261706 443336
rect 261942 443100 262026 443336
rect 262262 443100 262294 443336
rect 261674 443016 262294 443100
rect 261674 442780 261706 443016
rect 261942 442780 262026 443016
rect 262262 442780 262294 443016
rect 261674 407336 262294 442780
rect 261674 407100 261706 407336
rect 261942 407100 262026 407336
rect 262262 407100 262294 407336
rect 261674 407016 262294 407100
rect 261674 406780 261706 407016
rect 261942 406780 262026 407016
rect 262262 406780 262294 407016
rect 261674 371336 262294 406780
rect 261674 371100 261706 371336
rect 261942 371100 262026 371336
rect 262262 371100 262294 371336
rect 261674 371016 262294 371100
rect 261674 370780 261706 371016
rect 261942 370780 262026 371016
rect 262262 370780 262294 371016
rect 261674 335336 262294 370780
rect 261674 335100 261706 335336
rect 261942 335100 262026 335336
rect 262262 335100 262294 335336
rect 261674 335016 262294 335100
rect 261674 334780 261706 335016
rect 261942 334780 262026 335016
rect 262262 334780 262294 335016
rect 261674 299336 262294 334780
rect 261674 299100 261706 299336
rect 261942 299100 262026 299336
rect 262262 299100 262294 299336
rect 261674 299016 262294 299100
rect 261674 298780 261706 299016
rect 261942 298780 262026 299016
rect 262262 298780 262294 299016
rect 261674 263336 262294 298780
rect 261674 263100 261706 263336
rect 261942 263100 262026 263336
rect 262262 263100 262294 263336
rect 261674 263016 262294 263100
rect 261674 262780 261706 263016
rect 261942 262780 262026 263016
rect 262262 262780 262294 263016
rect 261674 227336 262294 262780
rect 261674 227100 261706 227336
rect 261942 227100 262026 227336
rect 262262 227100 262294 227336
rect 261674 227016 262294 227100
rect 261674 226780 261706 227016
rect 261942 226780 262026 227016
rect 262262 226780 262294 227016
rect 261674 191336 262294 226780
rect 261674 191100 261706 191336
rect 261942 191100 262026 191336
rect 262262 191100 262294 191336
rect 261674 191016 262294 191100
rect 261674 190780 261706 191016
rect 261942 190780 262026 191016
rect 262262 190780 262294 191016
rect 261674 155336 262294 190780
rect 261674 155100 261706 155336
rect 261942 155100 262026 155336
rect 262262 155100 262294 155336
rect 261674 155016 262294 155100
rect 261674 154780 261706 155016
rect 261942 154780 262026 155016
rect 262262 154780 262294 155016
rect 261674 119336 262294 154780
rect 261674 119100 261706 119336
rect 261942 119100 262026 119336
rect 262262 119100 262294 119336
rect 261674 119016 262294 119100
rect 261674 118780 261706 119016
rect 261942 118780 262026 119016
rect 262262 118780 262294 119016
rect 261674 83336 262294 118780
rect 261674 83100 261706 83336
rect 261942 83100 262026 83336
rect 262262 83100 262294 83336
rect 261674 83016 262294 83100
rect 261674 82780 261706 83016
rect 261942 82780 262026 83016
rect 262262 82780 262294 83016
rect 261674 47336 262294 82780
rect 261674 47100 261706 47336
rect 261942 47100 262026 47336
rect 262262 47100 262294 47336
rect 261674 47016 262294 47100
rect 261674 46780 261706 47016
rect 261942 46780 262026 47016
rect 262262 46780 262294 47016
rect 261674 11336 262294 46780
rect 261674 11100 261706 11336
rect 261942 11100 262026 11336
rect 262262 11100 262294 11336
rect 261674 11016 262294 11100
rect 261674 10780 261706 11016
rect 261942 10780 262026 11016
rect 262262 10780 262294 11016
rect 261674 -7064 262294 10780
rect 261674 -7300 261706 -7064
rect 261942 -7300 262026 -7064
rect 262262 -7300 262294 -7064
rect 261674 -7384 262294 -7300
rect 261674 -7620 261706 -7384
rect 261942 -7620 262026 -7384
rect 262262 -7620 262294 -7384
rect 261674 -7652 262294 -7620
rect 288994 704840 289614 711592
rect 288994 704604 289026 704840
rect 289262 704604 289346 704840
rect 289582 704604 289614 704840
rect 288994 704520 289614 704604
rect 288994 704284 289026 704520
rect 289262 704284 289346 704520
rect 289582 704284 289614 704520
rect 288994 686656 289614 704284
rect 288994 686420 289026 686656
rect 289262 686420 289346 686656
rect 289582 686420 289614 686656
rect 288994 686336 289614 686420
rect 288994 686100 289026 686336
rect 289262 686100 289346 686336
rect 289582 686100 289614 686336
rect 288994 650656 289614 686100
rect 288994 650420 289026 650656
rect 289262 650420 289346 650656
rect 289582 650420 289614 650656
rect 288994 650336 289614 650420
rect 288994 650100 289026 650336
rect 289262 650100 289346 650336
rect 289582 650100 289614 650336
rect 288994 614656 289614 650100
rect 288994 614420 289026 614656
rect 289262 614420 289346 614656
rect 289582 614420 289614 614656
rect 288994 614336 289614 614420
rect 288994 614100 289026 614336
rect 289262 614100 289346 614336
rect 289582 614100 289614 614336
rect 288994 578656 289614 614100
rect 288994 578420 289026 578656
rect 289262 578420 289346 578656
rect 289582 578420 289614 578656
rect 288994 578336 289614 578420
rect 288994 578100 289026 578336
rect 289262 578100 289346 578336
rect 289582 578100 289614 578336
rect 288994 542656 289614 578100
rect 288994 542420 289026 542656
rect 289262 542420 289346 542656
rect 289582 542420 289614 542656
rect 288994 542336 289614 542420
rect 288994 542100 289026 542336
rect 289262 542100 289346 542336
rect 289582 542100 289614 542336
rect 288994 506656 289614 542100
rect 288994 506420 289026 506656
rect 289262 506420 289346 506656
rect 289582 506420 289614 506656
rect 288994 506336 289614 506420
rect 288994 506100 289026 506336
rect 289262 506100 289346 506336
rect 289582 506100 289614 506336
rect 288994 470656 289614 506100
rect 288994 470420 289026 470656
rect 289262 470420 289346 470656
rect 289582 470420 289614 470656
rect 288994 470336 289614 470420
rect 288994 470100 289026 470336
rect 289262 470100 289346 470336
rect 289582 470100 289614 470336
rect 288994 434656 289614 470100
rect 288994 434420 289026 434656
rect 289262 434420 289346 434656
rect 289582 434420 289614 434656
rect 288994 434336 289614 434420
rect 288994 434100 289026 434336
rect 289262 434100 289346 434336
rect 289582 434100 289614 434336
rect 288994 398656 289614 434100
rect 288994 398420 289026 398656
rect 289262 398420 289346 398656
rect 289582 398420 289614 398656
rect 288994 398336 289614 398420
rect 288994 398100 289026 398336
rect 289262 398100 289346 398336
rect 289582 398100 289614 398336
rect 288994 362656 289614 398100
rect 288994 362420 289026 362656
rect 289262 362420 289346 362656
rect 289582 362420 289614 362656
rect 288994 362336 289614 362420
rect 288994 362100 289026 362336
rect 289262 362100 289346 362336
rect 289582 362100 289614 362336
rect 288994 326656 289614 362100
rect 288994 326420 289026 326656
rect 289262 326420 289346 326656
rect 289582 326420 289614 326656
rect 288994 326336 289614 326420
rect 288994 326100 289026 326336
rect 289262 326100 289346 326336
rect 289582 326100 289614 326336
rect 288994 290656 289614 326100
rect 288994 290420 289026 290656
rect 289262 290420 289346 290656
rect 289582 290420 289614 290656
rect 288994 290336 289614 290420
rect 288994 290100 289026 290336
rect 289262 290100 289346 290336
rect 289582 290100 289614 290336
rect 288994 254656 289614 290100
rect 288994 254420 289026 254656
rect 289262 254420 289346 254656
rect 289582 254420 289614 254656
rect 288994 254336 289614 254420
rect 288994 254100 289026 254336
rect 289262 254100 289346 254336
rect 289582 254100 289614 254336
rect 288994 218656 289614 254100
rect 288994 218420 289026 218656
rect 289262 218420 289346 218656
rect 289582 218420 289614 218656
rect 288994 218336 289614 218420
rect 288994 218100 289026 218336
rect 289262 218100 289346 218336
rect 289582 218100 289614 218336
rect 288994 182656 289614 218100
rect 288994 182420 289026 182656
rect 289262 182420 289346 182656
rect 289582 182420 289614 182656
rect 288994 182336 289614 182420
rect 288994 182100 289026 182336
rect 289262 182100 289346 182336
rect 289582 182100 289614 182336
rect 288994 146656 289614 182100
rect 288994 146420 289026 146656
rect 289262 146420 289346 146656
rect 289582 146420 289614 146656
rect 288994 146336 289614 146420
rect 288994 146100 289026 146336
rect 289262 146100 289346 146336
rect 289582 146100 289614 146336
rect 288994 110656 289614 146100
rect 288994 110420 289026 110656
rect 289262 110420 289346 110656
rect 289582 110420 289614 110656
rect 288994 110336 289614 110420
rect 288994 110100 289026 110336
rect 289262 110100 289346 110336
rect 289582 110100 289614 110336
rect 288994 74656 289614 110100
rect 288994 74420 289026 74656
rect 289262 74420 289346 74656
rect 289582 74420 289614 74656
rect 288994 74336 289614 74420
rect 288994 74100 289026 74336
rect 289262 74100 289346 74336
rect 289582 74100 289614 74336
rect 288994 38656 289614 74100
rect 288994 38420 289026 38656
rect 289262 38420 289346 38656
rect 289582 38420 289614 38656
rect 288994 38336 289614 38420
rect 288994 38100 289026 38336
rect 289262 38100 289346 38336
rect 289582 38100 289614 38336
rect 288994 2656 289614 38100
rect 288994 2420 289026 2656
rect 289262 2420 289346 2656
rect 289582 2420 289614 2656
rect 288994 2336 289614 2420
rect 288994 2100 289026 2336
rect 289262 2100 289346 2336
rect 289582 2100 289614 2336
rect 288994 -344 289614 2100
rect 288994 -580 289026 -344
rect 289262 -580 289346 -344
rect 289582 -580 289614 -344
rect 288994 -664 289614 -580
rect 288994 -900 289026 -664
rect 289262 -900 289346 -664
rect 289582 -900 289614 -664
rect 288994 -7652 289614 -900
rect 290234 705800 290854 711592
rect 290234 705564 290266 705800
rect 290502 705564 290586 705800
rect 290822 705564 290854 705800
rect 290234 705480 290854 705564
rect 290234 705244 290266 705480
rect 290502 705244 290586 705480
rect 290822 705244 290854 705480
rect 290234 687896 290854 705244
rect 290234 687660 290266 687896
rect 290502 687660 290586 687896
rect 290822 687660 290854 687896
rect 290234 687576 290854 687660
rect 290234 687340 290266 687576
rect 290502 687340 290586 687576
rect 290822 687340 290854 687576
rect 290234 651896 290854 687340
rect 290234 651660 290266 651896
rect 290502 651660 290586 651896
rect 290822 651660 290854 651896
rect 290234 651576 290854 651660
rect 290234 651340 290266 651576
rect 290502 651340 290586 651576
rect 290822 651340 290854 651576
rect 290234 615896 290854 651340
rect 290234 615660 290266 615896
rect 290502 615660 290586 615896
rect 290822 615660 290854 615896
rect 290234 615576 290854 615660
rect 290234 615340 290266 615576
rect 290502 615340 290586 615576
rect 290822 615340 290854 615576
rect 290234 579896 290854 615340
rect 290234 579660 290266 579896
rect 290502 579660 290586 579896
rect 290822 579660 290854 579896
rect 290234 579576 290854 579660
rect 290234 579340 290266 579576
rect 290502 579340 290586 579576
rect 290822 579340 290854 579576
rect 290234 543896 290854 579340
rect 290234 543660 290266 543896
rect 290502 543660 290586 543896
rect 290822 543660 290854 543896
rect 290234 543576 290854 543660
rect 290234 543340 290266 543576
rect 290502 543340 290586 543576
rect 290822 543340 290854 543576
rect 290234 507896 290854 543340
rect 290234 507660 290266 507896
rect 290502 507660 290586 507896
rect 290822 507660 290854 507896
rect 290234 507576 290854 507660
rect 290234 507340 290266 507576
rect 290502 507340 290586 507576
rect 290822 507340 290854 507576
rect 290234 471896 290854 507340
rect 290234 471660 290266 471896
rect 290502 471660 290586 471896
rect 290822 471660 290854 471896
rect 290234 471576 290854 471660
rect 290234 471340 290266 471576
rect 290502 471340 290586 471576
rect 290822 471340 290854 471576
rect 290234 435896 290854 471340
rect 290234 435660 290266 435896
rect 290502 435660 290586 435896
rect 290822 435660 290854 435896
rect 290234 435576 290854 435660
rect 290234 435340 290266 435576
rect 290502 435340 290586 435576
rect 290822 435340 290854 435576
rect 290234 399896 290854 435340
rect 290234 399660 290266 399896
rect 290502 399660 290586 399896
rect 290822 399660 290854 399896
rect 290234 399576 290854 399660
rect 290234 399340 290266 399576
rect 290502 399340 290586 399576
rect 290822 399340 290854 399576
rect 290234 363896 290854 399340
rect 290234 363660 290266 363896
rect 290502 363660 290586 363896
rect 290822 363660 290854 363896
rect 290234 363576 290854 363660
rect 290234 363340 290266 363576
rect 290502 363340 290586 363576
rect 290822 363340 290854 363576
rect 290234 327896 290854 363340
rect 290234 327660 290266 327896
rect 290502 327660 290586 327896
rect 290822 327660 290854 327896
rect 290234 327576 290854 327660
rect 290234 327340 290266 327576
rect 290502 327340 290586 327576
rect 290822 327340 290854 327576
rect 290234 291896 290854 327340
rect 290234 291660 290266 291896
rect 290502 291660 290586 291896
rect 290822 291660 290854 291896
rect 290234 291576 290854 291660
rect 290234 291340 290266 291576
rect 290502 291340 290586 291576
rect 290822 291340 290854 291576
rect 290234 255896 290854 291340
rect 290234 255660 290266 255896
rect 290502 255660 290586 255896
rect 290822 255660 290854 255896
rect 290234 255576 290854 255660
rect 290234 255340 290266 255576
rect 290502 255340 290586 255576
rect 290822 255340 290854 255576
rect 290234 219896 290854 255340
rect 290234 219660 290266 219896
rect 290502 219660 290586 219896
rect 290822 219660 290854 219896
rect 290234 219576 290854 219660
rect 290234 219340 290266 219576
rect 290502 219340 290586 219576
rect 290822 219340 290854 219576
rect 290234 183896 290854 219340
rect 290234 183660 290266 183896
rect 290502 183660 290586 183896
rect 290822 183660 290854 183896
rect 290234 183576 290854 183660
rect 290234 183340 290266 183576
rect 290502 183340 290586 183576
rect 290822 183340 290854 183576
rect 290234 147896 290854 183340
rect 290234 147660 290266 147896
rect 290502 147660 290586 147896
rect 290822 147660 290854 147896
rect 290234 147576 290854 147660
rect 290234 147340 290266 147576
rect 290502 147340 290586 147576
rect 290822 147340 290854 147576
rect 290234 111896 290854 147340
rect 290234 111660 290266 111896
rect 290502 111660 290586 111896
rect 290822 111660 290854 111896
rect 290234 111576 290854 111660
rect 290234 111340 290266 111576
rect 290502 111340 290586 111576
rect 290822 111340 290854 111576
rect 290234 75896 290854 111340
rect 290234 75660 290266 75896
rect 290502 75660 290586 75896
rect 290822 75660 290854 75896
rect 290234 75576 290854 75660
rect 290234 75340 290266 75576
rect 290502 75340 290586 75576
rect 290822 75340 290854 75576
rect 290234 39896 290854 75340
rect 290234 39660 290266 39896
rect 290502 39660 290586 39896
rect 290822 39660 290854 39896
rect 290234 39576 290854 39660
rect 290234 39340 290266 39576
rect 290502 39340 290586 39576
rect 290822 39340 290854 39576
rect 290234 3896 290854 39340
rect 290234 3660 290266 3896
rect 290502 3660 290586 3896
rect 290822 3660 290854 3896
rect 290234 3576 290854 3660
rect 290234 3340 290266 3576
rect 290502 3340 290586 3576
rect 290822 3340 290854 3576
rect 290234 -1304 290854 3340
rect 290234 -1540 290266 -1304
rect 290502 -1540 290586 -1304
rect 290822 -1540 290854 -1304
rect 290234 -1624 290854 -1540
rect 290234 -1860 290266 -1624
rect 290502 -1860 290586 -1624
rect 290822 -1860 290854 -1624
rect 290234 -7652 290854 -1860
rect 291474 706760 292094 711592
rect 291474 706524 291506 706760
rect 291742 706524 291826 706760
rect 292062 706524 292094 706760
rect 291474 706440 292094 706524
rect 291474 706204 291506 706440
rect 291742 706204 291826 706440
rect 292062 706204 292094 706440
rect 291474 689136 292094 706204
rect 291474 688900 291506 689136
rect 291742 688900 291826 689136
rect 292062 688900 292094 689136
rect 291474 688816 292094 688900
rect 291474 688580 291506 688816
rect 291742 688580 291826 688816
rect 292062 688580 292094 688816
rect 291474 653136 292094 688580
rect 291474 652900 291506 653136
rect 291742 652900 291826 653136
rect 292062 652900 292094 653136
rect 291474 652816 292094 652900
rect 291474 652580 291506 652816
rect 291742 652580 291826 652816
rect 292062 652580 292094 652816
rect 291474 617136 292094 652580
rect 291474 616900 291506 617136
rect 291742 616900 291826 617136
rect 292062 616900 292094 617136
rect 291474 616816 292094 616900
rect 291474 616580 291506 616816
rect 291742 616580 291826 616816
rect 292062 616580 292094 616816
rect 291474 581136 292094 616580
rect 291474 580900 291506 581136
rect 291742 580900 291826 581136
rect 292062 580900 292094 581136
rect 291474 580816 292094 580900
rect 291474 580580 291506 580816
rect 291742 580580 291826 580816
rect 292062 580580 292094 580816
rect 291474 545136 292094 580580
rect 291474 544900 291506 545136
rect 291742 544900 291826 545136
rect 292062 544900 292094 545136
rect 291474 544816 292094 544900
rect 291474 544580 291506 544816
rect 291742 544580 291826 544816
rect 292062 544580 292094 544816
rect 291474 509136 292094 544580
rect 291474 508900 291506 509136
rect 291742 508900 291826 509136
rect 292062 508900 292094 509136
rect 291474 508816 292094 508900
rect 291474 508580 291506 508816
rect 291742 508580 291826 508816
rect 292062 508580 292094 508816
rect 291474 473136 292094 508580
rect 291474 472900 291506 473136
rect 291742 472900 291826 473136
rect 292062 472900 292094 473136
rect 291474 472816 292094 472900
rect 291474 472580 291506 472816
rect 291742 472580 291826 472816
rect 292062 472580 292094 472816
rect 291474 437136 292094 472580
rect 291474 436900 291506 437136
rect 291742 436900 291826 437136
rect 292062 436900 292094 437136
rect 291474 436816 292094 436900
rect 291474 436580 291506 436816
rect 291742 436580 291826 436816
rect 292062 436580 292094 436816
rect 291474 401136 292094 436580
rect 291474 400900 291506 401136
rect 291742 400900 291826 401136
rect 292062 400900 292094 401136
rect 291474 400816 292094 400900
rect 291474 400580 291506 400816
rect 291742 400580 291826 400816
rect 292062 400580 292094 400816
rect 291474 365136 292094 400580
rect 291474 364900 291506 365136
rect 291742 364900 291826 365136
rect 292062 364900 292094 365136
rect 291474 364816 292094 364900
rect 291474 364580 291506 364816
rect 291742 364580 291826 364816
rect 292062 364580 292094 364816
rect 291474 329136 292094 364580
rect 291474 328900 291506 329136
rect 291742 328900 291826 329136
rect 292062 328900 292094 329136
rect 291474 328816 292094 328900
rect 291474 328580 291506 328816
rect 291742 328580 291826 328816
rect 292062 328580 292094 328816
rect 291474 293136 292094 328580
rect 291474 292900 291506 293136
rect 291742 292900 291826 293136
rect 292062 292900 292094 293136
rect 291474 292816 292094 292900
rect 291474 292580 291506 292816
rect 291742 292580 291826 292816
rect 292062 292580 292094 292816
rect 291474 257136 292094 292580
rect 291474 256900 291506 257136
rect 291742 256900 291826 257136
rect 292062 256900 292094 257136
rect 291474 256816 292094 256900
rect 291474 256580 291506 256816
rect 291742 256580 291826 256816
rect 292062 256580 292094 256816
rect 291474 221136 292094 256580
rect 291474 220900 291506 221136
rect 291742 220900 291826 221136
rect 292062 220900 292094 221136
rect 291474 220816 292094 220900
rect 291474 220580 291506 220816
rect 291742 220580 291826 220816
rect 292062 220580 292094 220816
rect 291474 185136 292094 220580
rect 291474 184900 291506 185136
rect 291742 184900 291826 185136
rect 292062 184900 292094 185136
rect 291474 184816 292094 184900
rect 291474 184580 291506 184816
rect 291742 184580 291826 184816
rect 292062 184580 292094 184816
rect 291474 149136 292094 184580
rect 291474 148900 291506 149136
rect 291742 148900 291826 149136
rect 292062 148900 292094 149136
rect 291474 148816 292094 148900
rect 291474 148580 291506 148816
rect 291742 148580 291826 148816
rect 292062 148580 292094 148816
rect 291474 113136 292094 148580
rect 291474 112900 291506 113136
rect 291742 112900 291826 113136
rect 292062 112900 292094 113136
rect 291474 112816 292094 112900
rect 291474 112580 291506 112816
rect 291742 112580 291826 112816
rect 292062 112580 292094 112816
rect 291474 77136 292094 112580
rect 291474 76900 291506 77136
rect 291742 76900 291826 77136
rect 292062 76900 292094 77136
rect 291474 76816 292094 76900
rect 291474 76580 291506 76816
rect 291742 76580 291826 76816
rect 292062 76580 292094 76816
rect 291474 41136 292094 76580
rect 291474 40900 291506 41136
rect 291742 40900 291826 41136
rect 292062 40900 292094 41136
rect 291474 40816 292094 40900
rect 291474 40580 291506 40816
rect 291742 40580 291826 40816
rect 292062 40580 292094 40816
rect 291474 5136 292094 40580
rect 291474 4900 291506 5136
rect 291742 4900 291826 5136
rect 292062 4900 292094 5136
rect 291474 4816 292094 4900
rect 291474 4580 291506 4816
rect 291742 4580 291826 4816
rect 292062 4580 292094 4816
rect 291474 -2264 292094 4580
rect 291474 -2500 291506 -2264
rect 291742 -2500 291826 -2264
rect 292062 -2500 292094 -2264
rect 291474 -2584 292094 -2500
rect 291474 -2820 291506 -2584
rect 291742 -2820 291826 -2584
rect 292062 -2820 292094 -2584
rect 291474 -7652 292094 -2820
rect 292714 707720 293334 711592
rect 292714 707484 292746 707720
rect 292982 707484 293066 707720
rect 293302 707484 293334 707720
rect 292714 707400 293334 707484
rect 292714 707164 292746 707400
rect 292982 707164 293066 707400
rect 293302 707164 293334 707400
rect 292714 690376 293334 707164
rect 292714 690140 292746 690376
rect 292982 690140 293066 690376
rect 293302 690140 293334 690376
rect 292714 690056 293334 690140
rect 292714 689820 292746 690056
rect 292982 689820 293066 690056
rect 293302 689820 293334 690056
rect 292714 654376 293334 689820
rect 292714 654140 292746 654376
rect 292982 654140 293066 654376
rect 293302 654140 293334 654376
rect 292714 654056 293334 654140
rect 292714 653820 292746 654056
rect 292982 653820 293066 654056
rect 293302 653820 293334 654056
rect 292714 618376 293334 653820
rect 292714 618140 292746 618376
rect 292982 618140 293066 618376
rect 293302 618140 293334 618376
rect 292714 618056 293334 618140
rect 292714 617820 292746 618056
rect 292982 617820 293066 618056
rect 293302 617820 293334 618056
rect 292714 582376 293334 617820
rect 292714 582140 292746 582376
rect 292982 582140 293066 582376
rect 293302 582140 293334 582376
rect 292714 582056 293334 582140
rect 292714 581820 292746 582056
rect 292982 581820 293066 582056
rect 293302 581820 293334 582056
rect 292714 546376 293334 581820
rect 292714 546140 292746 546376
rect 292982 546140 293066 546376
rect 293302 546140 293334 546376
rect 292714 546056 293334 546140
rect 292714 545820 292746 546056
rect 292982 545820 293066 546056
rect 293302 545820 293334 546056
rect 292714 510376 293334 545820
rect 292714 510140 292746 510376
rect 292982 510140 293066 510376
rect 293302 510140 293334 510376
rect 292714 510056 293334 510140
rect 292714 509820 292746 510056
rect 292982 509820 293066 510056
rect 293302 509820 293334 510056
rect 292714 474376 293334 509820
rect 292714 474140 292746 474376
rect 292982 474140 293066 474376
rect 293302 474140 293334 474376
rect 292714 474056 293334 474140
rect 292714 473820 292746 474056
rect 292982 473820 293066 474056
rect 293302 473820 293334 474056
rect 292714 438376 293334 473820
rect 292714 438140 292746 438376
rect 292982 438140 293066 438376
rect 293302 438140 293334 438376
rect 292714 438056 293334 438140
rect 292714 437820 292746 438056
rect 292982 437820 293066 438056
rect 293302 437820 293334 438056
rect 292714 402376 293334 437820
rect 292714 402140 292746 402376
rect 292982 402140 293066 402376
rect 293302 402140 293334 402376
rect 292714 402056 293334 402140
rect 292714 401820 292746 402056
rect 292982 401820 293066 402056
rect 293302 401820 293334 402056
rect 292714 366376 293334 401820
rect 292714 366140 292746 366376
rect 292982 366140 293066 366376
rect 293302 366140 293334 366376
rect 292714 366056 293334 366140
rect 292714 365820 292746 366056
rect 292982 365820 293066 366056
rect 293302 365820 293334 366056
rect 292714 330376 293334 365820
rect 292714 330140 292746 330376
rect 292982 330140 293066 330376
rect 293302 330140 293334 330376
rect 292714 330056 293334 330140
rect 292714 329820 292746 330056
rect 292982 329820 293066 330056
rect 293302 329820 293334 330056
rect 292714 294376 293334 329820
rect 292714 294140 292746 294376
rect 292982 294140 293066 294376
rect 293302 294140 293334 294376
rect 292714 294056 293334 294140
rect 292714 293820 292746 294056
rect 292982 293820 293066 294056
rect 293302 293820 293334 294056
rect 292714 258376 293334 293820
rect 292714 258140 292746 258376
rect 292982 258140 293066 258376
rect 293302 258140 293334 258376
rect 292714 258056 293334 258140
rect 292714 257820 292746 258056
rect 292982 257820 293066 258056
rect 293302 257820 293334 258056
rect 292714 222376 293334 257820
rect 292714 222140 292746 222376
rect 292982 222140 293066 222376
rect 293302 222140 293334 222376
rect 292714 222056 293334 222140
rect 292714 221820 292746 222056
rect 292982 221820 293066 222056
rect 293302 221820 293334 222056
rect 292714 186376 293334 221820
rect 292714 186140 292746 186376
rect 292982 186140 293066 186376
rect 293302 186140 293334 186376
rect 292714 186056 293334 186140
rect 292714 185820 292746 186056
rect 292982 185820 293066 186056
rect 293302 185820 293334 186056
rect 292714 150376 293334 185820
rect 292714 150140 292746 150376
rect 292982 150140 293066 150376
rect 293302 150140 293334 150376
rect 292714 150056 293334 150140
rect 292714 149820 292746 150056
rect 292982 149820 293066 150056
rect 293302 149820 293334 150056
rect 292714 114376 293334 149820
rect 292714 114140 292746 114376
rect 292982 114140 293066 114376
rect 293302 114140 293334 114376
rect 292714 114056 293334 114140
rect 292714 113820 292746 114056
rect 292982 113820 293066 114056
rect 293302 113820 293334 114056
rect 292714 78376 293334 113820
rect 292714 78140 292746 78376
rect 292982 78140 293066 78376
rect 293302 78140 293334 78376
rect 292714 78056 293334 78140
rect 292714 77820 292746 78056
rect 292982 77820 293066 78056
rect 293302 77820 293334 78056
rect 292714 42376 293334 77820
rect 292714 42140 292746 42376
rect 292982 42140 293066 42376
rect 293302 42140 293334 42376
rect 292714 42056 293334 42140
rect 292714 41820 292746 42056
rect 292982 41820 293066 42056
rect 293302 41820 293334 42056
rect 292714 6376 293334 41820
rect 292714 6140 292746 6376
rect 292982 6140 293066 6376
rect 293302 6140 293334 6376
rect 292714 6056 293334 6140
rect 292714 5820 292746 6056
rect 292982 5820 293066 6056
rect 293302 5820 293334 6056
rect 292714 -3224 293334 5820
rect 292714 -3460 292746 -3224
rect 292982 -3460 293066 -3224
rect 293302 -3460 293334 -3224
rect 292714 -3544 293334 -3460
rect 292714 -3780 292746 -3544
rect 292982 -3780 293066 -3544
rect 293302 -3780 293334 -3544
rect 292714 -7652 293334 -3780
rect 293954 708680 294574 711592
rect 293954 708444 293986 708680
rect 294222 708444 294306 708680
rect 294542 708444 294574 708680
rect 293954 708360 294574 708444
rect 293954 708124 293986 708360
rect 294222 708124 294306 708360
rect 294542 708124 294574 708360
rect 293954 691616 294574 708124
rect 293954 691380 293986 691616
rect 294222 691380 294306 691616
rect 294542 691380 294574 691616
rect 293954 691296 294574 691380
rect 293954 691060 293986 691296
rect 294222 691060 294306 691296
rect 294542 691060 294574 691296
rect 293954 655616 294574 691060
rect 293954 655380 293986 655616
rect 294222 655380 294306 655616
rect 294542 655380 294574 655616
rect 293954 655296 294574 655380
rect 293954 655060 293986 655296
rect 294222 655060 294306 655296
rect 294542 655060 294574 655296
rect 293954 619616 294574 655060
rect 293954 619380 293986 619616
rect 294222 619380 294306 619616
rect 294542 619380 294574 619616
rect 293954 619296 294574 619380
rect 293954 619060 293986 619296
rect 294222 619060 294306 619296
rect 294542 619060 294574 619296
rect 293954 583616 294574 619060
rect 293954 583380 293986 583616
rect 294222 583380 294306 583616
rect 294542 583380 294574 583616
rect 293954 583296 294574 583380
rect 293954 583060 293986 583296
rect 294222 583060 294306 583296
rect 294542 583060 294574 583296
rect 293954 547616 294574 583060
rect 293954 547380 293986 547616
rect 294222 547380 294306 547616
rect 294542 547380 294574 547616
rect 293954 547296 294574 547380
rect 293954 547060 293986 547296
rect 294222 547060 294306 547296
rect 294542 547060 294574 547296
rect 293954 511616 294574 547060
rect 293954 511380 293986 511616
rect 294222 511380 294306 511616
rect 294542 511380 294574 511616
rect 293954 511296 294574 511380
rect 293954 511060 293986 511296
rect 294222 511060 294306 511296
rect 294542 511060 294574 511296
rect 293954 475616 294574 511060
rect 293954 475380 293986 475616
rect 294222 475380 294306 475616
rect 294542 475380 294574 475616
rect 293954 475296 294574 475380
rect 293954 475060 293986 475296
rect 294222 475060 294306 475296
rect 294542 475060 294574 475296
rect 293954 439616 294574 475060
rect 293954 439380 293986 439616
rect 294222 439380 294306 439616
rect 294542 439380 294574 439616
rect 293954 439296 294574 439380
rect 293954 439060 293986 439296
rect 294222 439060 294306 439296
rect 294542 439060 294574 439296
rect 293954 403616 294574 439060
rect 293954 403380 293986 403616
rect 294222 403380 294306 403616
rect 294542 403380 294574 403616
rect 293954 403296 294574 403380
rect 293954 403060 293986 403296
rect 294222 403060 294306 403296
rect 294542 403060 294574 403296
rect 293954 367616 294574 403060
rect 293954 367380 293986 367616
rect 294222 367380 294306 367616
rect 294542 367380 294574 367616
rect 293954 367296 294574 367380
rect 293954 367060 293986 367296
rect 294222 367060 294306 367296
rect 294542 367060 294574 367296
rect 293954 331616 294574 367060
rect 293954 331380 293986 331616
rect 294222 331380 294306 331616
rect 294542 331380 294574 331616
rect 293954 331296 294574 331380
rect 293954 331060 293986 331296
rect 294222 331060 294306 331296
rect 294542 331060 294574 331296
rect 293954 295616 294574 331060
rect 293954 295380 293986 295616
rect 294222 295380 294306 295616
rect 294542 295380 294574 295616
rect 293954 295296 294574 295380
rect 293954 295060 293986 295296
rect 294222 295060 294306 295296
rect 294542 295060 294574 295296
rect 293954 259616 294574 295060
rect 293954 259380 293986 259616
rect 294222 259380 294306 259616
rect 294542 259380 294574 259616
rect 293954 259296 294574 259380
rect 293954 259060 293986 259296
rect 294222 259060 294306 259296
rect 294542 259060 294574 259296
rect 293954 223616 294574 259060
rect 293954 223380 293986 223616
rect 294222 223380 294306 223616
rect 294542 223380 294574 223616
rect 293954 223296 294574 223380
rect 293954 223060 293986 223296
rect 294222 223060 294306 223296
rect 294542 223060 294574 223296
rect 293954 187616 294574 223060
rect 293954 187380 293986 187616
rect 294222 187380 294306 187616
rect 294542 187380 294574 187616
rect 293954 187296 294574 187380
rect 293954 187060 293986 187296
rect 294222 187060 294306 187296
rect 294542 187060 294574 187296
rect 293954 151616 294574 187060
rect 293954 151380 293986 151616
rect 294222 151380 294306 151616
rect 294542 151380 294574 151616
rect 293954 151296 294574 151380
rect 293954 151060 293986 151296
rect 294222 151060 294306 151296
rect 294542 151060 294574 151296
rect 293954 115616 294574 151060
rect 293954 115380 293986 115616
rect 294222 115380 294306 115616
rect 294542 115380 294574 115616
rect 293954 115296 294574 115380
rect 293954 115060 293986 115296
rect 294222 115060 294306 115296
rect 294542 115060 294574 115296
rect 293954 79616 294574 115060
rect 293954 79380 293986 79616
rect 294222 79380 294306 79616
rect 294542 79380 294574 79616
rect 293954 79296 294574 79380
rect 293954 79060 293986 79296
rect 294222 79060 294306 79296
rect 294542 79060 294574 79296
rect 293954 43616 294574 79060
rect 293954 43380 293986 43616
rect 294222 43380 294306 43616
rect 294542 43380 294574 43616
rect 293954 43296 294574 43380
rect 293954 43060 293986 43296
rect 294222 43060 294306 43296
rect 294542 43060 294574 43296
rect 293954 7616 294574 43060
rect 293954 7380 293986 7616
rect 294222 7380 294306 7616
rect 294542 7380 294574 7616
rect 293954 7296 294574 7380
rect 293954 7060 293986 7296
rect 294222 7060 294306 7296
rect 294542 7060 294574 7296
rect 293954 -4184 294574 7060
rect 293954 -4420 293986 -4184
rect 294222 -4420 294306 -4184
rect 294542 -4420 294574 -4184
rect 293954 -4504 294574 -4420
rect 293954 -4740 293986 -4504
rect 294222 -4740 294306 -4504
rect 294542 -4740 294574 -4504
rect 293954 -7652 294574 -4740
rect 295194 709640 295814 711592
rect 295194 709404 295226 709640
rect 295462 709404 295546 709640
rect 295782 709404 295814 709640
rect 295194 709320 295814 709404
rect 295194 709084 295226 709320
rect 295462 709084 295546 709320
rect 295782 709084 295814 709320
rect 295194 692856 295814 709084
rect 295194 692620 295226 692856
rect 295462 692620 295546 692856
rect 295782 692620 295814 692856
rect 295194 692536 295814 692620
rect 295194 692300 295226 692536
rect 295462 692300 295546 692536
rect 295782 692300 295814 692536
rect 295194 656856 295814 692300
rect 295194 656620 295226 656856
rect 295462 656620 295546 656856
rect 295782 656620 295814 656856
rect 295194 656536 295814 656620
rect 295194 656300 295226 656536
rect 295462 656300 295546 656536
rect 295782 656300 295814 656536
rect 295194 620856 295814 656300
rect 295194 620620 295226 620856
rect 295462 620620 295546 620856
rect 295782 620620 295814 620856
rect 295194 620536 295814 620620
rect 295194 620300 295226 620536
rect 295462 620300 295546 620536
rect 295782 620300 295814 620536
rect 295194 584856 295814 620300
rect 295194 584620 295226 584856
rect 295462 584620 295546 584856
rect 295782 584620 295814 584856
rect 295194 584536 295814 584620
rect 295194 584300 295226 584536
rect 295462 584300 295546 584536
rect 295782 584300 295814 584536
rect 295194 548856 295814 584300
rect 295194 548620 295226 548856
rect 295462 548620 295546 548856
rect 295782 548620 295814 548856
rect 295194 548536 295814 548620
rect 295194 548300 295226 548536
rect 295462 548300 295546 548536
rect 295782 548300 295814 548536
rect 295194 512856 295814 548300
rect 295194 512620 295226 512856
rect 295462 512620 295546 512856
rect 295782 512620 295814 512856
rect 295194 512536 295814 512620
rect 295194 512300 295226 512536
rect 295462 512300 295546 512536
rect 295782 512300 295814 512536
rect 295194 476856 295814 512300
rect 295194 476620 295226 476856
rect 295462 476620 295546 476856
rect 295782 476620 295814 476856
rect 295194 476536 295814 476620
rect 295194 476300 295226 476536
rect 295462 476300 295546 476536
rect 295782 476300 295814 476536
rect 295194 440856 295814 476300
rect 295194 440620 295226 440856
rect 295462 440620 295546 440856
rect 295782 440620 295814 440856
rect 295194 440536 295814 440620
rect 295194 440300 295226 440536
rect 295462 440300 295546 440536
rect 295782 440300 295814 440536
rect 295194 404856 295814 440300
rect 295194 404620 295226 404856
rect 295462 404620 295546 404856
rect 295782 404620 295814 404856
rect 295194 404536 295814 404620
rect 295194 404300 295226 404536
rect 295462 404300 295546 404536
rect 295782 404300 295814 404536
rect 295194 368856 295814 404300
rect 295194 368620 295226 368856
rect 295462 368620 295546 368856
rect 295782 368620 295814 368856
rect 295194 368536 295814 368620
rect 295194 368300 295226 368536
rect 295462 368300 295546 368536
rect 295782 368300 295814 368536
rect 295194 332856 295814 368300
rect 295194 332620 295226 332856
rect 295462 332620 295546 332856
rect 295782 332620 295814 332856
rect 295194 332536 295814 332620
rect 295194 332300 295226 332536
rect 295462 332300 295546 332536
rect 295782 332300 295814 332536
rect 295194 296856 295814 332300
rect 295194 296620 295226 296856
rect 295462 296620 295546 296856
rect 295782 296620 295814 296856
rect 295194 296536 295814 296620
rect 295194 296300 295226 296536
rect 295462 296300 295546 296536
rect 295782 296300 295814 296536
rect 295194 260856 295814 296300
rect 295194 260620 295226 260856
rect 295462 260620 295546 260856
rect 295782 260620 295814 260856
rect 295194 260536 295814 260620
rect 295194 260300 295226 260536
rect 295462 260300 295546 260536
rect 295782 260300 295814 260536
rect 295194 224856 295814 260300
rect 295194 224620 295226 224856
rect 295462 224620 295546 224856
rect 295782 224620 295814 224856
rect 295194 224536 295814 224620
rect 295194 224300 295226 224536
rect 295462 224300 295546 224536
rect 295782 224300 295814 224536
rect 295194 188856 295814 224300
rect 295194 188620 295226 188856
rect 295462 188620 295546 188856
rect 295782 188620 295814 188856
rect 295194 188536 295814 188620
rect 295194 188300 295226 188536
rect 295462 188300 295546 188536
rect 295782 188300 295814 188536
rect 295194 152856 295814 188300
rect 295194 152620 295226 152856
rect 295462 152620 295546 152856
rect 295782 152620 295814 152856
rect 295194 152536 295814 152620
rect 295194 152300 295226 152536
rect 295462 152300 295546 152536
rect 295782 152300 295814 152536
rect 295194 116856 295814 152300
rect 295194 116620 295226 116856
rect 295462 116620 295546 116856
rect 295782 116620 295814 116856
rect 295194 116536 295814 116620
rect 295194 116300 295226 116536
rect 295462 116300 295546 116536
rect 295782 116300 295814 116536
rect 295194 80856 295814 116300
rect 295194 80620 295226 80856
rect 295462 80620 295546 80856
rect 295782 80620 295814 80856
rect 295194 80536 295814 80620
rect 295194 80300 295226 80536
rect 295462 80300 295546 80536
rect 295782 80300 295814 80536
rect 295194 44856 295814 80300
rect 295194 44620 295226 44856
rect 295462 44620 295546 44856
rect 295782 44620 295814 44856
rect 295194 44536 295814 44620
rect 295194 44300 295226 44536
rect 295462 44300 295546 44536
rect 295782 44300 295814 44536
rect 295194 8856 295814 44300
rect 295194 8620 295226 8856
rect 295462 8620 295546 8856
rect 295782 8620 295814 8856
rect 295194 8536 295814 8620
rect 295194 8300 295226 8536
rect 295462 8300 295546 8536
rect 295782 8300 295814 8536
rect 295194 -5144 295814 8300
rect 295194 -5380 295226 -5144
rect 295462 -5380 295546 -5144
rect 295782 -5380 295814 -5144
rect 295194 -5464 295814 -5380
rect 295194 -5700 295226 -5464
rect 295462 -5700 295546 -5464
rect 295782 -5700 295814 -5464
rect 295194 -7652 295814 -5700
rect 296434 710600 297054 711592
rect 296434 710364 296466 710600
rect 296702 710364 296786 710600
rect 297022 710364 297054 710600
rect 296434 710280 297054 710364
rect 296434 710044 296466 710280
rect 296702 710044 296786 710280
rect 297022 710044 297054 710280
rect 296434 694096 297054 710044
rect 296434 693860 296466 694096
rect 296702 693860 296786 694096
rect 297022 693860 297054 694096
rect 296434 693776 297054 693860
rect 296434 693540 296466 693776
rect 296702 693540 296786 693776
rect 297022 693540 297054 693776
rect 296434 658096 297054 693540
rect 296434 657860 296466 658096
rect 296702 657860 296786 658096
rect 297022 657860 297054 658096
rect 296434 657776 297054 657860
rect 296434 657540 296466 657776
rect 296702 657540 296786 657776
rect 297022 657540 297054 657776
rect 296434 622096 297054 657540
rect 296434 621860 296466 622096
rect 296702 621860 296786 622096
rect 297022 621860 297054 622096
rect 296434 621776 297054 621860
rect 296434 621540 296466 621776
rect 296702 621540 296786 621776
rect 297022 621540 297054 621776
rect 296434 586096 297054 621540
rect 296434 585860 296466 586096
rect 296702 585860 296786 586096
rect 297022 585860 297054 586096
rect 296434 585776 297054 585860
rect 296434 585540 296466 585776
rect 296702 585540 296786 585776
rect 297022 585540 297054 585776
rect 296434 550096 297054 585540
rect 296434 549860 296466 550096
rect 296702 549860 296786 550096
rect 297022 549860 297054 550096
rect 296434 549776 297054 549860
rect 296434 549540 296466 549776
rect 296702 549540 296786 549776
rect 297022 549540 297054 549776
rect 296434 514096 297054 549540
rect 296434 513860 296466 514096
rect 296702 513860 296786 514096
rect 297022 513860 297054 514096
rect 296434 513776 297054 513860
rect 296434 513540 296466 513776
rect 296702 513540 296786 513776
rect 297022 513540 297054 513776
rect 296434 478096 297054 513540
rect 296434 477860 296466 478096
rect 296702 477860 296786 478096
rect 297022 477860 297054 478096
rect 296434 477776 297054 477860
rect 296434 477540 296466 477776
rect 296702 477540 296786 477776
rect 297022 477540 297054 477776
rect 296434 442096 297054 477540
rect 296434 441860 296466 442096
rect 296702 441860 296786 442096
rect 297022 441860 297054 442096
rect 296434 441776 297054 441860
rect 296434 441540 296466 441776
rect 296702 441540 296786 441776
rect 297022 441540 297054 441776
rect 296434 406096 297054 441540
rect 296434 405860 296466 406096
rect 296702 405860 296786 406096
rect 297022 405860 297054 406096
rect 296434 405776 297054 405860
rect 296434 405540 296466 405776
rect 296702 405540 296786 405776
rect 297022 405540 297054 405776
rect 296434 370096 297054 405540
rect 296434 369860 296466 370096
rect 296702 369860 296786 370096
rect 297022 369860 297054 370096
rect 296434 369776 297054 369860
rect 296434 369540 296466 369776
rect 296702 369540 296786 369776
rect 297022 369540 297054 369776
rect 296434 334096 297054 369540
rect 296434 333860 296466 334096
rect 296702 333860 296786 334096
rect 297022 333860 297054 334096
rect 296434 333776 297054 333860
rect 296434 333540 296466 333776
rect 296702 333540 296786 333776
rect 297022 333540 297054 333776
rect 296434 298096 297054 333540
rect 296434 297860 296466 298096
rect 296702 297860 296786 298096
rect 297022 297860 297054 298096
rect 296434 297776 297054 297860
rect 296434 297540 296466 297776
rect 296702 297540 296786 297776
rect 297022 297540 297054 297776
rect 296434 262096 297054 297540
rect 296434 261860 296466 262096
rect 296702 261860 296786 262096
rect 297022 261860 297054 262096
rect 296434 261776 297054 261860
rect 296434 261540 296466 261776
rect 296702 261540 296786 261776
rect 297022 261540 297054 261776
rect 296434 226096 297054 261540
rect 296434 225860 296466 226096
rect 296702 225860 296786 226096
rect 297022 225860 297054 226096
rect 296434 225776 297054 225860
rect 296434 225540 296466 225776
rect 296702 225540 296786 225776
rect 297022 225540 297054 225776
rect 296434 190096 297054 225540
rect 296434 189860 296466 190096
rect 296702 189860 296786 190096
rect 297022 189860 297054 190096
rect 296434 189776 297054 189860
rect 296434 189540 296466 189776
rect 296702 189540 296786 189776
rect 297022 189540 297054 189776
rect 296434 154096 297054 189540
rect 296434 153860 296466 154096
rect 296702 153860 296786 154096
rect 297022 153860 297054 154096
rect 296434 153776 297054 153860
rect 296434 153540 296466 153776
rect 296702 153540 296786 153776
rect 297022 153540 297054 153776
rect 296434 118096 297054 153540
rect 296434 117860 296466 118096
rect 296702 117860 296786 118096
rect 297022 117860 297054 118096
rect 296434 117776 297054 117860
rect 296434 117540 296466 117776
rect 296702 117540 296786 117776
rect 297022 117540 297054 117776
rect 296434 82096 297054 117540
rect 296434 81860 296466 82096
rect 296702 81860 296786 82096
rect 297022 81860 297054 82096
rect 296434 81776 297054 81860
rect 296434 81540 296466 81776
rect 296702 81540 296786 81776
rect 297022 81540 297054 81776
rect 296434 46096 297054 81540
rect 296434 45860 296466 46096
rect 296702 45860 296786 46096
rect 297022 45860 297054 46096
rect 296434 45776 297054 45860
rect 296434 45540 296466 45776
rect 296702 45540 296786 45776
rect 297022 45540 297054 45776
rect 296434 10096 297054 45540
rect 296434 9860 296466 10096
rect 296702 9860 296786 10096
rect 297022 9860 297054 10096
rect 296434 9776 297054 9860
rect 296434 9540 296466 9776
rect 296702 9540 296786 9776
rect 297022 9540 297054 9776
rect 296434 -6104 297054 9540
rect 296434 -6340 296466 -6104
rect 296702 -6340 296786 -6104
rect 297022 -6340 297054 -6104
rect 296434 -6424 297054 -6340
rect 296434 -6660 296466 -6424
rect 296702 -6660 296786 -6424
rect 297022 -6660 297054 -6424
rect 296434 -7652 297054 -6660
rect 297674 711560 298294 711592
rect 297674 711324 297706 711560
rect 297942 711324 298026 711560
rect 298262 711324 298294 711560
rect 297674 711240 298294 711324
rect 297674 711004 297706 711240
rect 297942 711004 298026 711240
rect 298262 711004 298294 711240
rect 297674 695336 298294 711004
rect 297674 695100 297706 695336
rect 297942 695100 298026 695336
rect 298262 695100 298294 695336
rect 297674 695016 298294 695100
rect 297674 694780 297706 695016
rect 297942 694780 298026 695016
rect 298262 694780 298294 695016
rect 297674 659336 298294 694780
rect 297674 659100 297706 659336
rect 297942 659100 298026 659336
rect 298262 659100 298294 659336
rect 297674 659016 298294 659100
rect 297674 658780 297706 659016
rect 297942 658780 298026 659016
rect 298262 658780 298294 659016
rect 297674 623336 298294 658780
rect 297674 623100 297706 623336
rect 297942 623100 298026 623336
rect 298262 623100 298294 623336
rect 297674 623016 298294 623100
rect 297674 622780 297706 623016
rect 297942 622780 298026 623016
rect 298262 622780 298294 623016
rect 297674 587336 298294 622780
rect 297674 587100 297706 587336
rect 297942 587100 298026 587336
rect 298262 587100 298294 587336
rect 297674 587016 298294 587100
rect 297674 586780 297706 587016
rect 297942 586780 298026 587016
rect 298262 586780 298294 587016
rect 297674 551336 298294 586780
rect 297674 551100 297706 551336
rect 297942 551100 298026 551336
rect 298262 551100 298294 551336
rect 297674 551016 298294 551100
rect 297674 550780 297706 551016
rect 297942 550780 298026 551016
rect 298262 550780 298294 551016
rect 297674 515336 298294 550780
rect 297674 515100 297706 515336
rect 297942 515100 298026 515336
rect 298262 515100 298294 515336
rect 297674 515016 298294 515100
rect 297674 514780 297706 515016
rect 297942 514780 298026 515016
rect 298262 514780 298294 515016
rect 297674 479336 298294 514780
rect 297674 479100 297706 479336
rect 297942 479100 298026 479336
rect 298262 479100 298294 479336
rect 297674 479016 298294 479100
rect 297674 478780 297706 479016
rect 297942 478780 298026 479016
rect 298262 478780 298294 479016
rect 297674 443336 298294 478780
rect 297674 443100 297706 443336
rect 297942 443100 298026 443336
rect 298262 443100 298294 443336
rect 297674 443016 298294 443100
rect 297674 442780 297706 443016
rect 297942 442780 298026 443016
rect 298262 442780 298294 443016
rect 297674 407336 298294 442780
rect 297674 407100 297706 407336
rect 297942 407100 298026 407336
rect 298262 407100 298294 407336
rect 297674 407016 298294 407100
rect 297674 406780 297706 407016
rect 297942 406780 298026 407016
rect 298262 406780 298294 407016
rect 297674 371336 298294 406780
rect 297674 371100 297706 371336
rect 297942 371100 298026 371336
rect 298262 371100 298294 371336
rect 297674 371016 298294 371100
rect 297674 370780 297706 371016
rect 297942 370780 298026 371016
rect 298262 370780 298294 371016
rect 297674 335336 298294 370780
rect 297674 335100 297706 335336
rect 297942 335100 298026 335336
rect 298262 335100 298294 335336
rect 297674 335016 298294 335100
rect 297674 334780 297706 335016
rect 297942 334780 298026 335016
rect 298262 334780 298294 335016
rect 297674 299336 298294 334780
rect 297674 299100 297706 299336
rect 297942 299100 298026 299336
rect 298262 299100 298294 299336
rect 297674 299016 298294 299100
rect 297674 298780 297706 299016
rect 297942 298780 298026 299016
rect 298262 298780 298294 299016
rect 297674 263336 298294 298780
rect 297674 263100 297706 263336
rect 297942 263100 298026 263336
rect 298262 263100 298294 263336
rect 297674 263016 298294 263100
rect 297674 262780 297706 263016
rect 297942 262780 298026 263016
rect 298262 262780 298294 263016
rect 297674 227336 298294 262780
rect 297674 227100 297706 227336
rect 297942 227100 298026 227336
rect 298262 227100 298294 227336
rect 297674 227016 298294 227100
rect 297674 226780 297706 227016
rect 297942 226780 298026 227016
rect 298262 226780 298294 227016
rect 297674 191336 298294 226780
rect 297674 191100 297706 191336
rect 297942 191100 298026 191336
rect 298262 191100 298294 191336
rect 297674 191016 298294 191100
rect 297674 190780 297706 191016
rect 297942 190780 298026 191016
rect 298262 190780 298294 191016
rect 297674 155336 298294 190780
rect 297674 155100 297706 155336
rect 297942 155100 298026 155336
rect 298262 155100 298294 155336
rect 297674 155016 298294 155100
rect 297674 154780 297706 155016
rect 297942 154780 298026 155016
rect 298262 154780 298294 155016
rect 297674 119336 298294 154780
rect 297674 119100 297706 119336
rect 297942 119100 298026 119336
rect 298262 119100 298294 119336
rect 297674 119016 298294 119100
rect 297674 118780 297706 119016
rect 297942 118780 298026 119016
rect 298262 118780 298294 119016
rect 297674 83336 298294 118780
rect 297674 83100 297706 83336
rect 297942 83100 298026 83336
rect 298262 83100 298294 83336
rect 297674 83016 298294 83100
rect 297674 82780 297706 83016
rect 297942 82780 298026 83016
rect 298262 82780 298294 83016
rect 297674 47336 298294 82780
rect 297674 47100 297706 47336
rect 297942 47100 298026 47336
rect 298262 47100 298294 47336
rect 297674 47016 298294 47100
rect 297674 46780 297706 47016
rect 297942 46780 298026 47016
rect 298262 46780 298294 47016
rect 297674 11336 298294 46780
rect 297674 11100 297706 11336
rect 297942 11100 298026 11336
rect 298262 11100 298294 11336
rect 297674 11016 298294 11100
rect 297674 10780 297706 11016
rect 297942 10780 298026 11016
rect 298262 10780 298294 11016
rect 297674 -7064 298294 10780
rect 297674 -7300 297706 -7064
rect 297942 -7300 298026 -7064
rect 298262 -7300 298294 -7064
rect 297674 -7384 298294 -7300
rect 297674 -7620 297706 -7384
rect 297942 -7620 298026 -7384
rect 298262 -7620 298294 -7384
rect 297674 -7652 298294 -7620
rect 324994 704840 325614 711592
rect 324994 704604 325026 704840
rect 325262 704604 325346 704840
rect 325582 704604 325614 704840
rect 324994 704520 325614 704604
rect 324994 704284 325026 704520
rect 325262 704284 325346 704520
rect 325582 704284 325614 704520
rect 324994 702608 325614 704284
rect 324994 702544 325032 702608
rect 325096 702544 325112 702608
rect 325176 702544 325192 702608
rect 325256 702544 325272 702608
rect 325336 702544 325352 702608
rect 325416 702544 325432 702608
rect 325496 702544 325512 702608
rect 325576 702544 325614 702608
rect 324994 702528 325614 702544
rect 324994 702464 325032 702528
rect 325096 702464 325112 702528
rect 325176 702464 325192 702528
rect 325256 702464 325272 702528
rect 325336 702464 325352 702528
rect 325416 702464 325432 702528
rect 325496 702464 325512 702528
rect 325576 702464 325614 702528
rect 324994 702448 325614 702464
rect 324994 702384 325032 702448
rect 325096 702384 325112 702448
rect 325176 702384 325192 702448
rect 325256 702384 325272 702448
rect 325336 702384 325352 702448
rect 325416 702384 325432 702448
rect 325496 702384 325512 702448
rect 325576 702384 325614 702448
rect 324994 702368 325614 702384
rect 324994 702304 325032 702368
rect 325096 702304 325112 702368
rect 325176 702304 325192 702368
rect 325256 702304 325272 702368
rect 325336 702304 325352 702368
rect 325416 702304 325432 702368
rect 325496 702304 325512 702368
rect 325576 702304 325614 702368
rect 324994 686656 325614 702304
rect 324994 686420 325026 686656
rect 325262 686420 325346 686656
rect 325582 686420 325614 686656
rect 324994 686336 325614 686420
rect 324994 686100 325026 686336
rect 325262 686100 325346 686336
rect 325582 686100 325614 686336
rect 324994 650656 325614 686100
rect 324994 650420 325026 650656
rect 325262 650420 325346 650656
rect 325582 650420 325614 650656
rect 324994 650336 325614 650420
rect 324994 650100 325026 650336
rect 325262 650100 325346 650336
rect 325582 650100 325614 650336
rect 324994 614656 325614 650100
rect 324994 614420 325026 614656
rect 325262 614420 325346 614656
rect 325582 614420 325614 614656
rect 324994 614336 325614 614420
rect 324994 614100 325026 614336
rect 325262 614100 325346 614336
rect 325582 614100 325614 614336
rect 324994 578656 325614 614100
rect 324994 578420 325026 578656
rect 325262 578420 325346 578656
rect 325582 578420 325614 578656
rect 324994 578336 325614 578420
rect 324994 578100 325026 578336
rect 325262 578100 325346 578336
rect 325582 578100 325614 578336
rect 324994 542656 325614 578100
rect 324994 542420 325026 542656
rect 325262 542420 325346 542656
rect 325582 542420 325614 542656
rect 324994 542336 325614 542420
rect 324994 542100 325026 542336
rect 325262 542100 325346 542336
rect 325582 542100 325614 542336
rect 324994 506656 325614 542100
rect 324994 506420 325026 506656
rect 325262 506420 325346 506656
rect 325582 506420 325614 506656
rect 324994 506336 325614 506420
rect 324994 506100 325026 506336
rect 325262 506100 325346 506336
rect 325582 506100 325614 506336
rect 324994 470656 325614 506100
rect 324994 470420 325026 470656
rect 325262 470420 325346 470656
rect 325582 470420 325614 470656
rect 324994 470336 325614 470420
rect 324994 470100 325026 470336
rect 325262 470100 325346 470336
rect 325582 470100 325614 470336
rect 324994 434656 325614 470100
rect 324994 434420 325026 434656
rect 325262 434420 325346 434656
rect 325582 434420 325614 434656
rect 324994 434336 325614 434420
rect 324994 434100 325026 434336
rect 325262 434100 325346 434336
rect 325582 434100 325614 434336
rect 324994 398656 325614 434100
rect 324994 398420 325026 398656
rect 325262 398420 325346 398656
rect 325582 398420 325614 398656
rect 324994 398336 325614 398420
rect 324994 398100 325026 398336
rect 325262 398100 325346 398336
rect 325582 398100 325614 398336
rect 324994 362656 325614 398100
rect 324994 362420 325026 362656
rect 325262 362420 325346 362656
rect 325582 362420 325614 362656
rect 324994 362336 325614 362420
rect 324994 362100 325026 362336
rect 325262 362100 325346 362336
rect 325582 362100 325614 362336
rect 324994 326656 325614 362100
rect 324994 326420 325026 326656
rect 325262 326420 325346 326656
rect 325582 326420 325614 326656
rect 324994 326336 325614 326420
rect 324994 326100 325026 326336
rect 325262 326100 325346 326336
rect 325582 326100 325614 326336
rect 324994 290656 325614 326100
rect 324994 290420 325026 290656
rect 325262 290420 325346 290656
rect 325582 290420 325614 290656
rect 324994 290336 325614 290420
rect 324994 290100 325026 290336
rect 325262 290100 325346 290336
rect 325582 290100 325614 290336
rect 324994 254656 325614 290100
rect 324994 254420 325026 254656
rect 325262 254420 325346 254656
rect 325582 254420 325614 254656
rect 324994 254336 325614 254420
rect 324994 254100 325026 254336
rect 325262 254100 325346 254336
rect 325582 254100 325614 254336
rect 324994 218656 325614 254100
rect 324994 218420 325026 218656
rect 325262 218420 325346 218656
rect 325582 218420 325614 218656
rect 324994 218336 325614 218420
rect 324994 218100 325026 218336
rect 325262 218100 325346 218336
rect 325582 218100 325614 218336
rect 324994 182656 325614 218100
rect 324994 182420 325026 182656
rect 325262 182420 325346 182656
rect 325582 182420 325614 182656
rect 324994 182336 325614 182420
rect 324994 182100 325026 182336
rect 325262 182100 325346 182336
rect 325582 182100 325614 182336
rect 324994 146656 325614 182100
rect 324994 146420 325026 146656
rect 325262 146420 325346 146656
rect 325582 146420 325614 146656
rect 324994 146336 325614 146420
rect 324994 146100 325026 146336
rect 325262 146100 325346 146336
rect 325582 146100 325614 146336
rect 324994 110656 325614 146100
rect 324994 110420 325026 110656
rect 325262 110420 325346 110656
rect 325582 110420 325614 110656
rect 324994 110336 325614 110420
rect 324994 110100 325026 110336
rect 325262 110100 325346 110336
rect 325582 110100 325614 110336
rect 324994 74656 325614 110100
rect 324994 74420 325026 74656
rect 325262 74420 325346 74656
rect 325582 74420 325614 74656
rect 324994 74336 325614 74420
rect 324994 74100 325026 74336
rect 325262 74100 325346 74336
rect 325582 74100 325614 74336
rect 324994 38656 325614 74100
rect 324994 38420 325026 38656
rect 325262 38420 325346 38656
rect 325582 38420 325614 38656
rect 324994 38336 325614 38420
rect 324994 38100 325026 38336
rect 325262 38100 325346 38336
rect 325582 38100 325614 38336
rect 324994 2656 325614 38100
rect 324994 2420 325026 2656
rect 325262 2420 325346 2656
rect 325582 2420 325614 2656
rect 324994 2336 325614 2420
rect 324994 2100 325026 2336
rect 325262 2100 325346 2336
rect 325582 2100 325614 2336
rect 324994 -344 325614 2100
rect 324994 -580 325026 -344
rect 325262 -580 325346 -344
rect 325582 -580 325614 -344
rect 324994 -664 325614 -580
rect 324994 -900 325026 -664
rect 325262 -900 325346 -664
rect 325582 -900 325614 -664
rect 324994 -7652 325614 -900
rect 326234 705800 326854 711592
rect 326234 705564 326266 705800
rect 326502 705564 326586 705800
rect 326822 705564 326854 705800
rect 326234 705480 326854 705564
rect 326234 705244 326266 705480
rect 326502 705244 326586 705480
rect 326822 705244 326854 705480
rect 326234 703376 326854 705244
rect 326234 703312 326272 703376
rect 326336 703312 326352 703376
rect 326416 703312 326432 703376
rect 326496 703312 326512 703376
rect 326576 703312 326592 703376
rect 326656 703312 326672 703376
rect 326736 703312 326752 703376
rect 326816 703312 326854 703376
rect 326234 703296 326854 703312
rect 326234 703232 326272 703296
rect 326336 703232 326352 703296
rect 326416 703232 326432 703296
rect 326496 703232 326512 703296
rect 326576 703232 326592 703296
rect 326656 703232 326672 703296
rect 326736 703232 326752 703296
rect 326816 703232 326854 703296
rect 326234 703216 326854 703232
rect 326234 703152 326272 703216
rect 326336 703152 326352 703216
rect 326416 703152 326432 703216
rect 326496 703152 326512 703216
rect 326576 703152 326592 703216
rect 326656 703152 326672 703216
rect 326736 703152 326752 703216
rect 326816 703152 326854 703216
rect 326234 703136 326854 703152
rect 326234 703072 326272 703136
rect 326336 703072 326352 703136
rect 326416 703072 326432 703136
rect 326496 703072 326512 703136
rect 326576 703072 326592 703136
rect 326656 703072 326672 703136
rect 326736 703072 326752 703136
rect 326816 703072 326854 703136
rect 326234 687896 326854 703072
rect 326234 687660 326266 687896
rect 326502 687660 326586 687896
rect 326822 687660 326854 687896
rect 326234 687576 326854 687660
rect 326234 687340 326266 687576
rect 326502 687340 326586 687576
rect 326822 687340 326854 687576
rect 326234 651896 326854 687340
rect 326234 651660 326266 651896
rect 326502 651660 326586 651896
rect 326822 651660 326854 651896
rect 326234 651576 326854 651660
rect 326234 651340 326266 651576
rect 326502 651340 326586 651576
rect 326822 651340 326854 651576
rect 326234 615896 326854 651340
rect 326234 615660 326266 615896
rect 326502 615660 326586 615896
rect 326822 615660 326854 615896
rect 326234 615576 326854 615660
rect 326234 615340 326266 615576
rect 326502 615340 326586 615576
rect 326822 615340 326854 615576
rect 326234 579896 326854 615340
rect 326234 579660 326266 579896
rect 326502 579660 326586 579896
rect 326822 579660 326854 579896
rect 326234 579576 326854 579660
rect 326234 579340 326266 579576
rect 326502 579340 326586 579576
rect 326822 579340 326854 579576
rect 326234 543896 326854 579340
rect 326234 543660 326266 543896
rect 326502 543660 326586 543896
rect 326822 543660 326854 543896
rect 326234 543576 326854 543660
rect 326234 543340 326266 543576
rect 326502 543340 326586 543576
rect 326822 543340 326854 543576
rect 326234 507896 326854 543340
rect 326234 507660 326266 507896
rect 326502 507660 326586 507896
rect 326822 507660 326854 507896
rect 326234 507576 326854 507660
rect 326234 507340 326266 507576
rect 326502 507340 326586 507576
rect 326822 507340 326854 507576
rect 326234 471896 326854 507340
rect 326234 471660 326266 471896
rect 326502 471660 326586 471896
rect 326822 471660 326854 471896
rect 326234 471576 326854 471660
rect 326234 471340 326266 471576
rect 326502 471340 326586 471576
rect 326822 471340 326854 471576
rect 326234 435896 326854 471340
rect 326234 435660 326266 435896
rect 326502 435660 326586 435896
rect 326822 435660 326854 435896
rect 326234 435576 326854 435660
rect 326234 435340 326266 435576
rect 326502 435340 326586 435576
rect 326822 435340 326854 435576
rect 326234 399896 326854 435340
rect 326234 399660 326266 399896
rect 326502 399660 326586 399896
rect 326822 399660 326854 399896
rect 326234 399576 326854 399660
rect 326234 399340 326266 399576
rect 326502 399340 326586 399576
rect 326822 399340 326854 399576
rect 326234 363896 326854 399340
rect 326234 363660 326266 363896
rect 326502 363660 326586 363896
rect 326822 363660 326854 363896
rect 326234 363576 326854 363660
rect 326234 363340 326266 363576
rect 326502 363340 326586 363576
rect 326822 363340 326854 363576
rect 326234 327896 326854 363340
rect 326234 327660 326266 327896
rect 326502 327660 326586 327896
rect 326822 327660 326854 327896
rect 326234 327576 326854 327660
rect 326234 327340 326266 327576
rect 326502 327340 326586 327576
rect 326822 327340 326854 327576
rect 326234 291896 326854 327340
rect 326234 291660 326266 291896
rect 326502 291660 326586 291896
rect 326822 291660 326854 291896
rect 326234 291576 326854 291660
rect 326234 291340 326266 291576
rect 326502 291340 326586 291576
rect 326822 291340 326854 291576
rect 326234 255896 326854 291340
rect 326234 255660 326266 255896
rect 326502 255660 326586 255896
rect 326822 255660 326854 255896
rect 326234 255576 326854 255660
rect 326234 255340 326266 255576
rect 326502 255340 326586 255576
rect 326822 255340 326854 255576
rect 326234 219896 326854 255340
rect 326234 219660 326266 219896
rect 326502 219660 326586 219896
rect 326822 219660 326854 219896
rect 326234 219576 326854 219660
rect 326234 219340 326266 219576
rect 326502 219340 326586 219576
rect 326822 219340 326854 219576
rect 326234 183896 326854 219340
rect 326234 183660 326266 183896
rect 326502 183660 326586 183896
rect 326822 183660 326854 183896
rect 326234 183576 326854 183660
rect 326234 183340 326266 183576
rect 326502 183340 326586 183576
rect 326822 183340 326854 183576
rect 326234 147896 326854 183340
rect 326234 147660 326266 147896
rect 326502 147660 326586 147896
rect 326822 147660 326854 147896
rect 326234 147576 326854 147660
rect 326234 147340 326266 147576
rect 326502 147340 326586 147576
rect 326822 147340 326854 147576
rect 326234 111896 326854 147340
rect 326234 111660 326266 111896
rect 326502 111660 326586 111896
rect 326822 111660 326854 111896
rect 326234 111576 326854 111660
rect 326234 111340 326266 111576
rect 326502 111340 326586 111576
rect 326822 111340 326854 111576
rect 326234 75896 326854 111340
rect 326234 75660 326266 75896
rect 326502 75660 326586 75896
rect 326822 75660 326854 75896
rect 326234 75576 326854 75660
rect 326234 75340 326266 75576
rect 326502 75340 326586 75576
rect 326822 75340 326854 75576
rect 326234 39896 326854 75340
rect 326234 39660 326266 39896
rect 326502 39660 326586 39896
rect 326822 39660 326854 39896
rect 326234 39576 326854 39660
rect 326234 39340 326266 39576
rect 326502 39340 326586 39576
rect 326822 39340 326854 39576
rect 326234 3896 326854 39340
rect 326234 3660 326266 3896
rect 326502 3660 326586 3896
rect 326822 3660 326854 3896
rect 326234 3576 326854 3660
rect 326234 3340 326266 3576
rect 326502 3340 326586 3576
rect 326822 3340 326854 3576
rect 326234 -1304 326854 3340
rect 326234 -1540 326266 -1304
rect 326502 -1540 326586 -1304
rect 326822 -1540 326854 -1304
rect 326234 -1624 326854 -1540
rect 326234 -1860 326266 -1624
rect 326502 -1860 326586 -1624
rect 326822 -1860 326854 -1624
rect 326234 -7652 326854 -1860
rect 327474 706760 328094 711592
rect 327474 706524 327506 706760
rect 327742 706524 327826 706760
rect 328062 706524 328094 706760
rect 327474 706440 328094 706524
rect 327474 706204 327506 706440
rect 327742 706204 327826 706440
rect 328062 706204 328094 706440
rect 327474 689136 328094 706204
rect 327474 688900 327506 689136
rect 327742 688900 327826 689136
rect 328062 688900 328094 689136
rect 327474 688816 328094 688900
rect 327474 688580 327506 688816
rect 327742 688580 327826 688816
rect 328062 688580 328094 688816
rect 327474 653136 328094 688580
rect 327474 652900 327506 653136
rect 327742 652900 327826 653136
rect 328062 652900 328094 653136
rect 327474 652816 328094 652900
rect 327474 652580 327506 652816
rect 327742 652580 327826 652816
rect 328062 652580 328094 652816
rect 327474 617136 328094 652580
rect 327474 616900 327506 617136
rect 327742 616900 327826 617136
rect 328062 616900 328094 617136
rect 327474 616816 328094 616900
rect 327474 616580 327506 616816
rect 327742 616580 327826 616816
rect 328062 616580 328094 616816
rect 327474 581136 328094 616580
rect 327474 580900 327506 581136
rect 327742 580900 327826 581136
rect 328062 580900 328094 581136
rect 327474 580816 328094 580900
rect 327474 580580 327506 580816
rect 327742 580580 327826 580816
rect 328062 580580 328094 580816
rect 327474 545136 328094 580580
rect 327474 544900 327506 545136
rect 327742 544900 327826 545136
rect 328062 544900 328094 545136
rect 327474 544816 328094 544900
rect 327474 544580 327506 544816
rect 327742 544580 327826 544816
rect 328062 544580 328094 544816
rect 327474 509136 328094 544580
rect 327474 508900 327506 509136
rect 327742 508900 327826 509136
rect 328062 508900 328094 509136
rect 327474 508816 328094 508900
rect 327474 508580 327506 508816
rect 327742 508580 327826 508816
rect 328062 508580 328094 508816
rect 327474 473136 328094 508580
rect 327474 472900 327506 473136
rect 327742 472900 327826 473136
rect 328062 472900 328094 473136
rect 327474 472816 328094 472900
rect 327474 472580 327506 472816
rect 327742 472580 327826 472816
rect 328062 472580 328094 472816
rect 327474 437136 328094 472580
rect 327474 436900 327506 437136
rect 327742 436900 327826 437136
rect 328062 436900 328094 437136
rect 327474 436816 328094 436900
rect 327474 436580 327506 436816
rect 327742 436580 327826 436816
rect 328062 436580 328094 436816
rect 327474 401136 328094 436580
rect 327474 400900 327506 401136
rect 327742 400900 327826 401136
rect 328062 400900 328094 401136
rect 327474 400816 328094 400900
rect 327474 400580 327506 400816
rect 327742 400580 327826 400816
rect 328062 400580 328094 400816
rect 327474 365136 328094 400580
rect 327474 364900 327506 365136
rect 327742 364900 327826 365136
rect 328062 364900 328094 365136
rect 327474 364816 328094 364900
rect 327474 364580 327506 364816
rect 327742 364580 327826 364816
rect 328062 364580 328094 364816
rect 327474 329136 328094 364580
rect 327474 328900 327506 329136
rect 327742 328900 327826 329136
rect 328062 328900 328094 329136
rect 327474 328816 328094 328900
rect 327474 328580 327506 328816
rect 327742 328580 327826 328816
rect 328062 328580 328094 328816
rect 327474 293136 328094 328580
rect 327474 292900 327506 293136
rect 327742 292900 327826 293136
rect 328062 292900 328094 293136
rect 327474 292816 328094 292900
rect 327474 292580 327506 292816
rect 327742 292580 327826 292816
rect 328062 292580 328094 292816
rect 327474 257136 328094 292580
rect 327474 256900 327506 257136
rect 327742 256900 327826 257136
rect 328062 256900 328094 257136
rect 327474 256816 328094 256900
rect 327474 256580 327506 256816
rect 327742 256580 327826 256816
rect 328062 256580 328094 256816
rect 327474 221136 328094 256580
rect 327474 220900 327506 221136
rect 327742 220900 327826 221136
rect 328062 220900 328094 221136
rect 327474 220816 328094 220900
rect 327474 220580 327506 220816
rect 327742 220580 327826 220816
rect 328062 220580 328094 220816
rect 327474 185136 328094 220580
rect 327474 184900 327506 185136
rect 327742 184900 327826 185136
rect 328062 184900 328094 185136
rect 327474 184816 328094 184900
rect 327474 184580 327506 184816
rect 327742 184580 327826 184816
rect 328062 184580 328094 184816
rect 327474 149136 328094 184580
rect 327474 148900 327506 149136
rect 327742 148900 327826 149136
rect 328062 148900 328094 149136
rect 327474 148816 328094 148900
rect 327474 148580 327506 148816
rect 327742 148580 327826 148816
rect 328062 148580 328094 148816
rect 327474 113136 328094 148580
rect 327474 112900 327506 113136
rect 327742 112900 327826 113136
rect 328062 112900 328094 113136
rect 327474 112816 328094 112900
rect 327474 112580 327506 112816
rect 327742 112580 327826 112816
rect 328062 112580 328094 112816
rect 327474 77136 328094 112580
rect 327474 76900 327506 77136
rect 327742 76900 327826 77136
rect 328062 76900 328094 77136
rect 327474 76816 328094 76900
rect 327474 76580 327506 76816
rect 327742 76580 327826 76816
rect 328062 76580 328094 76816
rect 327474 41136 328094 76580
rect 327474 40900 327506 41136
rect 327742 40900 327826 41136
rect 328062 40900 328094 41136
rect 327474 40816 328094 40900
rect 327474 40580 327506 40816
rect 327742 40580 327826 40816
rect 328062 40580 328094 40816
rect 327474 5136 328094 40580
rect 327474 4900 327506 5136
rect 327742 4900 327826 5136
rect 328062 4900 328094 5136
rect 327474 4816 328094 4900
rect 327474 4580 327506 4816
rect 327742 4580 327826 4816
rect 328062 4580 328094 4816
rect 327474 -2264 328094 4580
rect 327474 -2500 327506 -2264
rect 327742 -2500 327826 -2264
rect 328062 -2500 328094 -2264
rect 327474 -2584 328094 -2500
rect 327474 -2820 327506 -2584
rect 327742 -2820 327826 -2584
rect 328062 -2820 328094 -2584
rect 327474 -7652 328094 -2820
rect 328714 707720 329334 711592
rect 328714 707484 328746 707720
rect 328982 707484 329066 707720
rect 329302 707484 329334 707720
rect 328714 707400 329334 707484
rect 328714 707164 328746 707400
rect 328982 707164 329066 707400
rect 329302 707164 329334 707400
rect 328714 690376 329334 707164
rect 328714 690140 328746 690376
rect 328982 690140 329066 690376
rect 329302 690140 329334 690376
rect 328714 690056 329334 690140
rect 328714 689820 328746 690056
rect 328982 689820 329066 690056
rect 329302 689820 329334 690056
rect 328714 654376 329334 689820
rect 328714 654140 328746 654376
rect 328982 654140 329066 654376
rect 329302 654140 329334 654376
rect 328714 654056 329334 654140
rect 328714 653820 328746 654056
rect 328982 653820 329066 654056
rect 329302 653820 329334 654056
rect 328714 618376 329334 653820
rect 328714 618140 328746 618376
rect 328982 618140 329066 618376
rect 329302 618140 329334 618376
rect 328714 618056 329334 618140
rect 328714 617820 328746 618056
rect 328982 617820 329066 618056
rect 329302 617820 329334 618056
rect 328714 582376 329334 617820
rect 328714 582140 328746 582376
rect 328982 582140 329066 582376
rect 329302 582140 329334 582376
rect 328714 582056 329334 582140
rect 328714 581820 328746 582056
rect 328982 581820 329066 582056
rect 329302 581820 329334 582056
rect 328714 546376 329334 581820
rect 328714 546140 328746 546376
rect 328982 546140 329066 546376
rect 329302 546140 329334 546376
rect 328714 546056 329334 546140
rect 328714 545820 328746 546056
rect 328982 545820 329066 546056
rect 329302 545820 329334 546056
rect 328714 510376 329334 545820
rect 328714 510140 328746 510376
rect 328982 510140 329066 510376
rect 329302 510140 329334 510376
rect 328714 510056 329334 510140
rect 328714 509820 328746 510056
rect 328982 509820 329066 510056
rect 329302 509820 329334 510056
rect 328714 474376 329334 509820
rect 328714 474140 328746 474376
rect 328982 474140 329066 474376
rect 329302 474140 329334 474376
rect 328714 474056 329334 474140
rect 328714 473820 328746 474056
rect 328982 473820 329066 474056
rect 329302 473820 329334 474056
rect 328714 438376 329334 473820
rect 328714 438140 328746 438376
rect 328982 438140 329066 438376
rect 329302 438140 329334 438376
rect 328714 438056 329334 438140
rect 328714 437820 328746 438056
rect 328982 437820 329066 438056
rect 329302 437820 329334 438056
rect 328714 402376 329334 437820
rect 328714 402140 328746 402376
rect 328982 402140 329066 402376
rect 329302 402140 329334 402376
rect 328714 402056 329334 402140
rect 328714 401820 328746 402056
rect 328982 401820 329066 402056
rect 329302 401820 329334 402056
rect 328714 366376 329334 401820
rect 328714 366140 328746 366376
rect 328982 366140 329066 366376
rect 329302 366140 329334 366376
rect 328714 366056 329334 366140
rect 328714 365820 328746 366056
rect 328982 365820 329066 366056
rect 329302 365820 329334 366056
rect 328714 330376 329334 365820
rect 328714 330140 328746 330376
rect 328982 330140 329066 330376
rect 329302 330140 329334 330376
rect 328714 330056 329334 330140
rect 328714 329820 328746 330056
rect 328982 329820 329066 330056
rect 329302 329820 329334 330056
rect 328714 294376 329334 329820
rect 328714 294140 328746 294376
rect 328982 294140 329066 294376
rect 329302 294140 329334 294376
rect 328714 294056 329334 294140
rect 328714 293820 328746 294056
rect 328982 293820 329066 294056
rect 329302 293820 329334 294056
rect 328714 258376 329334 293820
rect 328714 258140 328746 258376
rect 328982 258140 329066 258376
rect 329302 258140 329334 258376
rect 328714 258056 329334 258140
rect 328714 257820 328746 258056
rect 328982 257820 329066 258056
rect 329302 257820 329334 258056
rect 328714 222376 329334 257820
rect 328714 222140 328746 222376
rect 328982 222140 329066 222376
rect 329302 222140 329334 222376
rect 328714 222056 329334 222140
rect 328714 221820 328746 222056
rect 328982 221820 329066 222056
rect 329302 221820 329334 222056
rect 328714 186376 329334 221820
rect 328714 186140 328746 186376
rect 328982 186140 329066 186376
rect 329302 186140 329334 186376
rect 328714 186056 329334 186140
rect 328714 185820 328746 186056
rect 328982 185820 329066 186056
rect 329302 185820 329334 186056
rect 328714 150376 329334 185820
rect 328714 150140 328746 150376
rect 328982 150140 329066 150376
rect 329302 150140 329334 150376
rect 328714 150056 329334 150140
rect 328714 149820 328746 150056
rect 328982 149820 329066 150056
rect 329302 149820 329334 150056
rect 328714 114376 329334 149820
rect 328714 114140 328746 114376
rect 328982 114140 329066 114376
rect 329302 114140 329334 114376
rect 328714 114056 329334 114140
rect 328714 113820 328746 114056
rect 328982 113820 329066 114056
rect 329302 113820 329334 114056
rect 328714 78376 329334 113820
rect 328714 78140 328746 78376
rect 328982 78140 329066 78376
rect 329302 78140 329334 78376
rect 328714 78056 329334 78140
rect 328714 77820 328746 78056
rect 328982 77820 329066 78056
rect 329302 77820 329334 78056
rect 328714 42376 329334 77820
rect 328714 42140 328746 42376
rect 328982 42140 329066 42376
rect 329302 42140 329334 42376
rect 328714 42056 329334 42140
rect 328714 41820 328746 42056
rect 328982 41820 329066 42056
rect 329302 41820 329334 42056
rect 328714 6376 329334 41820
rect 328714 6140 328746 6376
rect 328982 6140 329066 6376
rect 329302 6140 329334 6376
rect 328714 6056 329334 6140
rect 328714 5820 328746 6056
rect 328982 5820 329066 6056
rect 329302 5820 329334 6056
rect 328714 -3224 329334 5820
rect 328714 -3460 328746 -3224
rect 328982 -3460 329066 -3224
rect 329302 -3460 329334 -3224
rect 328714 -3544 329334 -3460
rect 328714 -3780 328746 -3544
rect 328982 -3780 329066 -3544
rect 329302 -3780 329334 -3544
rect 328714 -7652 329334 -3780
rect 329954 708680 330574 711592
rect 329954 708444 329986 708680
rect 330222 708444 330306 708680
rect 330542 708444 330574 708680
rect 329954 708360 330574 708444
rect 329954 708124 329986 708360
rect 330222 708124 330306 708360
rect 330542 708124 330574 708360
rect 329954 691616 330574 708124
rect 329954 691380 329986 691616
rect 330222 691380 330306 691616
rect 330542 691380 330574 691616
rect 329954 691296 330574 691380
rect 329954 691060 329986 691296
rect 330222 691060 330306 691296
rect 330542 691060 330574 691296
rect 329954 655616 330574 691060
rect 329954 655380 329986 655616
rect 330222 655380 330306 655616
rect 330542 655380 330574 655616
rect 329954 655296 330574 655380
rect 329954 655060 329986 655296
rect 330222 655060 330306 655296
rect 330542 655060 330574 655296
rect 329954 619616 330574 655060
rect 329954 619380 329986 619616
rect 330222 619380 330306 619616
rect 330542 619380 330574 619616
rect 329954 619296 330574 619380
rect 329954 619060 329986 619296
rect 330222 619060 330306 619296
rect 330542 619060 330574 619296
rect 329954 583616 330574 619060
rect 329954 583380 329986 583616
rect 330222 583380 330306 583616
rect 330542 583380 330574 583616
rect 329954 583296 330574 583380
rect 329954 583060 329986 583296
rect 330222 583060 330306 583296
rect 330542 583060 330574 583296
rect 329954 547616 330574 583060
rect 329954 547380 329986 547616
rect 330222 547380 330306 547616
rect 330542 547380 330574 547616
rect 329954 547296 330574 547380
rect 329954 547060 329986 547296
rect 330222 547060 330306 547296
rect 330542 547060 330574 547296
rect 329954 511616 330574 547060
rect 329954 511380 329986 511616
rect 330222 511380 330306 511616
rect 330542 511380 330574 511616
rect 329954 511296 330574 511380
rect 329954 511060 329986 511296
rect 330222 511060 330306 511296
rect 330542 511060 330574 511296
rect 329954 475616 330574 511060
rect 329954 475380 329986 475616
rect 330222 475380 330306 475616
rect 330542 475380 330574 475616
rect 329954 475296 330574 475380
rect 329954 475060 329986 475296
rect 330222 475060 330306 475296
rect 330542 475060 330574 475296
rect 329954 439616 330574 475060
rect 329954 439380 329986 439616
rect 330222 439380 330306 439616
rect 330542 439380 330574 439616
rect 329954 439296 330574 439380
rect 329954 439060 329986 439296
rect 330222 439060 330306 439296
rect 330542 439060 330574 439296
rect 329954 403616 330574 439060
rect 329954 403380 329986 403616
rect 330222 403380 330306 403616
rect 330542 403380 330574 403616
rect 329954 403296 330574 403380
rect 329954 403060 329986 403296
rect 330222 403060 330306 403296
rect 330542 403060 330574 403296
rect 329954 367616 330574 403060
rect 329954 367380 329986 367616
rect 330222 367380 330306 367616
rect 330542 367380 330574 367616
rect 329954 367296 330574 367380
rect 329954 367060 329986 367296
rect 330222 367060 330306 367296
rect 330542 367060 330574 367296
rect 329954 331616 330574 367060
rect 329954 331380 329986 331616
rect 330222 331380 330306 331616
rect 330542 331380 330574 331616
rect 329954 331296 330574 331380
rect 329954 331060 329986 331296
rect 330222 331060 330306 331296
rect 330542 331060 330574 331296
rect 329954 295616 330574 331060
rect 329954 295380 329986 295616
rect 330222 295380 330306 295616
rect 330542 295380 330574 295616
rect 329954 295296 330574 295380
rect 329954 295060 329986 295296
rect 330222 295060 330306 295296
rect 330542 295060 330574 295296
rect 329954 259616 330574 295060
rect 329954 259380 329986 259616
rect 330222 259380 330306 259616
rect 330542 259380 330574 259616
rect 329954 259296 330574 259380
rect 329954 259060 329986 259296
rect 330222 259060 330306 259296
rect 330542 259060 330574 259296
rect 329954 223616 330574 259060
rect 329954 223380 329986 223616
rect 330222 223380 330306 223616
rect 330542 223380 330574 223616
rect 329954 223296 330574 223380
rect 329954 223060 329986 223296
rect 330222 223060 330306 223296
rect 330542 223060 330574 223296
rect 329954 187616 330574 223060
rect 329954 187380 329986 187616
rect 330222 187380 330306 187616
rect 330542 187380 330574 187616
rect 329954 187296 330574 187380
rect 329954 187060 329986 187296
rect 330222 187060 330306 187296
rect 330542 187060 330574 187296
rect 329954 151616 330574 187060
rect 329954 151380 329986 151616
rect 330222 151380 330306 151616
rect 330542 151380 330574 151616
rect 329954 151296 330574 151380
rect 329954 151060 329986 151296
rect 330222 151060 330306 151296
rect 330542 151060 330574 151296
rect 329954 115616 330574 151060
rect 329954 115380 329986 115616
rect 330222 115380 330306 115616
rect 330542 115380 330574 115616
rect 329954 115296 330574 115380
rect 329954 115060 329986 115296
rect 330222 115060 330306 115296
rect 330542 115060 330574 115296
rect 329954 79616 330574 115060
rect 329954 79380 329986 79616
rect 330222 79380 330306 79616
rect 330542 79380 330574 79616
rect 329954 79296 330574 79380
rect 329954 79060 329986 79296
rect 330222 79060 330306 79296
rect 330542 79060 330574 79296
rect 329954 43616 330574 79060
rect 329954 43380 329986 43616
rect 330222 43380 330306 43616
rect 330542 43380 330574 43616
rect 329954 43296 330574 43380
rect 329954 43060 329986 43296
rect 330222 43060 330306 43296
rect 330542 43060 330574 43296
rect 329954 7616 330574 43060
rect 329954 7380 329986 7616
rect 330222 7380 330306 7616
rect 330542 7380 330574 7616
rect 329954 7296 330574 7380
rect 329954 7060 329986 7296
rect 330222 7060 330306 7296
rect 330542 7060 330574 7296
rect 329954 -4184 330574 7060
rect 329954 -4420 329986 -4184
rect 330222 -4420 330306 -4184
rect 330542 -4420 330574 -4184
rect 329954 -4504 330574 -4420
rect 329954 -4740 329986 -4504
rect 330222 -4740 330306 -4504
rect 330542 -4740 330574 -4504
rect 329954 -7652 330574 -4740
rect 331194 709640 331814 711592
rect 331194 709404 331226 709640
rect 331462 709404 331546 709640
rect 331782 709404 331814 709640
rect 331194 709320 331814 709404
rect 331194 709084 331226 709320
rect 331462 709084 331546 709320
rect 331782 709084 331814 709320
rect 331194 692856 331814 709084
rect 331194 692620 331226 692856
rect 331462 692620 331546 692856
rect 331782 692620 331814 692856
rect 331194 692536 331814 692620
rect 331194 692300 331226 692536
rect 331462 692300 331546 692536
rect 331782 692300 331814 692536
rect 331194 656856 331814 692300
rect 331194 656620 331226 656856
rect 331462 656620 331546 656856
rect 331782 656620 331814 656856
rect 331194 656536 331814 656620
rect 331194 656300 331226 656536
rect 331462 656300 331546 656536
rect 331782 656300 331814 656536
rect 331194 620856 331814 656300
rect 331194 620620 331226 620856
rect 331462 620620 331546 620856
rect 331782 620620 331814 620856
rect 331194 620536 331814 620620
rect 331194 620300 331226 620536
rect 331462 620300 331546 620536
rect 331782 620300 331814 620536
rect 331194 584856 331814 620300
rect 331194 584620 331226 584856
rect 331462 584620 331546 584856
rect 331782 584620 331814 584856
rect 331194 584536 331814 584620
rect 331194 584300 331226 584536
rect 331462 584300 331546 584536
rect 331782 584300 331814 584536
rect 331194 548856 331814 584300
rect 331194 548620 331226 548856
rect 331462 548620 331546 548856
rect 331782 548620 331814 548856
rect 331194 548536 331814 548620
rect 331194 548300 331226 548536
rect 331462 548300 331546 548536
rect 331782 548300 331814 548536
rect 331194 512856 331814 548300
rect 331194 512620 331226 512856
rect 331462 512620 331546 512856
rect 331782 512620 331814 512856
rect 331194 512536 331814 512620
rect 331194 512300 331226 512536
rect 331462 512300 331546 512536
rect 331782 512300 331814 512536
rect 331194 476856 331814 512300
rect 331194 476620 331226 476856
rect 331462 476620 331546 476856
rect 331782 476620 331814 476856
rect 331194 476536 331814 476620
rect 331194 476300 331226 476536
rect 331462 476300 331546 476536
rect 331782 476300 331814 476536
rect 331194 440856 331814 476300
rect 331194 440620 331226 440856
rect 331462 440620 331546 440856
rect 331782 440620 331814 440856
rect 331194 440536 331814 440620
rect 331194 440300 331226 440536
rect 331462 440300 331546 440536
rect 331782 440300 331814 440536
rect 331194 404856 331814 440300
rect 331194 404620 331226 404856
rect 331462 404620 331546 404856
rect 331782 404620 331814 404856
rect 331194 404536 331814 404620
rect 331194 404300 331226 404536
rect 331462 404300 331546 404536
rect 331782 404300 331814 404536
rect 331194 368856 331814 404300
rect 331194 368620 331226 368856
rect 331462 368620 331546 368856
rect 331782 368620 331814 368856
rect 331194 368536 331814 368620
rect 331194 368300 331226 368536
rect 331462 368300 331546 368536
rect 331782 368300 331814 368536
rect 331194 332856 331814 368300
rect 331194 332620 331226 332856
rect 331462 332620 331546 332856
rect 331782 332620 331814 332856
rect 331194 332536 331814 332620
rect 331194 332300 331226 332536
rect 331462 332300 331546 332536
rect 331782 332300 331814 332536
rect 331194 296856 331814 332300
rect 331194 296620 331226 296856
rect 331462 296620 331546 296856
rect 331782 296620 331814 296856
rect 331194 296536 331814 296620
rect 331194 296300 331226 296536
rect 331462 296300 331546 296536
rect 331782 296300 331814 296536
rect 331194 260856 331814 296300
rect 331194 260620 331226 260856
rect 331462 260620 331546 260856
rect 331782 260620 331814 260856
rect 331194 260536 331814 260620
rect 331194 260300 331226 260536
rect 331462 260300 331546 260536
rect 331782 260300 331814 260536
rect 331194 224856 331814 260300
rect 331194 224620 331226 224856
rect 331462 224620 331546 224856
rect 331782 224620 331814 224856
rect 331194 224536 331814 224620
rect 331194 224300 331226 224536
rect 331462 224300 331546 224536
rect 331782 224300 331814 224536
rect 331194 188856 331814 224300
rect 331194 188620 331226 188856
rect 331462 188620 331546 188856
rect 331782 188620 331814 188856
rect 331194 188536 331814 188620
rect 331194 188300 331226 188536
rect 331462 188300 331546 188536
rect 331782 188300 331814 188536
rect 331194 152856 331814 188300
rect 331194 152620 331226 152856
rect 331462 152620 331546 152856
rect 331782 152620 331814 152856
rect 331194 152536 331814 152620
rect 331194 152300 331226 152536
rect 331462 152300 331546 152536
rect 331782 152300 331814 152536
rect 331194 116856 331814 152300
rect 331194 116620 331226 116856
rect 331462 116620 331546 116856
rect 331782 116620 331814 116856
rect 331194 116536 331814 116620
rect 331194 116300 331226 116536
rect 331462 116300 331546 116536
rect 331782 116300 331814 116536
rect 331194 80856 331814 116300
rect 331194 80620 331226 80856
rect 331462 80620 331546 80856
rect 331782 80620 331814 80856
rect 331194 80536 331814 80620
rect 331194 80300 331226 80536
rect 331462 80300 331546 80536
rect 331782 80300 331814 80536
rect 331194 44856 331814 80300
rect 331194 44620 331226 44856
rect 331462 44620 331546 44856
rect 331782 44620 331814 44856
rect 331194 44536 331814 44620
rect 331194 44300 331226 44536
rect 331462 44300 331546 44536
rect 331782 44300 331814 44536
rect 331194 8856 331814 44300
rect 331194 8620 331226 8856
rect 331462 8620 331546 8856
rect 331782 8620 331814 8856
rect 331194 8536 331814 8620
rect 331194 8300 331226 8536
rect 331462 8300 331546 8536
rect 331782 8300 331814 8536
rect 331194 -5144 331814 8300
rect 331194 -5380 331226 -5144
rect 331462 -5380 331546 -5144
rect 331782 -5380 331814 -5144
rect 331194 -5464 331814 -5380
rect 331194 -5700 331226 -5464
rect 331462 -5700 331546 -5464
rect 331782 -5700 331814 -5464
rect 331194 -7652 331814 -5700
rect 332434 710600 333054 711592
rect 332434 710364 332466 710600
rect 332702 710364 332786 710600
rect 333022 710364 333054 710600
rect 332434 710280 333054 710364
rect 332434 710044 332466 710280
rect 332702 710044 332786 710280
rect 333022 710044 333054 710280
rect 332434 694096 333054 710044
rect 332434 693860 332466 694096
rect 332702 693860 332786 694096
rect 333022 693860 333054 694096
rect 332434 693776 333054 693860
rect 332434 693540 332466 693776
rect 332702 693540 332786 693776
rect 333022 693540 333054 693776
rect 332434 658096 333054 693540
rect 332434 657860 332466 658096
rect 332702 657860 332786 658096
rect 333022 657860 333054 658096
rect 332434 657776 333054 657860
rect 332434 657540 332466 657776
rect 332702 657540 332786 657776
rect 333022 657540 333054 657776
rect 332434 622096 333054 657540
rect 332434 621860 332466 622096
rect 332702 621860 332786 622096
rect 333022 621860 333054 622096
rect 332434 621776 333054 621860
rect 332434 621540 332466 621776
rect 332702 621540 332786 621776
rect 333022 621540 333054 621776
rect 332434 586096 333054 621540
rect 332434 585860 332466 586096
rect 332702 585860 332786 586096
rect 333022 585860 333054 586096
rect 332434 585776 333054 585860
rect 332434 585540 332466 585776
rect 332702 585540 332786 585776
rect 333022 585540 333054 585776
rect 332434 550096 333054 585540
rect 332434 549860 332466 550096
rect 332702 549860 332786 550096
rect 333022 549860 333054 550096
rect 332434 549776 333054 549860
rect 332434 549540 332466 549776
rect 332702 549540 332786 549776
rect 333022 549540 333054 549776
rect 332434 514096 333054 549540
rect 332434 513860 332466 514096
rect 332702 513860 332786 514096
rect 333022 513860 333054 514096
rect 332434 513776 333054 513860
rect 332434 513540 332466 513776
rect 332702 513540 332786 513776
rect 333022 513540 333054 513776
rect 332434 478096 333054 513540
rect 332434 477860 332466 478096
rect 332702 477860 332786 478096
rect 333022 477860 333054 478096
rect 332434 477776 333054 477860
rect 332434 477540 332466 477776
rect 332702 477540 332786 477776
rect 333022 477540 333054 477776
rect 332434 442096 333054 477540
rect 332434 441860 332466 442096
rect 332702 441860 332786 442096
rect 333022 441860 333054 442096
rect 332434 441776 333054 441860
rect 332434 441540 332466 441776
rect 332702 441540 332786 441776
rect 333022 441540 333054 441776
rect 332434 406096 333054 441540
rect 332434 405860 332466 406096
rect 332702 405860 332786 406096
rect 333022 405860 333054 406096
rect 332434 405776 333054 405860
rect 332434 405540 332466 405776
rect 332702 405540 332786 405776
rect 333022 405540 333054 405776
rect 332434 370096 333054 405540
rect 332434 369860 332466 370096
rect 332702 369860 332786 370096
rect 333022 369860 333054 370096
rect 332434 369776 333054 369860
rect 332434 369540 332466 369776
rect 332702 369540 332786 369776
rect 333022 369540 333054 369776
rect 332434 334096 333054 369540
rect 332434 333860 332466 334096
rect 332702 333860 332786 334096
rect 333022 333860 333054 334096
rect 332434 333776 333054 333860
rect 332434 333540 332466 333776
rect 332702 333540 332786 333776
rect 333022 333540 333054 333776
rect 332434 298096 333054 333540
rect 332434 297860 332466 298096
rect 332702 297860 332786 298096
rect 333022 297860 333054 298096
rect 332434 297776 333054 297860
rect 332434 297540 332466 297776
rect 332702 297540 332786 297776
rect 333022 297540 333054 297776
rect 332434 262096 333054 297540
rect 332434 261860 332466 262096
rect 332702 261860 332786 262096
rect 333022 261860 333054 262096
rect 332434 261776 333054 261860
rect 332434 261540 332466 261776
rect 332702 261540 332786 261776
rect 333022 261540 333054 261776
rect 332434 226096 333054 261540
rect 332434 225860 332466 226096
rect 332702 225860 332786 226096
rect 333022 225860 333054 226096
rect 332434 225776 333054 225860
rect 332434 225540 332466 225776
rect 332702 225540 332786 225776
rect 333022 225540 333054 225776
rect 332434 190096 333054 225540
rect 332434 189860 332466 190096
rect 332702 189860 332786 190096
rect 333022 189860 333054 190096
rect 332434 189776 333054 189860
rect 332434 189540 332466 189776
rect 332702 189540 332786 189776
rect 333022 189540 333054 189776
rect 332434 154096 333054 189540
rect 332434 153860 332466 154096
rect 332702 153860 332786 154096
rect 333022 153860 333054 154096
rect 332434 153776 333054 153860
rect 332434 153540 332466 153776
rect 332702 153540 332786 153776
rect 333022 153540 333054 153776
rect 332434 118096 333054 153540
rect 332434 117860 332466 118096
rect 332702 117860 332786 118096
rect 333022 117860 333054 118096
rect 332434 117776 333054 117860
rect 332434 117540 332466 117776
rect 332702 117540 332786 117776
rect 333022 117540 333054 117776
rect 332434 82096 333054 117540
rect 332434 81860 332466 82096
rect 332702 81860 332786 82096
rect 333022 81860 333054 82096
rect 332434 81776 333054 81860
rect 332434 81540 332466 81776
rect 332702 81540 332786 81776
rect 333022 81540 333054 81776
rect 332434 46096 333054 81540
rect 332434 45860 332466 46096
rect 332702 45860 332786 46096
rect 333022 45860 333054 46096
rect 332434 45776 333054 45860
rect 332434 45540 332466 45776
rect 332702 45540 332786 45776
rect 333022 45540 333054 45776
rect 332434 10096 333054 45540
rect 332434 9860 332466 10096
rect 332702 9860 332786 10096
rect 333022 9860 333054 10096
rect 332434 9776 333054 9860
rect 332434 9540 332466 9776
rect 332702 9540 332786 9776
rect 333022 9540 333054 9776
rect 332434 -6104 333054 9540
rect 332434 -6340 332466 -6104
rect 332702 -6340 332786 -6104
rect 333022 -6340 333054 -6104
rect 332434 -6424 333054 -6340
rect 332434 -6660 332466 -6424
rect 332702 -6660 332786 -6424
rect 333022 -6660 333054 -6424
rect 332434 -7652 333054 -6660
rect 333674 711560 334294 711592
rect 333674 711324 333706 711560
rect 333942 711324 334026 711560
rect 334262 711324 334294 711560
rect 333674 711240 334294 711324
rect 333674 711004 333706 711240
rect 333942 711004 334026 711240
rect 334262 711004 334294 711240
rect 333674 695336 334294 711004
rect 333674 695100 333706 695336
rect 333942 695100 334026 695336
rect 334262 695100 334294 695336
rect 333674 695016 334294 695100
rect 333674 694780 333706 695016
rect 333942 694780 334026 695016
rect 334262 694780 334294 695016
rect 333674 659336 334294 694780
rect 333674 659100 333706 659336
rect 333942 659100 334026 659336
rect 334262 659100 334294 659336
rect 333674 659016 334294 659100
rect 333674 658780 333706 659016
rect 333942 658780 334026 659016
rect 334262 658780 334294 659016
rect 333674 623336 334294 658780
rect 333674 623100 333706 623336
rect 333942 623100 334026 623336
rect 334262 623100 334294 623336
rect 333674 623016 334294 623100
rect 333674 622780 333706 623016
rect 333942 622780 334026 623016
rect 334262 622780 334294 623016
rect 333674 587336 334294 622780
rect 333674 587100 333706 587336
rect 333942 587100 334026 587336
rect 334262 587100 334294 587336
rect 333674 587016 334294 587100
rect 333674 586780 333706 587016
rect 333942 586780 334026 587016
rect 334262 586780 334294 587016
rect 333674 551336 334294 586780
rect 333674 551100 333706 551336
rect 333942 551100 334026 551336
rect 334262 551100 334294 551336
rect 333674 551016 334294 551100
rect 333674 550780 333706 551016
rect 333942 550780 334026 551016
rect 334262 550780 334294 551016
rect 333674 515336 334294 550780
rect 333674 515100 333706 515336
rect 333942 515100 334026 515336
rect 334262 515100 334294 515336
rect 333674 515016 334294 515100
rect 333674 514780 333706 515016
rect 333942 514780 334026 515016
rect 334262 514780 334294 515016
rect 333674 479336 334294 514780
rect 333674 479100 333706 479336
rect 333942 479100 334026 479336
rect 334262 479100 334294 479336
rect 333674 479016 334294 479100
rect 333674 478780 333706 479016
rect 333942 478780 334026 479016
rect 334262 478780 334294 479016
rect 333674 443336 334294 478780
rect 333674 443100 333706 443336
rect 333942 443100 334026 443336
rect 334262 443100 334294 443336
rect 333674 443016 334294 443100
rect 333674 442780 333706 443016
rect 333942 442780 334026 443016
rect 334262 442780 334294 443016
rect 333674 407336 334294 442780
rect 333674 407100 333706 407336
rect 333942 407100 334026 407336
rect 334262 407100 334294 407336
rect 333674 407016 334294 407100
rect 333674 406780 333706 407016
rect 333942 406780 334026 407016
rect 334262 406780 334294 407016
rect 333674 371336 334294 406780
rect 333674 371100 333706 371336
rect 333942 371100 334026 371336
rect 334262 371100 334294 371336
rect 333674 371016 334294 371100
rect 333674 370780 333706 371016
rect 333942 370780 334026 371016
rect 334262 370780 334294 371016
rect 333674 335336 334294 370780
rect 333674 335100 333706 335336
rect 333942 335100 334026 335336
rect 334262 335100 334294 335336
rect 333674 335016 334294 335100
rect 333674 334780 333706 335016
rect 333942 334780 334026 335016
rect 334262 334780 334294 335016
rect 333674 299336 334294 334780
rect 333674 299100 333706 299336
rect 333942 299100 334026 299336
rect 334262 299100 334294 299336
rect 333674 299016 334294 299100
rect 333674 298780 333706 299016
rect 333942 298780 334026 299016
rect 334262 298780 334294 299016
rect 333674 263336 334294 298780
rect 333674 263100 333706 263336
rect 333942 263100 334026 263336
rect 334262 263100 334294 263336
rect 333674 263016 334294 263100
rect 333674 262780 333706 263016
rect 333942 262780 334026 263016
rect 334262 262780 334294 263016
rect 333674 227336 334294 262780
rect 333674 227100 333706 227336
rect 333942 227100 334026 227336
rect 334262 227100 334294 227336
rect 333674 227016 334294 227100
rect 333674 226780 333706 227016
rect 333942 226780 334026 227016
rect 334262 226780 334294 227016
rect 333674 191336 334294 226780
rect 333674 191100 333706 191336
rect 333942 191100 334026 191336
rect 334262 191100 334294 191336
rect 333674 191016 334294 191100
rect 333674 190780 333706 191016
rect 333942 190780 334026 191016
rect 334262 190780 334294 191016
rect 333674 155336 334294 190780
rect 333674 155100 333706 155336
rect 333942 155100 334026 155336
rect 334262 155100 334294 155336
rect 333674 155016 334294 155100
rect 333674 154780 333706 155016
rect 333942 154780 334026 155016
rect 334262 154780 334294 155016
rect 333674 119336 334294 154780
rect 333674 119100 333706 119336
rect 333942 119100 334026 119336
rect 334262 119100 334294 119336
rect 333674 119016 334294 119100
rect 333674 118780 333706 119016
rect 333942 118780 334026 119016
rect 334262 118780 334294 119016
rect 333674 83336 334294 118780
rect 333674 83100 333706 83336
rect 333942 83100 334026 83336
rect 334262 83100 334294 83336
rect 333674 83016 334294 83100
rect 333674 82780 333706 83016
rect 333942 82780 334026 83016
rect 334262 82780 334294 83016
rect 333674 47336 334294 82780
rect 333674 47100 333706 47336
rect 333942 47100 334026 47336
rect 334262 47100 334294 47336
rect 333674 47016 334294 47100
rect 333674 46780 333706 47016
rect 333942 46780 334026 47016
rect 334262 46780 334294 47016
rect 333674 11336 334294 46780
rect 333674 11100 333706 11336
rect 333942 11100 334026 11336
rect 334262 11100 334294 11336
rect 333674 11016 334294 11100
rect 333674 10780 333706 11016
rect 333942 10780 334026 11016
rect 334262 10780 334294 11016
rect 333674 -7064 334294 10780
rect 333674 -7300 333706 -7064
rect 333942 -7300 334026 -7064
rect 334262 -7300 334294 -7064
rect 333674 -7384 334294 -7300
rect 333674 -7620 333706 -7384
rect 333942 -7620 334026 -7384
rect 334262 -7620 334294 -7384
rect 333674 -7652 334294 -7620
rect 360994 704840 361614 711592
rect 360994 704604 361026 704840
rect 361262 704604 361346 704840
rect 361582 704604 361614 704840
rect 360994 704520 361614 704604
rect 360994 704284 361026 704520
rect 361262 704284 361346 704520
rect 361582 704284 361614 704520
rect 360994 702139 361614 704284
rect 360994 702075 361032 702139
rect 361096 702075 361112 702139
rect 361176 702075 361192 702139
rect 361256 702075 361272 702139
rect 361336 702075 361352 702139
rect 361416 702075 361432 702139
rect 361496 702075 361512 702139
rect 361576 702075 361614 702139
rect 360994 702059 361614 702075
rect 360994 701995 361032 702059
rect 361096 701995 361112 702059
rect 361176 701995 361192 702059
rect 361256 701995 361272 702059
rect 361336 701995 361352 702059
rect 361416 701995 361432 702059
rect 361496 701995 361512 702059
rect 361576 701995 361614 702059
rect 360994 701979 361614 701995
rect 360994 701915 361032 701979
rect 361096 701915 361112 701979
rect 361176 701915 361192 701979
rect 361256 701915 361272 701979
rect 361336 701915 361352 701979
rect 361416 701915 361432 701979
rect 361496 701915 361512 701979
rect 361576 701915 361614 701979
rect 360994 701899 361614 701915
rect 360994 701835 361032 701899
rect 361096 701835 361112 701899
rect 361176 701835 361192 701899
rect 361256 701835 361272 701899
rect 361336 701835 361352 701899
rect 361416 701835 361432 701899
rect 361496 701835 361512 701899
rect 361576 701835 361614 701899
rect 360994 686656 361614 701835
rect 360994 686420 361026 686656
rect 361262 686420 361346 686656
rect 361582 686420 361614 686656
rect 360994 686336 361614 686420
rect 360994 686100 361026 686336
rect 361262 686100 361346 686336
rect 361582 686100 361614 686336
rect 360994 650656 361614 686100
rect 360994 650420 361026 650656
rect 361262 650420 361346 650656
rect 361582 650420 361614 650656
rect 360994 650336 361614 650420
rect 360994 650100 361026 650336
rect 361262 650100 361346 650336
rect 361582 650100 361614 650336
rect 360994 614656 361614 650100
rect 360994 614420 361026 614656
rect 361262 614420 361346 614656
rect 361582 614420 361614 614656
rect 360994 614336 361614 614420
rect 360994 614100 361026 614336
rect 361262 614100 361346 614336
rect 361582 614100 361614 614336
rect 360994 578656 361614 614100
rect 360994 578420 361026 578656
rect 361262 578420 361346 578656
rect 361582 578420 361614 578656
rect 360994 578336 361614 578420
rect 360994 578100 361026 578336
rect 361262 578100 361346 578336
rect 361582 578100 361614 578336
rect 360994 542656 361614 578100
rect 360994 542420 361026 542656
rect 361262 542420 361346 542656
rect 361582 542420 361614 542656
rect 360994 542336 361614 542420
rect 360994 542100 361026 542336
rect 361262 542100 361346 542336
rect 361582 542100 361614 542336
rect 360994 506656 361614 542100
rect 360994 506420 361026 506656
rect 361262 506420 361346 506656
rect 361582 506420 361614 506656
rect 360994 506336 361614 506420
rect 360994 506100 361026 506336
rect 361262 506100 361346 506336
rect 361582 506100 361614 506336
rect 360994 470656 361614 506100
rect 360994 470420 361026 470656
rect 361262 470420 361346 470656
rect 361582 470420 361614 470656
rect 360994 470336 361614 470420
rect 360994 470100 361026 470336
rect 361262 470100 361346 470336
rect 361582 470100 361614 470336
rect 360994 434656 361614 470100
rect 360994 434420 361026 434656
rect 361262 434420 361346 434656
rect 361582 434420 361614 434656
rect 360994 434336 361614 434420
rect 360994 434100 361026 434336
rect 361262 434100 361346 434336
rect 361582 434100 361614 434336
rect 360994 398656 361614 434100
rect 360994 398420 361026 398656
rect 361262 398420 361346 398656
rect 361582 398420 361614 398656
rect 360994 398336 361614 398420
rect 360994 398100 361026 398336
rect 361262 398100 361346 398336
rect 361582 398100 361614 398336
rect 360994 362656 361614 398100
rect 360994 362420 361026 362656
rect 361262 362420 361346 362656
rect 361582 362420 361614 362656
rect 360994 362336 361614 362420
rect 360994 362100 361026 362336
rect 361262 362100 361346 362336
rect 361582 362100 361614 362336
rect 360994 326656 361614 362100
rect 360994 326420 361026 326656
rect 361262 326420 361346 326656
rect 361582 326420 361614 326656
rect 360994 326336 361614 326420
rect 360994 326100 361026 326336
rect 361262 326100 361346 326336
rect 361582 326100 361614 326336
rect 360994 290656 361614 326100
rect 360994 290420 361026 290656
rect 361262 290420 361346 290656
rect 361582 290420 361614 290656
rect 360994 290336 361614 290420
rect 360994 290100 361026 290336
rect 361262 290100 361346 290336
rect 361582 290100 361614 290336
rect 360994 254656 361614 290100
rect 360994 254420 361026 254656
rect 361262 254420 361346 254656
rect 361582 254420 361614 254656
rect 360994 254336 361614 254420
rect 360994 254100 361026 254336
rect 361262 254100 361346 254336
rect 361582 254100 361614 254336
rect 360994 218656 361614 254100
rect 360994 218420 361026 218656
rect 361262 218420 361346 218656
rect 361582 218420 361614 218656
rect 360994 218336 361614 218420
rect 360994 218100 361026 218336
rect 361262 218100 361346 218336
rect 361582 218100 361614 218336
rect 360994 182656 361614 218100
rect 360994 182420 361026 182656
rect 361262 182420 361346 182656
rect 361582 182420 361614 182656
rect 360994 182336 361614 182420
rect 360994 182100 361026 182336
rect 361262 182100 361346 182336
rect 361582 182100 361614 182336
rect 360994 146656 361614 182100
rect 360994 146420 361026 146656
rect 361262 146420 361346 146656
rect 361582 146420 361614 146656
rect 360994 146336 361614 146420
rect 360994 146100 361026 146336
rect 361262 146100 361346 146336
rect 361582 146100 361614 146336
rect 360994 110656 361614 146100
rect 360994 110420 361026 110656
rect 361262 110420 361346 110656
rect 361582 110420 361614 110656
rect 360994 110336 361614 110420
rect 360994 110100 361026 110336
rect 361262 110100 361346 110336
rect 361582 110100 361614 110336
rect 360994 74656 361614 110100
rect 360994 74420 361026 74656
rect 361262 74420 361346 74656
rect 361582 74420 361614 74656
rect 360994 74336 361614 74420
rect 360994 74100 361026 74336
rect 361262 74100 361346 74336
rect 361582 74100 361614 74336
rect 360994 38656 361614 74100
rect 360994 38420 361026 38656
rect 361262 38420 361346 38656
rect 361582 38420 361614 38656
rect 360994 38336 361614 38420
rect 360994 38100 361026 38336
rect 361262 38100 361346 38336
rect 361582 38100 361614 38336
rect 360994 2656 361614 38100
rect 360994 2420 361026 2656
rect 361262 2420 361346 2656
rect 361582 2420 361614 2656
rect 360994 2336 361614 2420
rect 360994 2100 361026 2336
rect 361262 2100 361346 2336
rect 361582 2100 361614 2336
rect 360994 -344 361614 2100
rect 360994 -580 361026 -344
rect 361262 -580 361346 -344
rect 361582 -580 361614 -344
rect 360994 -664 361614 -580
rect 360994 -900 361026 -664
rect 361262 -900 361346 -664
rect 361582 -900 361614 -664
rect 360994 -7652 361614 -900
rect 362234 705800 362854 711592
rect 362234 705564 362266 705800
rect 362502 705564 362586 705800
rect 362822 705564 362854 705800
rect 362234 705480 362854 705564
rect 362234 705244 362266 705480
rect 362502 705244 362586 705480
rect 362822 705244 362854 705480
rect 362234 702907 362854 705244
rect 362234 702843 362272 702907
rect 362336 702843 362352 702907
rect 362416 702843 362432 702907
rect 362496 702843 362512 702907
rect 362576 702843 362592 702907
rect 362656 702843 362672 702907
rect 362736 702843 362752 702907
rect 362816 702843 362854 702907
rect 362234 702827 362854 702843
rect 362234 702763 362272 702827
rect 362336 702763 362352 702827
rect 362416 702763 362432 702827
rect 362496 702763 362512 702827
rect 362576 702763 362592 702827
rect 362656 702763 362672 702827
rect 362736 702763 362752 702827
rect 362816 702763 362854 702827
rect 362234 702747 362854 702763
rect 362234 702683 362272 702747
rect 362336 702683 362352 702747
rect 362416 702683 362432 702747
rect 362496 702683 362512 702747
rect 362576 702683 362592 702747
rect 362656 702683 362672 702747
rect 362736 702683 362752 702747
rect 362816 702683 362854 702747
rect 362234 702667 362854 702683
rect 362234 702603 362272 702667
rect 362336 702603 362352 702667
rect 362416 702603 362432 702667
rect 362496 702603 362512 702667
rect 362576 702603 362592 702667
rect 362656 702603 362672 702667
rect 362736 702603 362752 702667
rect 362816 702603 362854 702667
rect 362234 687896 362854 702603
rect 362234 687660 362266 687896
rect 362502 687660 362586 687896
rect 362822 687660 362854 687896
rect 362234 687576 362854 687660
rect 362234 687340 362266 687576
rect 362502 687340 362586 687576
rect 362822 687340 362854 687576
rect 362234 651896 362854 687340
rect 362234 651660 362266 651896
rect 362502 651660 362586 651896
rect 362822 651660 362854 651896
rect 362234 651576 362854 651660
rect 362234 651340 362266 651576
rect 362502 651340 362586 651576
rect 362822 651340 362854 651576
rect 362234 615896 362854 651340
rect 362234 615660 362266 615896
rect 362502 615660 362586 615896
rect 362822 615660 362854 615896
rect 362234 615576 362854 615660
rect 362234 615340 362266 615576
rect 362502 615340 362586 615576
rect 362822 615340 362854 615576
rect 362234 579896 362854 615340
rect 362234 579660 362266 579896
rect 362502 579660 362586 579896
rect 362822 579660 362854 579896
rect 362234 579576 362854 579660
rect 362234 579340 362266 579576
rect 362502 579340 362586 579576
rect 362822 579340 362854 579576
rect 362234 543896 362854 579340
rect 362234 543660 362266 543896
rect 362502 543660 362586 543896
rect 362822 543660 362854 543896
rect 362234 543576 362854 543660
rect 362234 543340 362266 543576
rect 362502 543340 362586 543576
rect 362822 543340 362854 543576
rect 362234 507896 362854 543340
rect 362234 507660 362266 507896
rect 362502 507660 362586 507896
rect 362822 507660 362854 507896
rect 362234 507576 362854 507660
rect 362234 507340 362266 507576
rect 362502 507340 362586 507576
rect 362822 507340 362854 507576
rect 362234 471896 362854 507340
rect 362234 471660 362266 471896
rect 362502 471660 362586 471896
rect 362822 471660 362854 471896
rect 362234 471576 362854 471660
rect 362234 471340 362266 471576
rect 362502 471340 362586 471576
rect 362822 471340 362854 471576
rect 362234 435896 362854 471340
rect 362234 435660 362266 435896
rect 362502 435660 362586 435896
rect 362822 435660 362854 435896
rect 362234 435576 362854 435660
rect 362234 435340 362266 435576
rect 362502 435340 362586 435576
rect 362822 435340 362854 435576
rect 362234 399896 362854 435340
rect 362234 399660 362266 399896
rect 362502 399660 362586 399896
rect 362822 399660 362854 399896
rect 362234 399576 362854 399660
rect 362234 399340 362266 399576
rect 362502 399340 362586 399576
rect 362822 399340 362854 399576
rect 362234 363896 362854 399340
rect 362234 363660 362266 363896
rect 362502 363660 362586 363896
rect 362822 363660 362854 363896
rect 362234 363576 362854 363660
rect 362234 363340 362266 363576
rect 362502 363340 362586 363576
rect 362822 363340 362854 363576
rect 362234 327896 362854 363340
rect 362234 327660 362266 327896
rect 362502 327660 362586 327896
rect 362822 327660 362854 327896
rect 362234 327576 362854 327660
rect 362234 327340 362266 327576
rect 362502 327340 362586 327576
rect 362822 327340 362854 327576
rect 362234 291896 362854 327340
rect 362234 291660 362266 291896
rect 362502 291660 362586 291896
rect 362822 291660 362854 291896
rect 362234 291576 362854 291660
rect 362234 291340 362266 291576
rect 362502 291340 362586 291576
rect 362822 291340 362854 291576
rect 362234 255896 362854 291340
rect 362234 255660 362266 255896
rect 362502 255660 362586 255896
rect 362822 255660 362854 255896
rect 362234 255576 362854 255660
rect 362234 255340 362266 255576
rect 362502 255340 362586 255576
rect 362822 255340 362854 255576
rect 362234 219896 362854 255340
rect 362234 219660 362266 219896
rect 362502 219660 362586 219896
rect 362822 219660 362854 219896
rect 362234 219576 362854 219660
rect 362234 219340 362266 219576
rect 362502 219340 362586 219576
rect 362822 219340 362854 219576
rect 362234 183896 362854 219340
rect 362234 183660 362266 183896
rect 362502 183660 362586 183896
rect 362822 183660 362854 183896
rect 362234 183576 362854 183660
rect 362234 183340 362266 183576
rect 362502 183340 362586 183576
rect 362822 183340 362854 183576
rect 362234 147896 362854 183340
rect 362234 147660 362266 147896
rect 362502 147660 362586 147896
rect 362822 147660 362854 147896
rect 362234 147576 362854 147660
rect 362234 147340 362266 147576
rect 362502 147340 362586 147576
rect 362822 147340 362854 147576
rect 362234 111896 362854 147340
rect 362234 111660 362266 111896
rect 362502 111660 362586 111896
rect 362822 111660 362854 111896
rect 362234 111576 362854 111660
rect 362234 111340 362266 111576
rect 362502 111340 362586 111576
rect 362822 111340 362854 111576
rect 362234 75896 362854 111340
rect 362234 75660 362266 75896
rect 362502 75660 362586 75896
rect 362822 75660 362854 75896
rect 362234 75576 362854 75660
rect 362234 75340 362266 75576
rect 362502 75340 362586 75576
rect 362822 75340 362854 75576
rect 362234 39896 362854 75340
rect 362234 39660 362266 39896
rect 362502 39660 362586 39896
rect 362822 39660 362854 39896
rect 362234 39576 362854 39660
rect 362234 39340 362266 39576
rect 362502 39340 362586 39576
rect 362822 39340 362854 39576
rect 362234 3896 362854 39340
rect 362234 3660 362266 3896
rect 362502 3660 362586 3896
rect 362822 3660 362854 3896
rect 362234 3576 362854 3660
rect 362234 3340 362266 3576
rect 362502 3340 362586 3576
rect 362822 3340 362854 3576
rect 362234 -1304 362854 3340
rect 362234 -1540 362266 -1304
rect 362502 -1540 362586 -1304
rect 362822 -1540 362854 -1304
rect 362234 -1624 362854 -1540
rect 362234 -1860 362266 -1624
rect 362502 -1860 362586 -1624
rect 362822 -1860 362854 -1624
rect 362234 -7652 362854 -1860
rect 363474 706760 364094 711592
rect 363474 706524 363506 706760
rect 363742 706524 363826 706760
rect 364062 706524 364094 706760
rect 363474 706440 364094 706524
rect 363474 706204 363506 706440
rect 363742 706204 363826 706440
rect 364062 706204 364094 706440
rect 363474 689136 364094 706204
rect 363474 688900 363506 689136
rect 363742 688900 363826 689136
rect 364062 688900 364094 689136
rect 363474 688816 364094 688900
rect 363474 688580 363506 688816
rect 363742 688580 363826 688816
rect 364062 688580 364094 688816
rect 363474 653136 364094 688580
rect 363474 652900 363506 653136
rect 363742 652900 363826 653136
rect 364062 652900 364094 653136
rect 363474 652816 364094 652900
rect 363474 652580 363506 652816
rect 363742 652580 363826 652816
rect 364062 652580 364094 652816
rect 363474 617136 364094 652580
rect 363474 616900 363506 617136
rect 363742 616900 363826 617136
rect 364062 616900 364094 617136
rect 363474 616816 364094 616900
rect 363474 616580 363506 616816
rect 363742 616580 363826 616816
rect 364062 616580 364094 616816
rect 363474 581136 364094 616580
rect 363474 580900 363506 581136
rect 363742 580900 363826 581136
rect 364062 580900 364094 581136
rect 363474 580816 364094 580900
rect 363474 580580 363506 580816
rect 363742 580580 363826 580816
rect 364062 580580 364094 580816
rect 363474 545136 364094 580580
rect 363474 544900 363506 545136
rect 363742 544900 363826 545136
rect 364062 544900 364094 545136
rect 363474 544816 364094 544900
rect 363474 544580 363506 544816
rect 363742 544580 363826 544816
rect 364062 544580 364094 544816
rect 363474 509136 364094 544580
rect 363474 508900 363506 509136
rect 363742 508900 363826 509136
rect 364062 508900 364094 509136
rect 363474 508816 364094 508900
rect 363474 508580 363506 508816
rect 363742 508580 363826 508816
rect 364062 508580 364094 508816
rect 363474 473136 364094 508580
rect 363474 472900 363506 473136
rect 363742 472900 363826 473136
rect 364062 472900 364094 473136
rect 363474 472816 364094 472900
rect 363474 472580 363506 472816
rect 363742 472580 363826 472816
rect 364062 472580 364094 472816
rect 363474 437136 364094 472580
rect 363474 436900 363506 437136
rect 363742 436900 363826 437136
rect 364062 436900 364094 437136
rect 363474 436816 364094 436900
rect 363474 436580 363506 436816
rect 363742 436580 363826 436816
rect 364062 436580 364094 436816
rect 363474 401136 364094 436580
rect 363474 400900 363506 401136
rect 363742 400900 363826 401136
rect 364062 400900 364094 401136
rect 363474 400816 364094 400900
rect 363474 400580 363506 400816
rect 363742 400580 363826 400816
rect 364062 400580 364094 400816
rect 363474 365136 364094 400580
rect 363474 364900 363506 365136
rect 363742 364900 363826 365136
rect 364062 364900 364094 365136
rect 363474 364816 364094 364900
rect 363474 364580 363506 364816
rect 363742 364580 363826 364816
rect 364062 364580 364094 364816
rect 363474 329136 364094 364580
rect 363474 328900 363506 329136
rect 363742 328900 363826 329136
rect 364062 328900 364094 329136
rect 363474 328816 364094 328900
rect 363474 328580 363506 328816
rect 363742 328580 363826 328816
rect 364062 328580 364094 328816
rect 363474 293136 364094 328580
rect 363474 292900 363506 293136
rect 363742 292900 363826 293136
rect 364062 292900 364094 293136
rect 363474 292816 364094 292900
rect 363474 292580 363506 292816
rect 363742 292580 363826 292816
rect 364062 292580 364094 292816
rect 363474 257136 364094 292580
rect 363474 256900 363506 257136
rect 363742 256900 363826 257136
rect 364062 256900 364094 257136
rect 363474 256816 364094 256900
rect 363474 256580 363506 256816
rect 363742 256580 363826 256816
rect 364062 256580 364094 256816
rect 363474 221136 364094 256580
rect 363474 220900 363506 221136
rect 363742 220900 363826 221136
rect 364062 220900 364094 221136
rect 363474 220816 364094 220900
rect 363474 220580 363506 220816
rect 363742 220580 363826 220816
rect 364062 220580 364094 220816
rect 363474 185136 364094 220580
rect 363474 184900 363506 185136
rect 363742 184900 363826 185136
rect 364062 184900 364094 185136
rect 363474 184816 364094 184900
rect 363474 184580 363506 184816
rect 363742 184580 363826 184816
rect 364062 184580 364094 184816
rect 363474 149136 364094 184580
rect 363474 148900 363506 149136
rect 363742 148900 363826 149136
rect 364062 148900 364094 149136
rect 363474 148816 364094 148900
rect 363474 148580 363506 148816
rect 363742 148580 363826 148816
rect 364062 148580 364094 148816
rect 363474 113136 364094 148580
rect 363474 112900 363506 113136
rect 363742 112900 363826 113136
rect 364062 112900 364094 113136
rect 363474 112816 364094 112900
rect 363474 112580 363506 112816
rect 363742 112580 363826 112816
rect 364062 112580 364094 112816
rect 363474 77136 364094 112580
rect 363474 76900 363506 77136
rect 363742 76900 363826 77136
rect 364062 76900 364094 77136
rect 363474 76816 364094 76900
rect 363474 76580 363506 76816
rect 363742 76580 363826 76816
rect 364062 76580 364094 76816
rect 363474 41136 364094 76580
rect 363474 40900 363506 41136
rect 363742 40900 363826 41136
rect 364062 40900 364094 41136
rect 363474 40816 364094 40900
rect 363474 40580 363506 40816
rect 363742 40580 363826 40816
rect 364062 40580 364094 40816
rect 363474 5136 364094 40580
rect 363474 4900 363506 5136
rect 363742 4900 363826 5136
rect 364062 4900 364094 5136
rect 363474 4816 364094 4900
rect 363474 4580 363506 4816
rect 363742 4580 363826 4816
rect 364062 4580 364094 4816
rect 363474 -2264 364094 4580
rect 363474 -2500 363506 -2264
rect 363742 -2500 363826 -2264
rect 364062 -2500 364094 -2264
rect 363474 -2584 364094 -2500
rect 363474 -2820 363506 -2584
rect 363742 -2820 363826 -2584
rect 364062 -2820 364094 -2584
rect 363474 -7652 364094 -2820
rect 364714 707720 365334 711592
rect 364714 707484 364746 707720
rect 364982 707484 365066 707720
rect 365302 707484 365334 707720
rect 364714 707400 365334 707484
rect 364714 707164 364746 707400
rect 364982 707164 365066 707400
rect 365302 707164 365334 707400
rect 364714 690376 365334 707164
rect 364714 690140 364746 690376
rect 364982 690140 365066 690376
rect 365302 690140 365334 690376
rect 364714 690056 365334 690140
rect 364714 689820 364746 690056
rect 364982 689820 365066 690056
rect 365302 689820 365334 690056
rect 364714 654376 365334 689820
rect 364714 654140 364746 654376
rect 364982 654140 365066 654376
rect 365302 654140 365334 654376
rect 364714 654056 365334 654140
rect 364714 653820 364746 654056
rect 364982 653820 365066 654056
rect 365302 653820 365334 654056
rect 364714 618376 365334 653820
rect 364714 618140 364746 618376
rect 364982 618140 365066 618376
rect 365302 618140 365334 618376
rect 364714 618056 365334 618140
rect 364714 617820 364746 618056
rect 364982 617820 365066 618056
rect 365302 617820 365334 618056
rect 364714 582376 365334 617820
rect 364714 582140 364746 582376
rect 364982 582140 365066 582376
rect 365302 582140 365334 582376
rect 364714 582056 365334 582140
rect 364714 581820 364746 582056
rect 364982 581820 365066 582056
rect 365302 581820 365334 582056
rect 364714 546376 365334 581820
rect 364714 546140 364746 546376
rect 364982 546140 365066 546376
rect 365302 546140 365334 546376
rect 364714 546056 365334 546140
rect 364714 545820 364746 546056
rect 364982 545820 365066 546056
rect 365302 545820 365334 546056
rect 364714 510376 365334 545820
rect 364714 510140 364746 510376
rect 364982 510140 365066 510376
rect 365302 510140 365334 510376
rect 364714 510056 365334 510140
rect 364714 509820 364746 510056
rect 364982 509820 365066 510056
rect 365302 509820 365334 510056
rect 364714 474376 365334 509820
rect 364714 474140 364746 474376
rect 364982 474140 365066 474376
rect 365302 474140 365334 474376
rect 364714 474056 365334 474140
rect 364714 473820 364746 474056
rect 364982 473820 365066 474056
rect 365302 473820 365334 474056
rect 364714 438376 365334 473820
rect 364714 438140 364746 438376
rect 364982 438140 365066 438376
rect 365302 438140 365334 438376
rect 364714 438056 365334 438140
rect 364714 437820 364746 438056
rect 364982 437820 365066 438056
rect 365302 437820 365334 438056
rect 364714 402376 365334 437820
rect 364714 402140 364746 402376
rect 364982 402140 365066 402376
rect 365302 402140 365334 402376
rect 364714 402056 365334 402140
rect 364714 401820 364746 402056
rect 364982 401820 365066 402056
rect 365302 401820 365334 402056
rect 364714 366376 365334 401820
rect 364714 366140 364746 366376
rect 364982 366140 365066 366376
rect 365302 366140 365334 366376
rect 364714 366056 365334 366140
rect 364714 365820 364746 366056
rect 364982 365820 365066 366056
rect 365302 365820 365334 366056
rect 364714 330376 365334 365820
rect 364714 330140 364746 330376
rect 364982 330140 365066 330376
rect 365302 330140 365334 330376
rect 364714 330056 365334 330140
rect 364714 329820 364746 330056
rect 364982 329820 365066 330056
rect 365302 329820 365334 330056
rect 364714 294376 365334 329820
rect 364714 294140 364746 294376
rect 364982 294140 365066 294376
rect 365302 294140 365334 294376
rect 364714 294056 365334 294140
rect 364714 293820 364746 294056
rect 364982 293820 365066 294056
rect 365302 293820 365334 294056
rect 364714 258376 365334 293820
rect 364714 258140 364746 258376
rect 364982 258140 365066 258376
rect 365302 258140 365334 258376
rect 364714 258056 365334 258140
rect 364714 257820 364746 258056
rect 364982 257820 365066 258056
rect 365302 257820 365334 258056
rect 364714 222376 365334 257820
rect 364714 222140 364746 222376
rect 364982 222140 365066 222376
rect 365302 222140 365334 222376
rect 364714 222056 365334 222140
rect 364714 221820 364746 222056
rect 364982 221820 365066 222056
rect 365302 221820 365334 222056
rect 364714 186376 365334 221820
rect 364714 186140 364746 186376
rect 364982 186140 365066 186376
rect 365302 186140 365334 186376
rect 364714 186056 365334 186140
rect 364714 185820 364746 186056
rect 364982 185820 365066 186056
rect 365302 185820 365334 186056
rect 364714 150376 365334 185820
rect 364714 150140 364746 150376
rect 364982 150140 365066 150376
rect 365302 150140 365334 150376
rect 364714 150056 365334 150140
rect 364714 149820 364746 150056
rect 364982 149820 365066 150056
rect 365302 149820 365334 150056
rect 364714 114376 365334 149820
rect 364714 114140 364746 114376
rect 364982 114140 365066 114376
rect 365302 114140 365334 114376
rect 364714 114056 365334 114140
rect 364714 113820 364746 114056
rect 364982 113820 365066 114056
rect 365302 113820 365334 114056
rect 364714 78376 365334 113820
rect 364714 78140 364746 78376
rect 364982 78140 365066 78376
rect 365302 78140 365334 78376
rect 364714 78056 365334 78140
rect 364714 77820 364746 78056
rect 364982 77820 365066 78056
rect 365302 77820 365334 78056
rect 364714 42376 365334 77820
rect 364714 42140 364746 42376
rect 364982 42140 365066 42376
rect 365302 42140 365334 42376
rect 364714 42056 365334 42140
rect 364714 41820 364746 42056
rect 364982 41820 365066 42056
rect 365302 41820 365334 42056
rect 364714 6376 365334 41820
rect 364714 6140 364746 6376
rect 364982 6140 365066 6376
rect 365302 6140 365334 6376
rect 364714 6056 365334 6140
rect 364714 5820 364746 6056
rect 364982 5820 365066 6056
rect 365302 5820 365334 6056
rect 364714 -3224 365334 5820
rect 364714 -3460 364746 -3224
rect 364982 -3460 365066 -3224
rect 365302 -3460 365334 -3224
rect 364714 -3544 365334 -3460
rect 364714 -3780 364746 -3544
rect 364982 -3780 365066 -3544
rect 365302 -3780 365334 -3544
rect 364714 -7652 365334 -3780
rect 365954 708680 366574 711592
rect 365954 708444 365986 708680
rect 366222 708444 366306 708680
rect 366542 708444 366574 708680
rect 365954 708360 366574 708444
rect 365954 708124 365986 708360
rect 366222 708124 366306 708360
rect 366542 708124 366574 708360
rect 365954 691616 366574 708124
rect 365954 691380 365986 691616
rect 366222 691380 366306 691616
rect 366542 691380 366574 691616
rect 365954 691296 366574 691380
rect 365954 691060 365986 691296
rect 366222 691060 366306 691296
rect 366542 691060 366574 691296
rect 365954 655616 366574 691060
rect 365954 655380 365986 655616
rect 366222 655380 366306 655616
rect 366542 655380 366574 655616
rect 365954 655296 366574 655380
rect 365954 655060 365986 655296
rect 366222 655060 366306 655296
rect 366542 655060 366574 655296
rect 365954 619616 366574 655060
rect 365954 619380 365986 619616
rect 366222 619380 366306 619616
rect 366542 619380 366574 619616
rect 365954 619296 366574 619380
rect 365954 619060 365986 619296
rect 366222 619060 366306 619296
rect 366542 619060 366574 619296
rect 365954 583616 366574 619060
rect 365954 583380 365986 583616
rect 366222 583380 366306 583616
rect 366542 583380 366574 583616
rect 365954 583296 366574 583380
rect 365954 583060 365986 583296
rect 366222 583060 366306 583296
rect 366542 583060 366574 583296
rect 365954 547616 366574 583060
rect 365954 547380 365986 547616
rect 366222 547380 366306 547616
rect 366542 547380 366574 547616
rect 365954 547296 366574 547380
rect 365954 547060 365986 547296
rect 366222 547060 366306 547296
rect 366542 547060 366574 547296
rect 365954 511616 366574 547060
rect 365954 511380 365986 511616
rect 366222 511380 366306 511616
rect 366542 511380 366574 511616
rect 365954 511296 366574 511380
rect 365954 511060 365986 511296
rect 366222 511060 366306 511296
rect 366542 511060 366574 511296
rect 365954 475616 366574 511060
rect 365954 475380 365986 475616
rect 366222 475380 366306 475616
rect 366542 475380 366574 475616
rect 365954 475296 366574 475380
rect 365954 475060 365986 475296
rect 366222 475060 366306 475296
rect 366542 475060 366574 475296
rect 365954 439616 366574 475060
rect 365954 439380 365986 439616
rect 366222 439380 366306 439616
rect 366542 439380 366574 439616
rect 365954 439296 366574 439380
rect 365954 439060 365986 439296
rect 366222 439060 366306 439296
rect 366542 439060 366574 439296
rect 365954 403616 366574 439060
rect 365954 403380 365986 403616
rect 366222 403380 366306 403616
rect 366542 403380 366574 403616
rect 365954 403296 366574 403380
rect 365954 403060 365986 403296
rect 366222 403060 366306 403296
rect 366542 403060 366574 403296
rect 365954 367616 366574 403060
rect 365954 367380 365986 367616
rect 366222 367380 366306 367616
rect 366542 367380 366574 367616
rect 365954 367296 366574 367380
rect 365954 367060 365986 367296
rect 366222 367060 366306 367296
rect 366542 367060 366574 367296
rect 365954 331616 366574 367060
rect 365954 331380 365986 331616
rect 366222 331380 366306 331616
rect 366542 331380 366574 331616
rect 365954 331296 366574 331380
rect 365954 331060 365986 331296
rect 366222 331060 366306 331296
rect 366542 331060 366574 331296
rect 365954 295616 366574 331060
rect 365954 295380 365986 295616
rect 366222 295380 366306 295616
rect 366542 295380 366574 295616
rect 365954 295296 366574 295380
rect 365954 295060 365986 295296
rect 366222 295060 366306 295296
rect 366542 295060 366574 295296
rect 365954 259616 366574 295060
rect 365954 259380 365986 259616
rect 366222 259380 366306 259616
rect 366542 259380 366574 259616
rect 365954 259296 366574 259380
rect 365954 259060 365986 259296
rect 366222 259060 366306 259296
rect 366542 259060 366574 259296
rect 365954 223616 366574 259060
rect 365954 223380 365986 223616
rect 366222 223380 366306 223616
rect 366542 223380 366574 223616
rect 365954 223296 366574 223380
rect 365954 223060 365986 223296
rect 366222 223060 366306 223296
rect 366542 223060 366574 223296
rect 365954 187616 366574 223060
rect 365954 187380 365986 187616
rect 366222 187380 366306 187616
rect 366542 187380 366574 187616
rect 365954 187296 366574 187380
rect 365954 187060 365986 187296
rect 366222 187060 366306 187296
rect 366542 187060 366574 187296
rect 365954 151616 366574 187060
rect 365954 151380 365986 151616
rect 366222 151380 366306 151616
rect 366542 151380 366574 151616
rect 365954 151296 366574 151380
rect 365954 151060 365986 151296
rect 366222 151060 366306 151296
rect 366542 151060 366574 151296
rect 365954 115616 366574 151060
rect 365954 115380 365986 115616
rect 366222 115380 366306 115616
rect 366542 115380 366574 115616
rect 365954 115296 366574 115380
rect 365954 115060 365986 115296
rect 366222 115060 366306 115296
rect 366542 115060 366574 115296
rect 365954 79616 366574 115060
rect 365954 79380 365986 79616
rect 366222 79380 366306 79616
rect 366542 79380 366574 79616
rect 365954 79296 366574 79380
rect 365954 79060 365986 79296
rect 366222 79060 366306 79296
rect 366542 79060 366574 79296
rect 365954 43616 366574 79060
rect 365954 43380 365986 43616
rect 366222 43380 366306 43616
rect 366542 43380 366574 43616
rect 365954 43296 366574 43380
rect 365954 43060 365986 43296
rect 366222 43060 366306 43296
rect 366542 43060 366574 43296
rect 365954 7616 366574 43060
rect 365954 7380 365986 7616
rect 366222 7380 366306 7616
rect 366542 7380 366574 7616
rect 365954 7296 366574 7380
rect 365954 7060 365986 7296
rect 366222 7060 366306 7296
rect 366542 7060 366574 7296
rect 365954 -4184 366574 7060
rect 365954 -4420 365986 -4184
rect 366222 -4420 366306 -4184
rect 366542 -4420 366574 -4184
rect 365954 -4504 366574 -4420
rect 365954 -4740 365986 -4504
rect 366222 -4740 366306 -4504
rect 366542 -4740 366574 -4504
rect 365954 -7652 366574 -4740
rect 367194 709640 367814 711592
rect 367194 709404 367226 709640
rect 367462 709404 367546 709640
rect 367782 709404 367814 709640
rect 367194 709320 367814 709404
rect 367194 709084 367226 709320
rect 367462 709084 367546 709320
rect 367782 709084 367814 709320
rect 367194 692856 367814 709084
rect 367194 692620 367226 692856
rect 367462 692620 367546 692856
rect 367782 692620 367814 692856
rect 367194 692536 367814 692620
rect 367194 692300 367226 692536
rect 367462 692300 367546 692536
rect 367782 692300 367814 692536
rect 367194 656856 367814 692300
rect 367194 656620 367226 656856
rect 367462 656620 367546 656856
rect 367782 656620 367814 656856
rect 367194 656536 367814 656620
rect 367194 656300 367226 656536
rect 367462 656300 367546 656536
rect 367782 656300 367814 656536
rect 367194 620856 367814 656300
rect 367194 620620 367226 620856
rect 367462 620620 367546 620856
rect 367782 620620 367814 620856
rect 367194 620536 367814 620620
rect 367194 620300 367226 620536
rect 367462 620300 367546 620536
rect 367782 620300 367814 620536
rect 367194 584856 367814 620300
rect 367194 584620 367226 584856
rect 367462 584620 367546 584856
rect 367782 584620 367814 584856
rect 367194 584536 367814 584620
rect 367194 584300 367226 584536
rect 367462 584300 367546 584536
rect 367782 584300 367814 584536
rect 367194 548856 367814 584300
rect 367194 548620 367226 548856
rect 367462 548620 367546 548856
rect 367782 548620 367814 548856
rect 367194 548536 367814 548620
rect 367194 548300 367226 548536
rect 367462 548300 367546 548536
rect 367782 548300 367814 548536
rect 367194 512856 367814 548300
rect 367194 512620 367226 512856
rect 367462 512620 367546 512856
rect 367782 512620 367814 512856
rect 367194 512536 367814 512620
rect 367194 512300 367226 512536
rect 367462 512300 367546 512536
rect 367782 512300 367814 512536
rect 367194 476856 367814 512300
rect 367194 476620 367226 476856
rect 367462 476620 367546 476856
rect 367782 476620 367814 476856
rect 367194 476536 367814 476620
rect 367194 476300 367226 476536
rect 367462 476300 367546 476536
rect 367782 476300 367814 476536
rect 367194 440856 367814 476300
rect 367194 440620 367226 440856
rect 367462 440620 367546 440856
rect 367782 440620 367814 440856
rect 367194 440536 367814 440620
rect 367194 440300 367226 440536
rect 367462 440300 367546 440536
rect 367782 440300 367814 440536
rect 367194 404856 367814 440300
rect 367194 404620 367226 404856
rect 367462 404620 367546 404856
rect 367782 404620 367814 404856
rect 367194 404536 367814 404620
rect 367194 404300 367226 404536
rect 367462 404300 367546 404536
rect 367782 404300 367814 404536
rect 367194 368856 367814 404300
rect 367194 368620 367226 368856
rect 367462 368620 367546 368856
rect 367782 368620 367814 368856
rect 367194 368536 367814 368620
rect 367194 368300 367226 368536
rect 367462 368300 367546 368536
rect 367782 368300 367814 368536
rect 367194 332856 367814 368300
rect 367194 332620 367226 332856
rect 367462 332620 367546 332856
rect 367782 332620 367814 332856
rect 367194 332536 367814 332620
rect 367194 332300 367226 332536
rect 367462 332300 367546 332536
rect 367782 332300 367814 332536
rect 367194 296856 367814 332300
rect 367194 296620 367226 296856
rect 367462 296620 367546 296856
rect 367782 296620 367814 296856
rect 367194 296536 367814 296620
rect 367194 296300 367226 296536
rect 367462 296300 367546 296536
rect 367782 296300 367814 296536
rect 367194 260856 367814 296300
rect 367194 260620 367226 260856
rect 367462 260620 367546 260856
rect 367782 260620 367814 260856
rect 367194 260536 367814 260620
rect 367194 260300 367226 260536
rect 367462 260300 367546 260536
rect 367782 260300 367814 260536
rect 367194 224856 367814 260300
rect 367194 224620 367226 224856
rect 367462 224620 367546 224856
rect 367782 224620 367814 224856
rect 367194 224536 367814 224620
rect 367194 224300 367226 224536
rect 367462 224300 367546 224536
rect 367782 224300 367814 224536
rect 367194 188856 367814 224300
rect 367194 188620 367226 188856
rect 367462 188620 367546 188856
rect 367782 188620 367814 188856
rect 367194 188536 367814 188620
rect 367194 188300 367226 188536
rect 367462 188300 367546 188536
rect 367782 188300 367814 188536
rect 367194 152856 367814 188300
rect 367194 152620 367226 152856
rect 367462 152620 367546 152856
rect 367782 152620 367814 152856
rect 367194 152536 367814 152620
rect 367194 152300 367226 152536
rect 367462 152300 367546 152536
rect 367782 152300 367814 152536
rect 367194 116856 367814 152300
rect 367194 116620 367226 116856
rect 367462 116620 367546 116856
rect 367782 116620 367814 116856
rect 367194 116536 367814 116620
rect 367194 116300 367226 116536
rect 367462 116300 367546 116536
rect 367782 116300 367814 116536
rect 367194 80856 367814 116300
rect 367194 80620 367226 80856
rect 367462 80620 367546 80856
rect 367782 80620 367814 80856
rect 367194 80536 367814 80620
rect 367194 80300 367226 80536
rect 367462 80300 367546 80536
rect 367782 80300 367814 80536
rect 367194 44856 367814 80300
rect 367194 44620 367226 44856
rect 367462 44620 367546 44856
rect 367782 44620 367814 44856
rect 367194 44536 367814 44620
rect 367194 44300 367226 44536
rect 367462 44300 367546 44536
rect 367782 44300 367814 44536
rect 367194 8856 367814 44300
rect 367194 8620 367226 8856
rect 367462 8620 367546 8856
rect 367782 8620 367814 8856
rect 367194 8536 367814 8620
rect 367194 8300 367226 8536
rect 367462 8300 367546 8536
rect 367782 8300 367814 8536
rect 367194 -5144 367814 8300
rect 367194 -5380 367226 -5144
rect 367462 -5380 367546 -5144
rect 367782 -5380 367814 -5144
rect 367194 -5464 367814 -5380
rect 367194 -5700 367226 -5464
rect 367462 -5700 367546 -5464
rect 367782 -5700 367814 -5464
rect 367194 -7652 367814 -5700
rect 368434 710600 369054 711592
rect 368434 710364 368466 710600
rect 368702 710364 368786 710600
rect 369022 710364 369054 710600
rect 368434 710280 369054 710364
rect 368434 710044 368466 710280
rect 368702 710044 368786 710280
rect 369022 710044 369054 710280
rect 368434 694096 369054 710044
rect 368434 693860 368466 694096
rect 368702 693860 368786 694096
rect 369022 693860 369054 694096
rect 368434 693776 369054 693860
rect 368434 693540 368466 693776
rect 368702 693540 368786 693776
rect 369022 693540 369054 693776
rect 368434 658096 369054 693540
rect 368434 657860 368466 658096
rect 368702 657860 368786 658096
rect 369022 657860 369054 658096
rect 368434 657776 369054 657860
rect 368434 657540 368466 657776
rect 368702 657540 368786 657776
rect 369022 657540 369054 657776
rect 368434 622096 369054 657540
rect 368434 621860 368466 622096
rect 368702 621860 368786 622096
rect 369022 621860 369054 622096
rect 368434 621776 369054 621860
rect 368434 621540 368466 621776
rect 368702 621540 368786 621776
rect 369022 621540 369054 621776
rect 368434 586096 369054 621540
rect 368434 585860 368466 586096
rect 368702 585860 368786 586096
rect 369022 585860 369054 586096
rect 368434 585776 369054 585860
rect 368434 585540 368466 585776
rect 368702 585540 368786 585776
rect 369022 585540 369054 585776
rect 368434 550096 369054 585540
rect 368434 549860 368466 550096
rect 368702 549860 368786 550096
rect 369022 549860 369054 550096
rect 368434 549776 369054 549860
rect 368434 549540 368466 549776
rect 368702 549540 368786 549776
rect 369022 549540 369054 549776
rect 368434 514096 369054 549540
rect 368434 513860 368466 514096
rect 368702 513860 368786 514096
rect 369022 513860 369054 514096
rect 368434 513776 369054 513860
rect 368434 513540 368466 513776
rect 368702 513540 368786 513776
rect 369022 513540 369054 513776
rect 368434 478096 369054 513540
rect 368434 477860 368466 478096
rect 368702 477860 368786 478096
rect 369022 477860 369054 478096
rect 368434 477776 369054 477860
rect 368434 477540 368466 477776
rect 368702 477540 368786 477776
rect 369022 477540 369054 477776
rect 368434 442096 369054 477540
rect 368434 441860 368466 442096
rect 368702 441860 368786 442096
rect 369022 441860 369054 442096
rect 368434 441776 369054 441860
rect 368434 441540 368466 441776
rect 368702 441540 368786 441776
rect 369022 441540 369054 441776
rect 368434 406096 369054 441540
rect 368434 405860 368466 406096
rect 368702 405860 368786 406096
rect 369022 405860 369054 406096
rect 368434 405776 369054 405860
rect 368434 405540 368466 405776
rect 368702 405540 368786 405776
rect 369022 405540 369054 405776
rect 368434 370096 369054 405540
rect 368434 369860 368466 370096
rect 368702 369860 368786 370096
rect 369022 369860 369054 370096
rect 368434 369776 369054 369860
rect 368434 369540 368466 369776
rect 368702 369540 368786 369776
rect 369022 369540 369054 369776
rect 368434 334096 369054 369540
rect 368434 333860 368466 334096
rect 368702 333860 368786 334096
rect 369022 333860 369054 334096
rect 368434 333776 369054 333860
rect 368434 333540 368466 333776
rect 368702 333540 368786 333776
rect 369022 333540 369054 333776
rect 368434 298096 369054 333540
rect 368434 297860 368466 298096
rect 368702 297860 368786 298096
rect 369022 297860 369054 298096
rect 368434 297776 369054 297860
rect 368434 297540 368466 297776
rect 368702 297540 368786 297776
rect 369022 297540 369054 297776
rect 368434 262096 369054 297540
rect 368434 261860 368466 262096
rect 368702 261860 368786 262096
rect 369022 261860 369054 262096
rect 368434 261776 369054 261860
rect 368434 261540 368466 261776
rect 368702 261540 368786 261776
rect 369022 261540 369054 261776
rect 368434 226096 369054 261540
rect 368434 225860 368466 226096
rect 368702 225860 368786 226096
rect 369022 225860 369054 226096
rect 368434 225776 369054 225860
rect 368434 225540 368466 225776
rect 368702 225540 368786 225776
rect 369022 225540 369054 225776
rect 368434 190096 369054 225540
rect 368434 189860 368466 190096
rect 368702 189860 368786 190096
rect 369022 189860 369054 190096
rect 368434 189776 369054 189860
rect 368434 189540 368466 189776
rect 368702 189540 368786 189776
rect 369022 189540 369054 189776
rect 368434 154096 369054 189540
rect 368434 153860 368466 154096
rect 368702 153860 368786 154096
rect 369022 153860 369054 154096
rect 368434 153776 369054 153860
rect 368434 153540 368466 153776
rect 368702 153540 368786 153776
rect 369022 153540 369054 153776
rect 368434 118096 369054 153540
rect 368434 117860 368466 118096
rect 368702 117860 368786 118096
rect 369022 117860 369054 118096
rect 368434 117776 369054 117860
rect 368434 117540 368466 117776
rect 368702 117540 368786 117776
rect 369022 117540 369054 117776
rect 368434 82096 369054 117540
rect 368434 81860 368466 82096
rect 368702 81860 368786 82096
rect 369022 81860 369054 82096
rect 368434 81776 369054 81860
rect 368434 81540 368466 81776
rect 368702 81540 368786 81776
rect 369022 81540 369054 81776
rect 368434 46096 369054 81540
rect 368434 45860 368466 46096
rect 368702 45860 368786 46096
rect 369022 45860 369054 46096
rect 368434 45776 369054 45860
rect 368434 45540 368466 45776
rect 368702 45540 368786 45776
rect 369022 45540 369054 45776
rect 368434 10096 369054 45540
rect 368434 9860 368466 10096
rect 368702 9860 368786 10096
rect 369022 9860 369054 10096
rect 368434 9776 369054 9860
rect 368434 9540 368466 9776
rect 368702 9540 368786 9776
rect 369022 9540 369054 9776
rect 368434 -6104 369054 9540
rect 368434 -6340 368466 -6104
rect 368702 -6340 368786 -6104
rect 369022 -6340 369054 -6104
rect 368434 -6424 369054 -6340
rect 368434 -6660 368466 -6424
rect 368702 -6660 368786 -6424
rect 369022 -6660 369054 -6424
rect 368434 -7652 369054 -6660
rect 369674 711560 370294 711592
rect 369674 711324 369706 711560
rect 369942 711324 370026 711560
rect 370262 711324 370294 711560
rect 369674 711240 370294 711324
rect 369674 711004 369706 711240
rect 369942 711004 370026 711240
rect 370262 711004 370294 711240
rect 369674 695336 370294 711004
rect 369674 695100 369706 695336
rect 369942 695100 370026 695336
rect 370262 695100 370294 695336
rect 369674 695016 370294 695100
rect 369674 694780 369706 695016
rect 369942 694780 370026 695016
rect 370262 694780 370294 695016
rect 369674 659336 370294 694780
rect 369674 659100 369706 659336
rect 369942 659100 370026 659336
rect 370262 659100 370294 659336
rect 369674 659016 370294 659100
rect 369674 658780 369706 659016
rect 369942 658780 370026 659016
rect 370262 658780 370294 659016
rect 369674 623336 370294 658780
rect 369674 623100 369706 623336
rect 369942 623100 370026 623336
rect 370262 623100 370294 623336
rect 369674 623016 370294 623100
rect 369674 622780 369706 623016
rect 369942 622780 370026 623016
rect 370262 622780 370294 623016
rect 369674 587336 370294 622780
rect 369674 587100 369706 587336
rect 369942 587100 370026 587336
rect 370262 587100 370294 587336
rect 369674 587016 370294 587100
rect 369674 586780 369706 587016
rect 369942 586780 370026 587016
rect 370262 586780 370294 587016
rect 369674 551336 370294 586780
rect 369674 551100 369706 551336
rect 369942 551100 370026 551336
rect 370262 551100 370294 551336
rect 369674 551016 370294 551100
rect 369674 550780 369706 551016
rect 369942 550780 370026 551016
rect 370262 550780 370294 551016
rect 369674 515336 370294 550780
rect 369674 515100 369706 515336
rect 369942 515100 370026 515336
rect 370262 515100 370294 515336
rect 369674 515016 370294 515100
rect 369674 514780 369706 515016
rect 369942 514780 370026 515016
rect 370262 514780 370294 515016
rect 369674 479336 370294 514780
rect 369674 479100 369706 479336
rect 369942 479100 370026 479336
rect 370262 479100 370294 479336
rect 369674 479016 370294 479100
rect 369674 478780 369706 479016
rect 369942 478780 370026 479016
rect 370262 478780 370294 479016
rect 369674 443336 370294 478780
rect 369674 443100 369706 443336
rect 369942 443100 370026 443336
rect 370262 443100 370294 443336
rect 369674 443016 370294 443100
rect 369674 442780 369706 443016
rect 369942 442780 370026 443016
rect 370262 442780 370294 443016
rect 369674 407336 370294 442780
rect 369674 407100 369706 407336
rect 369942 407100 370026 407336
rect 370262 407100 370294 407336
rect 369674 407016 370294 407100
rect 369674 406780 369706 407016
rect 369942 406780 370026 407016
rect 370262 406780 370294 407016
rect 369674 371336 370294 406780
rect 369674 371100 369706 371336
rect 369942 371100 370026 371336
rect 370262 371100 370294 371336
rect 369674 371016 370294 371100
rect 369674 370780 369706 371016
rect 369942 370780 370026 371016
rect 370262 370780 370294 371016
rect 369674 335336 370294 370780
rect 369674 335100 369706 335336
rect 369942 335100 370026 335336
rect 370262 335100 370294 335336
rect 369674 335016 370294 335100
rect 369674 334780 369706 335016
rect 369942 334780 370026 335016
rect 370262 334780 370294 335016
rect 369674 299336 370294 334780
rect 369674 299100 369706 299336
rect 369942 299100 370026 299336
rect 370262 299100 370294 299336
rect 369674 299016 370294 299100
rect 369674 298780 369706 299016
rect 369942 298780 370026 299016
rect 370262 298780 370294 299016
rect 369674 263336 370294 298780
rect 369674 263100 369706 263336
rect 369942 263100 370026 263336
rect 370262 263100 370294 263336
rect 369674 263016 370294 263100
rect 369674 262780 369706 263016
rect 369942 262780 370026 263016
rect 370262 262780 370294 263016
rect 369674 227336 370294 262780
rect 369674 227100 369706 227336
rect 369942 227100 370026 227336
rect 370262 227100 370294 227336
rect 369674 227016 370294 227100
rect 369674 226780 369706 227016
rect 369942 226780 370026 227016
rect 370262 226780 370294 227016
rect 369674 191336 370294 226780
rect 369674 191100 369706 191336
rect 369942 191100 370026 191336
rect 370262 191100 370294 191336
rect 369674 191016 370294 191100
rect 369674 190780 369706 191016
rect 369942 190780 370026 191016
rect 370262 190780 370294 191016
rect 369674 155336 370294 190780
rect 369674 155100 369706 155336
rect 369942 155100 370026 155336
rect 370262 155100 370294 155336
rect 369674 155016 370294 155100
rect 369674 154780 369706 155016
rect 369942 154780 370026 155016
rect 370262 154780 370294 155016
rect 369674 119336 370294 154780
rect 369674 119100 369706 119336
rect 369942 119100 370026 119336
rect 370262 119100 370294 119336
rect 369674 119016 370294 119100
rect 369674 118780 369706 119016
rect 369942 118780 370026 119016
rect 370262 118780 370294 119016
rect 369674 83336 370294 118780
rect 369674 83100 369706 83336
rect 369942 83100 370026 83336
rect 370262 83100 370294 83336
rect 369674 83016 370294 83100
rect 369674 82780 369706 83016
rect 369942 82780 370026 83016
rect 370262 82780 370294 83016
rect 369674 47336 370294 82780
rect 369674 47100 369706 47336
rect 369942 47100 370026 47336
rect 370262 47100 370294 47336
rect 369674 47016 370294 47100
rect 369674 46780 369706 47016
rect 369942 46780 370026 47016
rect 370262 46780 370294 47016
rect 369674 11336 370294 46780
rect 369674 11100 369706 11336
rect 369942 11100 370026 11336
rect 370262 11100 370294 11336
rect 369674 11016 370294 11100
rect 369674 10780 369706 11016
rect 369942 10780 370026 11016
rect 370262 10780 370294 11016
rect 369674 -7064 370294 10780
rect 369674 -7300 369706 -7064
rect 369942 -7300 370026 -7064
rect 370262 -7300 370294 -7064
rect 369674 -7384 370294 -7300
rect 369674 -7620 369706 -7384
rect 369942 -7620 370026 -7384
rect 370262 -7620 370294 -7384
rect 369674 -7652 370294 -7620
rect 396994 704840 397614 711592
rect 396994 704604 397026 704840
rect 397262 704604 397346 704840
rect 397582 704604 397614 704840
rect 396994 704520 397614 704604
rect 396994 704284 397026 704520
rect 397262 704284 397346 704520
rect 397582 704284 397614 704520
rect 396994 686656 397614 704284
rect 396994 686420 397026 686656
rect 397262 686420 397346 686656
rect 397582 686420 397614 686656
rect 396994 686336 397614 686420
rect 396994 686100 397026 686336
rect 397262 686100 397346 686336
rect 397582 686100 397614 686336
rect 396994 650656 397614 686100
rect 396994 650420 397026 650656
rect 397262 650420 397346 650656
rect 397582 650420 397614 650656
rect 396994 650336 397614 650420
rect 396994 650100 397026 650336
rect 397262 650100 397346 650336
rect 397582 650100 397614 650336
rect 396994 614656 397614 650100
rect 396994 614420 397026 614656
rect 397262 614420 397346 614656
rect 397582 614420 397614 614656
rect 396994 614336 397614 614420
rect 396994 614100 397026 614336
rect 397262 614100 397346 614336
rect 397582 614100 397614 614336
rect 396994 578656 397614 614100
rect 396994 578420 397026 578656
rect 397262 578420 397346 578656
rect 397582 578420 397614 578656
rect 396994 578336 397614 578420
rect 396994 578100 397026 578336
rect 397262 578100 397346 578336
rect 397582 578100 397614 578336
rect 396994 542656 397614 578100
rect 396994 542420 397026 542656
rect 397262 542420 397346 542656
rect 397582 542420 397614 542656
rect 396994 542336 397614 542420
rect 396994 542100 397026 542336
rect 397262 542100 397346 542336
rect 397582 542100 397614 542336
rect 396994 506656 397614 542100
rect 396994 506420 397026 506656
rect 397262 506420 397346 506656
rect 397582 506420 397614 506656
rect 396994 506336 397614 506420
rect 396994 506100 397026 506336
rect 397262 506100 397346 506336
rect 397582 506100 397614 506336
rect 396994 470656 397614 506100
rect 396994 470420 397026 470656
rect 397262 470420 397346 470656
rect 397582 470420 397614 470656
rect 396994 470336 397614 470420
rect 396994 470100 397026 470336
rect 397262 470100 397346 470336
rect 397582 470100 397614 470336
rect 396994 434656 397614 470100
rect 396994 434420 397026 434656
rect 397262 434420 397346 434656
rect 397582 434420 397614 434656
rect 396994 434336 397614 434420
rect 396994 434100 397026 434336
rect 397262 434100 397346 434336
rect 397582 434100 397614 434336
rect 396994 398656 397614 434100
rect 396994 398420 397026 398656
rect 397262 398420 397346 398656
rect 397582 398420 397614 398656
rect 396994 398336 397614 398420
rect 396994 398100 397026 398336
rect 397262 398100 397346 398336
rect 397582 398100 397614 398336
rect 396994 362656 397614 398100
rect 396994 362420 397026 362656
rect 397262 362420 397346 362656
rect 397582 362420 397614 362656
rect 396994 362336 397614 362420
rect 396994 362100 397026 362336
rect 397262 362100 397346 362336
rect 397582 362100 397614 362336
rect 396994 326656 397614 362100
rect 396994 326420 397026 326656
rect 397262 326420 397346 326656
rect 397582 326420 397614 326656
rect 396994 326336 397614 326420
rect 396994 326100 397026 326336
rect 397262 326100 397346 326336
rect 397582 326100 397614 326336
rect 396994 290656 397614 326100
rect 396994 290420 397026 290656
rect 397262 290420 397346 290656
rect 397582 290420 397614 290656
rect 396994 290336 397614 290420
rect 396994 290100 397026 290336
rect 397262 290100 397346 290336
rect 397582 290100 397614 290336
rect 396994 254656 397614 290100
rect 396994 254420 397026 254656
rect 397262 254420 397346 254656
rect 397582 254420 397614 254656
rect 396994 254336 397614 254420
rect 396994 254100 397026 254336
rect 397262 254100 397346 254336
rect 397582 254100 397614 254336
rect 396994 218656 397614 254100
rect 396994 218420 397026 218656
rect 397262 218420 397346 218656
rect 397582 218420 397614 218656
rect 396994 218336 397614 218420
rect 396994 218100 397026 218336
rect 397262 218100 397346 218336
rect 397582 218100 397614 218336
rect 396994 182656 397614 218100
rect 396994 182420 397026 182656
rect 397262 182420 397346 182656
rect 397582 182420 397614 182656
rect 396994 182336 397614 182420
rect 396994 182100 397026 182336
rect 397262 182100 397346 182336
rect 397582 182100 397614 182336
rect 396994 146656 397614 182100
rect 396994 146420 397026 146656
rect 397262 146420 397346 146656
rect 397582 146420 397614 146656
rect 396994 146336 397614 146420
rect 396994 146100 397026 146336
rect 397262 146100 397346 146336
rect 397582 146100 397614 146336
rect 396994 110656 397614 146100
rect 396994 110420 397026 110656
rect 397262 110420 397346 110656
rect 397582 110420 397614 110656
rect 396994 110336 397614 110420
rect 396994 110100 397026 110336
rect 397262 110100 397346 110336
rect 397582 110100 397614 110336
rect 396994 74656 397614 110100
rect 396994 74420 397026 74656
rect 397262 74420 397346 74656
rect 397582 74420 397614 74656
rect 396994 74336 397614 74420
rect 396994 74100 397026 74336
rect 397262 74100 397346 74336
rect 397582 74100 397614 74336
rect 396994 38656 397614 74100
rect 396994 38420 397026 38656
rect 397262 38420 397346 38656
rect 397582 38420 397614 38656
rect 396994 38336 397614 38420
rect 396994 38100 397026 38336
rect 397262 38100 397346 38336
rect 397582 38100 397614 38336
rect 396994 2656 397614 38100
rect 396994 2420 397026 2656
rect 397262 2420 397346 2656
rect 397582 2420 397614 2656
rect 396994 2336 397614 2420
rect 396994 2100 397026 2336
rect 397262 2100 397346 2336
rect 397582 2100 397614 2336
rect 396994 -344 397614 2100
rect 396994 -580 397026 -344
rect 397262 -580 397346 -344
rect 397582 -580 397614 -344
rect 396994 -664 397614 -580
rect 396994 -900 397026 -664
rect 397262 -900 397346 -664
rect 397582 -900 397614 -664
rect 396994 -7652 397614 -900
rect 398234 705800 398854 711592
rect 398234 705564 398266 705800
rect 398502 705564 398586 705800
rect 398822 705564 398854 705800
rect 398234 705480 398854 705564
rect 398234 705244 398266 705480
rect 398502 705244 398586 705480
rect 398822 705244 398854 705480
rect 398234 687896 398854 705244
rect 398234 687660 398266 687896
rect 398502 687660 398586 687896
rect 398822 687660 398854 687896
rect 398234 687576 398854 687660
rect 398234 687340 398266 687576
rect 398502 687340 398586 687576
rect 398822 687340 398854 687576
rect 398234 651896 398854 687340
rect 398234 651660 398266 651896
rect 398502 651660 398586 651896
rect 398822 651660 398854 651896
rect 398234 651576 398854 651660
rect 398234 651340 398266 651576
rect 398502 651340 398586 651576
rect 398822 651340 398854 651576
rect 398234 615896 398854 651340
rect 398234 615660 398266 615896
rect 398502 615660 398586 615896
rect 398822 615660 398854 615896
rect 398234 615576 398854 615660
rect 398234 615340 398266 615576
rect 398502 615340 398586 615576
rect 398822 615340 398854 615576
rect 398234 579896 398854 615340
rect 398234 579660 398266 579896
rect 398502 579660 398586 579896
rect 398822 579660 398854 579896
rect 398234 579576 398854 579660
rect 398234 579340 398266 579576
rect 398502 579340 398586 579576
rect 398822 579340 398854 579576
rect 398234 543896 398854 579340
rect 398234 543660 398266 543896
rect 398502 543660 398586 543896
rect 398822 543660 398854 543896
rect 398234 543576 398854 543660
rect 398234 543340 398266 543576
rect 398502 543340 398586 543576
rect 398822 543340 398854 543576
rect 398234 507896 398854 543340
rect 398234 507660 398266 507896
rect 398502 507660 398586 507896
rect 398822 507660 398854 507896
rect 398234 507576 398854 507660
rect 398234 507340 398266 507576
rect 398502 507340 398586 507576
rect 398822 507340 398854 507576
rect 398234 471896 398854 507340
rect 398234 471660 398266 471896
rect 398502 471660 398586 471896
rect 398822 471660 398854 471896
rect 398234 471576 398854 471660
rect 398234 471340 398266 471576
rect 398502 471340 398586 471576
rect 398822 471340 398854 471576
rect 398234 435896 398854 471340
rect 398234 435660 398266 435896
rect 398502 435660 398586 435896
rect 398822 435660 398854 435896
rect 398234 435576 398854 435660
rect 398234 435340 398266 435576
rect 398502 435340 398586 435576
rect 398822 435340 398854 435576
rect 398234 399896 398854 435340
rect 398234 399660 398266 399896
rect 398502 399660 398586 399896
rect 398822 399660 398854 399896
rect 398234 399576 398854 399660
rect 398234 399340 398266 399576
rect 398502 399340 398586 399576
rect 398822 399340 398854 399576
rect 398234 363896 398854 399340
rect 398234 363660 398266 363896
rect 398502 363660 398586 363896
rect 398822 363660 398854 363896
rect 398234 363576 398854 363660
rect 398234 363340 398266 363576
rect 398502 363340 398586 363576
rect 398822 363340 398854 363576
rect 398234 327896 398854 363340
rect 398234 327660 398266 327896
rect 398502 327660 398586 327896
rect 398822 327660 398854 327896
rect 398234 327576 398854 327660
rect 398234 327340 398266 327576
rect 398502 327340 398586 327576
rect 398822 327340 398854 327576
rect 398234 291896 398854 327340
rect 398234 291660 398266 291896
rect 398502 291660 398586 291896
rect 398822 291660 398854 291896
rect 398234 291576 398854 291660
rect 398234 291340 398266 291576
rect 398502 291340 398586 291576
rect 398822 291340 398854 291576
rect 398234 255896 398854 291340
rect 398234 255660 398266 255896
rect 398502 255660 398586 255896
rect 398822 255660 398854 255896
rect 398234 255576 398854 255660
rect 398234 255340 398266 255576
rect 398502 255340 398586 255576
rect 398822 255340 398854 255576
rect 398234 219896 398854 255340
rect 398234 219660 398266 219896
rect 398502 219660 398586 219896
rect 398822 219660 398854 219896
rect 398234 219576 398854 219660
rect 398234 219340 398266 219576
rect 398502 219340 398586 219576
rect 398822 219340 398854 219576
rect 398234 183896 398854 219340
rect 398234 183660 398266 183896
rect 398502 183660 398586 183896
rect 398822 183660 398854 183896
rect 398234 183576 398854 183660
rect 398234 183340 398266 183576
rect 398502 183340 398586 183576
rect 398822 183340 398854 183576
rect 398234 147896 398854 183340
rect 398234 147660 398266 147896
rect 398502 147660 398586 147896
rect 398822 147660 398854 147896
rect 398234 147576 398854 147660
rect 398234 147340 398266 147576
rect 398502 147340 398586 147576
rect 398822 147340 398854 147576
rect 398234 111896 398854 147340
rect 398234 111660 398266 111896
rect 398502 111660 398586 111896
rect 398822 111660 398854 111896
rect 398234 111576 398854 111660
rect 398234 111340 398266 111576
rect 398502 111340 398586 111576
rect 398822 111340 398854 111576
rect 398234 75896 398854 111340
rect 398234 75660 398266 75896
rect 398502 75660 398586 75896
rect 398822 75660 398854 75896
rect 398234 75576 398854 75660
rect 398234 75340 398266 75576
rect 398502 75340 398586 75576
rect 398822 75340 398854 75576
rect 398234 39896 398854 75340
rect 398234 39660 398266 39896
rect 398502 39660 398586 39896
rect 398822 39660 398854 39896
rect 398234 39576 398854 39660
rect 398234 39340 398266 39576
rect 398502 39340 398586 39576
rect 398822 39340 398854 39576
rect 398234 3896 398854 39340
rect 398234 3660 398266 3896
rect 398502 3660 398586 3896
rect 398822 3660 398854 3896
rect 398234 3576 398854 3660
rect 398234 3340 398266 3576
rect 398502 3340 398586 3576
rect 398822 3340 398854 3576
rect 398234 -1304 398854 3340
rect 398234 -1540 398266 -1304
rect 398502 -1540 398586 -1304
rect 398822 -1540 398854 -1304
rect 398234 -1624 398854 -1540
rect 398234 -1860 398266 -1624
rect 398502 -1860 398586 -1624
rect 398822 -1860 398854 -1624
rect 398234 -7652 398854 -1860
rect 399474 706760 400094 711592
rect 399474 706524 399506 706760
rect 399742 706524 399826 706760
rect 400062 706524 400094 706760
rect 399474 706440 400094 706524
rect 399474 706204 399506 706440
rect 399742 706204 399826 706440
rect 400062 706204 400094 706440
rect 399474 689136 400094 706204
rect 399474 688900 399506 689136
rect 399742 688900 399826 689136
rect 400062 688900 400094 689136
rect 399474 688816 400094 688900
rect 399474 688580 399506 688816
rect 399742 688580 399826 688816
rect 400062 688580 400094 688816
rect 399474 653136 400094 688580
rect 399474 652900 399506 653136
rect 399742 652900 399826 653136
rect 400062 652900 400094 653136
rect 399474 652816 400094 652900
rect 399474 652580 399506 652816
rect 399742 652580 399826 652816
rect 400062 652580 400094 652816
rect 399474 617136 400094 652580
rect 399474 616900 399506 617136
rect 399742 616900 399826 617136
rect 400062 616900 400094 617136
rect 399474 616816 400094 616900
rect 399474 616580 399506 616816
rect 399742 616580 399826 616816
rect 400062 616580 400094 616816
rect 399474 581136 400094 616580
rect 399474 580900 399506 581136
rect 399742 580900 399826 581136
rect 400062 580900 400094 581136
rect 399474 580816 400094 580900
rect 399474 580580 399506 580816
rect 399742 580580 399826 580816
rect 400062 580580 400094 580816
rect 399474 545136 400094 580580
rect 399474 544900 399506 545136
rect 399742 544900 399826 545136
rect 400062 544900 400094 545136
rect 399474 544816 400094 544900
rect 399474 544580 399506 544816
rect 399742 544580 399826 544816
rect 400062 544580 400094 544816
rect 399474 509136 400094 544580
rect 399474 508900 399506 509136
rect 399742 508900 399826 509136
rect 400062 508900 400094 509136
rect 399474 508816 400094 508900
rect 399474 508580 399506 508816
rect 399742 508580 399826 508816
rect 400062 508580 400094 508816
rect 399474 473136 400094 508580
rect 399474 472900 399506 473136
rect 399742 472900 399826 473136
rect 400062 472900 400094 473136
rect 399474 472816 400094 472900
rect 399474 472580 399506 472816
rect 399742 472580 399826 472816
rect 400062 472580 400094 472816
rect 399474 437136 400094 472580
rect 399474 436900 399506 437136
rect 399742 436900 399826 437136
rect 400062 436900 400094 437136
rect 399474 436816 400094 436900
rect 399474 436580 399506 436816
rect 399742 436580 399826 436816
rect 400062 436580 400094 436816
rect 399474 401136 400094 436580
rect 399474 400900 399506 401136
rect 399742 400900 399826 401136
rect 400062 400900 400094 401136
rect 399474 400816 400094 400900
rect 399474 400580 399506 400816
rect 399742 400580 399826 400816
rect 400062 400580 400094 400816
rect 399474 365136 400094 400580
rect 399474 364900 399506 365136
rect 399742 364900 399826 365136
rect 400062 364900 400094 365136
rect 399474 364816 400094 364900
rect 399474 364580 399506 364816
rect 399742 364580 399826 364816
rect 400062 364580 400094 364816
rect 399474 329136 400094 364580
rect 399474 328900 399506 329136
rect 399742 328900 399826 329136
rect 400062 328900 400094 329136
rect 399474 328816 400094 328900
rect 399474 328580 399506 328816
rect 399742 328580 399826 328816
rect 400062 328580 400094 328816
rect 399474 293136 400094 328580
rect 399474 292900 399506 293136
rect 399742 292900 399826 293136
rect 400062 292900 400094 293136
rect 399474 292816 400094 292900
rect 399474 292580 399506 292816
rect 399742 292580 399826 292816
rect 400062 292580 400094 292816
rect 399474 257136 400094 292580
rect 399474 256900 399506 257136
rect 399742 256900 399826 257136
rect 400062 256900 400094 257136
rect 399474 256816 400094 256900
rect 399474 256580 399506 256816
rect 399742 256580 399826 256816
rect 400062 256580 400094 256816
rect 399474 221136 400094 256580
rect 399474 220900 399506 221136
rect 399742 220900 399826 221136
rect 400062 220900 400094 221136
rect 399474 220816 400094 220900
rect 399474 220580 399506 220816
rect 399742 220580 399826 220816
rect 400062 220580 400094 220816
rect 399474 185136 400094 220580
rect 399474 184900 399506 185136
rect 399742 184900 399826 185136
rect 400062 184900 400094 185136
rect 399474 184816 400094 184900
rect 399474 184580 399506 184816
rect 399742 184580 399826 184816
rect 400062 184580 400094 184816
rect 399474 149136 400094 184580
rect 399474 148900 399506 149136
rect 399742 148900 399826 149136
rect 400062 148900 400094 149136
rect 399474 148816 400094 148900
rect 399474 148580 399506 148816
rect 399742 148580 399826 148816
rect 400062 148580 400094 148816
rect 399474 113136 400094 148580
rect 399474 112900 399506 113136
rect 399742 112900 399826 113136
rect 400062 112900 400094 113136
rect 399474 112816 400094 112900
rect 399474 112580 399506 112816
rect 399742 112580 399826 112816
rect 400062 112580 400094 112816
rect 399474 77136 400094 112580
rect 399474 76900 399506 77136
rect 399742 76900 399826 77136
rect 400062 76900 400094 77136
rect 399474 76816 400094 76900
rect 399474 76580 399506 76816
rect 399742 76580 399826 76816
rect 400062 76580 400094 76816
rect 399474 41136 400094 76580
rect 399474 40900 399506 41136
rect 399742 40900 399826 41136
rect 400062 40900 400094 41136
rect 399474 40816 400094 40900
rect 399474 40580 399506 40816
rect 399742 40580 399826 40816
rect 400062 40580 400094 40816
rect 399474 5136 400094 40580
rect 399474 4900 399506 5136
rect 399742 4900 399826 5136
rect 400062 4900 400094 5136
rect 399474 4816 400094 4900
rect 399474 4580 399506 4816
rect 399742 4580 399826 4816
rect 400062 4580 400094 4816
rect 399474 -2264 400094 4580
rect 399474 -2500 399506 -2264
rect 399742 -2500 399826 -2264
rect 400062 -2500 400094 -2264
rect 399474 -2584 400094 -2500
rect 399474 -2820 399506 -2584
rect 399742 -2820 399826 -2584
rect 400062 -2820 400094 -2584
rect 399474 -7652 400094 -2820
rect 400714 707720 401334 711592
rect 400714 707484 400746 707720
rect 400982 707484 401066 707720
rect 401302 707484 401334 707720
rect 400714 707400 401334 707484
rect 400714 707164 400746 707400
rect 400982 707164 401066 707400
rect 401302 707164 401334 707400
rect 400714 690376 401334 707164
rect 400714 690140 400746 690376
rect 400982 690140 401066 690376
rect 401302 690140 401334 690376
rect 400714 690056 401334 690140
rect 400714 689820 400746 690056
rect 400982 689820 401066 690056
rect 401302 689820 401334 690056
rect 400714 654376 401334 689820
rect 400714 654140 400746 654376
rect 400982 654140 401066 654376
rect 401302 654140 401334 654376
rect 400714 654056 401334 654140
rect 400714 653820 400746 654056
rect 400982 653820 401066 654056
rect 401302 653820 401334 654056
rect 400714 618376 401334 653820
rect 400714 618140 400746 618376
rect 400982 618140 401066 618376
rect 401302 618140 401334 618376
rect 400714 618056 401334 618140
rect 400714 617820 400746 618056
rect 400982 617820 401066 618056
rect 401302 617820 401334 618056
rect 400714 582376 401334 617820
rect 400714 582140 400746 582376
rect 400982 582140 401066 582376
rect 401302 582140 401334 582376
rect 400714 582056 401334 582140
rect 400714 581820 400746 582056
rect 400982 581820 401066 582056
rect 401302 581820 401334 582056
rect 400714 546376 401334 581820
rect 400714 546140 400746 546376
rect 400982 546140 401066 546376
rect 401302 546140 401334 546376
rect 400714 546056 401334 546140
rect 400714 545820 400746 546056
rect 400982 545820 401066 546056
rect 401302 545820 401334 546056
rect 400714 510376 401334 545820
rect 400714 510140 400746 510376
rect 400982 510140 401066 510376
rect 401302 510140 401334 510376
rect 400714 510056 401334 510140
rect 400714 509820 400746 510056
rect 400982 509820 401066 510056
rect 401302 509820 401334 510056
rect 400714 474376 401334 509820
rect 400714 474140 400746 474376
rect 400982 474140 401066 474376
rect 401302 474140 401334 474376
rect 400714 474056 401334 474140
rect 400714 473820 400746 474056
rect 400982 473820 401066 474056
rect 401302 473820 401334 474056
rect 400714 438376 401334 473820
rect 400714 438140 400746 438376
rect 400982 438140 401066 438376
rect 401302 438140 401334 438376
rect 400714 438056 401334 438140
rect 400714 437820 400746 438056
rect 400982 437820 401066 438056
rect 401302 437820 401334 438056
rect 400714 402376 401334 437820
rect 400714 402140 400746 402376
rect 400982 402140 401066 402376
rect 401302 402140 401334 402376
rect 400714 402056 401334 402140
rect 400714 401820 400746 402056
rect 400982 401820 401066 402056
rect 401302 401820 401334 402056
rect 400714 366376 401334 401820
rect 400714 366140 400746 366376
rect 400982 366140 401066 366376
rect 401302 366140 401334 366376
rect 400714 366056 401334 366140
rect 400714 365820 400746 366056
rect 400982 365820 401066 366056
rect 401302 365820 401334 366056
rect 400714 330376 401334 365820
rect 400714 330140 400746 330376
rect 400982 330140 401066 330376
rect 401302 330140 401334 330376
rect 400714 330056 401334 330140
rect 400714 329820 400746 330056
rect 400982 329820 401066 330056
rect 401302 329820 401334 330056
rect 400714 294376 401334 329820
rect 400714 294140 400746 294376
rect 400982 294140 401066 294376
rect 401302 294140 401334 294376
rect 400714 294056 401334 294140
rect 400714 293820 400746 294056
rect 400982 293820 401066 294056
rect 401302 293820 401334 294056
rect 400714 258376 401334 293820
rect 400714 258140 400746 258376
rect 400982 258140 401066 258376
rect 401302 258140 401334 258376
rect 400714 258056 401334 258140
rect 400714 257820 400746 258056
rect 400982 257820 401066 258056
rect 401302 257820 401334 258056
rect 400714 222376 401334 257820
rect 400714 222140 400746 222376
rect 400982 222140 401066 222376
rect 401302 222140 401334 222376
rect 400714 222056 401334 222140
rect 400714 221820 400746 222056
rect 400982 221820 401066 222056
rect 401302 221820 401334 222056
rect 400714 186376 401334 221820
rect 400714 186140 400746 186376
rect 400982 186140 401066 186376
rect 401302 186140 401334 186376
rect 400714 186056 401334 186140
rect 400714 185820 400746 186056
rect 400982 185820 401066 186056
rect 401302 185820 401334 186056
rect 400714 150376 401334 185820
rect 400714 150140 400746 150376
rect 400982 150140 401066 150376
rect 401302 150140 401334 150376
rect 400714 150056 401334 150140
rect 400714 149820 400746 150056
rect 400982 149820 401066 150056
rect 401302 149820 401334 150056
rect 400714 114376 401334 149820
rect 400714 114140 400746 114376
rect 400982 114140 401066 114376
rect 401302 114140 401334 114376
rect 400714 114056 401334 114140
rect 400714 113820 400746 114056
rect 400982 113820 401066 114056
rect 401302 113820 401334 114056
rect 400714 78376 401334 113820
rect 400714 78140 400746 78376
rect 400982 78140 401066 78376
rect 401302 78140 401334 78376
rect 400714 78056 401334 78140
rect 400714 77820 400746 78056
rect 400982 77820 401066 78056
rect 401302 77820 401334 78056
rect 400714 42376 401334 77820
rect 400714 42140 400746 42376
rect 400982 42140 401066 42376
rect 401302 42140 401334 42376
rect 400714 42056 401334 42140
rect 400714 41820 400746 42056
rect 400982 41820 401066 42056
rect 401302 41820 401334 42056
rect 400714 6376 401334 41820
rect 400714 6140 400746 6376
rect 400982 6140 401066 6376
rect 401302 6140 401334 6376
rect 400714 6056 401334 6140
rect 400714 5820 400746 6056
rect 400982 5820 401066 6056
rect 401302 5820 401334 6056
rect 400714 -3224 401334 5820
rect 400714 -3460 400746 -3224
rect 400982 -3460 401066 -3224
rect 401302 -3460 401334 -3224
rect 400714 -3544 401334 -3460
rect 400714 -3780 400746 -3544
rect 400982 -3780 401066 -3544
rect 401302 -3780 401334 -3544
rect 400714 -7652 401334 -3780
rect 401954 708680 402574 711592
rect 401954 708444 401986 708680
rect 402222 708444 402306 708680
rect 402542 708444 402574 708680
rect 401954 708360 402574 708444
rect 401954 708124 401986 708360
rect 402222 708124 402306 708360
rect 402542 708124 402574 708360
rect 401954 691616 402574 708124
rect 401954 691380 401986 691616
rect 402222 691380 402306 691616
rect 402542 691380 402574 691616
rect 401954 691296 402574 691380
rect 401954 691060 401986 691296
rect 402222 691060 402306 691296
rect 402542 691060 402574 691296
rect 401954 655616 402574 691060
rect 401954 655380 401986 655616
rect 402222 655380 402306 655616
rect 402542 655380 402574 655616
rect 401954 655296 402574 655380
rect 401954 655060 401986 655296
rect 402222 655060 402306 655296
rect 402542 655060 402574 655296
rect 401954 619616 402574 655060
rect 401954 619380 401986 619616
rect 402222 619380 402306 619616
rect 402542 619380 402574 619616
rect 401954 619296 402574 619380
rect 401954 619060 401986 619296
rect 402222 619060 402306 619296
rect 402542 619060 402574 619296
rect 401954 583616 402574 619060
rect 401954 583380 401986 583616
rect 402222 583380 402306 583616
rect 402542 583380 402574 583616
rect 401954 583296 402574 583380
rect 401954 583060 401986 583296
rect 402222 583060 402306 583296
rect 402542 583060 402574 583296
rect 401954 547616 402574 583060
rect 401954 547380 401986 547616
rect 402222 547380 402306 547616
rect 402542 547380 402574 547616
rect 401954 547296 402574 547380
rect 401954 547060 401986 547296
rect 402222 547060 402306 547296
rect 402542 547060 402574 547296
rect 401954 511616 402574 547060
rect 401954 511380 401986 511616
rect 402222 511380 402306 511616
rect 402542 511380 402574 511616
rect 401954 511296 402574 511380
rect 401954 511060 401986 511296
rect 402222 511060 402306 511296
rect 402542 511060 402574 511296
rect 401954 475616 402574 511060
rect 401954 475380 401986 475616
rect 402222 475380 402306 475616
rect 402542 475380 402574 475616
rect 401954 475296 402574 475380
rect 401954 475060 401986 475296
rect 402222 475060 402306 475296
rect 402542 475060 402574 475296
rect 401954 439616 402574 475060
rect 401954 439380 401986 439616
rect 402222 439380 402306 439616
rect 402542 439380 402574 439616
rect 401954 439296 402574 439380
rect 401954 439060 401986 439296
rect 402222 439060 402306 439296
rect 402542 439060 402574 439296
rect 401954 403616 402574 439060
rect 401954 403380 401986 403616
rect 402222 403380 402306 403616
rect 402542 403380 402574 403616
rect 401954 403296 402574 403380
rect 401954 403060 401986 403296
rect 402222 403060 402306 403296
rect 402542 403060 402574 403296
rect 401954 367616 402574 403060
rect 401954 367380 401986 367616
rect 402222 367380 402306 367616
rect 402542 367380 402574 367616
rect 401954 367296 402574 367380
rect 401954 367060 401986 367296
rect 402222 367060 402306 367296
rect 402542 367060 402574 367296
rect 401954 331616 402574 367060
rect 401954 331380 401986 331616
rect 402222 331380 402306 331616
rect 402542 331380 402574 331616
rect 401954 331296 402574 331380
rect 401954 331060 401986 331296
rect 402222 331060 402306 331296
rect 402542 331060 402574 331296
rect 401954 295616 402574 331060
rect 401954 295380 401986 295616
rect 402222 295380 402306 295616
rect 402542 295380 402574 295616
rect 401954 295296 402574 295380
rect 401954 295060 401986 295296
rect 402222 295060 402306 295296
rect 402542 295060 402574 295296
rect 401954 259616 402574 295060
rect 401954 259380 401986 259616
rect 402222 259380 402306 259616
rect 402542 259380 402574 259616
rect 401954 259296 402574 259380
rect 401954 259060 401986 259296
rect 402222 259060 402306 259296
rect 402542 259060 402574 259296
rect 401954 223616 402574 259060
rect 401954 223380 401986 223616
rect 402222 223380 402306 223616
rect 402542 223380 402574 223616
rect 401954 223296 402574 223380
rect 401954 223060 401986 223296
rect 402222 223060 402306 223296
rect 402542 223060 402574 223296
rect 401954 187616 402574 223060
rect 401954 187380 401986 187616
rect 402222 187380 402306 187616
rect 402542 187380 402574 187616
rect 401954 187296 402574 187380
rect 401954 187060 401986 187296
rect 402222 187060 402306 187296
rect 402542 187060 402574 187296
rect 401954 151616 402574 187060
rect 401954 151380 401986 151616
rect 402222 151380 402306 151616
rect 402542 151380 402574 151616
rect 401954 151296 402574 151380
rect 401954 151060 401986 151296
rect 402222 151060 402306 151296
rect 402542 151060 402574 151296
rect 401954 115616 402574 151060
rect 401954 115380 401986 115616
rect 402222 115380 402306 115616
rect 402542 115380 402574 115616
rect 401954 115296 402574 115380
rect 401954 115060 401986 115296
rect 402222 115060 402306 115296
rect 402542 115060 402574 115296
rect 401954 79616 402574 115060
rect 401954 79380 401986 79616
rect 402222 79380 402306 79616
rect 402542 79380 402574 79616
rect 401954 79296 402574 79380
rect 401954 79060 401986 79296
rect 402222 79060 402306 79296
rect 402542 79060 402574 79296
rect 401954 43616 402574 79060
rect 401954 43380 401986 43616
rect 402222 43380 402306 43616
rect 402542 43380 402574 43616
rect 401954 43296 402574 43380
rect 401954 43060 401986 43296
rect 402222 43060 402306 43296
rect 402542 43060 402574 43296
rect 401954 7616 402574 43060
rect 401954 7380 401986 7616
rect 402222 7380 402306 7616
rect 402542 7380 402574 7616
rect 401954 7296 402574 7380
rect 401954 7060 401986 7296
rect 402222 7060 402306 7296
rect 402542 7060 402574 7296
rect 401954 -4184 402574 7060
rect 401954 -4420 401986 -4184
rect 402222 -4420 402306 -4184
rect 402542 -4420 402574 -4184
rect 401954 -4504 402574 -4420
rect 401954 -4740 401986 -4504
rect 402222 -4740 402306 -4504
rect 402542 -4740 402574 -4504
rect 401954 -7652 402574 -4740
rect 403194 709640 403814 711592
rect 403194 709404 403226 709640
rect 403462 709404 403546 709640
rect 403782 709404 403814 709640
rect 403194 709320 403814 709404
rect 403194 709084 403226 709320
rect 403462 709084 403546 709320
rect 403782 709084 403814 709320
rect 403194 692856 403814 709084
rect 403194 692620 403226 692856
rect 403462 692620 403546 692856
rect 403782 692620 403814 692856
rect 403194 692536 403814 692620
rect 403194 692300 403226 692536
rect 403462 692300 403546 692536
rect 403782 692300 403814 692536
rect 403194 656856 403814 692300
rect 403194 656620 403226 656856
rect 403462 656620 403546 656856
rect 403782 656620 403814 656856
rect 403194 656536 403814 656620
rect 403194 656300 403226 656536
rect 403462 656300 403546 656536
rect 403782 656300 403814 656536
rect 403194 620856 403814 656300
rect 403194 620620 403226 620856
rect 403462 620620 403546 620856
rect 403782 620620 403814 620856
rect 403194 620536 403814 620620
rect 403194 620300 403226 620536
rect 403462 620300 403546 620536
rect 403782 620300 403814 620536
rect 403194 584856 403814 620300
rect 403194 584620 403226 584856
rect 403462 584620 403546 584856
rect 403782 584620 403814 584856
rect 403194 584536 403814 584620
rect 403194 584300 403226 584536
rect 403462 584300 403546 584536
rect 403782 584300 403814 584536
rect 403194 548856 403814 584300
rect 403194 548620 403226 548856
rect 403462 548620 403546 548856
rect 403782 548620 403814 548856
rect 403194 548536 403814 548620
rect 403194 548300 403226 548536
rect 403462 548300 403546 548536
rect 403782 548300 403814 548536
rect 403194 512856 403814 548300
rect 403194 512620 403226 512856
rect 403462 512620 403546 512856
rect 403782 512620 403814 512856
rect 403194 512536 403814 512620
rect 403194 512300 403226 512536
rect 403462 512300 403546 512536
rect 403782 512300 403814 512536
rect 403194 476856 403814 512300
rect 403194 476620 403226 476856
rect 403462 476620 403546 476856
rect 403782 476620 403814 476856
rect 403194 476536 403814 476620
rect 403194 476300 403226 476536
rect 403462 476300 403546 476536
rect 403782 476300 403814 476536
rect 403194 440856 403814 476300
rect 403194 440620 403226 440856
rect 403462 440620 403546 440856
rect 403782 440620 403814 440856
rect 403194 440536 403814 440620
rect 403194 440300 403226 440536
rect 403462 440300 403546 440536
rect 403782 440300 403814 440536
rect 403194 404856 403814 440300
rect 403194 404620 403226 404856
rect 403462 404620 403546 404856
rect 403782 404620 403814 404856
rect 403194 404536 403814 404620
rect 403194 404300 403226 404536
rect 403462 404300 403546 404536
rect 403782 404300 403814 404536
rect 403194 368856 403814 404300
rect 403194 368620 403226 368856
rect 403462 368620 403546 368856
rect 403782 368620 403814 368856
rect 403194 368536 403814 368620
rect 403194 368300 403226 368536
rect 403462 368300 403546 368536
rect 403782 368300 403814 368536
rect 403194 332856 403814 368300
rect 403194 332620 403226 332856
rect 403462 332620 403546 332856
rect 403782 332620 403814 332856
rect 403194 332536 403814 332620
rect 403194 332300 403226 332536
rect 403462 332300 403546 332536
rect 403782 332300 403814 332536
rect 403194 296856 403814 332300
rect 403194 296620 403226 296856
rect 403462 296620 403546 296856
rect 403782 296620 403814 296856
rect 403194 296536 403814 296620
rect 403194 296300 403226 296536
rect 403462 296300 403546 296536
rect 403782 296300 403814 296536
rect 403194 260856 403814 296300
rect 403194 260620 403226 260856
rect 403462 260620 403546 260856
rect 403782 260620 403814 260856
rect 403194 260536 403814 260620
rect 403194 260300 403226 260536
rect 403462 260300 403546 260536
rect 403782 260300 403814 260536
rect 403194 224856 403814 260300
rect 403194 224620 403226 224856
rect 403462 224620 403546 224856
rect 403782 224620 403814 224856
rect 403194 224536 403814 224620
rect 403194 224300 403226 224536
rect 403462 224300 403546 224536
rect 403782 224300 403814 224536
rect 403194 188856 403814 224300
rect 403194 188620 403226 188856
rect 403462 188620 403546 188856
rect 403782 188620 403814 188856
rect 403194 188536 403814 188620
rect 403194 188300 403226 188536
rect 403462 188300 403546 188536
rect 403782 188300 403814 188536
rect 403194 152856 403814 188300
rect 403194 152620 403226 152856
rect 403462 152620 403546 152856
rect 403782 152620 403814 152856
rect 403194 152536 403814 152620
rect 403194 152300 403226 152536
rect 403462 152300 403546 152536
rect 403782 152300 403814 152536
rect 403194 116856 403814 152300
rect 403194 116620 403226 116856
rect 403462 116620 403546 116856
rect 403782 116620 403814 116856
rect 403194 116536 403814 116620
rect 403194 116300 403226 116536
rect 403462 116300 403546 116536
rect 403782 116300 403814 116536
rect 403194 80856 403814 116300
rect 403194 80620 403226 80856
rect 403462 80620 403546 80856
rect 403782 80620 403814 80856
rect 403194 80536 403814 80620
rect 403194 80300 403226 80536
rect 403462 80300 403546 80536
rect 403782 80300 403814 80536
rect 403194 44856 403814 80300
rect 403194 44620 403226 44856
rect 403462 44620 403546 44856
rect 403782 44620 403814 44856
rect 403194 44536 403814 44620
rect 403194 44300 403226 44536
rect 403462 44300 403546 44536
rect 403782 44300 403814 44536
rect 403194 8856 403814 44300
rect 403194 8620 403226 8856
rect 403462 8620 403546 8856
rect 403782 8620 403814 8856
rect 403194 8536 403814 8620
rect 403194 8300 403226 8536
rect 403462 8300 403546 8536
rect 403782 8300 403814 8536
rect 403194 -5144 403814 8300
rect 403194 -5380 403226 -5144
rect 403462 -5380 403546 -5144
rect 403782 -5380 403814 -5144
rect 403194 -5464 403814 -5380
rect 403194 -5700 403226 -5464
rect 403462 -5700 403546 -5464
rect 403782 -5700 403814 -5464
rect 403194 -7652 403814 -5700
rect 404434 710600 405054 711592
rect 404434 710364 404466 710600
rect 404702 710364 404786 710600
rect 405022 710364 405054 710600
rect 404434 710280 405054 710364
rect 404434 710044 404466 710280
rect 404702 710044 404786 710280
rect 405022 710044 405054 710280
rect 404434 694096 405054 710044
rect 404434 693860 404466 694096
rect 404702 693860 404786 694096
rect 405022 693860 405054 694096
rect 404434 693776 405054 693860
rect 404434 693540 404466 693776
rect 404702 693540 404786 693776
rect 405022 693540 405054 693776
rect 404434 658096 405054 693540
rect 404434 657860 404466 658096
rect 404702 657860 404786 658096
rect 405022 657860 405054 658096
rect 404434 657776 405054 657860
rect 404434 657540 404466 657776
rect 404702 657540 404786 657776
rect 405022 657540 405054 657776
rect 404434 622096 405054 657540
rect 404434 621860 404466 622096
rect 404702 621860 404786 622096
rect 405022 621860 405054 622096
rect 404434 621776 405054 621860
rect 404434 621540 404466 621776
rect 404702 621540 404786 621776
rect 405022 621540 405054 621776
rect 404434 586096 405054 621540
rect 404434 585860 404466 586096
rect 404702 585860 404786 586096
rect 405022 585860 405054 586096
rect 404434 585776 405054 585860
rect 404434 585540 404466 585776
rect 404702 585540 404786 585776
rect 405022 585540 405054 585776
rect 404434 550096 405054 585540
rect 404434 549860 404466 550096
rect 404702 549860 404786 550096
rect 405022 549860 405054 550096
rect 404434 549776 405054 549860
rect 404434 549540 404466 549776
rect 404702 549540 404786 549776
rect 405022 549540 405054 549776
rect 404434 514096 405054 549540
rect 404434 513860 404466 514096
rect 404702 513860 404786 514096
rect 405022 513860 405054 514096
rect 404434 513776 405054 513860
rect 404434 513540 404466 513776
rect 404702 513540 404786 513776
rect 405022 513540 405054 513776
rect 404434 478096 405054 513540
rect 404434 477860 404466 478096
rect 404702 477860 404786 478096
rect 405022 477860 405054 478096
rect 404434 477776 405054 477860
rect 404434 477540 404466 477776
rect 404702 477540 404786 477776
rect 405022 477540 405054 477776
rect 404434 442096 405054 477540
rect 404434 441860 404466 442096
rect 404702 441860 404786 442096
rect 405022 441860 405054 442096
rect 404434 441776 405054 441860
rect 404434 441540 404466 441776
rect 404702 441540 404786 441776
rect 405022 441540 405054 441776
rect 404434 406096 405054 441540
rect 404434 405860 404466 406096
rect 404702 405860 404786 406096
rect 405022 405860 405054 406096
rect 404434 405776 405054 405860
rect 404434 405540 404466 405776
rect 404702 405540 404786 405776
rect 405022 405540 405054 405776
rect 404434 370096 405054 405540
rect 404434 369860 404466 370096
rect 404702 369860 404786 370096
rect 405022 369860 405054 370096
rect 404434 369776 405054 369860
rect 404434 369540 404466 369776
rect 404702 369540 404786 369776
rect 405022 369540 405054 369776
rect 404434 334096 405054 369540
rect 404434 333860 404466 334096
rect 404702 333860 404786 334096
rect 405022 333860 405054 334096
rect 404434 333776 405054 333860
rect 404434 333540 404466 333776
rect 404702 333540 404786 333776
rect 405022 333540 405054 333776
rect 404434 298096 405054 333540
rect 404434 297860 404466 298096
rect 404702 297860 404786 298096
rect 405022 297860 405054 298096
rect 404434 297776 405054 297860
rect 404434 297540 404466 297776
rect 404702 297540 404786 297776
rect 405022 297540 405054 297776
rect 404434 262096 405054 297540
rect 404434 261860 404466 262096
rect 404702 261860 404786 262096
rect 405022 261860 405054 262096
rect 404434 261776 405054 261860
rect 404434 261540 404466 261776
rect 404702 261540 404786 261776
rect 405022 261540 405054 261776
rect 404434 226096 405054 261540
rect 404434 225860 404466 226096
rect 404702 225860 404786 226096
rect 405022 225860 405054 226096
rect 404434 225776 405054 225860
rect 404434 225540 404466 225776
rect 404702 225540 404786 225776
rect 405022 225540 405054 225776
rect 404434 190096 405054 225540
rect 404434 189860 404466 190096
rect 404702 189860 404786 190096
rect 405022 189860 405054 190096
rect 404434 189776 405054 189860
rect 404434 189540 404466 189776
rect 404702 189540 404786 189776
rect 405022 189540 405054 189776
rect 404434 154096 405054 189540
rect 404434 153860 404466 154096
rect 404702 153860 404786 154096
rect 405022 153860 405054 154096
rect 404434 153776 405054 153860
rect 404434 153540 404466 153776
rect 404702 153540 404786 153776
rect 405022 153540 405054 153776
rect 404434 118096 405054 153540
rect 404434 117860 404466 118096
rect 404702 117860 404786 118096
rect 405022 117860 405054 118096
rect 404434 117776 405054 117860
rect 404434 117540 404466 117776
rect 404702 117540 404786 117776
rect 405022 117540 405054 117776
rect 404434 82096 405054 117540
rect 404434 81860 404466 82096
rect 404702 81860 404786 82096
rect 405022 81860 405054 82096
rect 404434 81776 405054 81860
rect 404434 81540 404466 81776
rect 404702 81540 404786 81776
rect 405022 81540 405054 81776
rect 404434 46096 405054 81540
rect 404434 45860 404466 46096
rect 404702 45860 404786 46096
rect 405022 45860 405054 46096
rect 404434 45776 405054 45860
rect 404434 45540 404466 45776
rect 404702 45540 404786 45776
rect 405022 45540 405054 45776
rect 404434 10096 405054 45540
rect 404434 9860 404466 10096
rect 404702 9860 404786 10096
rect 405022 9860 405054 10096
rect 404434 9776 405054 9860
rect 404434 9540 404466 9776
rect 404702 9540 404786 9776
rect 405022 9540 405054 9776
rect 404434 -6104 405054 9540
rect 404434 -6340 404466 -6104
rect 404702 -6340 404786 -6104
rect 405022 -6340 405054 -6104
rect 404434 -6424 405054 -6340
rect 404434 -6660 404466 -6424
rect 404702 -6660 404786 -6424
rect 405022 -6660 405054 -6424
rect 404434 -7652 405054 -6660
rect 405674 711560 406294 711592
rect 405674 711324 405706 711560
rect 405942 711324 406026 711560
rect 406262 711324 406294 711560
rect 405674 711240 406294 711324
rect 405674 711004 405706 711240
rect 405942 711004 406026 711240
rect 406262 711004 406294 711240
rect 405674 695336 406294 711004
rect 405674 695100 405706 695336
rect 405942 695100 406026 695336
rect 406262 695100 406294 695336
rect 405674 695016 406294 695100
rect 405674 694780 405706 695016
rect 405942 694780 406026 695016
rect 406262 694780 406294 695016
rect 405674 659336 406294 694780
rect 405674 659100 405706 659336
rect 405942 659100 406026 659336
rect 406262 659100 406294 659336
rect 405674 659016 406294 659100
rect 405674 658780 405706 659016
rect 405942 658780 406026 659016
rect 406262 658780 406294 659016
rect 405674 623336 406294 658780
rect 405674 623100 405706 623336
rect 405942 623100 406026 623336
rect 406262 623100 406294 623336
rect 405674 623016 406294 623100
rect 405674 622780 405706 623016
rect 405942 622780 406026 623016
rect 406262 622780 406294 623016
rect 405674 587336 406294 622780
rect 405674 587100 405706 587336
rect 405942 587100 406026 587336
rect 406262 587100 406294 587336
rect 405674 587016 406294 587100
rect 405674 586780 405706 587016
rect 405942 586780 406026 587016
rect 406262 586780 406294 587016
rect 405674 551336 406294 586780
rect 405674 551100 405706 551336
rect 405942 551100 406026 551336
rect 406262 551100 406294 551336
rect 405674 551016 406294 551100
rect 405674 550780 405706 551016
rect 405942 550780 406026 551016
rect 406262 550780 406294 551016
rect 405674 515336 406294 550780
rect 405674 515100 405706 515336
rect 405942 515100 406026 515336
rect 406262 515100 406294 515336
rect 405674 515016 406294 515100
rect 405674 514780 405706 515016
rect 405942 514780 406026 515016
rect 406262 514780 406294 515016
rect 405674 479336 406294 514780
rect 405674 479100 405706 479336
rect 405942 479100 406026 479336
rect 406262 479100 406294 479336
rect 405674 479016 406294 479100
rect 405674 478780 405706 479016
rect 405942 478780 406026 479016
rect 406262 478780 406294 479016
rect 405674 443336 406294 478780
rect 405674 443100 405706 443336
rect 405942 443100 406026 443336
rect 406262 443100 406294 443336
rect 405674 443016 406294 443100
rect 405674 442780 405706 443016
rect 405942 442780 406026 443016
rect 406262 442780 406294 443016
rect 405674 407336 406294 442780
rect 405674 407100 405706 407336
rect 405942 407100 406026 407336
rect 406262 407100 406294 407336
rect 405674 407016 406294 407100
rect 405674 406780 405706 407016
rect 405942 406780 406026 407016
rect 406262 406780 406294 407016
rect 405674 371336 406294 406780
rect 405674 371100 405706 371336
rect 405942 371100 406026 371336
rect 406262 371100 406294 371336
rect 405674 371016 406294 371100
rect 405674 370780 405706 371016
rect 405942 370780 406026 371016
rect 406262 370780 406294 371016
rect 405674 335336 406294 370780
rect 405674 335100 405706 335336
rect 405942 335100 406026 335336
rect 406262 335100 406294 335336
rect 405674 335016 406294 335100
rect 405674 334780 405706 335016
rect 405942 334780 406026 335016
rect 406262 334780 406294 335016
rect 405674 299336 406294 334780
rect 405674 299100 405706 299336
rect 405942 299100 406026 299336
rect 406262 299100 406294 299336
rect 405674 299016 406294 299100
rect 405674 298780 405706 299016
rect 405942 298780 406026 299016
rect 406262 298780 406294 299016
rect 405674 263336 406294 298780
rect 405674 263100 405706 263336
rect 405942 263100 406026 263336
rect 406262 263100 406294 263336
rect 405674 263016 406294 263100
rect 405674 262780 405706 263016
rect 405942 262780 406026 263016
rect 406262 262780 406294 263016
rect 405674 227336 406294 262780
rect 405674 227100 405706 227336
rect 405942 227100 406026 227336
rect 406262 227100 406294 227336
rect 405674 227016 406294 227100
rect 405674 226780 405706 227016
rect 405942 226780 406026 227016
rect 406262 226780 406294 227016
rect 405674 191336 406294 226780
rect 405674 191100 405706 191336
rect 405942 191100 406026 191336
rect 406262 191100 406294 191336
rect 405674 191016 406294 191100
rect 405674 190780 405706 191016
rect 405942 190780 406026 191016
rect 406262 190780 406294 191016
rect 405674 155336 406294 190780
rect 405674 155100 405706 155336
rect 405942 155100 406026 155336
rect 406262 155100 406294 155336
rect 405674 155016 406294 155100
rect 405674 154780 405706 155016
rect 405942 154780 406026 155016
rect 406262 154780 406294 155016
rect 405674 119336 406294 154780
rect 405674 119100 405706 119336
rect 405942 119100 406026 119336
rect 406262 119100 406294 119336
rect 405674 119016 406294 119100
rect 405674 118780 405706 119016
rect 405942 118780 406026 119016
rect 406262 118780 406294 119016
rect 405674 83336 406294 118780
rect 405674 83100 405706 83336
rect 405942 83100 406026 83336
rect 406262 83100 406294 83336
rect 405674 83016 406294 83100
rect 405674 82780 405706 83016
rect 405942 82780 406026 83016
rect 406262 82780 406294 83016
rect 405674 47336 406294 82780
rect 405674 47100 405706 47336
rect 405942 47100 406026 47336
rect 406262 47100 406294 47336
rect 405674 47016 406294 47100
rect 405674 46780 405706 47016
rect 405942 46780 406026 47016
rect 406262 46780 406294 47016
rect 405674 11336 406294 46780
rect 405674 11100 405706 11336
rect 405942 11100 406026 11336
rect 406262 11100 406294 11336
rect 405674 11016 406294 11100
rect 405674 10780 405706 11016
rect 405942 10780 406026 11016
rect 406262 10780 406294 11016
rect 405674 -7064 406294 10780
rect 405674 -7300 405706 -7064
rect 405942 -7300 406026 -7064
rect 406262 -7300 406294 -7064
rect 405674 -7384 406294 -7300
rect 405674 -7620 405706 -7384
rect 405942 -7620 406026 -7384
rect 406262 -7620 406294 -7384
rect 405674 -7652 406294 -7620
rect 432994 704840 433614 711592
rect 432994 704604 433026 704840
rect 433262 704604 433346 704840
rect 433582 704604 433614 704840
rect 432994 704520 433614 704604
rect 432994 704284 433026 704520
rect 433262 704284 433346 704520
rect 433582 704284 433614 704520
rect 432994 702002 433614 704284
rect 432994 701938 433032 702002
rect 433096 701938 433112 702002
rect 433176 701938 433192 702002
rect 433256 701938 433272 702002
rect 433336 701938 433352 702002
rect 433416 701938 433432 702002
rect 433496 701938 433512 702002
rect 433576 701938 433614 702002
rect 432994 701922 433614 701938
rect 432994 701858 433032 701922
rect 433096 701858 433112 701922
rect 433176 701858 433192 701922
rect 433256 701858 433272 701922
rect 433336 701858 433352 701922
rect 433416 701858 433432 701922
rect 433496 701858 433512 701922
rect 433576 701858 433614 701922
rect 432994 701842 433614 701858
rect 432994 701778 433032 701842
rect 433096 701778 433112 701842
rect 433176 701778 433192 701842
rect 433256 701778 433272 701842
rect 433336 701778 433352 701842
rect 433416 701778 433432 701842
rect 433496 701778 433512 701842
rect 433576 701778 433614 701842
rect 432994 701762 433614 701778
rect 432994 701698 433032 701762
rect 433096 701698 433112 701762
rect 433176 701698 433192 701762
rect 433256 701698 433272 701762
rect 433336 701698 433352 701762
rect 433416 701698 433432 701762
rect 433496 701698 433512 701762
rect 433576 701698 433614 701762
rect 432994 686656 433614 701698
rect 432994 686420 433026 686656
rect 433262 686420 433346 686656
rect 433582 686420 433614 686656
rect 432994 686336 433614 686420
rect 432994 686100 433026 686336
rect 433262 686100 433346 686336
rect 433582 686100 433614 686336
rect 432994 650656 433614 686100
rect 432994 650420 433026 650656
rect 433262 650420 433346 650656
rect 433582 650420 433614 650656
rect 432994 650336 433614 650420
rect 432994 650100 433026 650336
rect 433262 650100 433346 650336
rect 433582 650100 433614 650336
rect 432994 614656 433614 650100
rect 432994 614420 433026 614656
rect 433262 614420 433346 614656
rect 433582 614420 433614 614656
rect 432994 614336 433614 614420
rect 432994 614100 433026 614336
rect 433262 614100 433346 614336
rect 433582 614100 433614 614336
rect 432994 578656 433614 614100
rect 432994 578420 433026 578656
rect 433262 578420 433346 578656
rect 433582 578420 433614 578656
rect 432994 578336 433614 578420
rect 432994 578100 433026 578336
rect 433262 578100 433346 578336
rect 433582 578100 433614 578336
rect 432994 542656 433614 578100
rect 432994 542420 433026 542656
rect 433262 542420 433346 542656
rect 433582 542420 433614 542656
rect 432994 542336 433614 542420
rect 432994 542100 433026 542336
rect 433262 542100 433346 542336
rect 433582 542100 433614 542336
rect 432994 506656 433614 542100
rect 432994 506420 433026 506656
rect 433262 506420 433346 506656
rect 433582 506420 433614 506656
rect 432994 506336 433614 506420
rect 432994 506100 433026 506336
rect 433262 506100 433346 506336
rect 433582 506100 433614 506336
rect 432994 470656 433614 506100
rect 432994 470420 433026 470656
rect 433262 470420 433346 470656
rect 433582 470420 433614 470656
rect 432994 470336 433614 470420
rect 432994 470100 433026 470336
rect 433262 470100 433346 470336
rect 433582 470100 433614 470336
rect 432994 434656 433614 470100
rect 432994 434420 433026 434656
rect 433262 434420 433346 434656
rect 433582 434420 433614 434656
rect 432994 434336 433614 434420
rect 432994 434100 433026 434336
rect 433262 434100 433346 434336
rect 433582 434100 433614 434336
rect 432994 398656 433614 434100
rect 432994 398420 433026 398656
rect 433262 398420 433346 398656
rect 433582 398420 433614 398656
rect 432994 398336 433614 398420
rect 432994 398100 433026 398336
rect 433262 398100 433346 398336
rect 433582 398100 433614 398336
rect 432994 362656 433614 398100
rect 432994 362420 433026 362656
rect 433262 362420 433346 362656
rect 433582 362420 433614 362656
rect 432994 362336 433614 362420
rect 432994 362100 433026 362336
rect 433262 362100 433346 362336
rect 433582 362100 433614 362336
rect 432994 326656 433614 362100
rect 432994 326420 433026 326656
rect 433262 326420 433346 326656
rect 433582 326420 433614 326656
rect 432994 326336 433614 326420
rect 432994 326100 433026 326336
rect 433262 326100 433346 326336
rect 433582 326100 433614 326336
rect 432994 290656 433614 326100
rect 432994 290420 433026 290656
rect 433262 290420 433346 290656
rect 433582 290420 433614 290656
rect 432994 290336 433614 290420
rect 432994 290100 433026 290336
rect 433262 290100 433346 290336
rect 433582 290100 433614 290336
rect 432994 254656 433614 290100
rect 432994 254420 433026 254656
rect 433262 254420 433346 254656
rect 433582 254420 433614 254656
rect 432994 254336 433614 254420
rect 432994 254100 433026 254336
rect 433262 254100 433346 254336
rect 433582 254100 433614 254336
rect 432994 218656 433614 254100
rect 432994 218420 433026 218656
rect 433262 218420 433346 218656
rect 433582 218420 433614 218656
rect 432994 218336 433614 218420
rect 432994 218100 433026 218336
rect 433262 218100 433346 218336
rect 433582 218100 433614 218336
rect 432994 182656 433614 218100
rect 432994 182420 433026 182656
rect 433262 182420 433346 182656
rect 433582 182420 433614 182656
rect 432994 182336 433614 182420
rect 432994 182100 433026 182336
rect 433262 182100 433346 182336
rect 433582 182100 433614 182336
rect 432994 146656 433614 182100
rect 432994 146420 433026 146656
rect 433262 146420 433346 146656
rect 433582 146420 433614 146656
rect 432994 146336 433614 146420
rect 432994 146100 433026 146336
rect 433262 146100 433346 146336
rect 433582 146100 433614 146336
rect 432994 110656 433614 146100
rect 432994 110420 433026 110656
rect 433262 110420 433346 110656
rect 433582 110420 433614 110656
rect 432994 110336 433614 110420
rect 432994 110100 433026 110336
rect 433262 110100 433346 110336
rect 433582 110100 433614 110336
rect 432994 74656 433614 110100
rect 432994 74420 433026 74656
rect 433262 74420 433346 74656
rect 433582 74420 433614 74656
rect 432994 74336 433614 74420
rect 432994 74100 433026 74336
rect 433262 74100 433346 74336
rect 433582 74100 433614 74336
rect 432994 38656 433614 74100
rect 432994 38420 433026 38656
rect 433262 38420 433346 38656
rect 433582 38420 433614 38656
rect 432994 38336 433614 38420
rect 432994 38100 433026 38336
rect 433262 38100 433346 38336
rect 433582 38100 433614 38336
rect 432994 2656 433614 38100
rect 432994 2420 433026 2656
rect 433262 2420 433346 2656
rect 433582 2420 433614 2656
rect 432994 2336 433614 2420
rect 432994 2100 433026 2336
rect 433262 2100 433346 2336
rect 433582 2100 433614 2336
rect 432994 -344 433614 2100
rect 432994 -580 433026 -344
rect 433262 -580 433346 -344
rect 433582 -580 433614 -344
rect 432994 -664 433614 -580
rect 432994 -900 433026 -664
rect 433262 -900 433346 -664
rect 433582 -900 433614 -664
rect 432994 -7652 433614 -900
rect 434234 705800 434854 711592
rect 434234 705564 434266 705800
rect 434502 705564 434586 705800
rect 434822 705564 434854 705800
rect 434234 705480 434854 705564
rect 434234 705244 434266 705480
rect 434502 705244 434586 705480
rect 434822 705244 434854 705480
rect 434234 702770 434854 705244
rect 434234 702706 434272 702770
rect 434336 702706 434352 702770
rect 434416 702706 434432 702770
rect 434496 702706 434512 702770
rect 434576 702706 434592 702770
rect 434656 702706 434672 702770
rect 434736 702706 434752 702770
rect 434816 702706 434854 702770
rect 434234 702690 434854 702706
rect 434234 702626 434272 702690
rect 434336 702626 434352 702690
rect 434416 702626 434432 702690
rect 434496 702626 434512 702690
rect 434576 702626 434592 702690
rect 434656 702626 434672 702690
rect 434736 702626 434752 702690
rect 434816 702626 434854 702690
rect 434234 702610 434854 702626
rect 434234 702546 434272 702610
rect 434336 702546 434352 702610
rect 434416 702546 434432 702610
rect 434496 702546 434512 702610
rect 434576 702546 434592 702610
rect 434656 702546 434672 702610
rect 434736 702546 434752 702610
rect 434816 702546 434854 702610
rect 434234 702530 434854 702546
rect 434234 702466 434272 702530
rect 434336 702466 434352 702530
rect 434416 702466 434432 702530
rect 434496 702466 434512 702530
rect 434576 702466 434592 702530
rect 434656 702466 434672 702530
rect 434736 702466 434752 702530
rect 434816 702466 434854 702530
rect 434234 687896 434854 702466
rect 434234 687660 434266 687896
rect 434502 687660 434586 687896
rect 434822 687660 434854 687896
rect 434234 687576 434854 687660
rect 434234 687340 434266 687576
rect 434502 687340 434586 687576
rect 434822 687340 434854 687576
rect 434234 651896 434854 687340
rect 434234 651660 434266 651896
rect 434502 651660 434586 651896
rect 434822 651660 434854 651896
rect 434234 651576 434854 651660
rect 434234 651340 434266 651576
rect 434502 651340 434586 651576
rect 434822 651340 434854 651576
rect 434234 615896 434854 651340
rect 434234 615660 434266 615896
rect 434502 615660 434586 615896
rect 434822 615660 434854 615896
rect 434234 615576 434854 615660
rect 434234 615340 434266 615576
rect 434502 615340 434586 615576
rect 434822 615340 434854 615576
rect 434234 579896 434854 615340
rect 434234 579660 434266 579896
rect 434502 579660 434586 579896
rect 434822 579660 434854 579896
rect 434234 579576 434854 579660
rect 434234 579340 434266 579576
rect 434502 579340 434586 579576
rect 434822 579340 434854 579576
rect 434234 543896 434854 579340
rect 434234 543660 434266 543896
rect 434502 543660 434586 543896
rect 434822 543660 434854 543896
rect 434234 543576 434854 543660
rect 434234 543340 434266 543576
rect 434502 543340 434586 543576
rect 434822 543340 434854 543576
rect 434234 507896 434854 543340
rect 434234 507660 434266 507896
rect 434502 507660 434586 507896
rect 434822 507660 434854 507896
rect 434234 507576 434854 507660
rect 434234 507340 434266 507576
rect 434502 507340 434586 507576
rect 434822 507340 434854 507576
rect 434234 471896 434854 507340
rect 434234 471660 434266 471896
rect 434502 471660 434586 471896
rect 434822 471660 434854 471896
rect 434234 471576 434854 471660
rect 434234 471340 434266 471576
rect 434502 471340 434586 471576
rect 434822 471340 434854 471576
rect 434234 435896 434854 471340
rect 434234 435660 434266 435896
rect 434502 435660 434586 435896
rect 434822 435660 434854 435896
rect 434234 435576 434854 435660
rect 434234 435340 434266 435576
rect 434502 435340 434586 435576
rect 434822 435340 434854 435576
rect 434234 399896 434854 435340
rect 434234 399660 434266 399896
rect 434502 399660 434586 399896
rect 434822 399660 434854 399896
rect 434234 399576 434854 399660
rect 434234 399340 434266 399576
rect 434502 399340 434586 399576
rect 434822 399340 434854 399576
rect 434234 363896 434854 399340
rect 434234 363660 434266 363896
rect 434502 363660 434586 363896
rect 434822 363660 434854 363896
rect 434234 363576 434854 363660
rect 434234 363340 434266 363576
rect 434502 363340 434586 363576
rect 434822 363340 434854 363576
rect 434234 327896 434854 363340
rect 434234 327660 434266 327896
rect 434502 327660 434586 327896
rect 434822 327660 434854 327896
rect 434234 327576 434854 327660
rect 434234 327340 434266 327576
rect 434502 327340 434586 327576
rect 434822 327340 434854 327576
rect 434234 291896 434854 327340
rect 434234 291660 434266 291896
rect 434502 291660 434586 291896
rect 434822 291660 434854 291896
rect 434234 291576 434854 291660
rect 434234 291340 434266 291576
rect 434502 291340 434586 291576
rect 434822 291340 434854 291576
rect 434234 255896 434854 291340
rect 434234 255660 434266 255896
rect 434502 255660 434586 255896
rect 434822 255660 434854 255896
rect 434234 255576 434854 255660
rect 434234 255340 434266 255576
rect 434502 255340 434586 255576
rect 434822 255340 434854 255576
rect 434234 219896 434854 255340
rect 434234 219660 434266 219896
rect 434502 219660 434586 219896
rect 434822 219660 434854 219896
rect 434234 219576 434854 219660
rect 434234 219340 434266 219576
rect 434502 219340 434586 219576
rect 434822 219340 434854 219576
rect 434234 183896 434854 219340
rect 434234 183660 434266 183896
rect 434502 183660 434586 183896
rect 434822 183660 434854 183896
rect 434234 183576 434854 183660
rect 434234 183340 434266 183576
rect 434502 183340 434586 183576
rect 434822 183340 434854 183576
rect 434234 147896 434854 183340
rect 434234 147660 434266 147896
rect 434502 147660 434586 147896
rect 434822 147660 434854 147896
rect 434234 147576 434854 147660
rect 434234 147340 434266 147576
rect 434502 147340 434586 147576
rect 434822 147340 434854 147576
rect 434234 111896 434854 147340
rect 434234 111660 434266 111896
rect 434502 111660 434586 111896
rect 434822 111660 434854 111896
rect 434234 111576 434854 111660
rect 434234 111340 434266 111576
rect 434502 111340 434586 111576
rect 434822 111340 434854 111576
rect 434234 75896 434854 111340
rect 434234 75660 434266 75896
rect 434502 75660 434586 75896
rect 434822 75660 434854 75896
rect 434234 75576 434854 75660
rect 434234 75340 434266 75576
rect 434502 75340 434586 75576
rect 434822 75340 434854 75576
rect 434234 39896 434854 75340
rect 434234 39660 434266 39896
rect 434502 39660 434586 39896
rect 434822 39660 434854 39896
rect 434234 39576 434854 39660
rect 434234 39340 434266 39576
rect 434502 39340 434586 39576
rect 434822 39340 434854 39576
rect 434234 3896 434854 39340
rect 434234 3660 434266 3896
rect 434502 3660 434586 3896
rect 434822 3660 434854 3896
rect 434234 3576 434854 3660
rect 434234 3340 434266 3576
rect 434502 3340 434586 3576
rect 434822 3340 434854 3576
rect 434234 -1304 434854 3340
rect 434234 -1540 434266 -1304
rect 434502 -1540 434586 -1304
rect 434822 -1540 434854 -1304
rect 434234 -1624 434854 -1540
rect 434234 -1860 434266 -1624
rect 434502 -1860 434586 -1624
rect 434822 -1860 434854 -1624
rect 434234 -7652 434854 -1860
rect 435474 706760 436094 711592
rect 435474 706524 435506 706760
rect 435742 706524 435826 706760
rect 436062 706524 436094 706760
rect 435474 706440 436094 706524
rect 435474 706204 435506 706440
rect 435742 706204 435826 706440
rect 436062 706204 436094 706440
rect 435474 689136 436094 706204
rect 435474 688900 435506 689136
rect 435742 688900 435826 689136
rect 436062 688900 436094 689136
rect 435474 688816 436094 688900
rect 435474 688580 435506 688816
rect 435742 688580 435826 688816
rect 436062 688580 436094 688816
rect 435474 653136 436094 688580
rect 435474 652900 435506 653136
rect 435742 652900 435826 653136
rect 436062 652900 436094 653136
rect 435474 652816 436094 652900
rect 435474 652580 435506 652816
rect 435742 652580 435826 652816
rect 436062 652580 436094 652816
rect 435474 617136 436094 652580
rect 435474 616900 435506 617136
rect 435742 616900 435826 617136
rect 436062 616900 436094 617136
rect 435474 616816 436094 616900
rect 435474 616580 435506 616816
rect 435742 616580 435826 616816
rect 436062 616580 436094 616816
rect 435474 581136 436094 616580
rect 435474 580900 435506 581136
rect 435742 580900 435826 581136
rect 436062 580900 436094 581136
rect 435474 580816 436094 580900
rect 435474 580580 435506 580816
rect 435742 580580 435826 580816
rect 436062 580580 436094 580816
rect 435474 545136 436094 580580
rect 435474 544900 435506 545136
rect 435742 544900 435826 545136
rect 436062 544900 436094 545136
rect 435474 544816 436094 544900
rect 435474 544580 435506 544816
rect 435742 544580 435826 544816
rect 436062 544580 436094 544816
rect 435474 509136 436094 544580
rect 435474 508900 435506 509136
rect 435742 508900 435826 509136
rect 436062 508900 436094 509136
rect 435474 508816 436094 508900
rect 435474 508580 435506 508816
rect 435742 508580 435826 508816
rect 436062 508580 436094 508816
rect 435474 473136 436094 508580
rect 435474 472900 435506 473136
rect 435742 472900 435826 473136
rect 436062 472900 436094 473136
rect 435474 472816 436094 472900
rect 435474 472580 435506 472816
rect 435742 472580 435826 472816
rect 436062 472580 436094 472816
rect 435474 437136 436094 472580
rect 435474 436900 435506 437136
rect 435742 436900 435826 437136
rect 436062 436900 436094 437136
rect 435474 436816 436094 436900
rect 435474 436580 435506 436816
rect 435742 436580 435826 436816
rect 436062 436580 436094 436816
rect 435474 401136 436094 436580
rect 435474 400900 435506 401136
rect 435742 400900 435826 401136
rect 436062 400900 436094 401136
rect 435474 400816 436094 400900
rect 435474 400580 435506 400816
rect 435742 400580 435826 400816
rect 436062 400580 436094 400816
rect 435474 365136 436094 400580
rect 435474 364900 435506 365136
rect 435742 364900 435826 365136
rect 436062 364900 436094 365136
rect 435474 364816 436094 364900
rect 435474 364580 435506 364816
rect 435742 364580 435826 364816
rect 436062 364580 436094 364816
rect 435474 329136 436094 364580
rect 435474 328900 435506 329136
rect 435742 328900 435826 329136
rect 436062 328900 436094 329136
rect 435474 328816 436094 328900
rect 435474 328580 435506 328816
rect 435742 328580 435826 328816
rect 436062 328580 436094 328816
rect 435474 293136 436094 328580
rect 435474 292900 435506 293136
rect 435742 292900 435826 293136
rect 436062 292900 436094 293136
rect 435474 292816 436094 292900
rect 435474 292580 435506 292816
rect 435742 292580 435826 292816
rect 436062 292580 436094 292816
rect 435474 257136 436094 292580
rect 435474 256900 435506 257136
rect 435742 256900 435826 257136
rect 436062 256900 436094 257136
rect 435474 256816 436094 256900
rect 435474 256580 435506 256816
rect 435742 256580 435826 256816
rect 436062 256580 436094 256816
rect 435474 221136 436094 256580
rect 435474 220900 435506 221136
rect 435742 220900 435826 221136
rect 436062 220900 436094 221136
rect 435474 220816 436094 220900
rect 435474 220580 435506 220816
rect 435742 220580 435826 220816
rect 436062 220580 436094 220816
rect 435474 185136 436094 220580
rect 435474 184900 435506 185136
rect 435742 184900 435826 185136
rect 436062 184900 436094 185136
rect 435474 184816 436094 184900
rect 435474 184580 435506 184816
rect 435742 184580 435826 184816
rect 436062 184580 436094 184816
rect 435474 149136 436094 184580
rect 435474 148900 435506 149136
rect 435742 148900 435826 149136
rect 436062 148900 436094 149136
rect 435474 148816 436094 148900
rect 435474 148580 435506 148816
rect 435742 148580 435826 148816
rect 436062 148580 436094 148816
rect 435474 113136 436094 148580
rect 435474 112900 435506 113136
rect 435742 112900 435826 113136
rect 436062 112900 436094 113136
rect 435474 112816 436094 112900
rect 435474 112580 435506 112816
rect 435742 112580 435826 112816
rect 436062 112580 436094 112816
rect 435474 77136 436094 112580
rect 435474 76900 435506 77136
rect 435742 76900 435826 77136
rect 436062 76900 436094 77136
rect 435474 76816 436094 76900
rect 435474 76580 435506 76816
rect 435742 76580 435826 76816
rect 436062 76580 436094 76816
rect 435474 41136 436094 76580
rect 435474 40900 435506 41136
rect 435742 40900 435826 41136
rect 436062 40900 436094 41136
rect 435474 40816 436094 40900
rect 435474 40580 435506 40816
rect 435742 40580 435826 40816
rect 436062 40580 436094 40816
rect 435474 5136 436094 40580
rect 435474 4900 435506 5136
rect 435742 4900 435826 5136
rect 436062 4900 436094 5136
rect 435474 4816 436094 4900
rect 435474 4580 435506 4816
rect 435742 4580 435826 4816
rect 436062 4580 436094 4816
rect 435474 -2264 436094 4580
rect 435474 -2500 435506 -2264
rect 435742 -2500 435826 -2264
rect 436062 -2500 436094 -2264
rect 435474 -2584 436094 -2500
rect 435474 -2820 435506 -2584
rect 435742 -2820 435826 -2584
rect 436062 -2820 436094 -2584
rect 435474 -7652 436094 -2820
rect 436714 707720 437334 711592
rect 436714 707484 436746 707720
rect 436982 707484 437066 707720
rect 437302 707484 437334 707720
rect 436714 707400 437334 707484
rect 436714 707164 436746 707400
rect 436982 707164 437066 707400
rect 437302 707164 437334 707400
rect 436714 690376 437334 707164
rect 436714 690140 436746 690376
rect 436982 690140 437066 690376
rect 437302 690140 437334 690376
rect 436714 690056 437334 690140
rect 436714 689820 436746 690056
rect 436982 689820 437066 690056
rect 437302 689820 437334 690056
rect 436714 654376 437334 689820
rect 436714 654140 436746 654376
rect 436982 654140 437066 654376
rect 437302 654140 437334 654376
rect 436714 654056 437334 654140
rect 436714 653820 436746 654056
rect 436982 653820 437066 654056
rect 437302 653820 437334 654056
rect 436714 618376 437334 653820
rect 436714 618140 436746 618376
rect 436982 618140 437066 618376
rect 437302 618140 437334 618376
rect 436714 618056 437334 618140
rect 436714 617820 436746 618056
rect 436982 617820 437066 618056
rect 437302 617820 437334 618056
rect 436714 582376 437334 617820
rect 436714 582140 436746 582376
rect 436982 582140 437066 582376
rect 437302 582140 437334 582376
rect 436714 582056 437334 582140
rect 436714 581820 436746 582056
rect 436982 581820 437066 582056
rect 437302 581820 437334 582056
rect 436714 546376 437334 581820
rect 436714 546140 436746 546376
rect 436982 546140 437066 546376
rect 437302 546140 437334 546376
rect 436714 546056 437334 546140
rect 436714 545820 436746 546056
rect 436982 545820 437066 546056
rect 437302 545820 437334 546056
rect 436714 510376 437334 545820
rect 436714 510140 436746 510376
rect 436982 510140 437066 510376
rect 437302 510140 437334 510376
rect 436714 510056 437334 510140
rect 436714 509820 436746 510056
rect 436982 509820 437066 510056
rect 437302 509820 437334 510056
rect 436714 474376 437334 509820
rect 436714 474140 436746 474376
rect 436982 474140 437066 474376
rect 437302 474140 437334 474376
rect 436714 474056 437334 474140
rect 436714 473820 436746 474056
rect 436982 473820 437066 474056
rect 437302 473820 437334 474056
rect 436714 438376 437334 473820
rect 436714 438140 436746 438376
rect 436982 438140 437066 438376
rect 437302 438140 437334 438376
rect 436714 438056 437334 438140
rect 436714 437820 436746 438056
rect 436982 437820 437066 438056
rect 437302 437820 437334 438056
rect 436714 402376 437334 437820
rect 436714 402140 436746 402376
rect 436982 402140 437066 402376
rect 437302 402140 437334 402376
rect 436714 402056 437334 402140
rect 436714 401820 436746 402056
rect 436982 401820 437066 402056
rect 437302 401820 437334 402056
rect 436714 366376 437334 401820
rect 436714 366140 436746 366376
rect 436982 366140 437066 366376
rect 437302 366140 437334 366376
rect 436714 366056 437334 366140
rect 436714 365820 436746 366056
rect 436982 365820 437066 366056
rect 437302 365820 437334 366056
rect 436714 330376 437334 365820
rect 436714 330140 436746 330376
rect 436982 330140 437066 330376
rect 437302 330140 437334 330376
rect 436714 330056 437334 330140
rect 436714 329820 436746 330056
rect 436982 329820 437066 330056
rect 437302 329820 437334 330056
rect 436714 294376 437334 329820
rect 436714 294140 436746 294376
rect 436982 294140 437066 294376
rect 437302 294140 437334 294376
rect 436714 294056 437334 294140
rect 436714 293820 436746 294056
rect 436982 293820 437066 294056
rect 437302 293820 437334 294056
rect 436714 258376 437334 293820
rect 436714 258140 436746 258376
rect 436982 258140 437066 258376
rect 437302 258140 437334 258376
rect 436714 258056 437334 258140
rect 436714 257820 436746 258056
rect 436982 257820 437066 258056
rect 437302 257820 437334 258056
rect 436714 222376 437334 257820
rect 436714 222140 436746 222376
rect 436982 222140 437066 222376
rect 437302 222140 437334 222376
rect 436714 222056 437334 222140
rect 436714 221820 436746 222056
rect 436982 221820 437066 222056
rect 437302 221820 437334 222056
rect 436714 186376 437334 221820
rect 436714 186140 436746 186376
rect 436982 186140 437066 186376
rect 437302 186140 437334 186376
rect 436714 186056 437334 186140
rect 436714 185820 436746 186056
rect 436982 185820 437066 186056
rect 437302 185820 437334 186056
rect 436714 150376 437334 185820
rect 436714 150140 436746 150376
rect 436982 150140 437066 150376
rect 437302 150140 437334 150376
rect 436714 150056 437334 150140
rect 436714 149820 436746 150056
rect 436982 149820 437066 150056
rect 437302 149820 437334 150056
rect 436714 114376 437334 149820
rect 436714 114140 436746 114376
rect 436982 114140 437066 114376
rect 437302 114140 437334 114376
rect 436714 114056 437334 114140
rect 436714 113820 436746 114056
rect 436982 113820 437066 114056
rect 437302 113820 437334 114056
rect 436714 78376 437334 113820
rect 436714 78140 436746 78376
rect 436982 78140 437066 78376
rect 437302 78140 437334 78376
rect 436714 78056 437334 78140
rect 436714 77820 436746 78056
rect 436982 77820 437066 78056
rect 437302 77820 437334 78056
rect 436714 42376 437334 77820
rect 436714 42140 436746 42376
rect 436982 42140 437066 42376
rect 437302 42140 437334 42376
rect 436714 42056 437334 42140
rect 436714 41820 436746 42056
rect 436982 41820 437066 42056
rect 437302 41820 437334 42056
rect 436714 6376 437334 41820
rect 436714 6140 436746 6376
rect 436982 6140 437066 6376
rect 437302 6140 437334 6376
rect 436714 6056 437334 6140
rect 436714 5820 436746 6056
rect 436982 5820 437066 6056
rect 437302 5820 437334 6056
rect 436714 -3224 437334 5820
rect 436714 -3460 436746 -3224
rect 436982 -3460 437066 -3224
rect 437302 -3460 437334 -3224
rect 436714 -3544 437334 -3460
rect 436714 -3780 436746 -3544
rect 436982 -3780 437066 -3544
rect 437302 -3780 437334 -3544
rect 436714 -7652 437334 -3780
rect 437954 708680 438574 711592
rect 437954 708444 437986 708680
rect 438222 708444 438306 708680
rect 438542 708444 438574 708680
rect 437954 708360 438574 708444
rect 437954 708124 437986 708360
rect 438222 708124 438306 708360
rect 438542 708124 438574 708360
rect 437954 691616 438574 708124
rect 437954 691380 437986 691616
rect 438222 691380 438306 691616
rect 438542 691380 438574 691616
rect 437954 691296 438574 691380
rect 437954 691060 437986 691296
rect 438222 691060 438306 691296
rect 438542 691060 438574 691296
rect 437954 655616 438574 691060
rect 437954 655380 437986 655616
rect 438222 655380 438306 655616
rect 438542 655380 438574 655616
rect 437954 655296 438574 655380
rect 437954 655060 437986 655296
rect 438222 655060 438306 655296
rect 438542 655060 438574 655296
rect 437954 619616 438574 655060
rect 437954 619380 437986 619616
rect 438222 619380 438306 619616
rect 438542 619380 438574 619616
rect 437954 619296 438574 619380
rect 437954 619060 437986 619296
rect 438222 619060 438306 619296
rect 438542 619060 438574 619296
rect 437954 583616 438574 619060
rect 437954 583380 437986 583616
rect 438222 583380 438306 583616
rect 438542 583380 438574 583616
rect 437954 583296 438574 583380
rect 437954 583060 437986 583296
rect 438222 583060 438306 583296
rect 438542 583060 438574 583296
rect 437954 547616 438574 583060
rect 437954 547380 437986 547616
rect 438222 547380 438306 547616
rect 438542 547380 438574 547616
rect 437954 547296 438574 547380
rect 437954 547060 437986 547296
rect 438222 547060 438306 547296
rect 438542 547060 438574 547296
rect 437954 511616 438574 547060
rect 437954 511380 437986 511616
rect 438222 511380 438306 511616
rect 438542 511380 438574 511616
rect 437954 511296 438574 511380
rect 437954 511060 437986 511296
rect 438222 511060 438306 511296
rect 438542 511060 438574 511296
rect 437954 475616 438574 511060
rect 437954 475380 437986 475616
rect 438222 475380 438306 475616
rect 438542 475380 438574 475616
rect 437954 475296 438574 475380
rect 437954 475060 437986 475296
rect 438222 475060 438306 475296
rect 438542 475060 438574 475296
rect 437954 439616 438574 475060
rect 437954 439380 437986 439616
rect 438222 439380 438306 439616
rect 438542 439380 438574 439616
rect 437954 439296 438574 439380
rect 437954 439060 437986 439296
rect 438222 439060 438306 439296
rect 438542 439060 438574 439296
rect 437954 403616 438574 439060
rect 437954 403380 437986 403616
rect 438222 403380 438306 403616
rect 438542 403380 438574 403616
rect 437954 403296 438574 403380
rect 437954 403060 437986 403296
rect 438222 403060 438306 403296
rect 438542 403060 438574 403296
rect 437954 367616 438574 403060
rect 437954 367380 437986 367616
rect 438222 367380 438306 367616
rect 438542 367380 438574 367616
rect 437954 367296 438574 367380
rect 437954 367060 437986 367296
rect 438222 367060 438306 367296
rect 438542 367060 438574 367296
rect 437954 331616 438574 367060
rect 437954 331380 437986 331616
rect 438222 331380 438306 331616
rect 438542 331380 438574 331616
rect 437954 331296 438574 331380
rect 437954 331060 437986 331296
rect 438222 331060 438306 331296
rect 438542 331060 438574 331296
rect 437954 295616 438574 331060
rect 437954 295380 437986 295616
rect 438222 295380 438306 295616
rect 438542 295380 438574 295616
rect 437954 295296 438574 295380
rect 437954 295060 437986 295296
rect 438222 295060 438306 295296
rect 438542 295060 438574 295296
rect 437954 259616 438574 295060
rect 437954 259380 437986 259616
rect 438222 259380 438306 259616
rect 438542 259380 438574 259616
rect 437954 259296 438574 259380
rect 437954 259060 437986 259296
rect 438222 259060 438306 259296
rect 438542 259060 438574 259296
rect 437954 223616 438574 259060
rect 437954 223380 437986 223616
rect 438222 223380 438306 223616
rect 438542 223380 438574 223616
rect 437954 223296 438574 223380
rect 437954 223060 437986 223296
rect 438222 223060 438306 223296
rect 438542 223060 438574 223296
rect 437954 187616 438574 223060
rect 437954 187380 437986 187616
rect 438222 187380 438306 187616
rect 438542 187380 438574 187616
rect 437954 187296 438574 187380
rect 437954 187060 437986 187296
rect 438222 187060 438306 187296
rect 438542 187060 438574 187296
rect 437954 151616 438574 187060
rect 437954 151380 437986 151616
rect 438222 151380 438306 151616
rect 438542 151380 438574 151616
rect 437954 151296 438574 151380
rect 437954 151060 437986 151296
rect 438222 151060 438306 151296
rect 438542 151060 438574 151296
rect 437954 115616 438574 151060
rect 437954 115380 437986 115616
rect 438222 115380 438306 115616
rect 438542 115380 438574 115616
rect 437954 115296 438574 115380
rect 437954 115060 437986 115296
rect 438222 115060 438306 115296
rect 438542 115060 438574 115296
rect 437954 79616 438574 115060
rect 437954 79380 437986 79616
rect 438222 79380 438306 79616
rect 438542 79380 438574 79616
rect 437954 79296 438574 79380
rect 437954 79060 437986 79296
rect 438222 79060 438306 79296
rect 438542 79060 438574 79296
rect 437954 43616 438574 79060
rect 437954 43380 437986 43616
rect 438222 43380 438306 43616
rect 438542 43380 438574 43616
rect 437954 43296 438574 43380
rect 437954 43060 437986 43296
rect 438222 43060 438306 43296
rect 438542 43060 438574 43296
rect 437954 7616 438574 43060
rect 437954 7380 437986 7616
rect 438222 7380 438306 7616
rect 438542 7380 438574 7616
rect 437954 7296 438574 7380
rect 437954 7060 437986 7296
rect 438222 7060 438306 7296
rect 438542 7060 438574 7296
rect 437954 -4184 438574 7060
rect 437954 -4420 437986 -4184
rect 438222 -4420 438306 -4184
rect 438542 -4420 438574 -4184
rect 437954 -4504 438574 -4420
rect 437954 -4740 437986 -4504
rect 438222 -4740 438306 -4504
rect 438542 -4740 438574 -4504
rect 437954 -7652 438574 -4740
rect 439194 709640 439814 711592
rect 439194 709404 439226 709640
rect 439462 709404 439546 709640
rect 439782 709404 439814 709640
rect 439194 709320 439814 709404
rect 439194 709084 439226 709320
rect 439462 709084 439546 709320
rect 439782 709084 439814 709320
rect 439194 692856 439814 709084
rect 439194 692620 439226 692856
rect 439462 692620 439546 692856
rect 439782 692620 439814 692856
rect 439194 692536 439814 692620
rect 439194 692300 439226 692536
rect 439462 692300 439546 692536
rect 439782 692300 439814 692536
rect 439194 656856 439814 692300
rect 439194 656620 439226 656856
rect 439462 656620 439546 656856
rect 439782 656620 439814 656856
rect 439194 656536 439814 656620
rect 439194 656300 439226 656536
rect 439462 656300 439546 656536
rect 439782 656300 439814 656536
rect 439194 620856 439814 656300
rect 439194 620620 439226 620856
rect 439462 620620 439546 620856
rect 439782 620620 439814 620856
rect 439194 620536 439814 620620
rect 439194 620300 439226 620536
rect 439462 620300 439546 620536
rect 439782 620300 439814 620536
rect 439194 584856 439814 620300
rect 439194 584620 439226 584856
rect 439462 584620 439546 584856
rect 439782 584620 439814 584856
rect 439194 584536 439814 584620
rect 439194 584300 439226 584536
rect 439462 584300 439546 584536
rect 439782 584300 439814 584536
rect 439194 548856 439814 584300
rect 439194 548620 439226 548856
rect 439462 548620 439546 548856
rect 439782 548620 439814 548856
rect 439194 548536 439814 548620
rect 439194 548300 439226 548536
rect 439462 548300 439546 548536
rect 439782 548300 439814 548536
rect 439194 512856 439814 548300
rect 439194 512620 439226 512856
rect 439462 512620 439546 512856
rect 439782 512620 439814 512856
rect 439194 512536 439814 512620
rect 439194 512300 439226 512536
rect 439462 512300 439546 512536
rect 439782 512300 439814 512536
rect 439194 476856 439814 512300
rect 439194 476620 439226 476856
rect 439462 476620 439546 476856
rect 439782 476620 439814 476856
rect 439194 476536 439814 476620
rect 439194 476300 439226 476536
rect 439462 476300 439546 476536
rect 439782 476300 439814 476536
rect 439194 440856 439814 476300
rect 439194 440620 439226 440856
rect 439462 440620 439546 440856
rect 439782 440620 439814 440856
rect 439194 440536 439814 440620
rect 439194 440300 439226 440536
rect 439462 440300 439546 440536
rect 439782 440300 439814 440536
rect 439194 404856 439814 440300
rect 439194 404620 439226 404856
rect 439462 404620 439546 404856
rect 439782 404620 439814 404856
rect 439194 404536 439814 404620
rect 439194 404300 439226 404536
rect 439462 404300 439546 404536
rect 439782 404300 439814 404536
rect 439194 368856 439814 404300
rect 439194 368620 439226 368856
rect 439462 368620 439546 368856
rect 439782 368620 439814 368856
rect 439194 368536 439814 368620
rect 439194 368300 439226 368536
rect 439462 368300 439546 368536
rect 439782 368300 439814 368536
rect 439194 332856 439814 368300
rect 439194 332620 439226 332856
rect 439462 332620 439546 332856
rect 439782 332620 439814 332856
rect 439194 332536 439814 332620
rect 439194 332300 439226 332536
rect 439462 332300 439546 332536
rect 439782 332300 439814 332536
rect 439194 296856 439814 332300
rect 439194 296620 439226 296856
rect 439462 296620 439546 296856
rect 439782 296620 439814 296856
rect 439194 296536 439814 296620
rect 439194 296300 439226 296536
rect 439462 296300 439546 296536
rect 439782 296300 439814 296536
rect 439194 260856 439814 296300
rect 439194 260620 439226 260856
rect 439462 260620 439546 260856
rect 439782 260620 439814 260856
rect 439194 260536 439814 260620
rect 439194 260300 439226 260536
rect 439462 260300 439546 260536
rect 439782 260300 439814 260536
rect 439194 224856 439814 260300
rect 439194 224620 439226 224856
rect 439462 224620 439546 224856
rect 439782 224620 439814 224856
rect 439194 224536 439814 224620
rect 439194 224300 439226 224536
rect 439462 224300 439546 224536
rect 439782 224300 439814 224536
rect 439194 188856 439814 224300
rect 439194 188620 439226 188856
rect 439462 188620 439546 188856
rect 439782 188620 439814 188856
rect 439194 188536 439814 188620
rect 439194 188300 439226 188536
rect 439462 188300 439546 188536
rect 439782 188300 439814 188536
rect 439194 152856 439814 188300
rect 439194 152620 439226 152856
rect 439462 152620 439546 152856
rect 439782 152620 439814 152856
rect 439194 152536 439814 152620
rect 439194 152300 439226 152536
rect 439462 152300 439546 152536
rect 439782 152300 439814 152536
rect 439194 116856 439814 152300
rect 439194 116620 439226 116856
rect 439462 116620 439546 116856
rect 439782 116620 439814 116856
rect 439194 116536 439814 116620
rect 439194 116300 439226 116536
rect 439462 116300 439546 116536
rect 439782 116300 439814 116536
rect 439194 80856 439814 116300
rect 439194 80620 439226 80856
rect 439462 80620 439546 80856
rect 439782 80620 439814 80856
rect 439194 80536 439814 80620
rect 439194 80300 439226 80536
rect 439462 80300 439546 80536
rect 439782 80300 439814 80536
rect 439194 44856 439814 80300
rect 439194 44620 439226 44856
rect 439462 44620 439546 44856
rect 439782 44620 439814 44856
rect 439194 44536 439814 44620
rect 439194 44300 439226 44536
rect 439462 44300 439546 44536
rect 439782 44300 439814 44536
rect 439194 8856 439814 44300
rect 439194 8620 439226 8856
rect 439462 8620 439546 8856
rect 439782 8620 439814 8856
rect 439194 8536 439814 8620
rect 439194 8300 439226 8536
rect 439462 8300 439546 8536
rect 439782 8300 439814 8536
rect 439194 -5144 439814 8300
rect 439194 -5380 439226 -5144
rect 439462 -5380 439546 -5144
rect 439782 -5380 439814 -5144
rect 439194 -5464 439814 -5380
rect 439194 -5700 439226 -5464
rect 439462 -5700 439546 -5464
rect 439782 -5700 439814 -5464
rect 439194 -7652 439814 -5700
rect 440434 710600 441054 711592
rect 440434 710364 440466 710600
rect 440702 710364 440786 710600
rect 441022 710364 441054 710600
rect 440434 710280 441054 710364
rect 440434 710044 440466 710280
rect 440702 710044 440786 710280
rect 441022 710044 441054 710280
rect 440434 694096 441054 710044
rect 440434 693860 440466 694096
rect 440702 693860 440786 694096
rect 441022 693860 441054 694096
rect 440434 693776 441054 693860
rect 440434 693540 440466 693776
rect 440702 693540 440786 693776
rect 441022 693540 441054 693776
rect 440434 658096 441054 693540
rect 440434 657860 440466 658096
rect 440702 657860 440786 658096
rect 441022 657860 441054 658096
rect 440434 657776 441054 657860
rect 440434 657540 440466 657776
rect 440702 657540 440786 657776
rect 441022 657540 441054 657776
rect 440434 622096 441054 657540
rect 440434 621860 440466 622096
rect 440702 621860 440786 622096
rect 441022 621860 441054 622096
rect 440434 621776 441054 621860
rect 440434 621540 440466 621776
rect 440702 621540 440786 621776
rect 441022 621540 441054 621776
rect 440434 586096 441054 621540
rect 440434 585860 440466 586096
rect 440702 585860 440786 586096
rect 441022 585860 441054 586096
rect 440434 585776 441054 585860
rect 440434 585540 440466 585776
rect 440702 585540 440786 585776
rect 441022 585540 441054 585776
rect 440434 550096 441054 585540
rect 440434 549860 440466 550096
rect 440702 549860 440786 550096
rect 441022 549860 441054 550096
rect 440434 549776 441054 549860
rect 440434 549540 440466 549776
rect 440702 549540 440786 549776
rect 441022 549540 441054 549776
rect 440434 514096 441054 549540
rect 440434 513860 440466 514096
rect 440702 513860 440786 514096
rect 441022 513860 441054 514096
rect 440434 513776 441054 513860
rect 440434 513540 440466 513776
rect 440702 513540 440786 513776
rect 441022 513540 441054 513776
rect 440434 478096 441054 513540
rect 440434 477860 440466 478096
rect 440702 477860 440786 478096
rect 441022 477860 441054 478096
rect 440434 477776 441054 477860
rect 440434 477540 440466 477776
rect 440702 477540 440786 477776
rect 441022 477540 441054 477776
rect 440434 442096 441054 477540
rect 440434 441860 440466 442096
rect 440702 441860 440786 442096
rect 441022 441860 441054 442096
rect 440434 441776 441054 441860
rect 440434 441540 440466 441776
rect 440702 441540 440786 441776
rect 441022 441540 441054 441776
rect 440434 406096 441054 441540
rect 440434 405860 440466 406096
rect 440702 405860 440786 406096
rect 441022 405860 441054 406096
rect 440434 405776 441054 405860
rect 440434 405540 440466 405776
rect 440702 405540 440786 405776
rect 441022 405540 441054 405776
rect 440434 370096 441054 405540
rect 440434 369860 440466 370096
rect 440702 369860 440786 370096
rect 441022 369860 441054 370096
rect 440434 369776 441054 369860
rect 440434 369540 440466 369776
rect 440702 369540 440786 369776
rect 441022 369540 441054 369776
rect 440434 334096 441054 369540
rect 440434 333860 440466 334096
rect 440702 333860 440786 334096
rect 441022 333860 441054 334096
rect 440434 333776 441054 333860
rect 440434 333540 440466 333776
rect 440702 333540 440786 333776
rect 441022 333540 441054 333776
rect 440434 298096 441054 333540
rect 440434 297860 440466 298096
rect 440702 297860 440786 298096
rect 441022 297860 441054 298096
rect 440434 297776 441054 297860
rect 440434 297540 440466 297776
rect 440702 297540 440786 297776
rect 441022 297540 441054 297776
rect 440434 262096 441054 297540
rect 440434 261860 440466 262096
rect 440702 261860 440786 262096
rect 441022 261860 441054 262096
rect 440434 261776 441054 261860
rect 440434 261540 440466 261776
rect 440702 261540 440786 261776
rect 441022 261540 441054 261776
rect 440434 226096 441054 261540
rect 440434 225860 440466 226096
rect 440702 225860 440786 226096
rect 441022 225860 441054 226096
rect 440434 225776 441054 225860
rect 440434 225540 440466 225776
rect 440702 225540 440786 225776
rect 441022 225540 441054 225776
rect 440434 190096 441054 225540
rect 440434 189860 440466 190096
rect 440702 189860 440786 190096
rect 441022 189860 441054 190096
rect 440434 189776 441054 189860
rect 440434 189540 440466 189776
rect 440702 189540 440786 189776
rect 441022 189540 441054 189776
rect 440434 154096 441054 189540
rect 440434 153860 440466 154096
rect 440702 153860 440786 154096
rect 441022 153860 441054 154096
rect 440434 153776 441054 153860
rect 440434 153540 440466 153776
rect 440702 153540 440786 153776
rect 441022 153540 441054 153776
rect 440434 118096 441054 153540
rect 440434 117860 440466 118096
rect 440702 117860 440786 118096
rect 441022 117860 441054 118096
rect 440434 117776 441054 117860
rect 440434 117540 440466 117776
rect 440702 117540 440786 117776
rect 441022 117540 441054 117776
rect 440434 82096 441054 117540
rect 440434 81860 440466 82096
rect 440702 81860 440786 82096
rect 441022 81860 441054 82096
rect 440434 81776 441054 81860
rect 440434 81540 440466 81776
rect 440702 81540 440786 81776
rect 441022 81540 441054 81776
rect 440434 46096 441054 81540
rect 440434 45860 440466 46096
rect 440702 45860 440786 46096
rect 441022 45860 441054 46096
rect 440434 45776 441054 45860
rect 440434 45540 440466 45776
rect 440702 45540 440786 45776
rect 441022 45540 441054 45776
rect 440434 10096 441054 45540
rect 440434 9860 440466 10096
rect 440702 9860 440786 10096
rect 441022 9860 441054 10096
rect 440434 9776 441054 9860
rect 440434 9540 440466 9776
rect 440702 9540 440786 9776
rect 441022 9540 441054 9776
rect 440434 -6104 441054 9540
rect 440434 -6340 440466 -6104
rect 440702 -6340 440786 -6104
rect 441022 -6340 441054 -6104
rect 440434 -6424 441054 -6340
rect 440434 -6660 440466 -6424
rect 440702 -6660 440786 -6424
rect 441022 -6660 441054 -6424
rect 440434 -7652 441054 -6660
rect 441674 711560 442294 711592
rect 441674 711324 441706 711560
rect 441942 711324 442026 711560
rect 442262 711324 442294 711560
rect 441674 711240 442294 711324
rect 441674 711004 441706 711240
rect 441942 711004 442026 711240
rect 442262 711004 442294 711240
rect 441674 695336 442294 711004
rect 441674 695100 441706 695336
rect 441942 695100 442026 695336
rect 442262 695100 442294 695336
rect 441674 695016 442294 695100
rect 441674 694780 441706 695016
rect 441942 694780 442026 695016
rect 442262 694780 442294 695016
rect 441674 659336 442294 694780
rect 441674 659100 441706 659336
rect 441942 659100 442026 659336
rect 442262 659100 442294 659336
rect 441674 659016 442294 659100
rect 441674 658780 441706 659016
rect 441942 658780 442026 659016
rect 442262 658780 442294 659016
rect 441674 623336 442294 658780
rect 441674 623100 441706 623336
rect 441942 623100 442026 623336
rect 442262 623100 442294 623336
rect 441674 623016 442294 623100
rect 441674 622780 441706 623016
rect 441942 622780 442026 623016
rect 442262 622780 442294 623016
rect 441674 587336 442294 622780
rect 441674 587100 441706 587336
rect 441942 587100 442026 587336
rect 442262 587100 442294 587336
rect 441674 587016 442294 587100
rect 441674 586780 441706 587016
rect 441942 586780 442026 587016
rect 442262 586780 442294 587016
rect 441674 551336 442294 586780
rect 441674 551100 441706 551336
rect 441942 551100 442026 551336
rect 442262 551100 442294 551336
rect 441674 551016 442294 551100
rect 441674 550780 441706 551016
rect 441942 550780 442026 551016
rect 442262 550780 442294 551016
rect 441674 515336 442294 550780
rect 441674 515100 441706 515336
rect 441942 515100 442026 515336
rect 442262 515100 442294 515336
rect 441674 515016 442294 515100
rect 441674 514780 441706 515016
rect 441942 514780 442026 515016
rect 442262 514780 442294 515016
rect 441674 479336 442294 514780
rect 441674 479100 441706 479336
rect 441942 479100 442026 479336
rect 442262 479100 442294 479336
rect 441674 479016 442294 479100
rect 441674 478780 441706 479016
rect 441942 478780 442026 479016
rect 442262 478780 442294 479016
rect 441674 443336 442294 478780
rect 441674 443100 441706 443336
rect 441942 443100 442026 443336
rect 442262 443100 442294 443336
rect 441674 443016 442294 443100
rect 441674 442780 441706 443016
rect 441942 442780 442026 443016
rect 442262 442780 442294 443016
rect 441674 407336 442294 442780
rect 441674 407100 441706 407336
rect 441942 407100 442026 407336
rect 442262 407100 442294 407336
rect 441674 407016 442294 407100
rect 441674 406780 441706 407016
rect 441942 406780 442026 407016
rect 442262 406780 442294 407016
rect 441674 371336 442294 406780
rect 441674 371100 441706 371336
rect 441942 371100 442026 371336
rect 442262 371100 442294 371336
rect 441674 371016 442294 371100
rect 441674 370780 441706 371016
rect 441942 370780 442026 371016
rect 442262 370780 442294 371016
rect 441674 335336 442294 370780
rect 441674 335100 441706 335336
rect 441942 335100 442026 335336
rect 442262 335100 442294 335336
rect 441674 335016 442294 335100
rect 441674 334780 441706 335016
rect 441942 334780 442026 335016
rect 442262 334780 442294 335016
rect 441674 299336 442294 334780
rect 441674 299100 441706 299336
rect 441942 299100 442026 299336
rect 442262 299100 442294 299336
rect 441674 299016 442294 299100
rect 441674 298780 441706 299016
rect 441942 298780 442026 299016
rect 442262 298780 442294 299016
rect 441674 263336 442294 298780
rect 441674 263100 441706 263336
rect 441942 263100 442026 263336
rect 442262 263100 442294 263336
rect 441674 263016 442294 263100
rect 441674 262780 441706 263016
rect 441942 262780 442026 263016
rect 442262 262780 442294 263016
rect 441674 227336 442294 262780
rect 441674 227100 441706 227336
rect 441942 227100 442026 227336
rect 442262 227100 442294 227336
rect 441674 227016 442294 227100
rect 441674 226780 441706 227016
rect 441942 226780 442026 227016
rect 442262 226780 442294 227016
rect 441674 191336 442294 226780
rect 441674 191100 441706 191336
rect 441942 191100 442026 191336
rect 442262 191100 442294 191336
rect 441674 191016 442294 191100
rect 441674 190780 441706 191016
rect 441942 190780 442026 191016
rect 442262 190780 442294 191016
rect 441674 155336 442294 190780
rect 441674 155100 441706 155336
rect 441942 155100 442026 155336
rect 442262 155100 442294 155336
rect 441674 155016 442294 155100
rect 441674 154780 441706 155016
rect 441942 154780 442026 155016
rect 442262 154780 442294 155016
rect 441674 119336 442294 154780
rect 441674 119100 441706 119336
rect 441942 119100 442026 119336
rect 442262 119100 442294 119336
rect 441674 119016 442294 119100
rect 441674 118780 441706 119016
rect 441942 118780 442026 119016
rect 442262 118780 442294 119016
rect 441674 83336 442294 118780
rect 441674 83100 441706 83336
rect 441942 83100 442026 83336
rect 442262 83100 442294 83336
rect 441674 83016 442294 83100
rect 441674 82780 441706 83016
rect 441942 82780 442026 83016
rect 442262 82780 442294 83016
rect 441674 47336 442294 82780
rect 441674 47100 441706 47336
rect 441942 47100 442026 47336
rect 442262 47100 442294 47336
rect 441674 47016 442294 47100
rect 441674 46780 441706 47016
rect 441942 46780 442026 47016
rect 442262 46780 442294 47016
rect 441674 11336 442294 46780
rect 441674 11100 441706 11336
rect 441942 11100 442026 11336
rect 442262 11100 442294 11336
rect 441674 11016 442294 11100
rect 441674 10780 441706 11016
rect 441942 10780 442026 11016
rect 442262 10780 442294 11016
rect 441674 -7064 442294 10780
rect 441674 -7300 441706 -7064
rect 441942 -7300 442026 -7064
rect 442262 -7300 442294 -7064
rect 441674 -7384 442294 -7300
rect 441674 -7620 441706 -7384
rect 441942 -7620 442026 -7384
rect 442262 -7620 442294 -7384
rect 441674 -7652 442294 -7620
rect 468994 704840 469614 711592
rect 468994 704604 469026 704840
rect 469262 704604 469346 704840
rect 469582 704604 469614 704840
rect 468994 704520 469614 704604
rect 468994 704284 469026 704520
rect 469262 704284 469346 704520
rect 469582 704284 469614 704520
rect 468994 686656 469614 704284
rect 468994 686420 469026 686656
rect 469262 686420 469346 686656
rect 469582 686420 469614 686656
rect 468994 686336 469614 686420
rect 468994 686100 469026 686336
rect 469262 686100 469346 686336
rect 469582 686100 469614 686336
rect 468994 650656 469614 686100
rect 468994 650420 469026 650656
rect 469262 650420 469346 650656
rect 469582 650420 469614 650656
rect 468994 650336 469614 650420
rect 468994 650100 469026 650336
rect 469262 650100 469346 650336
rect 469582 650100 469614 650336
rect 468994 614656 469614 650100
rect 468994 614420 469026 614656
rect 469262 614420 469346 614656
rect 469582 614420 469614 614656
rect 468994 614336 469614 614420
rect 468994 614100 469026 614336
rect 469262 614100 469346 614336
rect 469582 614100 469614 614336
rect 468994 578656 469614 614100
rect 468994 578420 469026 578656
rect 469262 578420 469346 578656
rect 469582 578420 469614 578656
rect 468994 578336 469614 578420
rect 468994 578100 469026 578336
rect 469262 578100 469346 578336
rect 469582 578100 469614 578336
rect 468994 542656 469614 578100
rect 468994 542420 469026 542656
rect 469262 542420 469346 542656
rect 469582 542420 469614 542656
rect 468994 542336 469614 542420
rect 468994 542100 469026 542336
rect 469262 542100 469346 542336
rect 469582 542100 469614 542336
rect 468994 506656 469614 542100
rect 468994 506420 469026 506656
rect 469262 506420 469346 506656
rect 469582 506420 469614 506656
rect 468994 506336 469614 506420
rect 468994 506100 469026 506336
rect 469262 506100 469346 506336
rect 469582 506100 469614 506336
rect 468994 470656 469614 506100
rect 468994 470420 469026 470656
rect 469262 470420 469346 470656
rect 469582 470420 469614 470656
rect 468994 470336 469614 470420
rect 468994 470100 469026 470336
rect 469262 470100 469346 470336
rect 469582 470100 469614 470336
rect 468994 450399 469614 470100
rect 468994 450335 469032 450399
rect 469096 450335 469112 450399
rect 469176 450335 469192 450399
rect 469256 450335 469272 450399
rect 469336 450335 469352 450399
rect 469416 450335 469432 450399
rect 469496 450335 469512 450399
rect 469576 450335 469614 450399
rect 468994 450319 469614 450335
rect 468994 450255 469032 450319
rect 469096 450255 469112 450319
rect 469176 450255 469192 450319
rect 469256 450255 469272 450319
rect 469336 450255 469352 450319
rect 469416 450255 469432 450319
rect 469496 450255 469512 450319
rect 469576 450255 469614 450319
rect 468994 450239 469614 450255
rect 468994 450175 469032 450239
rect 469096 450175 469112 450239
rect 469176 450175 469192 450239
rect 469256 450175 469272 450239
rect 469336 450175 469352 450239
rect 469416 450175 469432 450239
rect 469496 450175 469512 450239
rect 469576 450175 469614 450239
rect 468994 450159 469614 450175
rect 468994 450095 469032 450159
rect 469096 450095 469112 450159
rect 469176 450095 469192 450159
rect 469256 450095 469272 450159
rect 469336 450095 469352 450159
rect 469416 450095 469432 450159
rect 469496 450095 469512 450159
rect 469576 450095 469614 450159
rect 468994 434656 469614 450095
rect 468994 434420 469026 434656
rect 469262 434420 469346 434656
rect 469582 434420 469614 434656
rect 468994 434336 469614 434420
rect 468994 434100 469026 434336
rect 469262 434100 469346 434336
rect 469582 434100 469614 434336
rect 468994 431999 469614 434100
rect 468994 431935 469032 431999
rect 469096 431935 469112 431999
rect 469176 431935 469192 431999
rect 469256 431935 469272 431999
rect 469336 431935 469352 431999
rect 469416 431935 469432 431999
rect 469496 431935 469512 431999
rect 469576 431935 469614 431999
rect 468994 431919 469614 431935
rect 468994 431855 469032 431919
rect 469096 431855 469112 431919
rect 469176 431855 469192 431919
rect 469256 431855 469272 431919
rect 469336 431855 469352 431919
rect 469416 431855 469432 431919
rect 469496 431855 469512 431919
rect 469576 431855 469614 431919
rect 468994 431839 469614 431855
rect 468994 431775 469032 431839
rect 469096 431775 469112 431839
rect 469176 431775 469192 431839
rect 469256 431775 469272 431839
rect 469336 431775 469352 431839
rect 469416 431775 469432 431839
rect 469496 431775 469512 431839
rect 469576 431775 469614 431839
rect 468994 431759 469614 431775
rect 468994 431695 469032 431759
rect 469096 431695 469112 431759
rect 469176 431695 469192 431759
rect 469256 431695 469272 431759
rect 469336 431695 469352 431759
rect 469416 431695 469432 431759
rect 469496 431695 469512 431759
rect 469576 431695 469614 431759
rect 468994 411000 469614 431695
rect 468994 410936 469032 411000
rect 469096 410936 469112 411000
rect 469176 410936 469192 411000
rect 469256 410936 469272 411000
rect 469336 410936 469352 411000
rect 469416 410936 469432 411000
rect 469496 410936 469512 411000
rect 469576 410936 469614 411000
rect 468994 410920 469614 410936
rect 468994 410856 469032 410920
rect 469096 410856 469112 410920
rect 469176 410856 469192 410920
rect 469256 410856 469272 410920
rect 469336 410856 469352 410920
rect 469416 410856 469432 410920
rect 469496 410856 469512 410920
rect 469576 410856 469614 410920
rect 468994 410840 469614 410856
rect 468994 410776 469032 410840
rect 469096 410776 469112 410840
rect 469176 410776 469192 410840
rect 469256 410776 469272 410840
rect 469336 410776 469352 410840
rect 469416 410776 469432 410840
rect 469496 410776 469512 410840
rect 469576 410776 469614 410840
rect 468994 410760 469614 410776
rect 468994 410696 469032 410760
rect 469096 410696 469112 410760
rect 469176 410696 469192 410760
rect 469256 410696 469272 410760
rect 469336 410696 469352 410760
rect 469416 410696 469432 410760
rect 469496 410696 469512 410760
rect 469576 410696 469614 410760
rect 468994 398656 469614 410696
rect 468994 398420 469026 398656
rect 469262 398420 469346 398656
rect 469582 398420 469614 398656
rect 468994 398336 469614 398420
rect 468994 398100 469026 398336
rect 469262 398100 469346 398336
rect 469582 398100 469614 398336
rect 468994 390004 469614 398100
rect 468994 389940 469032 390004
rect 469096 389940 469112 390004
rect 469176 389940 469192 390004
rect 469256 389940 469272 390004
rect 469336 389940 469352 390004
rect 469416 389940 469432 390004
rect 469496 389940 469512 390004
rect 469576 389940 469614 390004
rect 468994 389924 469614 389940
rect 468994 389860 469032 389924
rect 469096 389860 469112 389924
rect 469176 389860 469192 389924
rect 469256 389860 469272 389924
rect 469336 389860 469352 389924
rect 469416 389860 469432 389924
rect 469496 389860 469512 389924
rect 469576 389860 469614 389924
rect 468994 389844 469614 389860
rect 468994 389780 469032 389844
rect 469096 389780 469112 389844
rect 469176 389780 469192 389844
rect 469256 389780 469272 389844
rect 469336 389780 469352 389844
rect 469416 389780 469432 389844
rect 469496 389780 469512 389844
rect 469576 389780 469614 389844
rect 468994 389764 469614 389780
rect 468994 389700 469032 389764
rect 469096 389700 469112 389764
rect 469176 389700 469192 389764
rect 469256 389700 469272 389764
rect 469336 389700 469352 389764
rect 469416 389700 469432 389764
rect 469496 389700 469512 389764
rect 469576 389700 469614 389764
rect 468994 362656 469614 389700
rect 468994 362420 469026 362656
rect 469262 362420 469346 362656
rect 469582 362420 469614 362656
rect 468994 362336 469614 362420
rect 468994 362100 469026 362336
rect 469262 362100 469346 362336
rect 469582 362100 469614 362336
rect 468994 357401 469614 362100
rect 468994 357337 469032 357401
rect 469096 357337 469112 357401
rect 469176 357337 469192 357401
rect 469256 357337 469272 357401
rect 469336 357337 469352 357401
rect 469416 357337 469432 357401
rect 469496 357337 469512 357401
rect 469576 357337 469614 357401
rect 468994 357321 469614 357337
rect 468994 357257 469032 357321
rect 469096 357257 469112 357321
rect 469176 357257 469192 357321
rect 469256 357257 469272 357321
rect 469336 357257 469352 357321
rect 469416 357257 469432 357321
rect 469496 357257 469512 357321
rect 469576 357257 469614 357321
rect 468994 357241 469614 357257
rect 468994 357177 469032 357241
rect 469096 357177 469112 357241
rect 469176 357177 469192 357241
rect 469256 357177 469272 357241
rect 469336 357177 469352 357241
rect 469416 357177 469432 357241
rect 469496 357177 469512 357241
rect 469576 357177 469614 357241
rect 468994 357161 469614 357177
rect 468994 357097 469032 357161
rect 469096 357097 469112 357161
rect 469176 357097 469192 357161
rect 469256 357097 469272 357161
rect 469336 357097 469352 357161
rect 469416 357097 469432 357161
rect 469496 357097 469512 357161
rect 469576 357097 469614 357161
rect 468994 341399 469614 357097
rect 468994 341335 469032 341399
rect 469096 341335 469112 341399
rect 469176 341335 469192 341399
rect 469256 341335 469272 341399
rect 469336 341335 469352 341399
rect 469416 341335 469432 341399
rect 469496 341335 469512 341399
rect 469576 341335 469614 341399
rect 468994 341319 469614 341335
rect 468994 341255 469032 341319
rect 469096 341255 469112 341319
rect 469176 341255 469192 341319
rect 469256 341255 469272 341319
rect 469336 341255 469352 341319
rect 469416 341255 469432 341319
rect 469496 341255 469512 341319
rect 469576 341255 469614 341319
rect 468994 341239 469614 341255
rect 468994 341175 469032 341239
rect 469096 341175 469112 341239
rect 469176 341175 469192 341239
rect 469256 341175 469272 341239
rect 469336 341175 469352 341239
rect 469416 341175 469432 341239
rect 469496 341175 469512 341239
rect 469576 341175 469614 341239
rect 468994 341159 469614 341175
rect 468994 341095 469032 341159
rect 469096 341095 469112 341159
rect 469176 341095 469192 341159
rect 469256 341095 469272 341159
rect 469336 341095 469352 341159
rect 469416 341095 469432 341159
rect 469496 341095 469512 341159
rect 469576 341095 469614 341159
rect 468994 326656 469614 341095
rect 468994 326420 469026 326656
rect 469262 326420 469346 326656
rect 469582 326420 469614 326656
rect 468994 326336 469614 326420
rect 468994 326100 469026 326336
rect 469262 326100 469346 326336
rect 469582 326100 469614 326336
rect 468994 321399 469614 326100
rect 468994 321335 469032 321399
rect 469096 321335 469112 321399
rect 469176 321335 469192 321399
rect 469256 321335 469272 321399
rect 469336 321335 469352 321399
rect 469416 321335 469432 321399
rect 469496 321335 469512 321399
rect 469576 321335 469614 321399
rect 468994 321319 469614 321335
rect 468994 321255 469032 321319
rect 469096 321255 469112 321319
rect 469176 321255 469192 321319
rect 469256 321255 469272 321319
rect 469336 321255 469352 321319
rect 469416 321255 469432 321319
rect 469496 321255 469512 321319
rect 469576 321255 469614 321319
rect 468994 321239 469614 321255
rect 468994 321175 469032 321239
rect 469096 321175 469112 321239
rect 469176 321175 469192 321239
rect 469256 321175 469272 321239
rect 469336 321175 469352 321239
rect 469416 321175 469432 321239
rect 469496 321175 469512 321239
rect 469576 321175 469614 321239
rect 468994 321159 469614 321175
rect 468994 321095 469032 321159
rect 469096 321095 469112 321159
rect 469176 321095 469192 321159
rect 469256 321095 469272 321159
rect 469336 321095 469352 321159
rect 469416 321095 469432 321159
rect 469496 321095 469512 321159
rect 469576 321095 469614 321159
rect 468994 306001 469614 321095
rect 468994 305937 469032 306001
rect 469096 305937 469112 306001
rect 469176 305937 469192 306001
rect 469256 305937 469272 306001
rect 469336 305937 469352 306001
rect 469416 305937 469432 306001
rect 469496 305937 469512 306001
rect 469576 305937 469614 306001
rect 468994 305921 469614 305937
rect 468994 305857 469032 305921
rect 469096 305857 469112 305921
rect 469176 305857 469192 305921
rect 469256 305857 469272 305921
rect 469336 305857 469352 305921
rect 469416 305857 469432 305921
rect 469496 305857 469512 305921
rect 469576 305857 469614 305921
rect 468994 305841 469614 305857
rect 468994 305777 469032 305841
rect 469096 305777 469112 305841
rect 469176 305777 469192 305841
rect 469256 305777 469272 305841
rect 469336 305777 469352 305841
rect 469416 305777 469432 305841
rect 469496 305777 469512 305841
rect 469576 305777 469614 305841
rect 468994 305761 469614 305777
rect 468994 305697 469032 305761
rect 469096 305697 469112 305761
rect 469176 305697 469192 305761
rect 469256 305697 469272 305761
rect 469336 305697 469352 305761
rect 469416 305697 469432 305761
rect 469496 305697 469512 305761
rect 469576 305697 469614 305761
rect 468994 290656 469614 305697
rect 468994 290420 469026 290656
rect 469262 290420 469346 290656
rect 469582 290420 469614 290656
rect 468994 290336 469614 290420
rect 468994 290100 469026 290336
rect 469262 290100 469346 290336
rect 469582 290100 469614 290336
rect 468994 286402 469614 290100
rect 468994 286338 469032 286402
rect 469096 286338 469112 286402
rect 469176 286338 469192 286402
rect 469256 286338 469272 286402
rect 469336 286338 469352 286402
rect 469416 286338 469432 286402
rect 469496 286338 469512 286402
rect 469576 286338 469614 286402
rect 468994 286322 469614 286338
rect 468994 286258 469032 286322
rect 469096 286258 469112 286322
rect 469176 286258 469192 286322
rect 469256 286258 469272 286322
rect 469336 286258 469352 286322
rect 469416 286258 469432 286322
rect 469496 286258 469512 286322
rect 469576 286258 469614 286322
rect 468994 286242 469614 286258
rect 468994 286178 469032 286242
rect 469096 286178 469112 286242
rect 469176 286178 469192 286242
rect 469256 286178 469272 286242
rect 469336 286178 469352 286242
rect 469416 286178 469432 286242
rect 469496 286178 469512 286242
rect 469576 286178 469614 286242
rect 468994 286162 469614 286178
rect 468994 286098 469032 286162
rect 469096 286098 469112 286162
rect 469176 286098 469192 286162
rect 469256 286098 469272 286162
rect 469336 286098 469352 286162
rect 469416 286098 469432 286162
rect 469496 286098 469512 286162
rect 469576 286098 469614 286162
rect 468994 266401 469614 286098
rect 468994 266337 469032 266401
rect 469096 266337 469112 266401
rect 469176 266337 469192 266401
rect 469256 266337 469272 266401
rect 469336 266337 469352 266401
rect 469416 266337 469432 266401
rect 469496 266337 469512 266401
rect 469576 266337 469614 266401
rect 468994 266321 469614 266337
rect 468994 266257 469032 266321
rect 469096 266257 469112 266321
rect 469176 266257 469192 266321
rect 469256 266257 469272 266321
rect 469336 266257 469352 266321
rect 469416 266257 469432 266321
rect 469496 266257 469512 266321
rect 469576 266257 469614 266321
rect 468994 266241 469614 266257
rect 468994 266177 469032 266241
rect 469096 266177 469112 266241
rect 469176 266177 469192 266241
rect 469256 266177 469272 266241
rect 469336 266177 469352 266241
rect 469416 266177 469432 266241
rect 469496 266177 469512 266241
rect 469576 266177 469614 266241
rect 468994 266161 469614 266177
rect 468994 266097 469032 266161
rect 469096 266097 469112 266161
rect 469176 266097 469192 266161
rect 469256 266097 469272 266161
rect 469336 266097 469352 266161
rect 469416 266097 469432 266161
rect 469496 266097 469512 266161
rect 469576 266097 469614 266161
rect 468994 254656 469614 266097
rect 468994 254420 469026 254656
rect 469262 254420 469346 254656
rect 469582 254420 469614 254656
rect 468994 254336 469614 254420
rect 468994 254100 469026 254336
rect 469262 254100 469346 254336
rect 469582 254100 469614 254336
rect 468994 218656 469614 254100
rect 468994 218420 469026 218656
rect 469262 218420 469346 218656
rect 469582 218420 469614 218656
rect 468994 218336 469614 218420
rect 468994 218100 469026 218336
rect 469262 218100 469346 218336
rect 469582 218100 469614 218336
rect 468994 182656 469614 218100
rect 468994 182420 469026 182656
rect 469262 182420 469346 182656
rect 469582 182420 469614 182656
rect 468994 182336 469614 182420
rect 468994 182100 469026 182336
rect 469262 182100 469346 182336
rect 469582 182100 469614 182336
rect 468994 146656 469614 182100
rect 468994 146420 469026 146656
rect 469262 146420 469346 146656
rect 469582 146420 469614 146656
rect 468994 146336 469614 146420
rect 468994 146100 469026 146336
rect 469262 146100 469346 146336
rect 469582 146100 469614 146336
rect 468994 110656 469614 146100
rect 468994 110420 469026 110656
rect 469262 110420 469346 110656
rect 469582 110420 469614 110656
rect 468994 110336 469614 110420
rect 468994 110100 469026 110336
rect 469262 110100 469346 110336
rect 469582 110100 469614 110336
rect 468994 74656 469614 110100
rect 468994 74420 469026 74656
rect 469262 74420 469346 74656
rect 469582 74420 469614 74656
rect 468994 74336 469614 74420
rect 468994 74100 469026 74336
rect 469262 74100 469346 74336
rect 469582 74100 469614 74336
rect 468994 38656 469614 74100
rect 468994 38420 469026 38656
rect 469262 38420 469346 38656
rect 469582 38420 469614 38656
rect 468994 38336 469614 38420
rect 468994 38100 469026 38336
rect 469262 38100 469346 38336
rect 469582 38100 469614 38336
rect 468994 2656 469614 38100
rect 468994 2420 469026 2656
rect 469262 2420 469346 2656
rect 469582 2420 469614 2656
rect 468994 2336 469614 2420
rect 468994 2100 469026 2336
rect 469262 2100 469346 2336
rect 469582 2100 469614 2336
rect 468994 -344 469614 2100
rect 468994 -580 469026 -344
rect 469262 -580 469346 -344
rect 469582 -580 469614 -344
rect 468994 -664 469614 -580
rect 468994 -900 469026 -664
rect 469262 -900 469346 -664
rect 469582 -900 469614 -664
rect 468994 -7652 469614 -900
rect 470234 705800 470854 711592
rect 470234 705564 470266 705800
rect 470502 705564 470586 705800
rect 470822 705564 470854 705800
rect 470234 705480 470854 705564
rect 470234 705244 470266 705480
rect 470502 705244 470586 705480
rect 470822 705244 470854 705480
rect 470234 687896 470854 705244
rect 470234 687660 470266 687896
rect 470502 687660 470586 687896
rect 470822 687660 470854 687896
rect 470234 687576 470854 687660
rect 470234 687340 470266 687576
rect 470502 687340 470586 687576
rect 470822 687340 470854 687576
rect 470234 651896 470854 687340
rect 470234 651660 470266 651896
rect 470502 651660 470586 651896
rect 470822 651660 470854 651896
rect 470234 651576 470854 651660
rect 470234 651340 470266 651576
rect 470502 651340 470586 651576
rect 470822 651340 470854 651576
rect 470234 615896 470854 651340
rect 470234 615660 470266 615896
rect 470502 615660 470586 615896
rect 470822 615660 470854 615896
rect 470234 615576 470854 615660
rect 470234 615340 470266 615576
rect 470502 615340 470586 615576
rect 470822 615340 470854 615576
rect 470234 579896 470854 615340
rect 470234 579660 470266 579896
rect 470502 579660 470586 579896
rect 470822 579660 470854 579896
rect 470234 579576 470854 579660
rect 470234 579340 470266 579576
rect 470502 579340 470586 579576
rect 470822 579340 470854 579576
rect 470234 543896 470854 579340
rect 470234 543660 470266 543896
rect 470502 543660 470586 543896
rect 470822 543660 470854 543896
rect 470234 543576 470854 543660
rect 470234 543340 470266 543576
rect 470502 543340 470586 543576
rect 470822 543340 470854 543576
rect 470234 507896 470854 543340
rect 470234 507660 470266 507896
rect 470502 507660 470586 507896
rect 470822 507660 470854 507896
rect 470234 507576 470854 507660
rect 470234 507340 470266 507576
rect 470502 507340 470586 507576
rect 470822 507340 470854 507576
rect 470234 471896 470854 507340
rect 470234 471660 470266 471896
rect 470502 471660 470586 471896
rect 470822 471660 470854 471896
rect 470234 471576 470854 471660
rect 470234 471340 470266 471576
rect 470502 471340 470586 471576
rect 470822 471340 470854 471576
rect 470234 451485 470854 471340
rect 470234 451421 470272 451485
rect 470336 451421 470352 451485
rect 470416 451421 470432 451485
rect 470496 451421 470512 451485
rect 470576 451421 470592 451485
rect 470656 451421 470672 451485
rect 470736 451421 470752 451485
rect 470816 451421 470854 451485
rect 470234 451405 470854 451421
rect 470234 451341 470272 451405
rect 470336 451341 470352 451405
rect 470416 451341 470432 451405
rect 470496 451341 470512 451405
rect 470576 451341 470592 451405
rect 470656 451341 470672 451405
rect 470736 451341 470752 451405
rect 470816 451341 470854 451405
rect 470234 451325 470854 451341
rect 470234 451261 470272 451325
rect 470336 451261 470352 451325
rect 470416 451261 470432 451325
rect 470496 451261 470512 451325
rect 470576 451261 470592 451325
rect 470656 451261 470672 451325
rect 470736 451261 470752 451325
rect 470816 451261 470854 451325
rect 470234 451245 470854 451261
rect 470234 451181 470272 451245
rect 470336 451181 470352 451245
rect 470416 451181 470432 451245
rect 470496 451181 470512 451245
rect 470576 451181 470592 451245
rect 470656 451181 470672 451245
rect 470736 451181 470752 451245
rect 470816 451181 470854 451245
rect 470234 449314 470854 451181
rect 470234 449250 470272 449314
rect 470336 449250 470352 449314
rect 470416 449250 470432 449314
rect 470496 449250 470512 449314
rect 470576 449250 470592 449314
rect 470656 449250 470672 449314
rect 470736 449250 470752 449314
rect 470816 449250 470854 449314
rect 470234 449234 470854 449250
rect 470234 449170 470272 449234
rect 470336 449170 470352 449234
rect 470416 449170 470432 449234
rect 470496 449170 470512 449234
rect 470576 449170 470592 449234
rect 470656 449170 470672 449234
rect 470736 449170 470752 449234
rect 470816 449170 470854 449234
rect 470234 449154 470854 449170
rect 470234 449090 470272 449154
rect 470336 449090 470352 449154
rect 470416 449090 470432 449154
rect 470496 449090 470512 449154
rect 470576 449090 470592 449154
rect 470656 449090 470672 449154
rect 470736 449090 470752 449154
rect 470816 449090 470854 449154
rect 470234 449074 470854 449090
rect 470234 449010 470272 449074
rect 470336 449010 470352 449074
rect 470416 449010 470432 449074
rect 470496 449010 470512 449074
rect 470576 449010 470592 449074
rect 470656 449010 470672 449074
rect 470736 449010 470752 449074
rect 470816 449010 470854 449074
rect 470234 435896 470854 449010
rect 470234 435660 470266 435896
rect 470502 435660 470586 435896
rect 470822 435660 470854 435896
rect 470234 435576 470854 435660
rect 470234 435340 470266 435576
rect 470502 435340 470586 435576
rect 470822 435340 470854 435576
rect 470234 433086 470854 435340
rect 470234 433022 470272 433086
rect 470336 433022 470352 433086
rect 470416 433022 470432 433086
rect 470496 433022 470512 433086
rect 470576 433022 470592 433086
rect 470656 433022 470672 433086
rect 470736 433022 470752 433086
rect 470816 433022 470854 433086
rect 470234 433006 470854 433022
rect 470234 432942 470272 433006
rect 470336 432942 470352 433006
rect 470416 432942 470432 433006
rect 470496 432942 470512 433006
rect 470576 432942 470592 433006
rect 470656 432942 470672 433006
rect 470736 432942 470752 433006
rect 470816 432942 470854 433006
rect 470234 432926 470854 432942
rect 470234 432862 470272 432926
rect 470336 432862 470352 432926
rect 470416 432862 470432 432926
rect 470496 432862 470512 432926
rect 470576 432862 470592 432926
rect 470656 432862 470672 432926
rect 470736 432862 470752 432926
rect 470816 432862 470854 432926
rect 470234 432846 470854 432862
rect 470234 432782 470272 432846
rect 470336 432782 470352 432846
rect 470416 432782 470432 432846
rect 470496 432782 470512 432846
rect 470576 432782 470592 432846
rect 470656 432782 470672 432846
rect 470736 432782 470752 432846
rect 470816 432782 470854 432846
rect 470234 430914 470854 432782
rect 470234 430850 470272 430914
rect 470336 430850 470352 430914
rect 470416 430850 470432 430914
rect 470496 430850 470512 430914
rect 470576 430850 470592 430914
rect 470656 430850 470672 430914
rect 470736 430850 470752 430914
rect 470816 430850 470854 430914
rect 470234 430834 470854 430850
rect 470234 430770 470272 430834
rect 470336 430770 470352 430834
rect 470416 430770 470432 430834
rect 470496 430770 470512 430834
rect 470576 430770 470592 430834
rect 470656 430770 470672 430834
rect 470736 430770 470752 430834
rect 470816 430770 470854 430834
rect 470234 430754 470854 430770
rect 470234 430690 470272 430754
rect 470336 430690 470352 430754
rect 470416 430690 470432 430754
rect 470496 430690 470512 430754
rect 470576 430690 470592 430754
rect 470656 430690 470672 430754
rect 470736 430690 470752 430754
rect 470816 430690 470854 430754
rect 470234 430674 470854 430690
rect 470234 430610 470272 430674
rect 470336 430610 470352 430674
rect 470416 430610 470432 430674
rect 470496 430610 470512 430674
rect 470576 430610 470592 430674
rect 470656 430610 470672 430674
rect 470736 430610 470752 430674
rect 470816 430610 470854 430674
rect 470234 412086 470854 430610
rect 470234 412022 470272 412086
rect 470336 412022 470352 412086
rect 470416 412022 470432 412086
rect 470496 412022 470512 412086
rect 470576 412022 470592 412086
rect 470656 412022 470672 412086
rect 470736 412022 470752 412086
rect 470816 412022 470854 412086
rect 470234 412006 470854 412022
rect 470234 411942 470272 412006
rect 470336 411942 470352 412006
rect 470416 411942 470432 412006
rect 470496 411942 470512 412006
rect 470576 411942 470592 412006
rect 470656 411942 470672 412006
rect 470736 411942 470752 412006
rect 470816 411942 470854 412006
rect 470234 411926 470854 411942
rect 470234 411862 470272 411926
rect 470336 411862 470352 411926
rect 470416 411862 470432 411926
rect 470496 411862 470512 411926
rect 470576 411862 470592 411926
rect 470656 411862 470672 411926
rect 470736 411862 470752 411926
rect 470816 411862 470854 411926
rect 470234 411846 470854 411862
rect 470234 411782 470272 411846
rect 470336 411782 470352 411846
rect 470416 411782 470432 411846
rect 470496 411782 470512 411846
rect 470576 411782 470592 411846
rect 470656 411782 470672 411846
rect 470736 411782 470752 411846
rect 470816 411782 470854 411846
rect 470234 409914 470854 411782
rect 470234 409850 470272 409914
rect 470336 409850 470352 409914
rect 470416 409850 470432 409914
rect 470496 409850 470512 409914
rect 470576 409850 470592 409914
rect 470656 409850 470672 409914
rect 470736 409850 470752 409914
rect 470816 409850 470854 409914
rect 470234 409834 470854 409850
rect 470234 409770 470272 409834
rect 470336 409770 470352 409834
rect 470416 409770 470432 409834
rect 470496 409770 470512 409834
rect 470576 409770 470592 409834
rect 470656 409770 470672 409834
rect 470736 409770 470752 409834
rect 470816 409770 470854 409834
rect 470234 409754 470854 409770
rect 470234 409690 470272 409754
rect 470336 409690 470352 409754
rect 470416 409690 470432 409754
rect 470496 409690 470512 409754
rect 470576 409690 470592 409754
rect 470656 409690 470672 409754
rect 470736 409690 470752 409754
rect 470816 409690 470854 409754
rect 470234 409674 470854 409690
rect 470234 409610 470272 409674
rect 470336 409610 470352 409674
rect 470416 409610 470432 409674
rect 470496 409610 470512 409674
rect 470576 409610 470592 409674
rect 470656 409610 470672 409674
rect 470736 409610 470752 409674
rect 470816 409610 470854 409674
rect 470234 399896 470854 409610
rect 470234 399660 470266 399896
rect 470502 399660 470586 399896
rect 470822 399660 470854 399896
rect 470234 399576 470854 399660
rect 470234 399340 470266 399576
rect 470502 399340 470586 399576
rect 470822 399340 470854 399576
rect 470234 391087 470854 399340
rect 470234 391023 470272 391087
rect 470336 391023 470352 391087
rect 470416 391023 470432 391087
rect 470496 391023 470512 391087
rect 470576 391023 470592 391087
rect 470656 391023 470672 391087
rect 470736 391023 470752 391087
rect 470816 391023 470854 391087
rect 470234 391007 470854 391023
rect 470234 390943 470272 391007
rect 470336 390943 470352 391007
rect 470416 390943 470432 391007
rect 470496 390943 470512 391007
rect 470576 390943 470592 391007
rect 470656 390943 470672 391007
rect 470736 390943 470752 391007
rect 470816 390943 470854 391007
rect 470234 390927 470854 390943
rect 470234 390863 470272 390927
rect 470336 390863 470352 390927
rect 470416 390863 470432 390927
rect 470496 390863 470512 390927
rect 470576 390863 470592 390927
rect 470656 390863 470672 390927
rect 470736 390863 470752 390927
rect 470816 390863 470854 390927
rect 470234 390847 470854 390863
rect 470234 390783 470272 390847
rect 470336 390783 470352 390847
rect 470416 390783 470432 390847
rect 470496 390783 470512 390847
rect 470576 390783 470592 390847
rect 470656 390783 470672 390847
rect 470736 390783 470752 390847
rect 470816 390783 470854 390847
rect 470234 388914 470854 390783
rect 470234 388850 470272 388914
rect 470336 388850 470352 388914
rect 470416 388850 470432 388914
rect 470496 388850 470512 388914
rect 470576 388850 470592 388914
rect 470656 388850 470672 388914
rect 470736 388850 470752 388914
rect 470816 388850 470854 388914
rect 470234 388834 470854 388850
rect 470234 388770 470272 388834
rect 470336 388770 470352 388834
rect 470416 388770 470432 388834
rect 470496 388770 470512 388834
rect 470576 388770 470592 388834
rect 470656 388770 470672 388834
rect 470736 388770 470752 388834
rect 470816 388770 470854 388834
rect 470234 388754 470854 388770
rect 470234 388690 470272 388754
rect 470336 388690 470352 388754
rect 470416 388690 470432 388754
rect 470496 388690 470512 388754
rect 470576 388690 470592 388754
rect 470656 388690 470672 388754
rect 470736 388690 470752 388754
rect 470816 388690 470854 388754
rect 470234 388674 470854 388690
rect 470234 388610 470272 388674
rect 470336 388610 470352 388674
rect 470416 388610 470432 388674
rect 470496 388610 470512 388674
rect 470576 388610 470592 388674
rect 470656 388610 470672 388674
rect 470736 388610 470752 388674
rect 470816 388610 470854 388674
rect 470234 363896 470854 388610
rect 470234 363660 470266 363896
rect 470502 363660 470586 363896
rect 470822 363660 470854 363896
rect 470234 363576 470854 363660
rect 470234 363340 470266 363576
rect 470502 363340 470586 363576
rect 470822 363340 470854 363576
rect 470234 358487 470854 363340
rect 470234 358423 470272 358487
rect 470336 358423 470352 358487
rect 470416 358423 470432 358487
rect 470496 358423 470512 358487
rect 470576 358423 470592 358487
rect 470656 358423 470672 358487
rect 470736 358423 470752 358487
rect 470816 358423 470854 358487
rect 470234 358407 470854 358423
rect 470234 358343 470272 358407
rect 470336 358343 470352 358407
rect 470416 358343 470432 358407
rect 470496 358343 470512 358407
rect 470576 358343 470592 358407
rect 470656 358343 470672 358407
rect 470736 358343 470752 358407
rect 470816 358343 470854 358407
rect 470234 358327 470854 358343
rect 470234 358263 470272 358327
rect 470336 358263 470352 358327
rect 470416 358263 470432 358327
rect 470496 358263 470512 358327
rect 470576 358263 470592 358327
rect 470656 358263 470672 358327
rect 470736 358263 470752 358327
rect 470816 358263 470854 358327
rect 470234 358247 470854 358263
rect 470234 358183 470272 358247
rect 470336 358183 470352 358247
rect 470416 358183 470432 358247
rect 470496 358183 470512 358247
rect 470576 358183 470592 358247
rect 470656 358183 470672 358247
rect 470736 358183 470752 358247
rect 470816 358183 470854 358247
rect 470234 356314 470854 358183
rect 470234 356250 470272 356314
rect 470336 356250 470352 356314
rect 470416 356250 470432 356314
rect 470496 356250 470512 356314
rect 470576 356250 470592 356314
rect 470656 356250 470672 356314
rect 470736 356250 470752 356314
rect 470816 356250 470854 356314
rect 470234 356234 470854 356250
rect 470234 356170 470272 356234
rect 470336 356170 470352 356234
rect 470416 356170 470432 356234
rect 470496 356170 470512 356234
rect 470576 356170 470592 356234
rect 470656 356170 470672 356234
rect 470736 356170 470752 356234
rect 470816 356170 470854 356234
rect 470234 356154 470854 356170
rect 470234 356090 470272 356154
rect 470336 356090 470352 356154
rect 470416 356090 470432 356154
rect 470496 356090 470512 356154
rect 470576 356090 470592 356154
rect 470656 356090 470672 356154
rect 470736 356090 470752 356154
rect 470816 356090 470854 356154
rect 470234 356074 470854 356090
rect 470234 356010 470272 356074
rect 470336 356010 470352 356074
rect 470416 356010 470432 356074
rect 470496 356010 470512 356074
rect 470576 356010 470592 356074
rect 470656 356010 470672 356074
rect 470736 356010 470752 356074
rect 470816 356010 470854 356074
rect 470234 342486 470854 356010
rect 470234 342422 470272 342486
rect 470336 342422 470352 342486
rect 470416 342422 470432 342486
rect 470496 342422 470512 342486
rect 470576 342422 470592 342486
rect 470656 342422 470672 342486
rect 470736 342422 470752 342486
rect 470816 342422 470854 342486
rect 470234 342406 470854 342422
rect 470234 342342 470272 342406
rect 470336 342342 470352 342406
rect 470416 342342 470432 342406
rect 470496 342342 470512 342406
rect 470576 342342 470592 342406
rect 470656 342342 470672 342406
rect 470736 342342 470752 342406
rect 470816 342342 470854 342406
rect 470234 342326 470854 342342
rect 470234 342262 470272 342326
rect 470336 342262 470352 342326
rect 470416 342262 470432 342326
rect 470496 342262 470512 342326
rect 470576 342262 470592 342326
rect 470656 342262 470672 342326
rect 470736 342262 470752 342326
rect 470816 342262 470854 342326
rect 470234 342246 470854 342262
rect 470234 342182 470272 342246
rect 470336 342182 470352 342246
rect 470416 342182 470432 342246
rect 470496 342182 470512 342246
rect 470576 342182 470592 342246
rect 470656 342182 470672 342246
rect 470736 342182 470752 342246
rect 470816 342182 470854 342246
rect 470234 340314 470854 342182
rect 470234 340250 470272 340314
rect 470336 340250 470352 340314
rect 470416 340250 470432 340314
rect 470496 340250 470512 340314
rect 470576 340250 470592 340314
rect 470656 340250 470672 340314
rect 470736 340250 470752 340314
rect 470816 340250 470854 340314
rect 470234 340234 470854 340250
rect 470234 340170 470272 340234
rect 470336 340170 470352 340234
rect 470416 340170 470432 340234
rect 470496 340170 470512 340234
rect 470576 340170 470592 340234
rect 470656 340170 470672 340234
rect 470736 340170 470752 340234
rect 470816 340170 470854 340234
rect 470234 340154 470854 340170
rect 470234 340090 470272 340154
rect 470336 340090 470352 340154
rect 470416 340090 470432 340154
rect 470496 340090 470512 340154
rect 470576 340090 470592 340154
rect 470656 340090 470672 340154
rect 470736 340090 470752 340154
rect 470816 340090 470854 340154
rect 470234 340074 470854 340090
rect 470234 340010 470272 340074
rect 470336 340010 470352 340074
rect 470416 340010 470432 340074
rect 470496 340010 470512 340074
rect 470576 340010 470592 340074
rect 470656 340010 470672 340074
rect 470736 340010 470752 340074
rect 470816 340010 470854 340074
rect 470234 327896 470854 340010
rect 470234 327660 470266 327896
rect 470502 327660 470586 327896
rect 470822 327660 470854 327896
rect 470234 327576 470854 327660
rect 470234 327340 470266 327576
rect 470502 327340 470586 327576
rect 470822 327340 470854 327576
rect 470234 322486 470854 327340
rect 470234 322422 470272 322486
rect 470336 322422 470352 322486
rect 470416 322422 470432 322486
rect 470496 322422 470512 322486
rect 470576 322422 470592 322486
rect 470656 322422 470672 322486
rect 470736 322422 470752 322486
rect 470816 322422 470854 322486
rect 470234 322406 470854 322422
rect 470234 322342 470272 322406
rect 470336 322342 470352 322406
rect 470416 322342 470432 322406
rect 470496 322342 470512 322406
rect 470576 322342 470592 322406
rect 470656 322342 470672 322406
rect 470736 322342 470752 322406
rect 470816 322342 470854 322406
rect 470234 322326 470854 322342
rect 470234 322262 470272 322326
rect 470336 322262 470352 322326
rect 470416 322262 470432 322326
rect 470496 322262 470512 322326
rect 470576 322262 470592 322326
rect 470656 322262 470672 322326
rect 470736 322262 470752 322326
rect 470816 322262 470854 322326
rect 470234 322246 470854 322262
rect 470234 322182 470272 322246
rect 470336 322182 470352 322246
rect 470416 322182 470432 322246
rect 470496 322182 470512 322246
rect 470576 322182 470592 322246
rect 470656 322182 470672 322246
rect 470736 322182 470752 322246
rect 470816 322182 470854 322246
rect 470234 320314 470854 322182
rect 470234 320250 470272 320314
rect 470336 320250 470352 320314
rect 470416 320250 470432 320314
rect 470496 320250 470512 320314
rect 470576 320250 470592 320314
rect 470656 320250 470672 320314
rect 470736 320250 470752 320314
rect 470816 320250 470854 320314
rect 470234 320234 470854 320250
rect 470234 320170 470272 320234
rect 470336 320170 470352 320234
rect 470416 320170 470432 320234
rect 470496 320170 470512 320234
rect 470576 320170 470592 320234
rect 470656 320170 470672 320234
rect 470736 320170 470752 320234
rect 470816 320170 470854 320234
rect 470234 320154 470854 320170
rect 470234 320090 470272 320154
rect 470336 320090 470352 320154
rect 470416 320090 470432 320154
rect 470496 320090 470512 320154
rect 470576 320090 470592 320154
rect 470656 320090 470672 320154
rect 470736 320090 470752 320154
rect 470816 320090 470854 320154
rect 470234 320074 470854 320090
rect 470234 320010 470272 320074
rect 470336 320010 470352 320074
rect 470416 320010 470432 320074
rect 470496 320010 470512 320074
rect 470576 320010 470592 320074
rect 470656 320010 470672 320074
rect 470736 320010 470752 320074
rect 470816 320010 470854 320074
rect 470234 307086 470854 320010
rect 470234 307022 470272 307086
rect 470336 307022 470352 307086
rect 470416 307022 470432 307086
rect 470496 307022 470512 307086
rect 470576 307022 470592 307086
rect 470656 307022 470672 307086
rect 470736 307022 470752 307086
rect 470816 307022 470854 307086
rect 470234 307006 470854 307022
rect 470234 306942 470272 307006
rect 470336 306942 470352 307006
rect 470416 306942 470432 307006
rect 470496 306942 470512 307006
rect 470576 306942 470592 307006
rect 470656 306942 470672 307006
rect 470736 306942 470752 307006
rect 470816 306942 470854 307006
rect 470234 306926 470854 306942
rect 470234 306862 470272 306926
rect 470336 306862 470352 306926
rect 470416 306862 470432 306926
rect 470496 306862 470512 306926
rect 470576 306862 470592 306926
rect 470656 306862 470672 306926
rect 470736 306862 470752 306926
rect 470816 306862 470854 306926
rect 470234 306846 470854 306862
rect 470234 306782 470272 306846
rect 470336 306782 470352 306846
rect 470416 306782 470432 306846
rect 470496 306782 470512 306846
rect 470576 306782 470592 306846
rect 470656 306782 470672 306846
rect 470736 306782 470752 306846
rect 470816 306782 470854 306846
rect 470234 304914 470854 306782
rect 470234 304850 470272 304914
rect 470336 304850 470352 304914
rect 470416 304850 470432 304914
rect 470496 304850 470512 304914
rect 470576 304850 470592 304914
rect 470656 304850 470672 304914
rect 470736 304850 470752 304914
rect 470816 304850 470854 304914
rect 470234 304834 470854 304850
rect 470234 304770 470272 304834
rect 470336 304770 470352 304834
rect 470416 304770 470432 304834
rect 470496 304770 470512 304834
rect 470576 304770 470592 304834
rect 470656 304770 470672 304834
rect 470736 304770 470752 304834
rect 470816 304770 470854 304834
rect 470234 304754 470854 304770
rect 470234 304690 470272 304754
rect 470336 304690 470352 304754
rect 470416 304690 470432 304754
rect 470496 304690 470512 304754
rect 470576 304690 470592 304754
rect 470656 304690 470672 304754
rect 470736 304690 470752 304754
rect 470816 304690 470854 304754
rect 470234 304674 470854 304690
rect 470234 304610 470272 304674
rect 470336 304610 470352 304674
rect 470416 304610 470432 304674
rect 470496 304610 470512 304674
rect 470576 304610 470592 304674
rect 470656 304610 470672 304674
rect 470736 304610 470752 304674
rect 470816 304610 470854 304674
rect 470234 291896 470854 304610
rect 470234 291660 470266 291896
rect 470502 291660 470586 291896
rect 470822 291660 470854 291896
rect 470234 291576 470854 291660
rect 470234 291340 470266 291576
rect 470502 291340 470586 291576
rect 470822 291340 470854 291576
rect 470234 287487 470854 291340
rect 470234 287423 470272 287487
rect 470336 287423 470352 287487
rect 470416 287423 470432 287487
rect 470496 287423 470512 287487
rect 470576 287423 470592 287487
rect 470656 287423 470672 287487
rect 470736 287423 470752 287487
rect 470816 287423 470854 287487
rect 470234 287407 470854 287423
rect 470234 287343 470272 287407
rect 470336 287343 470352 287407
rect 470416 287343 470432 287407
rect 470496 287343 470512 287407
rect 470576 287343 470592 287407
rect 470656 287343 470672 287407
rect 470736 287343 470752 287407
rect 470816 287343 470854 287407
rect 470234 287327 470854 287343
rect 470234 287263 470272 287327
rect 470336 287263 470352 287327
rect 470416 287263 470432 287327
rect 470496 287263 470512 287327
rect 470576 287263 470592 287327
rect 470656 287263 470672 287327
rect 470736 287263 470752 287327
rect 470816 287263 470854 287327
rect 470234 287247 470854 287263
rect 470234 287183 470272 287247
rect 470336 287183 470352 287247
rect 470416 287183 470432 287247
rect 470496 287183 470512 287247
rect 470576 287183 470592 287247
rect 470656 287183 470672 287247
rect 470736 287183 470752 287247
rect 470816 287183 470854 287247
rect 470234 285314 470854 287183
rect 470234 285250 470272 285314
rect 470336 285250 470352 285314
rect 470416 285250 470432 285314
rect 470496 285250 470512 285314
rect 470576 285250 470592 285314
rect 470656 285250 470672 285314
rect 470736 285250 470752 285314
rect 470816 285250 470854 285314
rect 470234 285234 470854 285250
rect 470234 285170 470272 285234
rect 470336 285170 470352 285234
rect 470416 285170 470432 285234
rect 470496 285170 470512 285234
rect 470576 285170 470592 285234
rect 470656 285170 470672 285234
rect 470736 285170 470752 285234
rect 470816 285170 470854 285234
rect 470234 285154 470854 285170
rect 470234 285090 470272 285154
rect 470336 285090 470352 285154
rect 470416 285090 470432 285154
rect 470496 285090 470512 285154
rect 470576 285090 470592 285154
rect 470656 285090 470672 285154
rect 470736 285090 470752 285154
rect 470816 285090 470854 285154
rect 470234 285074 470854 285090
rect 470234 285010 470272 285074
rect 470336 285010 470352 285074
rect 470416 285010 470432 285074
rect 470496 285010 470512 285074
rect 470576 285010 470592 285074
rect 470656 285010 470672 285074
rect 470736 285010 470752 285074
rect 470816 285010 470854 285074
rect 470234 267487 470854 285010
rect 470234 267423 470272 267487
rect 470336 267423 470352 267487
rect 470416 267423 470432 267487
rect 470496 267423 470512 267487
rect 470576 267423 470592 267487
rect 470656 267423 470672 267487
rect 470736 267423 470752 267487
rect 470816 267423 470854 267487
rect 470234 267407 470854 267423
rect 470234 267343 470272 267407
rect 470336 267343 470352 267407
rect 470416 267343 470432 267407
rect 470496 267343 470512 267407
rect 470576 267343 470592 267407
rect 470656 267343 470672 267407
rect 470736 267343 470752 267407
rect 470816 267343 470854 267407
rect 470234 267327 470854 267343
rect 470234 267263 470272 267327
rect 470336 267263 470352 267327
rect 470416 267263 470432 267327
rect 470496 267263 470512 267327
rect 470576 267263 470592 267327
rect 470656 267263 470672 267327
rect 470736 267263 470752 267327
rect 470816 267263 470854 267327
rect 470234 267247 470854 267263
rect 470234 267183 470272 267247
rect 470336 267183 470352 267247
rect 470416 267183 470432 267247
rect 470496 267183 470512 267247
rect 470576 267183 470592 267247
rect 470656 267183 470672 267247
rect 470736 267183 470752 267247
rect 470816 267183 470854 267247
rect 470234 265314 470854 267183
rect 470234 265250 470272 265314
rect 470336 265250 470352 265314
rect 470416 265250 470432 265314
rect 470496 265250 470512 265314
rect 470576 265250 470592 265314
rect 470656 265250 470672 265314
rect 470736 265250 470752 265314
rect 470816 265250 470854 265314
rect 470234 265234 470854 265250
rect 470234 265170 470272 265234
rect 470336 265170 470352 265234
rect 470416 265170 470432 265234
rect 470496 265170 470512 265234
rect 470576 265170 470592 265234
rect 470656 265170 470672 265234
rect 470736 265170 470752 265234
rect 470816 265170 470854 265234
rect 470234 265154 470854 265170
rect 470234 265090 470272 265154
rect 470336 265090 470352 265154
rect 470416 265090 470432 265154
rect 470496 265090 470512 265154
rect 470576 265090 470592 265154
rect 470656 265090 470672 265154
rect 470736 265090 470752 265154
rect 470816 265090 470854 265154
rect 470234 265074 470854 265090
rect 470234 265010 470272 265074
rect 470336 265010 470352 265074
rect 470416 265010 470432 265074
rect 470496 265010 470512 265074
rect 470576 265010 470592 265074
rect 470656 265010 470672 265074
rect 470736 265010 470752 265074
rect 470816 265010 470854 265074
rect 470234 255896 470854 265010
rect 470234 255660 470266 255896
rect 470502 255660 470586 255896
rect 470822 255660 470854 255896
rect 470234 255576 470854 255660
rect 470234 255340 470266 255576
rect 470502 255340 470586 255576
rect 470822 255340 470854 255576
rect 470234 219896 470854 255340
rect 470234 219660 470266 219896
rect 470502 219660 470586 219896
rect 470822 219660 470854 219896
rect 470234 219576 470854 219660
rect 470234 219340 470266 219576
rect 470502 219340 470586 219576
rect 470822 219340 470854 219576
rect 470234 183896 470854 219340
rect 470234 183660 470266 183896
rect 470502 183660 470586 183896
rect 470822 183660 470854 183896
rect 470234 183576 470854 183660
rect 470234 183340 470266 183576
rect 470502 183340 470586 183576
rect 470822 183340 470854 183576
rect 470234 147896 470854 183340
rect 470234 147660 470266 147896
rect 470502 147660 470586 147896
rect 470822 147660 470854 147896
rect 470234 147576 470854 147660
rect 470234 147340 470266 147576
rect 470502 147340 470586 147576
rect 470822 147340 470854 147576
rect 470234 111896 470854 147340
rect 470234 111660 470266 111896
rect 470502 111660 470586 111896
rect 470822 111660 470854 111896
rect 470234 111576 470854 111660
rect 470234 111340 470266 111576
rect 470502 111340 470586 111576
rect 470822 111340 470854 111576
rect 470234 75896 470854 111340
rect 470234 75660 470266 75896
rect 470502 75660 470586 75896
rect 470822 75660 470854 75896
rect 470234 75576 470854 75660
rect 470234 75340 470266 75576
rect 470502 75340 470586 75576
rect 470822 75340 470854 75576
rect 470234 39896 470854 75340
rect 470234 39660 470266 39896
rect 470502 39660 470586 39896
rect 470822 39660 470854 39896
rect 470234 39576 470854 39660
rect 470234 39340 470266 39576
rect 470502 39340 470586 39576
rect 470822 39340 470854 39576
rect 470234 3896 470854 39340
rect 470234 3660 470266 3896
rect 470502 3660 470586 3896
rect 470822 3660 470854 3896
rect 470234 3576 470854 3660
rect 470234 3340 470266 3576
rect 470502 3340 470586 3576
rect 470822 3340 470854 3576
rect 470234 -1304 470854 3340
rect 470234 -1540 470266 -1304
rect 470502 -1540 470586 -1304
rect 470822 -1540 470854 -1304
rect 470234 -1624 470854 -1540
rect 470234 -1860 470266 -1624
rect 470502 -1860 470586 -1624
rect 470822 -1860 470854 -1624
rect 470234 -7652 470854 -1860
rect 471474 706760 472094 711592
rect 471474 706524 471506 706760
rect 471742 706524 471826 706760
rect 472062 706524 472094 706760
rect 471474 706440 472094 706524
rect 471474 706204 471506 706440
rect 471742 706204 471826 706440
rect 472062 706204 472094 706440
rect 471474 689136 472094 706204
rect 471474 688900 471506 689136
rect 471742 688900 471826 689136
rect 472062 688900 472094 689136
rect 471474 688816 472094 688900
rect 471474 688580 471506 688816
rect 471742 688580 471826 688816
rect 472062 688580 472094 688816
rect 471474 653136 472094 688580
rect 471474 652900 471506 653136
rect 471742 652900 471826 653136
rect 472062 652900 472094 653136
rect 471474 652816 472094 652900
rect 471474 652580 471506 652816
rect 471742 652580 471826 652816
rect 472062 652580 472094 652816
rect 471474 617136 472094 652580
rect 471474 616900 471506 617136
rect 471742 616900 471826 617136
rect 472062 616900 472094 617136
rect 471474 616816 472094 616900
rect 471474 616580 471506 616816
rect 471742 616580 471826 616816
rect 472062 616580 472094 616816
rect 471474 581136 472094 616580
rect 471474 580900 471506 581136
rect 471742 580900 471826 581136
rect 472062 580900 472094 581136
rect 471474 580816 472094 580900
rect 471474 580580 471506 580816
rect 471742 580580 471826 580816
rect 472062 580580 472094 580816
rect 471474 545136 472094 580580
rect 471474 544900 471506 545136
rect 471742 544900 471826 545136
rect 472062 544900 472094 545136
rect 471474 544816 472094 544900
rect 471474 544580 471506 544816
rect 471742 544580 471826 544816
rect 472062 544580 472094 544816
rect 471474 509136 472094 544580
rect 471474 508900 471506 509136
rect 471742 508900 471826 509136
rect 472062 508900 472094 509136
rect 471474 508816 472094 508900
rect 471474 508580 471506 508816
rect 471742 508580 471826 508816
rect 472062 508580 472094 508816
rect 471474 473136 472094 508580
rect 471474 472900 471506 473136
rect 471742 472900 471826 473136
rect 472062 472900 472094 473136
rect 471474 472816 472094 472900
rect 471474 472580 471506 472816
rect 471742 472580 471826 472816
rect 472062 472580 472094 472816
rect 471474 437136 472094 472580
rect 471474 436900 471506 437136
rect 471742 436900 471826 437136
rect 472062 436900 472094 437136
rect 471474 436816 472094 436900
rect 471474 436580 471506 436816
rect 471742 436580 471826 436816
rect 472062 436580 472094 436816
rect 471474 401136 472094 436580
rect 471474 400900 471506 401136
rect 471742 400900 471826 401136
rect 472062 400900 472094 401136
rect 471474 400816 472094 400900
rect 471474 400580 471506 400816
rect 471742 400580 471826 400816
rect 472062 400580 472094 400816
rect 471474 365136 472094 400580
rect 471474 364900 471506 365136
rect 471742 364900 471826 365136
rect 472062 364900 472094 365136
rect 471474 364816 472094 364900
rect 471474 364580 471506 364816
rect 471742 364580 471826 364816
rect 472062 364580 472094 364816
rect 471474 329136 472094 364580
rect 472714 707720 473334 711592
rect 472714 707484 472746 707720
rect 472982 707484 473066 707720
rect 473302 707484 473334 707720
rect 472714 707400 473334 707484
rect 472714 707164 472746 707400
rect 472982 707164 473066 707400
rect 473302 707164 473334 707400
rect 472714 690376 473334 707164
rect 472714 690140 472746 690376
rect 472982 690140 473066 690376
rect 473302 690140 473334 690376
rect 472714 690056 473334 690140
rect 472714 689820 472746 690056
rect 472982 689820 473066 690056
rect 473302 689820 473334 690056
rect 472714 654376 473334 689820
rect 472714 654140 472746 654376
rect 472982 654140 473066 654376
rect 473302 654140 473334 654376
rect 472714 654056 473334 654140
rect 472714 653820 472746 654056
rect 472982 653820 473066 654056
rect 473302 653820 473334 654056
rect 472714 618376 473334 653820
rect 472714 618140 472746 618376
rect 472982 618140 473066 618376
rect 473302 618140 473334 618376
rect 472714 618056 473334 618140
rect 472714 617820 472746 618056
rect 472982 617820 473066 618056
rect 473302 617820 473334 618056
rect 472714 582376 473334 617820
rect 472714 582140 472746 582376
rect 472982 582140 473066 582376
rect 473302 582140 473334 582376
rect 472714 582056 473334 582140
rect 472714 581820 472746 582056
rect 472982 581820 473066 582056
rect 473302 581820 473334 582056
rect 472714 546376 473334 581820
rect 472714 546140 472746 546376
rect 472982 546140 473066 546376
rect 473302 546140 473334 546376
rect 472714 546056 473334 546140
rect 472714 545820 472746 546056
rect 472982 545820 473066 546056
rect 473302 545820 473334 546056
rect 472714 510376 473334 545820
rect 472714 510140 472746 510376
rect 472982 510140 473066 510376
rect 473302 510140 473334 510376
rect 472714 510056 473334 510140
rect 472714 509820 472746 510056
rect 472982 509820 473066 510056
rect 473302 509820 473334 510056
rect 472714 474376 473334 509820
rect 472714 474140 472746 474376
rect 472982 474140 473066 474376
rect 473302 474140 473334 474376
rect 472714 474056 473334 474140
rect 472714 473820 472746 474056
rect 472982 473820 473066 474056
rect 473302 473820 473334 474056
rect 472714 438376 473334 473820
rect 473954 708680 474574 711592
rect 473954 708444 473986 708680
rect 474222 708444 474306 708680
rect 474542 708444 474574 708680
rect 473954 708360 474574 708444
rect 473954 708124 473986 708360
rect 474222 708124 474306 708360
rect 474542 708124 474574 708360
rect 473954 691616 474574 708124
rect 473954 691380 473986 691616
rect 474222 691380 474306 691616
rect 474542 691380 474574 691616
rect 473954 691296 474574 691380
rect 473954 691060 473986 691296
rect 474222 691060 474306 691296
rect 474542 691060 474574 691296
rect 473954 655616 474574 691060
rect 473954 655380 473986 655616
rect 474222 655380 474306 655616
rect 474542 655380 474574 655616
rect 473954 655296 474574 655380
rect 473954 655060 473986 655296
rect 474222 655060 474306 655296
rect 474542 655060 474574 655296
rect 473954 619616 474574 655060
rect 473954 619380 473986 619616
rect 474222 619380 474306 619616
rect 474542 619380 474574 619616
rect 473954 619296 474574 619380
rect 473954 619060 473986 619296
rect 474222 619060 474306 619296
rect 474542 619060 474574 619296
rect 473954 583616 474574 619060
rect 473954 583380 473986 583616
rect 474222 583380 474306 583616
rect 474542 583380 474574 583616
rect 473954 583296 474574 583380
rect 473954 583060 473986 583296
rect 474222 583060 474306 583296
rect 474542 583060 474574 583296
rect 473954 547616 474574 583060
rect 473954 547380 473986 547616
rect 474222 547380 474306 547616
rect 474542 547380 474574 547616
rect 473954 547296 474574 547380
rect 473954 547060 473986 547296
rect 474222 547060 474306 547296
rect 474542 547060 474574 547296
rect 473954 511616 474574 547060
rect 473954 511380 473986 511616
rect 474222 511380 474306 511616
rect 474542 511380 474574 511616
rect 473954 511296 474574 511380
rect 473954 511060 473986 511296
rect 474222 511060 474306 511296
rect 474542 511060 474574 511296
rect 473954 475616 474574 511060
rect 473954 475380 473986 475616
rect 474222 475380 474306 475616
rect 474542 475380 474574 475616
rect 473954 475296 474574 475380
rect 473954 475060 473986 475296
rect 474222 475060 474306 475296
rect 474542 475060 474574 475296
rect 473675 449718 473741 449719
rect 473675 449654 473676 449718
rect 473740 449654 473741 449718
rect 473675 449653 473741 449654
rect 472714 438140 472746 438376
rect 472982 438140 473066 438376
rect 473302 438140 473334 438376
rect 472714 438056 473334 438140
rect 472714 437820 472746 438056
rect 472982 437820 473066 438056
rect 473302 437820 473334 438056
rect 472714 402376 473334 437820
rect 473678 431903 473738 449653
rect 473954 439616 474574 475060
rect 473954 439380 473986 439616
rect 474222 439380 474306 439616
rect 474542 439380 474574 439616
rect 473954 439296 474574 439380
rect 473954 439060 473986 439296
rect 474222 439060 474306 439296
rect 474542 439060 474574 439296
rect 473675 431902 473741 431903
rect 473675 431838 473676 431902
rect 473740 431838 473741 431902
rect 473675 431837 473741 431838
rect 473678 410959 473738 431837
rect 473675 410958 473741 410959
rect 473675 410894 473676 410958
rect 473740 410894 473741 410958
rect 473675 410893 473741 410894
rect 472714 402140 472746 402376
rect 472982 402140 473066 402376
rect 473302 402140 473334 402376
rect 472714 402056 473334 402140
rect 472714 401820 472746 402056
rect 472982 401820 473066 402056
rect 473302 401820 473334 402056
rect 472714 366376 473334 401820
rect 473678 392055 473738 410893
rect 473954 403616 474574 439060
rect 473954 403380 473986 403616
rect 474222 403380 474306 403616
rect 474542 403380 474574 403616
rect 473954 403296 474574 403380
rect 473954 403060 473986 403296
rect 474222 403060 474306 403296
rect 474542 403060 474574 403296
rect 473675 392054 473741 392055
rect 473675 391990 473676 392054
rect 473740 391990 473741 392054
rect 473675 391989 473741 391990
rect 472714 366140 472746 366376
rect 472982 366140 473066 366376
rect 473302 366140 473334 366376
rect 472714 366056 473334 366140
rect 472714 365820 472746 366056
rect 472982 365820 473066 366056
rect 473302 365820 473334 366056
rect 472714 359062 473334 365820
rect 473954 367616 474574 403060
rect 475194 709640 475814 711592
rect 475194 709404 475226 709640
rect 475462 709404 475546 709640
rect 475782 709404 475814 709640
rect 475194 709320 475814 709404
rect 475194 709084 475226 709320
rect 475462 709084 475546 709320
rect 475782 709084 475814 709320
rect 475194 692856 475814 709084
rect 475194 692620 475226 692856
rect 475462 692620 475546 692856
rect 475782 692620 475814 692856
rect 475194 692536 475814 692620
rect 475194 692300 475226 692536
rect 475462 692300 475546 692536
rect 475782 692300 475814 692536
rect 475194 656856 475814 692300
rect 475194 656620 475226 656856
rect 475462 656620 475546 656856
rect 475782 656620 475814 656856
rect 475194 656536 475814 656620
rect 475194 656300 475226 656536
rect 475462 656300 475546 656536
rect 475782 656300 475814 656536
rect 475194 620856 475814 656300
rect 475194 620620 475226 620856
rect 475462 620620 475546 620856
rect 475782 620620 475814 620856
rect 475194 620536 475814 620620
rect 475194 620300 475226 620536
rect 475462 620300 475546 620536
rect 475782 620300 475814 620536
rect 475194 584856 475814 620300
rect 475194 584620 475226 584856
rect 475462 584620 475546 584856
rect 475782 584620 475814 584856
rect 475194 584536 475814 584620
rect 475194 584300 475226 584536
rect 475462 584300 475546 584536
rect 475782 584300 475814 584536
rect 475194 548856 475814 584300
rect 475194 548620 475226 548856
rect 475462 548620 475546 548856
rect 475782 548620 475814 548856
rect 475194 548536 475814 548620
rect 475194 548300 475226 548536
rect 475462 548300 475546 548536
rect 475782 548300 475814 548536
rect 475194 512856 475814 548300
rect 475194 512620 475226 512856
rect 475462 512620 475546 512856
rect 475782 512620 475814 512856
rect 475194 512536 475814 512620
rect 475194 512300 475226 512536
rect 475462 512300 475546 512536
rect 475782 512300 475814 512536
rect 475194 476856 475814 512300
rect 475194 476620 475226 476856
rect 475462 476620 475546 476856
rect 475782 476620 475814 476856
rect 475194 476536 475814 476620
rect 475194 476300 475226 476536
rect 475462 476300 475546 476536
rect 475782 476300 475814 476536
rect 475194 440856 475814 476300
rect 475194 440620 475226 440856
rect 475462 440620 475546 440856
rect 475782 440620 475814 440856
rect 475194 440536 475814 440620
rect 475194 440300 475226 440536
rect 475462 440300 475546 440536
rect 475782 440300 475814 440536
rect 475194 404856 475814 440300
rect 475194 404620 475226 404856
rect 475462 404620 475546 404856
rect 475782 404620 475814 404856
rect 475194 404536 475814 404620
rect 475194 404300 475226 404536
rect 475462 404300 475546 404536
rect 475782 404300 475814 404536
rect 474963 392054 475029 392055
rect 474963 391990 474964 392054
rect 475028 391990 475029 392054
rect 474963 391989 475029 391990
rect 474966 389335 475026 391989
rect 474963 389334 475029 389335
rect 474963 389270 474964 389334
rect 475028 389270 475029 389334
rect 474963 389269 475029 389270
rect 473954 367380 473986 367616
rect 474222 367380 474306 367616
rect 474542 367380 474574 367616
rect 473954 367296 474574 367380
rect 473954 367060 473986 367296
rect 474222 367060 474306 367296
rect 474542 367060 474574 367296
rect 473954 359062 474574 367060
rect 474966 357511 475026 389269
rect 475194 368856 475814 404300
rect 475194 368620 475226 368856
rect 475462 368620 475546 368856
rect 475782 368620 475814 368856
rect 475194 368536 475814 368620
rect 475194 368300 475226 368536
rect 475462 368300 475546 368536
rect 475782 368300 475814 368536
rect 475194 359062 475814 368300
rect 476434 710600 477054 711592
rect 476434 710364 476466 710600
rect 476702 710364 476786 710600
rect 477022 710364 477054 710600
rect 476434 710280 477054 710364
rect 476434 710044 476466 710280
rect 476702 710044 476786 710280
rect 477022 710044 477054 710280
rect 476434 694096 477054 710044
rect 476434 693860 476466 694096
rect 476702 693860 476786 694096
rect 477022 693860 477054 694096
rect 476434 693776 477054 693860
rect 476434 693540 476466 693776
rect 476702 693540 476786 693776
rect 477022 693540 477054 693776
rect 476434 658096 477054 693540
rect 476434 657860 476466 658096
rect 476702 657860 476786 658096
rect 477022 657860 477054 658096
rect 476434 657776 477054 657860
rect 476434 657540 476466 657776
rect 476702 657540 476786 657776
rect 477022 657540 477054 657776
rect 476434 622096 477054 657540
rect 476434 621860 476466 622096
rect 476702 621860 476786 622096
rect 477022 621860 477054 622096
rect 476434 621776 477054 621860
rect 476434 621540 476466 621776
rect 476702 621540 476786 621776
rect 477022 621540 477054 621776
rect 476434 586096 477054 621540
rect 476434 585860 476466 586096
rect 476702 585860 476786 586096
rect 477022 585860 477054 586096
rect 476434 585776 477054 585860
rect 476434 585540 476466 585776
rect 476702 585540 476786 585776
rect 477022 585540 477054 585776
rect 476434 550096 477054 585540
rect 476434 549860 476466 550096
rect 476702 549860 476786 550096
rect 477022 549860 477054 550096
rect 476434 549776 477054 549860
rect 476434 549540 476466 549776
rect 476702 549540 476786 549776
rect 477022 549540 477054 549776
rect 476434 514096 477054 549540
rect 476434 513860 476466 514096
rect 476702 513860 476786 514096
rect 477022 513860 477054 514096
rect 476434 513776 477054 513860
rect 476434 513540 476466 513776
rect 476702 513540 476786 513776
rect 477022 513540 477054 513776
rect 476434 478096 477054 513540
rect 476434 477860 476466 478096
rect 476702 477860 476786 478096
rect 477022 477860 477054 478096
rect 476434 477776 477054 477860
rect 476434 477540 476466 477776
rect 476702 477540 476786 477776
rect 477022 477540 477054 477776
rect 476434 442096 477054 477540
rect 476434 441860 476466 442096
rect 476702 441860 476786 442096
rect 477022 441860 477054 442096
rect 476434 441776 477054 441860
rect 476434 441540 476466 441776
rect 476702 441540 476786 441776
rect 477022 441540 477054 441776
rect 476434 406096 477054 441540
rect 476434 405860 476466 406096
rect 476702 405860 476786 406096
rect 477022 405860 477054 406096
rect 476434 405776 477054 405860
rect 476434 405540 476466 405776
rect 476702 405540 476786 405776
rect 477022 405540 477054 405776
rect 476434 370096 477054 405540
rect 476434 369860 476466 370096
rect 476702 369860 476786 370096
rect 477022 369860 477054 370096
rect 476434 369776 477054 369860
rect 476434 369540 476466 369776
rect 476702 369540 476786 369776
rect 477022 369540 477054 369776
rect 476434 359062 477054 369540
rect 477674 711560 478294 711592
rect 477674 711324 477706 711560
rect 477942 711324 478026 711560
rect 478262 711324 478294 711560
rect 477674 711240 478294 711324
rect 477674 711004 477706 711240
rect 477942 711004 478026 711240
rect 478262 711004 478294 711240
rect 477674 695336 478294 711004
rect 477674 695100 477706 695336
rect 477942 695100 478026 695336
rect 478262 695100 478294 695336
rect 477674 695016 478294 695100
rect 477674 694780 477706 695016
rect 477942 694780 478026 695016
rect 478262 694780 478294 695016
rect 477674 659336 478294 694780
rect 477674 659100 477706 659336
rect 477942 659100 478026 659336
rect 478262 659100 478294 659336
rect 477674 659016 478294 659100
rect 477674 658780 477706 659016
rect 477942 658780 478026 659016
rect 478262 658780 478294 659016
rect 477674 623336 478294 658780
rect 477674 623100 477706 623336
rect 477942 623100 478026 623336
rect 478262 623100 478294 623336
rect 477674 623016 478294 623100
rect 477674 622780 477706 623016
rect 477942 622780 478026 623016
rect 478262 622780 478294 623016
rect 477674 587336 478294 622780
rect 477674 587100 477706 587336
rect 477942 587100 478026 587336
rect 478262 587100 478294 587336
rect 477674 587016 478294 587100
rect 477674 586780 477706 587016
rect 477942 586780 478026 587016
rect 478262 586780 478294 587016
rect 477674 551336 478294 586780
rect 477674 551100 477706 551336
rect 477942 551100 478026 551336
rect 478262 551100 478294 551336
rect 477674 551016 478294 551100
rect 477674 550780 477706 551016
rect 477942 550780 478026 551016
rect 478262 550780 478294 551016
rect 477674 515336 478294 550780
rect 477674 515100 477706 515336
rect 477942 515100 478026 515336
rect 478262 515100 478294 515336
rect 477674 515016 478294 515100
rect 477674 514780 477706 515016
rect 477942 514780 478026 515016
rect 478262 514780 478294 515016
rect 477674 479336 478294 514780
rect 477674 479100 477706 479336
rect 477942 479100 478026 479336
rect 478262 479100 478294 479336
rect 477674 479016 478294 479100
rect 477674 478780 477706 479016
rect 477942 478780 478026 479016
rect 478262 478780 478294 479016
rect 477674 443336 478294 478780
rect 504994 704840 505614 711592
rect 504994 704604 505026 704840
rect 505262 704604 505346 704840
rect 505582 704604 505614 704840
rect 504994 704520 505614 704604
rect 504994 704284 505026 704520
rect 505262 704284 505346 704520
rect 505582 704284 505614 704520
rect 504994 701756 505614 704284
rect 504994 701692 505032 701756
rect 505096 701692 505112 701756
rect 505176 701692 505192 701756
rect 505256 701692 505272 701756
rect 505336 701692 505352 701756
rect 505416 701692 505432 701756
rect 505496 701692 505512 701756
rect 505576 701692 505614 701756
rect 504994 701676 505614 701692
rect 504994 701612 505032 701676
rect 505096 701612 505112 701676
rect 505176 701612 505192 701676
rect 505256 701612 505272 701676
rect 505336 701612 505352 701676
rect 505416 701612 505432 701676
rect 505496 701612 505512 701676
rect 505576 701612 505614 701676
rect 504994 701596 505614 701612
rect 504994 701532 505032 701596
rect 505096 701532 505112 701596
rect 505176 701532 505192 701596
rect 505256 701532 505272 701596
rect 505336 701532 505352 701596
rect 505416 701532 505432 701596
rect 505496 701532 505512 701596
rect 505576 701532 505614 701596
rect 504994 701516 505614 701532
rect 504994 701452 505032 701516
rect 505096 701452 505112 701516
rect 505176 701452 505192 701516
rect 505256 701452 505272 701516
rect 505336 701452 505352 701516
rect 505416 701452 505432 701516
rect 505496 701452 505512 701516
rect 505576 701452 505614 701516
rect 504994 686656 505614 701452
rect 504994 686420 505026 686656
rect 505262 686420 505346 686656
rect 505582 686420 505614 686656
rect 504994 686336 505614 686420
rect 504994 686100 505026 686336
rect 505262 686100 505346 686336
rect 505582 686100 505614 686336
rect 504994 650656 505614 686100
rect 504994 650420 505026 650656
rect 505262 650420 505346 650656
rect 505582 650420 505614 650656
rect 504994 650336 505614 650420
rect 504994 650100 505026 650336
rect 505262 650100 505346 650336
rect 505582 650100 505614 650336
rect 504994 614656 505614 650100
rect 504994 614420 505026 614656
rect 505262 614420 505346 614656
rect 505582 614420 505614 614656
rect 504994 614336 505614 614420
rect 504994 614100 505026 614336
rect 505262 614100 505346 614336
rect 505582 614100 505614 614336
rect 504994 578656 505614 614100
rect 504994 578420 505026 578656
rect 505262 578420 505346 578656
rect 505582 578420 505614 578656
rect 504994 578336 505614 578420
rect 504994 578100 505026 578336
rect 505262 578100 505346 578336
rect 505582 578100 505614 578336
rect 504994 554602 505614 578100
rect 504994 554538 505032 554602
rect 505096 554538 505112 554602
rect 505176 554538 505192 554602
rect 505256 554538 505272 554602
rect 505336 554538 505352 554602
rect 505416 554538 505432 554602
rect 505496 554538 505512 554602
rect 505576 554538 505614 554602
rect 504994 554522 505614 554538
rect 504994 554458 505032 554522
rect 505096 554458 505112 554522
rect 505176 554458 505192 554522
rect 505256 554458 505272 554522
rect 505336 554458 505352 554522
rect 505416 554458 505432 554522
rect 505496 554458 505512 554522
rect 505576 554458 505614 554522
rect 504994 554442 505614 554458
rect 504994 554378 505032 554442
rect 505096 554378 505112 554442
rect 505176 554378 505192 554442
rect 505256 554378 505272 554442
rect 505336 554378 505352 554442
rect 505416 554378 505432 554442
rect 505496 554378 505512 554442
rect 505576 554378 505614 554442
rect 504994 554362 505614 554378
rect 504994 554298 505032 554362
rect 505096 554298 505112 554362
rect 505176 554298 505192 554362
rect 505256 554298 505272 554362
rect 505336 554298 505352 554362
rect 505416 554298 505432 554362
rect 505496 554298 505512 554362
rect 505576 554298 505614 554362
rect 504994 542656 505614 554298
rect 504994 542420 505026 542656
rect 505262 542420 505346 542656
rect 505582 542420 505614 542656
rect 504994 542336 505614 542420
rect 504994 542100 505026 542336
rect 505262 542100 505346 542336
rect 505582 542100 505614 542336
rect 504994 506656 505614 542100
rect 504994 506420 505026 506656
rect 505262 506420 505346 506656
rect 505582 506420 505614 506656
rect 504994 506336 505614 506420
rect 504994 506100 505026 506336
rect 505262 506100 505346 506336
rect 505582 506100 505614 506336
rect 504994 470656 505614 506100
rect 504994 470420 505026 470656
rect 505262 470420 505346 470656
rect 505582 470420 505614 470656
rect 504994 470336 505614 470420
rect 504994 470100 505026 470336
rect 505262 470100 505346 470336
rect 505582 470100 505614 470336
rect 478459 450262 478525 450263
rect 478459 450198 478460 450262
rect 478524 450198 478525 450262
rect 478459 450197 478525 450198
rect 481219 450262 481285 450263
rect 481219 450198 481220 450262
rect 481284 450198 481285 450262
rect 481219 450197 481285 450198
rect 487843 450262 487909 450263
rect 487843 450198 487844 450262
rect 487908 450198 487909 450262
rect 487843 450197 487909 450198
rect 477674 443100 477706 443336
rect 477942 443100 478026 443336
rect 478262 443100 478294 443336
rect 477674 443016 478294 443100
rect 477674 442780 477706 443016
rect 477942 442780 478026 443016
rect 478262 442780 478294 443016
rect 477674 407336 478294 442780
rect 478462 431631 478522 450197
rect 481222 432175 481282 450197
rect 487846 441632 487906 450197
rect 487846 441572 488458 441632
rect 483611 432854 483677 432855
rect 483611 432790 483612 432854
rect 483676 432790 483677 432854
rect 483611 432789 483677 432790
rect 483614 432311 483674 432789
rect 483611 432310 483677 432311
rect 483611 432246 483612 432310
rect 483676 432246 483677 432310
rect 483611 432245 483677 432246
rect 481219 432174 481285 432175
rect 481219 432110 481220 432174
rect 481284 432110 481285 432174
rect 481219 432109 481285 432110
rect 481222 431972 481282 432109
rect 481038 431912 481282 431972
rect 483614 431972 483674 432245
rect 483614 431912 484226 431972
rect 478459 431630 478525 431631
rect 478459 431566 478460 431630
rect 478524 431566 478525 431630
rect 478459 431565 478525 431566
rect 478462 410143 478522 431565
rect 480115 427958 480181 427959
rect 480115 427894 480116 427958
rect 480180 427894 480181 427958
rect 480115 427893 480181 427894
rect 478459 410142 478525 410143
rect 478459 410078 478460 410142
rect 478524 410078 478525 410142
rect 478459 410077 478525 410078
rect 477674 407100 477706 407336
rect 477942 407100 478026 407336
rect 478262 407100 478294 407336
rect 477674 407016 478294 407100
rect 477674 406780 477706 407016
rect 477942 406780 478026 407016
rect 478262 406780 478294 407016
rect 477674 371336 478294 406780
rect 478462 402992 478522 410077
rect 480118 407559 480178 427893
rect 481038 422312 481098 431912
rect 481038 422252 481466 422312
rect 481406 410143 481466 422252
rect 484166 410415 484226 431912
rect 488398 431631 488458 441572
rect 504994 434656 505614 470100
rect 504994 434420 505026 434656
rect 505262 434420 505346 434656
rect 505582 434420 505614 434656
rect 504994 434336 505614 434420
rect 504994 434100 505026 434336
rect 505262 434100 505346 434336
rect 505582 434100 505614 434336
rect 488395 431630 488461 431631
rect 488395 431566 488396 431630
rect 488460 431566 488461 431630
rect 488395 431565 488461 431566
rect 486555 427958 486621 427959
rect 486555 427894 486556 427958
rect 486620 427894 486621 427958
rect 486555 427893 486621 427894
rect 484163 410414 484229 410415
rect 484163 410350 484164 410414
rect 484228 410350 484229 410414
rect 484163 410349 484229 410350
rect 481403 410142 481469 410143
rect 481403 410078 481404 410142
rect 481468 410078 481469 410142
rect 481403 410077 481469 410078
rect 480115 407558 480181 407559
rect 480115 407494 480116 407558
rect 480180 407494 480181 407558
rect 480115 407493 480181 407494
rect 478462 402932 478706 402992
rect 478646 389335 478706 402932
rect 481406 393332 481466 410077
rect 482875 407150 482941 407151
rect 482875 407086 482876 407150
rect 482940 407086 482941 407150
rect 482875 407085 482941 407086
rect 481406 393272 481834 393332
rect 481774 389471 481834 393272
rect 481771 389470 481837 389471
rect 481771 389406 481772 389470
rect 481836 389406 481837 389470
rect 481771 389405 481837 389406
rect 478643 389334 478709 389335
rect 478643 389270 478644 389334
rect 478708 389270 478709 389334
rect 478643 389269 478709 389270
rect 477674 371100 477706 371336
rect 477942 371100 478026 371336
rect 478262 371100 478294 371336
rect 477674 371016 478294 371100
rect 477674 370780 477706 371016
rect 477942 370780 478026 371016
rect 478262 370780 478294 371016
rect 477674 359062 478294 370780
rect 478646 358055 478706 389269
rect 481774 358055 481834 389405
rect 482878 370159 482938 407085
rect 484166 393332 484226 410349
rect 485635 407150 485701 407151
rect 485635 407086 485636 407150
rect 485700 407086 485701 407150
rect 485635 407085 485701 407086
rect 484166 393272 484962 393332
rect 484902 390300 484962 393272
rect 484899 390299 484965 390300
rect 484899 390235 484900 390299
rect 484964 390235 484965 390299
rect 484899 390234 484965 390235
rect 482875 370158 482941 370159
rect 482875 370094 482876 370158
rect 482940 370094 482941 370158
rect 482875 370093 482941 370094
rect 484902 358055 484962 390234
rect 478643 358054 478709 358055
rect 478643 357990 478644 358054
rect 478708 357990 478709 358054
rect 478643 357989 478709 357990
rect 481771 358054 481837 358055
rect 481771 357990 481772 358054
rect 481836 357990 481837 358054
rect 481771 357989 481837 357990
rect 484899 358054 484965 358055
rect 484899 357990 484900 358054
rect 484964 357990 484965 358054
rect 484899 357989 484965 357990
rect 474963 357510 475029 357511
rect 474963 357446 474964 357510
rect 475028 357446 475029 357510
rect 474963 357445 475029 357446
rect 474966 357372 475026 357445
rect 474966 357312 475394 357372
rect 475334 356692 475394 357312
rect 474966 356632 475394 356692
rect 471474 328900 471506 329136
rect 471742 328900 471826 329136
rect 472062 328900 472094 329136
rect 471474 328816 472094 328900
rect 471474 328580 471506 328816
rect 471742 328580 471826 328816
rect 472062 328580 472094 328816
rect 471474 293136 472094 328580
rect 471474 292900 471506 293136
rect 471742 292900 471826 293136
rect 472062 292900 472094 293136
rect 471474 292816 472094 292900
rect 471474 292580 471506 292816
rect 471742 292580 471826 292816
rect 472062 292580 472094 292816
rect 471474 257136 472094 292580
rect 472714 330376 473334 354617
rect 473675 343774 473741 343775
rect 473675 343710 473676 343774
rect 473740 343710 473741 343774
rect 473675 343709 473741 343710
rect 473678 340511 473738 343709
rect 473675 340510 473741 340511
rect 473675 340446 473676 340510
rect 473740 340446 473741 340510
rect 473675 340445 473741 340446
rect 472714 330140 472746 330376
rect 472982 330140 473066 330376
rect 473302 330140 473334 330376
rect 472714 330056 473334 330140
rect 472714 329820 472746 330056
rect 472982 329820 473066 330056
rect 473302 329820 473334 330056
rect 472714 294376 473334 329820
rect 473678 321335 473738 340445
rect 473954 331616 474574 354617
rect 474966 343775 475026 356632
rect 474963 343774 475029 343775
rect 474963 343710 474964 343774
rect 475028 343710 475029 343774
rect 474963 343709 475029 343710
rect 473954 331380 473986 331616
rect 474222 331380 474306 331616
rect 474542 331380 474574 331616
rect 473954 331296 474574 331380
rect 473954 331060 473986 331296
rect 474222 331060 474306 331296
rect 474542 331060 474574 331296
rect 473675 321334 473741 321335
rect 473675 321270 473676 321334
rect 473740 321270 473741 321334
rect 473675 321269 473741 321270
rect 473678 305967 473738 321269
rect 473675 305966 473741 305967
rect 473675 305902 473676 305966
rect 473740 305902 473741 305966
rect 473675 305901 473741 305902
rect 472714 294140 472746 294376
rect 472982 294140 473066 294376
rect 473302 294140 473334 294376
rect 472714 294056 473334 294140
rect 472714 293820 472746 294056
rect 472982 293820 473066 294056
rect 473302 293820 473334 294056
rect 472714 268062 473334 293820
rect 473678 289783 473738 305901
rect 473954 295616 474574 331060
rect 473954 295380 473986 295616
rect 474222 295380 474306 295616
rect 474542 295380 474574 295616
rect 473954 295296 474574 295380
rect 473954 295060 473986 295296
rect 474222 295060 474306 295296
rect 474542 295060 474574 295296
rect 473675 289782 473741 289783
rect 473675 289718 473676 289782
rect 473740 289718 473741 289782
rect 473675 289717 473741 289718
rect 473954 268062 474574 295060
rect 475194 332856 475814 354617
rect 475194 332620 475226 332856
rect 475462 332620 475546 332856
rect 475782 332620 475814 332856
rect 475194 332536 475814 332620
rect 475194 332300 475226 332536
rect 475462 332300 475546 332536
rect 475782 332300 475814 332536
rect 475194 296856 475814 332300
rect 475194 296620 475226 296856
rect 475462 296620 475546 296856
rect 475782 296620 475814 296856
rect 475194 296536 475814 296620
rect 475194 296300 475226 296536
rect 475462 296300 475546 296536
rect 475782 296300 475814 296536
rect 475194 268062 475814 296300
rect 476434 334096 477054 354617
rect 476434 333860 476466 334096
rect 476702 333860 476786 334096
rect 477022 333860 477054 334096
rect 476434 333776 477054 333860
rect 476434 333540 476466 333776
rect 476702 333540 476786 333776
rect 477022 333540 477054 333776
rect 476434 298096 477054 333540
rect 476434 297860 476466 298096
rect 476702 297860 476786 298096
rect 477022 297860 477054 298096
rect 476434 297776 477054 297860
rect 476434 297540 476466 297776
rect 476702 297540 476786 297776
rect 477022 297540 477054 297776
rect 476067 289782 476133 289783
rect 476067 289718 476068 289782
rect 476132 289718 476133 289782
rect 476067 289717 476133 289718
rect 476070 286655 476130 289717
rect 476067 286654 476133 286655
rect 476067 286590 476068 286654
rect 476132 286590 476133 286654
rect 476067 286589 476133 286590
rect 476070 267752 476130 286589
rect 476434 268062 477054 297540
rect 477674 335336 478294 354617
rect 478646 345032 478706 357989
rect 481774 354692 481834 357989
rect 481590 354632 481834 354692
rect 484902 354692 484962 357989
rect 484902 354632 485514 354692
rect 481590 345032 481650 354632
rect 485454 351935 485514 354632
rect 485451 351934 485517 351935
rect 485451 351870 485452 351934
rect 485516 351870 485517 351934
rect 485451 351869 485517 351870
rect 478462 344972 478706 345032
rect 481406 344972 481650 345032
rect 478462 341055 478522 344972
rect 481406 341055 481466 344972
rect 478459 341054 478525 341055
rect 478459 340990 478460 341054
rect 478524 340990 478525 341054
rect 478459 340989 478525 340990
rect 481403 341054 481469 341055
rect 481403 340990 481404 341054
rect 481468 340990 481469 341054
rect 481403 340989 481469 340990
rect 477674 335100 477706 335336
rect 477942 335100 478026 335336
rect 478262 335100 478294 335336
rect 477674 335016 478294 335100
rect 477674 334780 477706 335016
rect 477942 334780 478026 335016
rect 478262 334780 478294 335016
rect 477674 299336 478294 334780
rect 478462 325712 478522 340989
rect 481406 325712 481466 340989
rect 485638 334119 485698 407085
rect 486558 335479 486618 427893
rect 488398 413951 488458 431565
rect 488395 413950 488461 413951
rect 488395 413886 488396 413950
rect 488460 413886 488461 413950
rect 488395 413885 488461 413886
rect 504994 398656 505614 434100
rect 504994 398420 505026 398656
rect 505262 398420 505346 398656
rect 505582 398420 505614 398656
rect 504994 398336 505614 398420
rect 504994 398100 505026 398336
rect 505262 398100 505346 398336
rect 505582 398100 505614 398336
rect 489315 392054 489381 392055
rect 489315 391990 489316 392054
rect 489380 391990 489381 392054
rect 489315 391989 489381 391990
rect 489318 389471 489378 391989
rect 489315 389470 489381 389471
rect 489315 389406 489316 389470
rect 489380 389406 489381 389470
rect 489315 389405 489381 389406
rect 486739 386478 486805 386479
rect 486739 386414 486740 386478
rect 486804 386414 486805 386478
rect 486739 386413 486805 386414
rect 486555 335478 486621 335479
rect 486555 335414 486556 335478
rect 486620 335414 486621 335478
rect 486555 335413 486621 335414
rect 485635 334118 485701 334119
rect 485635 334054 485636 334118
rect 485700 334054 485701 334118
rect 485635 334053 485701 334054
rect 486742 332759 486802 386413
rect 489318 358055 489378 389405
rect 504994 362656 505614 398100
rect 504994 362420 505026 362656
rect 505262 362420 505346 362656
rect 505582 362420 505614 362656
rect 504994 362336 505614 362420
rect 504994 362100 505026 362336
rect 505262 362100 505346 362336
rect 505582 362100 505614 362336
rect 488395 358054 488461 358055
rect 488395 357990 488396 358054
rect 488460 357990 488461 358054
rect 488395 357989 488461 357990
rect 489315 358054 489381 358055
rect 489315 357990 489316 358054
rect 489380 357990 489381 358054
rect 489315 357989 489381 357990
rect 488398 345032 488458 357989
rect 488030 344972 488458 345032
rect 488030 341055 488090 344972
rect 488027 341054 488093 341055
rect 488027 340990 488028 341054
rect 488092 340990 488093 341054
rect 488027 340989 488093 340990
rect 486739 332758 486805 332759
rect 486739 332694 486740 332758
rect 486804 332694 486805 332758
rect 486739 332693 486805 332694
rect 478462 325652 478706 325712
rect 478646 320927 478706 325652
rect 481038 325652 481466 325712
rect 481038 321063 481098 325652
rect 483611 322150 483677 322151
rect 483611 322086 483612 322150
rect 483676 322086 483677 322150
rect 483611 322085 483677 322086
rect 483614 321607 483674 322085
rect 483611 321606 483677 321607
rect 483611 321542 483612 321606
rect 483676 321542 483677 321606
rect 483611 321541 483677 321542
rect 481035 321062 481101 321063
rect 481035 320998 481036 321062
rect 481100 320998 481101 321062
rect 481035 320997 481101 320998
rect 478643 320926 478709 320927
rect 478643 320862 478644 320926
rect 478708 320862 478709 320926
rect 478643 320861 478709 320862
rect 478646 306392 478706 320861
rect 481038 316052 481098 320997
rect 480854 315992 481098 316052
rect 483614 316052 483674 321541
rect 488030 321063 488090 340989
rect 504994 326656 505614 362100
rect 504994 326420 505026 326656
rect 505262 326420 505346 326656
rect 505582 326420 505614 326656
rect 504994 326336 505614 326420
rect 504994 326100 505026 326336
rect 505262 326100 505346 326336
rect 505582 326100 505614 326336
rect 488027 321062 488093 321063
rect 488027 320998 488028 321062
rect 488092 320998 488093 321062
rect 488027 320997 488093 320998
rect 488030 316052 488090 320997
rect 483614 315992 484226 316052
rect 480854 306511 480914 315992
rect 480851 306510 480917 306511
rect 480851 306446 480852 306510
rect 480916 306446 480917 306510
rect 480851 306445 480917 306446
rect 478646 306332 478890 306392
rect 478830 305695 478890 306332
rect 478827 305694 478893 305695
rect 478827 305630 478828 305694
rect 478892 305630 478893 305694
rect 478827 305629 478893 305630
rect 477674 299100 477706 299336
rect 477942 299100 478026 299336
rect 478262 299100 478294 299336
rect 477674 299016 478294 299100
rect 477674 298780 477706 299016
rect 477942 298780 478026 299016
rect 478262 298780 478294 299016
rect 477674 268062 478294 298780
rect 478830 287072 478890 305629
rect 480854 302295 480914 306445
rect 484166 305559 484226 315992
rect 487662 315992 488090 316052
rect 487662 306392 487722 315992
rect 487662 306375 488458 306392
rect 487659 306374 488458 306375
rect 487659 306310 487660 306374
rect 487724 306332 488458 306374
rect 487724 306310 487725 306332
rect 487659 306309 487725 306310
rect 484163 305558 484229 305559
rect 484163 305494 484164 305558
rect 484228 305494 484229 305558
rect 484163 305493 484229 305494
rect 480851 302294 480917 302295
rect 480851 302230 480852 302294
rect 480916 302230 480917 302294
rect 480851 302229 480917 302230
rect 482139 288422 482205 288423
rect 482139 288358 482140 288422
rect 482204 288358 482205 288422
rect 482139 288357 482205 288358
rect 478830 287012 479074 287072
rect 478830 286927 478890 287012
rect 478827 286926 478893 286927
rect 478827 286862 478828 286926
rect 478892 286862 478893 286926
rect 478827 286861 478893 286862
rect 476070 267692 476498 267752
rect 476438 265031 476498 267692
rect 479014 265983 479074 287012
rect 482142 285703 482202 288357
rect 484166 286655 484226 305493
rect 488398 286791 488458 306332
rect 504994 290656 505614 326100
rect 504994 290420 505026 290656
rect 505262 290420 505346 290656
rect 505582 290420 505614 290656
rect 504994 290336 505614 290420
rect 504994 290100 505026 290336
rect 505262 290100 505346 290336
rect 505582 290100 505614 290336
rect 488395 286790 488461 286791
rect 488395 286726 488396 286790
rect 488460 286726 488461 286790
rect 488395 286725 488461 286726
rect 484163 286654 484229 286655
rect 484163 286590 484164 286654
rect 484228 286590 484229 286654
rect 484163 286589 484229 286590
rect 482139 285702 482205 285703
rect 482139 285638 482140 285702
rect 482204 285638 482205 285702
rect 482139 285637 482205 285638
rect 482142 273327 482202 285637
rect 482139 273326 482205 273327
rect 482139 273262 482140 273326
rect 482204 273262 482205 273326
rect 482139 273261 482205 273262
rect 484166 272647 484226 286589
rect 484163 272646 484229 272647
rect 484163 272582 484164 272646
rect 484228 272582 484229 272646
rect 484163 272581 484229 272582
rect 488398 267071 488458 286725
rect 488395 267070 488461 267071
rect 488395 267006 488396 267070
rect 488460 267006 488461 267070
rect 488395 267005 488461 267006
rect 479011 265982 479077 265983
rect 479011 265918 479012 265982
rect 479076 265918 479077 265982
rect 479011 265917 479077 265918
rect 476435 265030 476501 265031
rect 476435 264966 476436 265030
rect 476500 264966 476501 265030
rect 476435 264965 476501 264966
rect 477355 265030 477421 265031
rect 477355 264966 477356 265030
rect 477420 264966 477421 265030
rect 477355 264965 477421 264966
rect 480115 265030 480181 265031
rect 480115 264966 480116 265030
rect 480180 264966 480181 265030
rect 480115 264965 480181 264966
rect 471474 256900 471506 257136
rect 471742 256900 471826 257136
rect 472062 256900 472094 257136
rect 471474 256816 472094 256900
rect 471474 256580 471506 256816
rect 471742 256580 471826 256816
rect 472062 256580 472094 256816
rect 471474 221136 472094 256580
rect 471474 220900 471506 221136
rect 471742 220900 471826 221136
rect 472062 220900 472094 221136
rect 471474 220816 472094 220900
rect 471474 220580 471506 220816
rect 471742 220580 471826 220816
rect 472062 220580 472094 220816
rect 471474 185136 472094 220580
rect 471474 184900 471506 185136
rect 471742 184900 471826 185136
rect 472062 184900 472094 185136
rect 471474 184816 472094 184900
rect 471474 184580 471506 184816
rect 471742 184580 471826 184816
rect 472062 184580 472094 184816
rect 471474 149136 472094 184580
rect 471474 148900 471506 149136
rect 471742 148900 471826 149136
rect 472062 148900 472094 149136
rect 471474 148816 472094 148900
rect 471474 148580 471506 148816
rect 471742 148580 471826 148816
rect 472062 148580 472094 148816
rect 471474 113136 472094 148580
rect 471474 112900 471506 113136
rect 471742 112900 471826 113136
rect 472062 112900 472094 113136
rect 471474 112816 472094 112900
rect 471474 112580 471506 112816
rect 471742 112580 471826 112816
rect 472062 112580 472094 112816
rect 471474 77136 472094 112580
rect 471474 76900 471506 77136
rect 471742 76900 471826 77136
rect 472062 76900 472094 77136
rect 471474 76816 472094 76900
rect 471474 76580 471506 76816
rect 471742 76580 471826 76816
rect 472062 76580 472094 76816
rect 471474 41136 472094 76580
rect 471474 40900 471506 41136
rect 471742 40900 471826 41136
rect 472062 40900 472094 41136
rect 471474 40816 472094 40900
rect 471474 40580 471506 40816
rect 471742 40580 471826 40816
rect 472062 40580 472094 40816
rect 471474 5136 472094 40580
rect 471474 4900 471506 5136
rect 471742 4900 471826 5136
rect 472062 4900 472094 5136
rect 471474 4816 472094 4900
rect 471474 4580 471506 4816
rect 471742 4580 471826 4816
rect 472062 4580 472094 4816
rect 471474 -2264 472094 4580
rect 471474 -2500 471506 -2264
rect 471742 -2500 471826 -2264
rect 472062 -2500 472094 -2264
rect 471474 -2584 472094 -2500
rect 471474 -2820 471506 -2584
rect 471742 -2820 471826 -2584
rect 472062 -2820 472094 -2584
rect 471474 -7652 472094 -2820
rect 472714 258376 473334 263617
rect 472714 258140 472746 258376
rect 472982 258140 473066 258376
rect 473302 258140 473334 258376
rect 472714 258056 473334 258140
rect 472714 257820 472746 258056
rect 472982 257820 473066 258056
rect 473302 257820 473334 258056
rect 472714 222376 473334 257820
rect 472714 222140 472746 222376
rect 472982 222140 473066 222376
rect 473302 222140 473334 222376
rect 472714 222056 473334 222140
rect 472714 221820 472746 222056
rect 472982 221820 473066 222056
rect 473302 221820 473334 222056
rect 472714 186376 473334 221820
rect 472714 186140 472746 186376
rect 472982 186140 473066 186376
rect 473302 186140 473334 186376
rect 472714 186056 473334 186140
rect 472714 185820 472746 186056
rect 472982 185820 473066 186056
rect 473302 185820 473334 186056
rect 472714 150376 473334 185820
rect 472714 150140 472746 150376
rect 472982 150140 473066 150376
rect 473302 150140 473334 150376
rect 472714 150056 473334 150140
rect 472714 149820 472746 150056
rect 472982 149820 473066 150056
rect 473302 149820 473334 150056
rect 472714 114376 473334 149820
rect 472714 114140 472746 114376
rect 472982 114140 473066 114376
rect 473302 114140 473334 114376
rect 472714 114056 473334 114140
rect 472714 113820 472746 114056
rect 472982 113820 473066 114056
rect 473302 113820 473334 114056
rect 472714 78376 473334 113820
rect 472714 78140 472746 78376
rect 472982 78140 473066 78376
rect 473302 78140 473334 78376
rect 472714 78056 473334 78140
rect 472714 77820 472746 78056
rect 472982 77820 473066 78056
rect 473302 77820 473334 78056
rect 472714 42376 473334 77820
rect 472714 42140 472746 42376
rect 472982 42140 473066 42376
rect 473302 42140 473334 42376
rect 472714 42056 473334 42140
rect 472714 41820 472746 42056
rect 472982 41820 473066 42056
rect 473302 41820 473334 42056
rect 472714 6376 473334 41820
rect 472714 6140 472746 6376
rect 472982 6140 473066 6376
rect 473302 6140 473334 6376
rect 472714 6056 473334 6140
rect 472714 5820 472746 6056
rect 472982 5820 473066 6056
rect 473302 5820 473334 6056
rect 472714 -3224 473334 5820
rect 472714 -3460 472746 -3224
rect 472982 -3460 473066 -3224
rect 473302 -3460 473334 -3224
rect 472714 -3544 473334 -3460
rect 472714 -3780 472746 -3544
rect 472982 -3780 473066 -3544
rect 473302 -3780 473334 -3544
rect 472714 -7652 473334 -3780
rect 473954 259616 474574 263617
rect 473954 259380 473986 259616
rect 474222 259380 474306 259616
rect 474542 259380 474574 259616
rect 473954 259296 474574 259380
rect 473954 259060 473986 259296
rect 474222 259060 474306 259296
rect 474542 259060 474574 259296
rect 473954 223616 474574 259060
rect 473954 223380 473986 223616
rect 474222 223380 474306 223616
rect 474542 223380 474574 223616
rect 473954 223296 474574 223380
rect 473954 223060 473986 223296
rect 474222 223060 474306 223296
rect 474542 223060 474574 223296
rect 473954 187616 474574 223060
rect 473954 187380 473986 187616
rect 474222 187380 474306 187616
rect 474542 187380 474574 187616
rect 473954 187296 474574 187380
rect 473954 187060 473986 187296
rect 474222 187060 474306 187296
rect 474542 187060 474574 187296
rect 473954 151616 474574 187060
rect 473954 151380 473986 151616
rect 474222 151380 474306 151616
rect 474542 151380 474574 151616
rect 473954 151296 474574 151380
rect 473954 151060 473986 151296
rect 474222 151060 474306 151296
rect 474542 151060 474574 151296
rect 473954 115616 474574 151060
rect 473954 115380 473986 115616
rect 474222 115380 474306 115616
rect 474542 115380 474574 115616
rect 473954 115296 474574 115380
rect 473954 115060 473986 115296
rect 474222 115060 474306 115296
rect 474542 115060 474574 115296
rect 473954 79616 474574 115060
rect 473954 79380 473986 79616
rect 474222 79380 474306 79616
rect 474542 79380 474574 79616
rect 473954 79296 474574 79380
rect 473954 79060 473986 79296
rect 474222 79060 474306 79296
rect 474542 79060 474574 79296
rect 473954 43616 474574 79060
rect 473954 43380 473986 43616
rect 474222 43380 474306 43616
rect 474542 43380 474574 43616
rect 473954 43296 474574 43380
rect 473954 43060 473986 43296
rect 474222 43060 474306 43296
rect 474542 43060 474574 43296
rect 473954 7616 474574 43060
rect 473954 7380 473986 7616
rect 474222 7380 474306 7616
rect 474542 7380 474574 7616
rect 473954 7296 474574 7380
rect 473954 7060 473986 7296
rect 474222 7060 474306 7296
rect 474542 7060 474574 7296
rect 473954 -4184 474574 7060
rect 473954 -4420 473986 -4184
rect 474222 -4420 474306 -4184
rect 474542 -4420 474574 -4184
rect 473954 -4504 474574 -4420
rect 473954 -4740 473986 -4504
rect 474222 -4740 474306 -4504
rect 474542 -4740 474574 -4504
rect 473954 -7652 474574 -4740
rect 475194 260856 475814 263617
rect 475194 260620 475226 260856
rect 475462 260620 475546 260856
rect 475782 260620 475814 260856
rect 475194 260536 475814 260620
rect 475194 260300 475226 260536
rect 475462 260300 475546 260536
rect 475782 260300 475814 260536
rect 475194 224856 475814 260300
rect 475194 224620 475226 224856
rect 475462 224620 475546 224856
rect 475782 224620 475814 224856
rect 475194 224536 475814 224620
rect 475194 224300 475226 224536
rect 475462 224300 475546 224536
rect 475782 224300 475814 224536
rect 475194 188856 475814 224300
rect 475194 188620 475226 188856
rect 475462 188620 475546 188856
rect 475782 188620 475814 188856
rect 475194 188536 475814 188620
rect 475194 188300 475226 188536
rect 475462 188300 475546 188536
rect 475782 188300 475814 188536
rect 475194 152856 475814 188300
rect 475194 152620 475226 152856
rect 475462 152620 475546 152856
rect 475782 152620 475814 152856
rect 475194 152536 475814 152620
rect 475194 152300 475226 152536
rect 475462 152300 475546 152536
rect 475782 152300 475814 152536
rect 475194 116856 475814 152300
rect 475194 116620 475226 116856
rect 475462 116620 475546 116856
rect 475782 116620 475814 116856
rect 475194 116536 475814 116620
rect 475194 116300 475226 116536
rect 475462 116300 475546 116536
rect 475782 116300 475814 116536
rect 475194 80856 475814 116300
rect 475194 80620 475226 80856
rect 475462 80620 475546 80856
rect 475782 80620 475814 80856
rect 475194 80536 475814 80620
rect 475194 80300 475226 80536
rect 475462 80300 475546 80536
rect 475782 80300 475814 80536
rect 475194 44856 475814 80300
rect 475194 44620 475226 44856
rect 475462 44620 475546 44856
rect 475782 44620 475814 44856
rect 475194 44536 475814 44620
rect 475194 44300 475226 44536
rect 475462 44300 475546 44536
rect 475782 44300 475814 44536
rect 475194 8856 475814 44300
rect 475194 8620 475226 8856
rect 475462 8620 475546 8856
rect 475782 8620 475814 8856
rect 475194 8536 475814 8620
rect 475194 8300 475226 8536
rect 475462 8300 475546 8536
rect 475782 8300 475814 8536
rect 475194 -5144 475814 8300
rect 475194 -5380 475226 -5144
rect 475462 -5380 475546 -5144
rect 475782 -5380 475814 -5144
rect 475194 -5464 475814 -5380
rect 475194 -5700 475226 -5464
rect 475462 -5700 475546 -5464
rect 475782 -5700 475814 -5464
rect 475194 -7652 475814 -5700
rect 476434 262096 477054 263617
rect 476434 261860 476466 262096
rect 476702 261860 476786 262096
rect 477022 261860 477054 262096
rect 476434 261776 477054 261860
rect 476434 261540 476466 261776
rect 476702 261540 476786 261776
rect 477022 261540 477054 261776
rect 476434 226096 477054 261540
rect 476434 225860 476466 226096
rect 476702 225860 476786 226096
rect 477022 225860 477054 226096
rect 476434 225776 477054 225860
rect 476434 225540 476466 225776
rect 476702 225540 476786 225776
rect 477022 225540 477054 225776
rect 476434 190096 477054 225540
rect 477358 205735 477418 264965
rect 477674 263336 478294 263617
rect 477674 263100 477706 263336
rect 477942 263100 478026 263336
rect 478262 263100 478294 263336
rect 477674 263016 478294 263100
rect 477674 262780 477706 263016
rect 477942 262780 478026 263016
rect 478262 262780 478294 263016
rect 477674 227336 478294 262780
rect 480118 245583 480178 264965
rect 504994 254656 505614 290100
rect 504994 254420 505026 254656
rect 505262 254420 505346 254656
rect 505582 254420 505614 254656
rect 504994 254336 505614 254420
rect 504994 254100 505026 254336
rect 505262 254100 505346 254336
rect 505582 254100 505614 254336
rect 480115 245582 480181 245583
rect 480115 245518 480116 245582
rect 480180 245518 480181 245582
rect 480115 245517 480181 245518
rect 477674 227100 477706 227336
rect 477942 227100 478026 227336
rect 478262 227100 478294 227336
rect 477674 227016 478294 227100
rect 477674 226780 477706 227016
rect 477942 226780 478026 227016
rect 478262 226780 478294 227016
rect 477355 205734 477421 205735
rect 477355 205670 477356 205734
rect 477420 205670 477421 205734
rect 477355 205669 477421 205670
rect 476434 189860 476466 190096
rect 476702 189860 476786 190096
rect 477022 189860 477054 190096
rect 476434 189776 477054 189860
rect 476434 189540 476466 189776
rect 476702 189540 476786 189776
rect 477022 189540 477054 189776
rect 476434 154096 477054 189540
rect 476434 153860 476466 154096
rect 476702 153860 476786 154096
rect 477022 153860 477054 154096
rect 476434 153776 477054 153860
rect 476434 153540 476466 153776
rect 476702 153540 476786 153776
rect 477022 153540 477054 153776
rect 476434 118096 477054 153540
rect 476434 117860 476466 118096
rect 476702 117860 476786 118096
rect 477022 117860 477054 118096
rect 476434 117776 477054 117860
rect 476434 117540 476466 117776
rect 476702 117540 476786 117776
rect 477022 117540 477054 117776
rect 476434 82096 477054 117540
rect 476434 81860 476466 82096
rect 476702 81860 476786 82096
rect 477022 81860 477054 82096
rect 476434 81776 477054 81860
rect 476434 81540 476466 81776
rect 476702 81540 476786 81776
rect 477022 81540 477054 81776
rect 476434 46096 477054 81540
rect 476434 45860 476466 46096
rect 476702 45860 476786 46096
rect 477022 45860 477054 46096
rect 476434 45776 477054 45860
rect 476434 45540 476466 45776
rect 476702 45540 476786 45776
rect 477022 45540 477054 45776
rect 476434 10096 477054 45540
rect 476434 9860 476466 10096
rect 476702 9860 476786 10096
rect 477022 9860 477054 10096
rect 476434 9776 477054 9860
rect 476434 9540 476466 9776
rect 476702 9540 476786 9776
rect 477022 9540 477054 9776
rect 476434 -6104 477054 9540
rect 476434 -6340 476466 -6104
rect 476702 -6340 476786 -6104
rect 477022 -6340 477054 -6104
rect 476434 -6424 477054 -6340
rect 476434 -6660 476466 -6424
rect 476702 -6660 476786 -6424
rect 477022 -6660 477054 -6424
rect 476434 -7652 477054 -6660
rect 477674 191336 478294 226780
rect 477674 191100 477706 191336
rect 477942 191100 478026 191336
rect 478262 191100 478294 191336
rect 477674 191016 478294 191100
rect 477674 190780 477706 191016
rect 477942 190780 478026 191016
rect 478262 190780 478294 191016
rect 477674 155336 478294 190780
rect 477674 155100 477706 155336
rect 477942 155100 478026 155336
rect 478262 155100 478294 155336
rect 477674 155016 478294 155100
rect 477674 154780 477706 155016
rect 477942 154780 478026 155016
rect 478262 154780 478294 155016
rect 477674 119336 478294 154780
rect 477674 119100 477706 119336
rect 477942 119100 478026 119336
rect 478262 119100 478294 119336
rect 477674 119016 478294 119100
rect 477674 118780 477706 119016
rect 477942 118780 478026 119016
rect 478262 118780 478294 119016
rect 477674 83336 478294 118780
rect 477674 83100 477706 83336
rect 477942 83100 478026 83336
rect 478262 83100 478294 83336
rect 477674 83016 478294 83100
rect 477674 82780 477706 83016
rect 477942 82780 478026 83016
rect 478262 82780 478294 83016
rect 477674 47336 478294 82780
rect 477674 47100 477706 47336
rect 477942 47100 478026 47336
rect 478262 47100 478294 47336
rect 477674 47016 478294 47100
rect 477674 46780 477706 47016
rect 477942 46780 478026 47016
rect 478262 46780 478294 47016
rect 477674 11336 478294 46780
rect 477674 11100 477706 11336
rect 477942 11100 478026 11336
rect 478262 11100 478294 11336
rect 477674 11016 478294 11100
rect 477674 10780 477706 11016
rect 477942 10780 478026 11016
rect 478262 10780 478294 11016
rect 477674 -7064 478294 10780
rect 477674 -7300 477706 -7064
rect 477942 -7300 478026 -7064
rect 478262 -7300 478294 -7064
rect 477674 -7384 478294 -7300
rect 477674 -7620 477706 -7384
rect 477942 -7620 478026 -7384
rect 478262 -7620 478294 -7384
rect 477674 -7652 478294 -7620
rect 504994 218656 505614 254100
rect 504994 218420 505026 218656
rect 505262 218420 505346 218656
rect 505582 218420 505614 218656
rect 504994 218336 505614 218420
rect 504994 218100 505026 218336
rect 505262 218100 505346 218336
rect 505582 218100 505614 218336
rect 504994 182656 505614 218100
rect 504994 182420 505026 182656
rect 505262 182420 505346 182656
rect 505582 182420 505614 182656
rect 504994 182336 505614 182420
rect 504994 182100 505026 182336
rect 505262 182100 505346 182336
rect 505582 182100 505614 182336
rect 504994 146656 505614 182100
rect 504994 146420 505026 146656
rect 505262 146420 505346 146656
rect 505582 146420 505614 146656
rect 504994 146336 505614 146420
rect 504994 146100 505026 146336
rect 505262 146100 505346 146336
rect 505582 146100 505614 146336
rect 504994 110656 505614 146100
rect 504994 110420 505026 110656
rect 505262 110420 505346 110656
rect 505582 110420 505614 110656
rect 504994 110336 505614 110420
rect 504994 110100 505026 110336
rect 505262 110100 505346 110336
rect 505582 110100 505614 110336
rect 504994 74656 505614 110100
rect 504994 74420 505026 74656
rect 505262 74420 505346 74656
rect 505582 74420 505614 74656
rect 504994 74336 505614 74420
rect 504994 74100 505026 74336
rect 505262 74100 505346 74336
rect 505582 74100 505614 74336
rect 504994 38656 505614 74100
rect 504994 38420 505026 38656
rect 505262 38420 505346 38656
rect 505582 38420 505614 38656
rect 504994 38336 505614 38420
rect 504994 38100 505026 38336
rect 505262 38100 505346 38336
rect 505582 38100 505614 38336
rect 504994 2656 505614 38100
rect 504994 2420 505026 2656
rect 505262 2420 505346 2656
rect 505582 2420 505614 2656
rect 504994 2336 505614 2420
rect 504994 2100 505026 2336
rect 505262 2100 505346 2336
rect 505582 2100 505614 2336
rect 504994 -344 505614 2100
rect 504994 -580 505026 -344
rect 505262 -580 505346 -344
rect 505582 -580 505614 -344
rect 504994 -664 505614 -580
rect 504994 -900 505026 -664
rect 505262 -900 505346 -664
rect 505582 -900 505614 -664
rect 504994 -7652 505614 -900
rect 506234 705800 506854 711592
rect 506234 705564 506266 705800
rect 506502 705564 506586 705800
rect 506822 705564 506854 705800
rect 506234 705480 506854 705564
rect 506234 705244 506266 705480
rect 506502 705244 506586 705480
rect 506822 705244 506854 705480
rect 506234 702524 506854 705244
rect 506234 702460 506272 702524
rect 506336 702460 506352 702524
rect 506416 702460 506432 702524
rect 506496 702460 506512 702524
rect 506576 702460 506592 702524
rect 506656 702460 506672 702524
rect 506736 702460 506752 702524
rect 506816 702460 506854 702524
rect 506234 702444 506854 702460
rect 506234 702380 506272 702444
rect 506336 702380 506352 702444
rect 506416 702380 506432 702444
rect 506496 702380 506512 702444
rect 506576 702380 506592 702444
rect 506656 702380 506672 702444
rect 506736 702380 506752 702444
rect 506816 702380 506854 702444
rect 506234 702364 506854 702380
rect 506234 702300 506272 702364
rect 506336 702300 506352 702364
rect 506416 702300 506432 702364
rect 506496 702300 506512 702364
rect 506576 702300 506592 702364
rect 506656 702300 506672 702364
rect 506736 702300 506752 702364
rect 506816 702300 506854 702364
rect 506234 702284 506854 702300
rect 506234 702220 506272 702284
rect 506336 702220 506352 702284
rect 506416 702220 506432 702284
rect 506496 702220 506512 702284
rect 506576 702220 506592 702284
rect 506656 702220 506672 702284
rect 506736 702220 506752 702284
rect 506816 702220 506854 702284
rect 506234 687896 506854 702220
rect 506234 687660 506266 687896
rect 506502 687660 506586 687896
rect 506822 687660 506854 687896
rect 506234 687576 506854 687660
rect 506234 687340 506266 687576
rect 506502 687340 506586 687576
rect 506822 687340 506854 687576
rect 506234 651896 506854 687340
rect 506234 651660 506266 651896
rect 506502 651660 506586 651896
rect 506822 651660 506854 651896
rect 506234 651576 506854 651660
rect 506234 651340 506266 651576
rect 506502 651340 506586 651576
rect 506822 651340 506854 651576
rect 506234 615896 506854 651340
rect 506234 615660 506266 615896
rect 506502 615660 506586 615896
rect 506822 615660 506854 615896
rect 506234 615576 506854 615660
rect 506234 615340 506266 615576
rect 506502 615340 506586 615576
rect 506822 615340 506854 615576
rect 506234 579896 506854 615340
rect 506234 579660 506266 579896
rect 506502 579660 506586 579896
rect 506822 579660 506854 579896
rect 506234 579576 506854 579660
rect 506234 579340 506266 579576
rect 506502 579340 506586 579576
rect 506822 579340 506854 579576
rect 506234 553807 506854 579340
rect 506234 553743 506272 553807
rect 506336 553743 506352 553807
rect 506416 553743 506432 553807
rect 506496 553743 506512 553807
rect 506576 553743 506592 553807
rect 506656 553743 506672 553807
rect 506736 553743 506752 553807
rect 506816 553743 506854 553807
rect 506234 553727 506854 553743
rect 506234 553663 506272 553727
rect 506336 553663 506352 553727
rect 506416 553663 506432 553727
rect 506496 553663 506512 553727
rect 506576 553663 506592 553727
rect 506656 553663 506672 553727
rect 506736 553663 506752 553727
rect 506816 553663 506854 553727
rect 506234 553647 506854 553663
rect 506234 553583 506272 553647
rect 506336 553583 506352 553647
rect 506416 553583 506432 553647
rect 506496 553583 506512 553647
rect 506576 553583 506592 553647
rect 506656 553583 506672 553647
rect 506736 553583 506752 553647
rect 506816 553583 506854 553647
rect 506234 553567 506854 553583
rect 506234 553503 506272 553567
rect 506336 553503 506352 553567
rect 506416 553503 506432 553567
rect 506496 553503 506512 553567
rect 506576 553503 506592 553567
rect 506656 553503 506672 553567
rect 506736 553503 506752 553567
rect 506816 553503 506854 553567
rect 506234 543896 506854 553503
rect 506234 543660 506266 543896
rect 506502 543660 506586 543896
rect 506822 543660 506854 543896
rect 506234 543576 506854 543660
rect 506234 543340 506266 543576
rect 506502 543340 506586 543576
rect 506822 543340 506854 543576
rect 506234 507896 506854 543340
rect 506234 507660 506266 507896
rect 506502 507660 506586 507896
rect 506822 507660 506854 507896
rect 506234 507576 506854 507660
rect 506234 507340 506266 507576
rect 506502 507340 506586 507576
rect 506822 507340 506854 507576
rect 506234 471896 506854 507340
rect 506234 471660 506266 471896
rect 506502 471660 506586 471896
rect 506822 471660 506854 471896
rect 506234 471576 506854 471660
rect 506234 471340 506266 471576
rect 506502 471340 506586 471576
rect 506822 471340 506854 471576
rect 506234 435896 506854 471340
rect 506234 435660 506266 435896
rect 506502 435660 506586 435896
rect 506822 435660 506854 435896
rect 506234 435576 506854 435660
rect 506234 435340 506266 435576
rect 506502 435340 506586 435576
rect 506822 435340 506854 435576
rect 506234 399896 506854 435340
rect 506234 399660 506266 399896
rect 506502 399660 506586 399896
rect 506822 399660 506854 399896
rect 506234 399576 506854 399660
rect 506234 399340 506266 399576
rect 506502 399340 506586 399576
rect 506822 399340 506854 399576
rect 506234 363896 506854 399340
rect 506234 363660 506266 363896
rect 506502 363660 506586 363896
rect 506822 363660 506854 363896
rect 506234 363576 506854 363660
rect 506234 363340 506266 363576
rect 506502 363340 506586 363576
rect 506822 363340 506854 363576
rect 506234 327896 506854 363340
rect 506234 327660 506266 327896
rect 506502 327660 506586 327896
rect 506822 327660 506854 327896
rect 506234 327576 506854 327660
rect 506234 327340 506266 327576
rect 506502 327340 506586 327576
rect 506822 327340 506854 327576
rect 506234 291896 506854 327340
rect 506234 291660 506266 291896
rect 506502 291660 506586 291896
rect 506822 291660 506854 291896
rect 506234 291576 506854 291660
rect 506234 291340 506266 291576
rect 506502 291340 506586 291576
rect 506822 291340 506854 291576
rect 506234 255896 506854 291340
rect 506234 255660 506266 255896
rect 506502 255660 506586 255896
rect 506822 255660 506854 255896
rect 506234 255576 506854 255660
rect 506234 255340 506266 255576
rect 506502 255340 506586 255576
rect 506822 255340 506854 255576
rect 506234 219896 506854 255340
rect 506234 219660 506266 219896
rect 506502 219660 506586 219896
rect 506822 219660 506854 219896
rect 506234 219576 506854 219660
rect 506234 219340 506266 219576
rect 506502 219340 506586 219576
rect 506822 219340 506854 219576
rect 506234 183896 506854 219340
rect 506234 183660 506266 183896
rect 506502 183660 506586 183896
rect 506822 183660 506854 183896
rect 506234 183576 506854 183660
rect 506234 183340 506266 183576
rect 506502 183340 506586 183576
rect 506822 183340 506854 183576
rect 506234 147896 506854 183340
rect 506234 147660 506266 147896
rect 506502 147660 506586 147896
rect 506822 147660 506854 147896
rect 506234 147576 506854 147660
rect 506234 147340 506266 147576
rect 506502 147340 506586 147576
rect 506822 147340 506854 147576
rect 506234 111896 506854 147340
rect 506234 111660 506266 111896
rect 506502 111660 506586 111896
rect 506822 111660 506854 111896
rect 506234 111576 506854 111660
rect 506234 111340 506266 111576
rect 506502 111340 506586 111576
rect 506822 111340 506854 111576
rect 506234 75896 506854 111340
rect 506234 75660 506266 75896
rect 506502 75660 506586 75896
rect 506822 75660 506854 75896
rect 506234 75576 506854 75660
rect 506234 75340 506266 75576
rect 506502 75340 506586 75576
rect 506822 75340 506854 75576
rect 506234 39896 506854 75340
rect 506234 39660 506266 39896
rect 506502 39660 506586 39896
rect 506822 39660 506854 39896
rect 506234 39576 506854 39660
rect 506234 39340 506266 39576
rect 506502 39340 506586 39576
rect 506822 39340 506854 39576
rect 506234 3896 506854 39340
rect 506234 3660 506266 3896
rect 506502 3660 506586 3896
rect 506822 3660 506854 3896
rect 506234 3576 506854 3660
rect 506234 3340 506266 3576
rect 506502 3340 506586 3576
rect 506822 3340 506854 3576
rect 506234 -1304 506854 3340
rect 506234 -1540 506266 -1304
rect 506502 -1540 506586 -1304
rect 506822 -1540 506854 -1304
rect 506234 -1624 506854 -1540
rect 506234 -1860 506266 -1624
rect 506502 -1860 506586 -1624
rect 506822 -1860 506854 -1624
rect 506234 -7652 506854 -1860
rect 507474 706760 508094 711592
rect 507474 706524 507506 706760
rect 507742 706524 507826 706760
rect 508062 706524 508094 706760
rect 507474 706440 508094 706524
rect 507474 706204 507506 706440
rect 507742 706204 507826 706440
rect 508062 706204 508094 706440
rect 507474 689136 508094 706204
rect 507474 688900 507506 689136
rect 507742 688900 507826 689136
rect 508062 688900 508094 689136
rect 507474 688816 508094 688900
rect 507474 688580 507506 688816
rect 507742 688580 507826 688816
rect 508062 688580 508094 688816
rect 507474 653136 508094 688580
rect 507474 652900 507506 653136
rect 507742 652900 507826 653136
rect 508062 652900 508094 653136
rect 507474 652816 508094 652900
rect 507474 652580 507506 652816
rect 507742 652580 507826 652816
rect 508062 652580 508094 652816
rect 507474 617136 508094 652580
rect 507474 616900 507506 617136
rect 507742 616900 507826 617136
rect 508062 616900 508094 617136
rect 507474 616816 508094 616900
rect 507474 616580 507506 616816
rect 507742 616580 507826 616816
rect 508062 616580 508094 616816
rect 507474 581136 508094 616580
rect 507474 580900 507506 581136
rect 507742 580900 507826 581136
rect 508062 580900 508094 581136
rect 507474 580816 508094 580900
rect 507474 580580 507506 580816
rect 507742 580580 507826 580816
rect 508062 580580 508094 580816
rect 507474 545136 508094 580580
rect 507474 544900 507506 545136
rect 507742 544900 507826 545136
rect 508062 544900 508094 545136
rect 507474 544816 508094 544900
rect 507474 544580 507506 544816
rect 507742 544580 507826 544816
rect 508062 544580 508094 544816
rect 507474 509136 508094 544580
rect 507474 508900 507506 509136
rect 507742 508900 507826 509136
rect 508062 508900 508094 509136
rect 507474 508816 508094 508900
rect 507474 508580 507506 508816
rect 507742 508580 507826 508816
rect 508062 508580 508094 508816
rect 507474 473136 508094 508580
rect 507474 472900 507506 473136
rect 507742 472900 507826 473136
rect 508062 472900 508094 473136
rect 507474 472816 508094 472900
rect 507474 472580 507506 472816
rect 507742 472580 507826 472816
rect 508062 472580 508094 472816
rect 507474 437136 508094 472580
rect 507474 436900 507506 437136
rect 507742 436900 507826 437136
rect 508062 436900 508094 437136
rect 507474 436816 508094 436900
rect 507474 436580 507506 436816
rect 507742 436580 507826 436816
rect 508062 436580 508094 436816
rect 507474 401136 508094 436580
rect 507474 400900 507506 401136
rect 507742 400900 507826 401136
rect 508062 400900 508094 401136
rect 507474 400816 508094 400900
rect 507474 400580 507506 400816
rect 507742 400580 507826 400816
rect 508062 400580 508094 400816
rect 507474 365136 508094 400580
rect 507474 364900 507506 365136
rect 507742 364900 507826 365136
rect 508062 364900 508094 365136
rect 507474 364816 508094 364900
rect 507474 364580 507506 364816
rect 507742 364580 507826 364816
rect 508062 364580 508094 364816
rect 507474 329136 508094 364580
rect 507474 328900 507506 329136
rect 507742 328900 507826 329136
rect 508062 328900 508094 329136
rect 507474 328816 508094 328900
rect 507474 328580 507506 328816
rect 507742 328580 507826 328816
rect 508062 328580 508094 328816
rect 507474 293136 508094 328580
rect 507474 292900 507506 293136
rect 507742 292900 507826 293136
rect 508062 292900 508094 293136
rect 507474 292816 508094 292900
rect 507474 292580 507506 292816
rect 507742 292580 507826 292816
rect 508062 292580 508094 292816
rect 507474 257136 508094 292580
rect 507474 256900 507506 257136
rect 507742 256900 507826 257136
rect 508062 256900 508094 257136
rect 507474 256816 508094 256900
rect 507474 256580 507506 256816
rect 507742 256580 507826 256816
rect 508062 256580 508094 256816
rect 507474 221136 508094 256580
rect 507474 220900 507506 221136
rect 507742 220900 507826 221136
rect 508062 220900 508094 221136
rect 507474 220816 508094 220900
rect 507474 220580 507506 220816
rect 507742 220580 507826 220816
rect 508062 220580 508094 220816
rect 507474 185136 508094 220580
rect 507474 184900 507506 185136
rect 507742 184900 507826 185136
rect 508062 184900 508094 185136
rect 507474 184816 508094 184900
rect 507474 184580 507506 184816
rect 507742 184580 507826 184816
rect 508062 184580 508094 184816
rect 507474 149136 508094 184580
rect 507474 148900 507506 149136
rect 507742 148900 507826 149136
rect 508062 148900 508094 149136
rect 507474 148816 508094 148900
rect 507474 148580 507506 148816
rect 507742 148580 507826 148816
rect 508062 148580 508094 148816
rect 507474 113136 508094 148580
rect 507474 112900 507506 113136
rect 507742 112900 507826 113136
rect 508062 112900 508094 113136
rect 507474 112816 508094 112900
rect 507474 112580 507506 112816
rect 507742 112580 507826 112816
rect 508062 112580 508094 112816
rect 507474 77136 508094 112580
rect 507474 76900 507506 77136
rect 507742 76900 507826 77136
rect 508062 76900 508094 77136
rect 507474 76816 508094 76900
rect 507474 76580 507506 76816
rect 507742 76580 507826 76816
rect 508062 76580 508094 76816
rect 507474 41136 508094 76580
rect 507474 40900 507506 41136
rect 507742 40900 507826 41136
rect 508062 40900 508094 41136
rect 507474 40816 508094 40900
rect 507474 40580 507506 40816
rect 507742 40580 507826 40816
rect 508062 40580 508094 40816
rect 507474 5136 508094 40580
rect 507474 4900 507506 5136
rect 507742 4900 507826 5136
rect 508062 4900 508094 5136
rect 507474 4816 508094 4900
rect 507474 4580 507506 4816
rect 507742 4580 507826 4816
rect 508062 4580 508094 4816
rect 507474 -2264 508094 4580
rect 507474 -2500 507506 -2264
rect 507742 -2500 507826 -2264
rect 508062 -2500 508094 -2264
rect 507474 -2584 508094 -2500
rect 507474 -2820 507506 -2584
rect 507742 -2820 507826 -2584
rect 508062 -2820 508094 -2584
rect 507474 -7652 508094 -2820
rect 508714 707720 509334 711592
rect 508714 707484 508746 707720
rect 508982 707484 509066 707720
rect 509302 707484 509334 707720
rect 508714 707400 509334 707484
rect 508714 707164 508746 707400
rect 508982 707164 509066 707400
rect 509302 707164 509334 707400
rect 508714 690376 509334 707164
rect 508714 690140 508746 690376
rect 508982 690140 509066 690376
rect 509302 690140 509334 690376
rect 508714 690056 509334 690140
rect 508714 689820 508746 690056
rect 508982 689820 509066 690056
rect 509302 689820 509334 690056
rect 508714 654376 509334 689820
rect 508714 654140 508746 654376
rect 508982 654140 509066 654376
rect 509302 654140 509334 654376
rect 508714 654056 509334 654140
rect 508714 653820 508746 654056
rect 508982 653820 509066 654056
rect 509302 653820 509334 654056
rect 508714 618376 509334 653820
rect 508714 618140 508746 618376
rect 508982 618140 509066 618376
rect 509302 618140 509334 618376
rect 508714 618056 509334 618140
rect 508714 617820 508746 618056
rect 508982 617820 509066 618056
rect 509302 617820 509334 618056
rect 508714 582376 509334 617820
rect 508714 582140 508746 582376
rect 508982 582140 509066 582376
rect 509302 582140 509334 582376
rect 508714 582056 509334 582140
rect 508714 581820 508746 582056
rect 508982 581820 509066 582056
rect 509302 581820 509334 582056
rect 508714 546376 509334 581820
rect 508714 546140 508746 546376
rect 508982 546140 509066 546376
rect 509302 546140 509334 546376
rect 508714 546056 509334 546140
rect 508714 545820 508746 546056
rect 508982 545820 509066 546056
rect 509302 545820 509334 546056
rect 508714 510376 509334 545820
rect 508714 510140 508746 510376
rect 508982 510140 509066 510376
rect 509302 510140 509334 510376
rect 508714 510056 509334 510140
rect 508714 509820 508746 510056
rect 508982 509820 509066 510056
rect 509302 509820 509334 510056
rect 508714 474376 509334 509820
rect 508714 474140 508746 474376
rect 508982 474140 509066 474376
rect 509302 474140 509334 474376
rect 508714 474056 509334 474140
rect 508714 473820 508746 474056
rect 508982 473820 509066 474056
rect 509302 473820 509334 474056
rect 508714 438376 509334 473820
rect 508714 438140 508746 438376
rect 508982 438140 509066 438376
rect 509302 438140 509334 438376
rect 508714 438056 509334 438140
rect 508714 437820 508746 438056
rect 508982 437820 509066 438056
rect 509302 437820 509334 438056
rect 508714 402376 509334 437820
rect 508714 402140 508746 402376
rect 508982 402140 509066 402376
rect 509302 402140 509334 402376
rect 508714 402056 509334 402140
rect 508714 401820 508746 402056
rect 508982 401820 509066 402056
rect 509302 401820 509334 402056
rect 508714 366376 509334 401820
rect 508714 366140 508746 366376
rect 508982 366140 509066 366376
rect 509302 366140 509334 366376
rect 508714 366056 509334 366140
rect 508714 365820 508746 366056
rect 508982 365820 509066 366056
rect 509302 365820 509334 366056
rect 508714 330376 509334 365820
rect 508714 330140 508746 330376
rect 508982 330140 509066 330376
rect 509302 330140 509334 330376
rect 508714 330056 509334 330140
rect 508714 329820 508746 330056
rect 508982 329820 509066 330056
rect 509302 329820 509334 330056
rect 508714 294376 509334 329820
rect 508714 294140 508746 294376
rect 508982 294140 509066 294376
rect 509302 294140 509334 294376
rect 508714 294056 509334 294140
rect 508714 293820 508746 294056
rect 508982 293820 509066 294056
rect 509302 293820 509334 294056
rect 508714 258376 509334 293820
rect 508714 258140 508746 258376
rect 508982 258140 509066 258376
rect 509302 258140 509334 258376
rect 508714 258056 509334 258140
rect 508714 257820 508746 258056
rect 508982 257820 509066 258056
rect 509302 257820 509334 258056
rect 508714 222376 509334 257820
rect 508714 222140 508746 222376
rect 508982 222140 509066 222376
rect 509302 222140 509334 222376
rect 508714 222056 509334 222140
rect 508714 221820 508746 222056
rect 508982 221820 509066 222056
rect 509302 221820 509334 222056
rect 508714 186376 509334 221820
rect 508714 186140 508746 186376
rect 508982 186140 509066 186376
rect 509302 186140 509334 186376
rect 508714 186056 509334 186140
rect 508714 185820 508746 186056
rect 508982 185820 509066 186056
rect 509302 185820 509334 186056
rect 508714 150376 509334 185820
rect 508714 150140 508746 150376
rect 508982 150140 509066 150376
rect 509302 150140 509334 150376
rect 508714 150056 509334 150140
rect 508714 149820 508746 150056
rect 508982 149820 509066 150056
rect 509302 149820 509334 150056
rect 508714 114376 509334 149820
rect 508714 114140 508746 114376
rect 508982 114140 509066 114376
rect 509302 114140 509334 114376
rect 508714 114056 509334 114140
rect 508714 113820 508746 114056
rect 508982 113820 509066 114056
rect 509302 113820 509334 114056
rect 508714 78376 509334 113820
rect 508714 78140 508746 78376
rect 508982 78140 509066 78376
rect 509302 78140 509334 78376
rect 508714 78056 509334 78140
rect 508714 77820 508746 78056
rect 508982 77820 509066 78056
rect 509302 77820 509334 78056
rect 508714 42376 509334 77820
rect 508714 42140 508746 42376
rect 508982 42140 509066 42376
rect 509302 42140 509334 42376
rect 508714 42056 509334 42140
rect 508714 41820 508746 42056
rect 508982 41820 509066 42056
rect 509302 41820 509334 42056
rect 508714 6376 509334 41820
rect 508714 6140 508746 6376
rect 508982 6140 509066 6376
rect 509302 6140 509334 6376
rect 508714 6056 509334 6140
rect 508714 5820 508746 6056
rect 508982 5820 509066 6056
rect 509302 5820 509334 6056
rect 508714 -3224 509334 5820
rect 508714 -3460 508746 -3224
rect 508982 -3460 509066 -3224
rect 509302 -3460 509334 -3224
rect 508714 -3544 509334 -3460
rect 508714 -3780 508746 -3544
rect 508982 -3780 509066 -3544
rect 509302 -3780 509334 -3544
rect 508714 -7652 509334 -3780
rect 509954 708680 510574 711592
rect 509954 708444 509986 708680
rect 510222 708444 510306 708680
rect 510542 708444 510574 708680
rect 509954 708360 510574 708444
rect 509954 708124 509986 708360
rect 510222 708124 510306 708360
rect 510542 708124 510574 708360
rect 509954 691616 510574 708124
rect 509954 691380 509986 691616
rect 510222 691380 510306 691616
rect 510542 691380 510574 691616
rect 509954 691296 510574 691380
rect 509954 691060 509986 691296
rect 510222 691060 510306 691296
rect 510542 691060 510574 691296
rect 509954 655616 510574 691060
rect 509954 655380 509986 655616
rect 510222 655380 510306 655616
rect 510542 655380 510574 655616
rect 509954 655296 510574 655380
rect 509954 655060 509986 655296
rect 510222 655060 510306 655296
rect 510542 655060 510574 655296
rect 509954 619616 510574 655060
rect 509954 619380 509986 619616
rect 510222 619380 510306 619616
rect 510542 619380 510574 619616
rect 509954 619296 510574 619380
rect 509954 619060 509986 619296
rect 510222 619060 510306 619296
rect 510542 619060 510574 619296
rect 509954 583616 510574 619060
rect 509954 583380 509986 583616
rect 510222 583380 510306 583616
rect 510542 583380 510574 583616
rect 509954 583296 510574 583380
rect 509954 583060 509986 583296
rect 510222 583060 510306 583296
rect 510542 583060 510574 583296
rect 509954 547616 510574 583060
rect 509954 547380 509986 547616
rect 510222 547380 510306 547616
rect 510542 547380 510574 547616
rect 509954 547296 510574 547380
rect 509954 547060 509986 547296
rect 510222 547060 510306 547296
rect 510542 547060 510574 547296
rect 509954 511616 510574 547060
rect 509954 511380 509986 511616
rect 510222 511380 510306 511616
rect 510542 511380 510574 511616
rect 509954 511296 510574 511380
rect 509954 511060 509986 511296
rect 510222 511060 510306 511296
rect 510542 511060 510574 511296
rect 509954 475616 510574 511060
rect 509954 475380 509986 475616
rect 510222 475380 510306 475616
rect 510542 475380 510574 475616
rect 509954 475296 510574 475380
rect 509954 475060 509986 475296
rect 510222 475060 510306 475296
rect 510542 475060 510574 475296
rect 509954 439616 510574 475060
rect 509954 439380 509986 439616
rect 510222 439380 510306 439616
rect 510542 439380 510574 439616
rect 509954 439296 510574 439380
rect 509954 439060 509986 439296
rect 510222 439060 510306 439296
rect 510542 439060 510574 439296
rect 509954 403616 510574 439060
rect 509954 403380 509986 403616
rect 510222 403380 510306 403616
rect 510542 403380 510574 403616
rect 509954 403296 510574 403380
rect 509954 403060 509986 403296
rect 510222 403060 510306 403296
rect 510542 403060 510574 403296
rect 509954 367616 510574 403060
rect 509954 367380 509986 367616
rect 510222 367380 510306 367616
rect 510542 367380 510574 367616
rect 509954 367296 510574 367380
rect 509954 367060 509986 367296
rect 510222 367060 510306 367296
rect 510542 367060 510574 367296
rect 509954 331616 510574 367060
rect 509954 331380 509986 331616
rect 510222 331380 510306 331616
rect 510542 331380 510574 331616
rect 509954 331296 510574 331380
rect 509954 331060 509986 331296
rect 510222 331060 510306 331296
rect 510542 331060 510574 331296
rect 509954 295616 510574 331060
rect 509954 295380 509986 295616
rect 510222 295380 510306 295616
rect 510542 295380 510574 295616
rect 509954 295296 510574 295380
rect 509954 295060 509986 295296
rect 510222 295060 510306 295296
rect 510542 295060 510574 295296
rect 509954 259616 510574 295060
rect 509954 259380 509986 259616
rect 510222 259380 510306 259616
rect 510542 259380 510574 259616
rect 509954 259296 510574 259380
rect 509954 259060 509986 259296
rect 510222 259060 510306 259296
rect 510542 259060 510574 259296
rect 509954 223616 510574 259060
rect 509954 223380 509986 223616
rect 510222 223380 510306 223616
rect 510542 223380 510574 223616
rect 509954 223296 510574 223380
rect 509954 223060 509986 223296
rect 510222 223060 510306 223296
rect 510542 223060 510574 223296
rect 509954 187616 510574 223060
rect 509954 187380 509986 187616
rect 510222 187380 510306 187616
rect 510542 187380 510574 187616
rect 509954 187296 510574 187380
rect 509954 187060 509986 187296
rect 510222 187060 510306 187296
rect 510542 187060 510574 187296
rect 509954 151616 510574 187060
rect 509954 151380 509986 151616
rect 510222 151380 510306 151616
rect 510542 151380 510574 151616
rect 509954 151296 510574 151380
rect 509954 151060 509986 151296
rect 510222 151060 510306 151296
rect 510542 151060 510574 151296
rect 509954 115616 510574 151060
rect 509954 115380 509986 115616
rect 510222 115380 510306 115616
rect 510542 115380 510574 115616
rect 509954 115296 510574 115380
rect 509954 115060 509986 115296
rect 510222 115060 510306 115296
rect 510542 115060 510574 115296
rect 509954 79616 510574 115060
rect 509954 79380 509986 79616
rect 510222 79380 510306 79616
rect 510542 79380 510574 79616
rect 509954 79296 510574 79380
rect 509954 79060 509986 79296
rect 510222 79060 510306 79296
rect 510542 79060 510574 79296
rect 509954 43616 510574 79060
rect 509954 43380 509986 43616
rect 510222 43380 510306 43616
rect 510542 43380 510574 43616
rect 509954 43296 510574 43380
rect 509954 43060 509986 43296
rect 510222 43060 510306 43296
rect 510542 43060 510574 43296
rect 509954 7616 510574 43060
rect 509954 7380 509986 7616
rect 510222 7380 510306 7616
rect 510542 7380 510574 7616
rect 509954 7296 510574 7380
rect 509954 7060 509986 7296
rect 510222 7060 510306 7296
rect 510542 7060 510574 7296
rect 509954 -4184 510574 7060
rect 509954 -4420 509986 -4184
rect 510222 -4420 510306 -4184
rect 510542 -4420 510574 -4184
rect 509954 -4504 510574 -4420
rect 509954 -4740 509986 -4504
rect 510222 -4740 510306 -4504
rect 510542 -4740 510574 -4504
rect 509954 -7652 510574 -4740
rect 511194 709640 511814 711592
rect 511194 709404 511226 709640
rect 511462 709404 511546 709640
rect 511782 709404 511814 709640
rect 511194 709320 511814 709404
rect 511194 709084 511226 709320
rect 511462 709084 511546 709320
rect 511782 709084 511814 709320
rect 511194 692856 511814 709084
rect 511194 692620 511226 692856
rect 511462 692620 511546 692856
rect 511782 692620 511814 692856
rect 511194 692536 511814 692620
rect 511194 692300 511226 692536
rect 511462 692300 511546 692536
rect 511782 692300 511814 692536
rect 511194 656856 511814 692300
rect 511194 656620 511226 656856
rect 511462 656620 511546 656856
rect 511782 656620 511814 656856
rect 511194 656536 511814 656620
rect 511194 656300 511226 656536
rect 511462 656300 511546 656536
rect 511782 656300 511814 656536
rect 511194 620856 511814 656300
rect 511194 620620 511226 620856
rect 511462 620620 511546 620856
rect 511782 620620 511814 620856
rect 511194 620536 511814 620620
rect 511194 620300 511226 620536
rect 511462 620300 511546 620536
rect 511782 620300 511814 620536
rect 511194 584856 511814 620300
rect 511194 584620 511226 584856
rect 511462 584620 511546 584856
rect 511782 584620 511814 584856
rect 511194 584536 511814 584620
rect 511194 584300 511226 584536
rect 511462 584300 511546 584536
rect 511782 584300 511814 584536
rect 511194 548856 511814 584300
rect 511194 548620 511226 548856
rect 511462 548620 511546 548856
rect 511782 548620 511814 548856
rect 511194 548536 511814 548620
rect 511194 548300 511226 548536
rect 511462 548300 511546 548536
rect 511782 548300 511814 548536
rect 511194 512856 511814 548300
rect 511194 512620 511226 512856
rect 511462 512620 511546 512856
rect 511782 512620 511814 512856
rect 511194 512536 511814 512620
rect 511194 512300 511226 512536
rect 511462 512300 511546 512536
rect 511782 512300 511814 512536
rect 511194 476856 511814 512300
rect 511194 476620 511226 476856
rect 511462 476620 511546 476856
rect 511782 476620 511814 476856
rect 511194 476536 511814 476620
rect 511194 476300 511226 476536
rect 511462 476300 511546 476536
rect 511782 476300 511814 476536
rect 511194 440856 511814 476300
rect 511194 440620 511226 440856
rect 511462 440620 511546 440856
rect 511782 440620 511814 440856
rect 511194 440536 511814 440620
rect 511194 440300 511226 440536
rect 511462 440300 511546 440536
rect 511782 440300 511814 440536
rect 511194 404856 511814 440300
rect 511194 404620 511226 404856
rect 511462 404620 511546 404856
rect 511782 404620 511814 404856
rect 511194 404536 511814 404620
rect 511194 404300 511226 404536
rect 511462 404300 511546 404536
rect 511782 404300 511814 404536
rect 511194 368856 511814 404300
rect 511194 368620 511226 368856
rect 511462 368620 511546 368856
rect 511782 368620 511814 368856
rect 511194 368536 511814 368620
rect 511194 368300 511226 368536
rect 511462 368300 511546 368536
rect 511782 368300 511814 368536
rect 511194 332856 511814 368300
rect 511194 332620 511226 332856
rect 511462 332620 511546 332856
rect 511782 332620 511814 332856
rect 511194 332536 511814 332620
rect 511194 332300 511226 332536
rect 511462 332300 511546 332536
rect 511782 332300 511814 332536
rect 511194 296856 511814 332300
rect 511194 296620 511226 296856
rect 511462 296620 511546 296856
rect 511782 296620 511814 296856
rect 511194 296536 511814 296620
rect 511194 296300 511226 296536
rect 511462 296300 511546 296536
rect 511782 296300 511814 296536
rect 511194 260856 511814 296300
rect 511194 260620 511226 260856
rect 511462 260620 511546 260856
rect 511782 260620 511814 260856
rect 511194 260536 511814 260620
rect 511194 260300 511226 260536
rect 511462 260300 511546 260536
rect 511782 260300 511814 260536
rect 511194 224856 511814 260300
rect 511194 224620 511226 224856
rect 511462 224620 511546 224856
rect 511782 224620 511814 224856
rect 511194 224536 511814 224620
rect 511194 224300 511226 224536
rect 511462 224300 511546 224536
rect 511782 224300 511814 224536
rect 511194 188856 511814 224300
rect 511194 188620 511226 188856
rect 511462 188620 511546 188856
rect 511782 188620 511814 188856
rect 511194 188536 511814 188620
rect 511194 188300 511226 188536
rect 511462 188300 511546 188536
rect 511782 188300 511814 188536
rect 511194 152856 511814 188300
rect 511194 152620 511226 152856
rect 511462 152620 511546 152856
rect 511782 152620 511814 152856
rect 511194 152536 511814 152620
rect 511194 152300 511226 152536
rect 511462 152300 511546 152536
rect 511782 152300 511814 152536
rect 511194 116856 511814 152300
rect 511194 116620 511226 116856
rect 511462 116620 511546 116856
rect 511782 116620 511814 116856
rect 511194 116536 511814 116620
rect 511194 116300 511226 116536
rect 511462 116300 511546 116536
rect 511782 116300 511814 116536
rect 511194 80856 511814 116300
rect 511194 80620 511226 80856
rect 511462 80620 511546 80856
rect 511782 80620 511814 80856
rect 511194 80536 511814 80620
rect 511194 80300 511226 80536
rect 511462 80300 511546 80536
rect 511782 80300 511814 80536
rect 511194 44856 511814 80300
rect 511194 44620 511226 44856
rect 511462 44620 511546 44856
rect 511782 44620 511814 44856
rect 511194 44536 511814 44620
rect 511194 44300 511226 44536
rect 511462 44300 511546 44536
rect 511782 44300 511814 44536
rect 511194 8856 511814 44300
rect 511194 8620 511226 8856
rect 511462 8620 511546 8856
rect 511782 8620 511814 8856
rect 511194 8536 511814 8620
rect 511194 8300 511226 8536
rect 511462 8300 511546 8536
rect 511782 8300 511814 8536
rect 511194 -5144 511814 8300
rect 511194 -5380 511226 -5144
rect 511462 -5380 511546 -5144
rect 511782 -5380 511814 -5144
rect 511194 -5464 511814 -5380
rect 511194 -5700 511226 -5464
rect 511462 -5700 511546 -5464
rect 511782 -5700 511814 -5464
rect 511194 -7652 511814 -5700
rect 512434 710600 513054 711592
rect 512434 710364 512466 710600
rect 512702 710364 512786 710600
rect 513022 710364 513054 710600
rect 512434 710280 513054 710364
rect 512434 710044 512466 710280
rect 512702 710044 512786 710280
rect 513022 710044 513054 710280
rect 512434 694096 513054 710044
rect 512434 693860 512466 694096
rect 512702 693860 512786 694096
rect 513022 693860 513054 694096
rect 512434 693776 513054 693860
rect 512434 693540 512466 693776
rect 512702 693540 512786 693776
rect 513022 693540 513054 693776
rect 512434 658096 513054 693540
rect 512434 657860 512466 658096
rect 512702 657860 512786 658096
rect 513022 657860 513054 658096
rect 512434 657776 513054 657860
rect 512434 657540 512466 657776
rect 512702 657540 512786 657776
rect 513022 657540 513054 657776
rect 512434 622096 513054 657540
rect 512434 621860 512466 622096
rect 512702 621860 512786 622096
rect 513022 621860 513054 622096
rect 512434 621776 513054 621860
rect 512434 621540 512466 621776
rect 512702 621540 512786 621776
rect 513022 621540 513054 621776
rect 512434 586096 513054 621540
rect 512434 585860 512466 586096
rect 512702 585860 512786 586096
rect 513022 585860 513054 586096
rect 512434 585776 513054 585860
rect 512434 585540 512466 585776
rect 512702 585540 512786 585776
rect 513022 585540 513054 585776
rect 512434 550096 513054 585540
rect 512434 549860 512466 550096
rect 512702 549860 512786 550096
rect 513022 549860 513054 550096
rect 512434 549776 513054 549860
rect 512434 549540 512466 549776
rect 512702 549540 512786 549776
rect 513022 549540 513054 549776
rect 512434 514096 513054 549540
rect 512434 513860 512466 514096
rect 512702 513860 512786 514096
rect 513022 513860 513054 514096
rect 512434 513776 513054 513860
rect 512434 513540 512466 513776
rect 512702 513540 512786 513776
rect 513022 513540 513054 513776
rect 512434 478096 513054 513540
rect 512434 477860 512466 478096
rect 512702 477860 512786 478096
rect 513022 477860 513054 478096
rect 512434 477776 513054 477860
rect 512434 477540 512466 477776
rect 512702 477540 512786 477776
rect 513022 477540 513054 477776
rect 512434 442096 513054 477540
rect 512434 441860 512466 442096
rect 512702 441860 512786 442096
rect 513022 441860 513054 442096
rect 512434 441776 513054 441860
rect 512434 441540 512466 441776
rect 512702 441540 512786 441776
rect 513022 441540 513054 441776
rect 512434 406096 513054 441540
rect 512434 405860 512466 406096
rect 512702 405860 512786 406096
rect 513022 405860 513054 406096
rect 512434 405776 513054 405860
rect 512434 405540 512466 405776
rect 512702 405540 512786 405776
rect 513022 405540 513054 405776
rect 512434 370096 513054 405540
rect 512434 369860 512466 370096
rect 512702 369860 512786 370096
rect 513022 369860 513054 370096
rect 512434 369776 513054 369860
rect 512434 369540 512466 369776
rect 512702 369540 512786 369776
rect 513022 369540 513054 369776
rect 512434 334096 513054 369540
rect 512434 333860 512466 334096
rect 512702 333860 512786 334096
rect 513022 333860 513054 334096
rect 512434 333776 513054 333860
rect 512434 333540 512466 333776
rect 512702 333540 512786 333776
rect 513022 333540 513054 333776
rect 512434 298096 513054 333540
rect 512434 297860 512466 298096
rect 512702 297860 512786 298096
rect 513022 297860 513054 298096
rect 512434 297776 513054 297860
rect 512434 297540 512466 297776
rect 512702 297540 512786 297776
rect 513022 297540 513054 297776
rect 512434 262096 513054 297540
rect 512434 261860 512466 262096
rect 512702 261860 512786 262096
rect 513022 261860 513054 262096
rect 512434 261776 513054 261860
rect 512434 261540 512466 261776
rect 512702 261540 512786 261776
rect 513022 261540 513054 261776
rect 512434 226096 513054 261540
rect 512434 225860 512466 226096
rect 512702 225860 512786 226096
rect 513022 225860 513054 226096
rect 512434 225776 513054 225860
rect 512434 225540 512466 225776
rect 512702 225540 512786 225776
rect 513022 225540 513054 225776
rect 512434 190096 513054 225540
rect 512434 189860 512466 190096
rect 512702 189860 512786 190096
rect 513022 189860 513054 190096
rect 512434 189776 513054 189860
rect 512434 189540 512466 189776
rect 512702 189540 512786 189776
rect 513022 189540 513054 189776
rect 512434 154096 513054 189540
rect 512434 153860 512466 154096
rect 512702 153860 512786 154096
rect 513022 153860 513054 154096
rect 512434 153776 513054 153860
rect 512434 153540 512466 153776
rect 512702 153540 512786 153776
rect 513022 153540 513054 153776
rect 512434 118096 513054 153540
rect 512434 117860 512466 118096
rect 512702 117860 512786 118096
rect 513022 117860 513054 118096
rect 512434 117776 513054 117860
rect 512434 117540 512466 117776
rect 512702 117540 512786 117776
rect 513022 117540 513054 117776
rect 512434 82096 513054 117540
rect 512434 81860 512466 82096
rect 512702 81860 512786 82096
rect 513022 81860 513054 82096
rect 512434 81776 513054 81860
rect 512434 81540 512466 81776
rect 512702 81540 512786 81776
rect 513022 81540 513054 81776
rect 512434 46096 513054 81540
rect 512434 45860 512466 46096
rect 512702 45860 512786 46096
rect 513022 45860 513054 46096
rect 512434 45776 513054 45860
rect 512434 45540 512466 45776
rect 512702 45540 512786 45776
rect 513022 45540 513054 45776
rect 512434 10096 513054 45540
rect 512434 9860 512466 10096
rect 512702 9860 512786 10096
rect 513022 9860 513054 10096
rect 512434 9776 513054 9860
rect 512434 9540 512466 9776
rect 512702 9540 512786 9776
rect 513022 9540 513054 9776
rect 512434 -6104 513054 9540
rect 512434 -6340 512466 -6104
rect 512702 -6340 512786 -6104
rect 513022 -6340 513054 -6104
rect 512434 -6424 513054 -6340
rect 512434 -6660 512466 -6424
rect 512702 -6660 512786 -6424
rect 513022 -6660 513054 -6424
rect 512434 -7652 513054 -6660
rect 513674 711560 514294 711592
rect 513674 711324 513706 711560
rect 513942 711324 514026 711560
rect 514262 711324 514294 711560
rect 513674 711240 514294 711324
rect 513674 711004 513706 711240
rect 513942 711004 514026 711240
rect 514262 711004 514294 711240
rect 513674 695336 514294 711004
rect 513674 695100 513706 695336
rect 513942 695100 514026 695336
rect 514262 695100 514294 695336
rect 513674 695016 514294 695100
rect 513674 694780 513706 695016
rect 513942 694780 514026 695016
rect 514262 694780 514294 695016
rect 513674 659336 514294 694780
rect 513674 659100 513706 659336
rect 513942 659100 514026 659336
rect 514262 659100 514294 659336
rect 513674 659016 514294 659100
rect 513674 658780 513706 659016
rect 513942 658780 514026 659016
rect 514262 658780 514294 659016
rect 513674 623336 514294 658780
rect 513674 623100 513706 623336
rect 513942 623100 514026 623336
rect 514262 623100 514294 623336
rect 513674 623016 514294 623100
rect 513674 622780 513706 623016
rect 513942 622780 514026 623016
rect 514262 622780 514294 623016
rect 513674 587336 514294 622780
rect 513674 587100 513706 587336
rect 513942 587100 514026 587336
rect 514262 587100 514294 587336
rect 513674 587016 514294 587100
rect 513674 586780 513706 587016
rect 513942 586780 514026 587016
rect 514262 586780 514294 587016
rect 513674 551336 514294 586780
rect 513674 551100 513706 551336
rect 513942 551100 514026 551336
rect 514262 551100 514294 551336
rect 513674 551016 514294 551100
rect 513674 550780 513706 551016
rect 513942 550780 514026 551016
rect 514262 550780 514294 551016
rect 513674 515336 514294 550780
rect 513674 515100 513706 515336
rect 513942 515100 514026 515336
rect 514262 515100 514294 515336
rect 513674 515016 514294 515100
rect 513674 514780 513706 515016
rect 513942 514780 514026 515016
rect 514262 514780 514294 515016
rect 513674 479336 514294 514780
rect 513674 479100 513706 479336
rect 513942 479100 514026 479336
rect 514262 479100 514294 479336
rect 513674 479016 514294 479100
rect 513674 478780 513706 479016
rect 513942 478780 514026 479016
rect 514262 478780 514294 479016
rect 513674 443336 514294 478780
rect 540994 704840 541614 711592
rect 540994 704604 541026 704840
rect 541262 704604 541346 704840
rect 541582 704604 541614 704840
rect 540994 704520 541614 704604
rect 540994 704284 541026 704520
rect 541262 704284 541346 704520
rect 541582 704284 541614 704520
rect 540994 686656 541614 704284
rect 540994 686420 541026 686656
rect 541262 686420 541346 686656
rect 541582 686420 541614 686656
rect 540994 686336 541614 686420
rect 540994 686100 541026 686336
rect 541262 686100 541346 686336
rect 541582 686100 541614 686336
rect 540994 650656 541614 686100
rect 540994 650420 541026 650656
rect 541262 650420 541346 650656
rect 541582 650420 541614 650656
rect 540994 650336 541614 650420
rect 540994 650100 541026 650336
rect 541262 650100 541346 650336
rect 541582 650100 541614 650336
rect 540994 614656 541614 650100
rect 540994 614420 541026 614656
rect 541262 614420 541346 614656
rect 541582 614420 541614 614656
rect 540994 614336 541614 614420
rect 540994 614100 541026 614336
rect 541262 614100 541346 614336
rect 541582 614100 541614 614336
rect 540994 578656 541614 614100
rect 540994 578420 541026 578656
rect 541262 578420 541346 578656
rect 541582 578420 541614 578656
rect 540994 578336 541614 578420
rect 540994 578100 541026 578336
rect 541262 578100 541346 578336
rect 541582 578100 541614 578336
rect 540994 542656 541614 578100
rect 540994 542420 541026 542656
rect 541262 542420 541346 542656
rect 541582 542420 541614 542656
rect 540994 542336 541614 542420
rect 540994 542100 541026 542336
rect 541262 542100 541346 542336
rect 541582 542100 541614 542336
rect 540994 506656 541614 542100
rect 540994 506420 541026 506656
rect 541262 506420 541346 506656
rect 541582 506420 541614 506656
rect 540994 506336 541614 506420
rect 540994 506100 541026 506336
rect 541262 506100 541346 506336
rect 541582 506100 541614 506336
rect 540994 470656 541614 506100
rect 540994 470420 541026 470656
rect 541262 470420 541346 470656
rect 541582 470420 541614 470656
rect 540994 470336 541614 470420
rect 540994 470100 541026 470336
rect 541262 470100 541346 470336
rect 541582 470100 541614 470336
rect 540994 445574 541614 470100
rect 542234 705800 542854 711592
rect 542234 705564 542266 705800
rect 542502 705564 542586 705800
rect 542822 705564 542854 705800
rect 542234 705480 542854 705564
rect 542234 705244 542266 705480
rect 542502 705244 542586 705480
rect 542822 705244 542854 705480
rect 542234 687896 542854 705244
rect 542234 687660 542266 687896
rect 542502 687660 542586 687896
rect 542822 687660 542854 687896
rect 542234 687576 542854 687660
rect 542234 687340 542266 687576
rect 542502 687340 542586 687576
rect 542822 687340 542854 687576
rect 542234 651896 542854 687340
rect 542234 651660 542266 651896
rect 542502 651660 542586 651896
rect 542822 651660 542854 651896
rect 542234 651576 542854 651660
rect 542234 651340 542266 651576
rect 542502 651340 542586 651576
rect 542822 651340 542854 651576
rect 542234 615896 542854 651340
rect 542234 615660 542266 615896
rect 542502 615660 542586 615896
rect 542822 615660 542854 615896
rect 542234 615576 542854 615660
rect 542234 615340 542266 615576
rect 542502 615340 542586 615576
rect 542822 615340 542854 615576
rect 542234 579896 542854 615340
rect 542234 579660 542266 579896
rect 542502 579660 542586 579896
rect 542822 579660 542854 579896
rect 542234 579576 542854 579660
rect 542234 579340 542266 579576
rect 542502 579340 542586 579576
rect 542822 579340 542854 579576
rect 542234 543896 542854 579340
rect 542234 543660 542266 543896
rect 542502 543660 542586 543896
rect 542822 543660 542854 543896
rect 542234 543576 542854 543660
rect 542234 543340 542266 543576
rect 542502 543340 542586 543576
rect 542822 543340 542854 543576
rect 542234 507896 542854 543340
rect 542234 507660 542266 507896
rect 542502 507660 542586 507896
rect 542822 507660 542854 507896
rect 542234 507576 542854 507660
rect 542234 507340 542266 507576
rect 542502 507340 542586 507576
rect 542822 507340 542854 507576
rect 542234 471896 542854 507340
rect 542234 471660 542266 471896
rect 542502 471660 542586 471896
rect 542822 471660 542854 471896
rect 542234 471576 542854 471660
rect 542234 471340 542266 471576
rect 542502 471340 542586 471576
rect 542822 471340 542854 471576
rect 542234 445574 542854 471340
rect 543474 706760 544094 711592
rect 543474 706524 543506 706760
rect 543742 706524 543826 706760
rect 544062 706524 544094 706760
rect 543474 706440 544094 706524
rect 543474 706204 543506 706440
rect 543742 706204 543826 706440
rect 544062 706204 544094 706440
rect 543474 689136 544094 706204
rect 543474 688900 543506 689136
rect 543742 688900 543826 689136
rect 544062 688900 544094 689136
rect 543474 688816 544094 688900
rect 543474 688580 543506 688816
rect 543742 688580 543826 688816
rect 544062 688580 544094 688816
rect 543474 653136 544094 688580
rect 543474 652900 543506 653136
rect 543742 652900 543826 653136
rect 544062 652900 544094 653136
rect 543474 652816 544094 652900
rect 543474 652580 543506 652816
rect 543742 652580 543826 652816
rect 544062 652580 544094 652816
rect 543474 617136 544094 652580
rect 543474 616900 543506 617136
rect 543742 616900 543826 617136
rect 544062 616900 544094 617136
rect 543474 616816 544094 616900
rect 543474 616580 543506 616816
rect 543742 616580 543826 616816
rect 544062 616580 544094 616816
rect 543474 581136 544094 616580
rect 543474 580900 543506 581136
rect 543742 580900 543826 581136
rect 544062 580900 544094 581136
rect 543474 580816 544094 580900
rect 543474 580580 543506 580816
rect 543742 580580 543826 580816
rect 544062 580580 544094 580816
rect 543474 545136 544094 580580
rect 543474 544900 543506 545136
rect 543742 544900 543826 545136
rect 544062 544900 544094 545136
rect 543474 544816 544094 544900
rect 543474 544580 543506 544816
rect 543742 544580 543826 544816
rect 544062 544580 544094 544816
rect 543474 509136 544094 544580
rect 543474 508900 543506 509136
rect 543742 508900 543826 509136
rect 544062 508900 544094 509136
rect 543474 508816 544094 508900
rect 543474 508580 543506 508816
rect 543742 508580 543826 508816
rect 544062 508580 544094 508816
rect 543474 473136 544094 508580
rect 543474 472900 543506 473136
rect 543742 472900 543826 473136
rect 544062 472900 544094 473136
rect 543474 472816 544094 472900
rect 543474 472580 543506 472816
rect 543742 472580 543826 472816
rect 544062 472580 544094 472816
rect 543474 445574 544094 472580
rect 544714 707720 545334 711592
rect 544714 707484 544746 707720
rect 544982 707484 545066 707720
rect 545302 707484 545334 707720
rect 544714 707400 545334 707484
rect 544714 707164 544746 707400
rect 544982 707164 545066 707400
rect 545302 707164 545334 707400
rect 544714 690376 545334 707164
rect 544714 690140 544746 690376
rect 544982 690140 545066 690376
rect 545302 690140 545334 690376
rect 544714 690056 545334 690140
rect 544714 689820 544746 690056
rect 544982 689820 545066 690056
rect 545302 689820 545334 690056
rect 544714 654376 545334 689820
rect 544714 654140 544746 654376
rect 544982 654140 545066 654376
rect 545302 654140 545334 654376
rect 544714 654056 545334 654140
rect 544714 653820 544746 654056
rect 544982 653820 545066 654056
rect 545302 653820 545334 654056
rect 544714 618376 545334 653820
rect 544714 618140 544746 618376
rect 544982 618140 545066 618376
rect 545302 618140 545334 618376
rect 544714 618056 545334 618140
rect 544714 617820 544746 618056
rect 544982 617820 545066 618056
rect 545302 617820 545334 618056
rect 544714 582376 545334 617820
rect 544714 582140 544746 582376
rect 544982 582140 545066 582376
rect 545302 582140 545334 582376
rect 544714 582056 545334 582140
rect 544714 581820 544746 582056
rect 544982 581820 545066 582056
rect 545302 581820 545334 582056
rect 544714 546376 545334 581820
rect 544714 546140 544746 546376
rect 544982 546140 545066 546376
rect 545302 546140 545334 546376
rect 544714 546056 545334 546140
rect 544714 545820 544746 546056
rect 544982 545820 545066 546056
rect 545302 545820 545334 546056
rect 544714 510376 545334 545820
rect 544714 510140 544746 510376
rect 544982 510140 545066 510376
rect 545302 510140 545334 510376
rect 544714 510056 545334 510140
rect 544714 509820 544746 510056
rect 544982 509820 545066 510056
rect 545302 509820 545334 510056
rect 544714 474376 545334 509820
rect 544714 474140 544746 474376
rect 544982 474140 545066 474376
rect 545302 474140 545334 474376
rect 544714 474056 545334 474140
rect 544714 473820 544746 474056
rect 544982 473820 545066 474056
rect 545302 473820 545334 474056
rect 544331 445774 544397 445775
rect 544331 445710 544332 445774
rect 544396 445710 544397 445774
rect 544331 445709 544397 445710
rect 541571 445366 541637 445367
rect 541571 445302 541572 445366
rect 541636 445302 541637 445366
rect 541571 445301 541637 445302
rect 513674 443100 513706 443336
rect 513942 443100 514026 443336
rect 514262 443100 514294 443336
rect 513674 443016 514294 443100
rect 513674 442780 513706 443016
rect 513942 442780 514026 443016
rect 514262 442780 514294 443016
rect 513674 407336 514294 442780
rect 540876 435896 541196 435928
rect 540876 435660 540918 435896
rect 541154 435660 541196 435896
rect 540876 435576 541196 435660
rect 540876 435340 540918 435576
rect 541154 435340 541196 435576
rect 540876 435308 541196 435340
rect 539910 434656 540230 434688
rect 539910 434420 539952 434656
rect 540188 434420 540230 434656
rect 539910 434336 540230 434420
rect 539910 434100 539952 434336
rect 540188 434100 540230 434336
rect 539910 434068 540230 434100
rect 541574 409327 541634 445301
rect 542808 435896 543128 435928
rect 542808 435660 542850 435896
rect 543086 435660 543128 435896
rect 542808 435576 543128 435660
rect 542808 435340 542850 435576
rect 543086 435340 543128 435576
rect 542808 435308 543128 435340
rect 541842 434656 542162 434688
rect 541842 434420 541884 434656
rect 542120 434420 542162 434656
rect 541842 434336 542162 434420
rect 541842 434100 541884 434336
rect 542120 434100 542162 434336
rect 541842 434068 542162 434100
rect 543774 434656 544094 434688
rect 543774 434420 543816 434656
rect 544052 434420 544094 434656
rect 543774 434336 544094 434420
rect 543774 434100 543816 434336
rect 544052 434100 544094 434336
rect 543774 434068 544094 434100
rect 544334 409327 544394 445709
rect 544714 445574 545334 473820
rect 545954 708680 546574 711592
rect 545954 708444 545986 708680
rect 546222 708444 546306 708680
rect 546542 708444 546574 708680
rect 545954 708360 546574 708444
rect 545954 708124 545986 708360
rect 546222 708124 546306 708360
rect 546542 708124 546574 708360
rect 545954 691616 546574 708124
rect 545954 691380 545986 691616
rect 546222 691380 546306 691616
rect 546542 691380 546574 691616
rect 545954 691296 546574 691380
rect 545954 691060 545986 691296
rect 546222 691060 546306 691296
rect 546542 691060 546574 691296
rect 545954 655616 546574 691060
rect 545954 655380 545986 655616
rect 546222 655380 546306 655616
rect 546542 655380 546574 655616
rect 545954 655296 546574 655380
rect 545954 655060 545986 655296
rect 546222 655060 546306 655296
rect 546542 655060 546574 655296
rect 545954 619616 546574 655060
rect 545954 619380 545986 619616
rect 546222 619380 546306 619616
rect 546542 619380 546574 619616
rect 545954 619296 546574 619380
rect 545954 619060 545986 619296
rect 546222 619060 546306 619296
rect 546542 619060 546574 619296
rect 545954 583616 546574 619060
rect 545954 583380 545986 583616
rect 546222 583380 546306 583616
rect 546542 583380 546574 583616
rect 545954 583296 546574 583380
rect 545954 583060 545986 583296
rect 546222 583060 546306 583296
rect 546542 583060 546574 583296
rect 545954 547616 546574 583060
rect 545954 547380 545986 547616
rect 546222 547380 546306 547616
rect 546542 547380 546574 547616
rect 545954 547296 546574 547380
rect 545954 547060 545986 547296
rect 546222 547060 546306 547296
rect 546542 547060 546574 547296
rect 545954 511616 546574 547060
rect 545954 511380 545986 511616
rect 546222 511380 546306 511616
rect 546542 511380 546574 511616
rect 545954 511296 546574 511380
rect 545954 511060 545986 511296
rect 546222 511060 546306 511296
rect 546542 511060 546574 511296
rect 545954 475616 546574 511060
rect 545954 475380 545986 475616
rect 546222 475380 546306 475616
rect 546542 475380 546574 475616
rect 545954 475296 546574 475380
rect 545954 475060 545986 475296
rect 546222 475060 546306 475296
rect 546542 475060 546574 475296
rect 545954 445574 546574 475060
rect 547194 709640 547814 711592
rect 547194 709404 547226 709640
rect 547462 709404 547546 709640
rect 547782 709404 547814 709640
rect 547194 709320 547814 709404
rect 547194 709084 547226 709320
rect 547462 709084 547546 709320
rect 547782 709084 547814 709320
rect 547194 692856 547814 709084
rect 547194 692620 547226 692856
rect 547462 692620 547546 692856
rect 547782 692620 547814 692856
rect 547194 692536 547814 692620
rect 547194 692300 547226 692536
rect 547462 692300 547546 692536
rect 547782 692300 547814 692536
rect 547194 656856 547814 692300
rect 547194 656620 547226 656856
rect 547462 656620 547546 656856
rect 547782 656620 547814 656856
rect 547194 656536 547814 656620
rect 547194 656300 547226 656536
rect 547462 656300 547546 656536
rect 547782 656300 547814 656536
rect 547194 620856 547814 656300
rect 547194 620620 547226 620856
rect 547462 620620 547546 620856
rect 547782 620620 547814 620856
rect 547194 620536 547814 620620
rect 547194 620300 547226 620536
rect 547462 620300 547546 620536
rect 547782 620300 547814 620536
rect 547194 584856 547814 620300
rect 547194 584620 547226 584856
rect 547462 584620 547546 584856
rect 547782 584620 547814 584856
rect 547194 584536 547814 584620
rect 547194 584300 547226 584536
rect 547462 584300 547546 584536
rect 547782 584300 547814 584536
rect 547194 548856 547814 584300
rect 547194 548620 547226 548856
rect 547462 548620 547546 548856
rect 547782 548620 547814 548856
rect 547194 548536 547814 548620
rect 547194 548300 547226 548536
rect 547462 548300 547546 548536
rect 547782 548300 547814 548536
rect 547194 512856 547814 548300
rect 547194 512620 547226 512856
rect 547462 512620 547546 512856
rect 547782 512620 547814 512856
rect 547194 512536 547814 512620
rect 547194 512300 547226 512536
rect 547462 512300 547546 512536
rect 547782 512300 547814 512536
rect 547194 476856 547814 512300
rect 547194 476620 547226 476856
rect 547462 476620 547546 476856
rect 547782 476620 547814 476856
rect 547194 476536 547814 476620
rect 547194 476300 547226 476536
rect 547462 476300 547546 476536
rect 547782 476300 547814 476536
rect 547194 440856 547814 476300
rect 547194 440620 547226 440856
rect 547462 440620 547546 440856
rect 547782 440620 547814 440856
rect 547194 440536 547814 440620
rect 547194 440300 547226 440536
rect 547462 440300 547546 440536
rect 547782 440300 547814 440536
rect 544740 435896 545060 435928
rect 544740 435660 544782 435896
rect 545018 435660 545060 435896
rect 544740 435576 545060 435660
rect 544740 435340 544782 435576
rect 545018 435340 545060 435576
rect 544740 435308 545060 435340
rect 546672 435896 546992 435928
rect 546672 435660 546714 435896
rect 546950 435660 546992 435896
rect 546672 435576 546992 435660
rect 546672 435340 546714 435576
rect 546950 435340 546992 435576
rect 546672 435308 546992 435340
rect 545706 434656 546026 434688
rect 545706 434420 545748 434656
rect 545984 434420 546026 434656
rect 545706 434336 546026 434420
rect 545706 434100 545748 434336
rect 545984 434100 546026 434336
rect 545706 434068 546026 434100
rect 541571 409326 541637 409327
rect 541571 409262 541572 409326
rect 541636 409262 541637 409326
rect 541571 409261 541637 409262
rect 544331 409326 544397 409327
rect 544331 409262 544332 409326
rect 544396 409262 544397 409326
rect 544331 409261 544397 409262
rect 513674 407100 513706 407336
rect 513942 407100 514026 407336
rect 514262 407100 514294 407336
rect 513674 407016 514294 407100
rect 513674 406780 513706 407016
rect 513942 406780 514026 407016
rect 514262 406780 514294 407016
rect 513674 371336 514294 406780
rect 540876 399896 541196 399928
rect 540876 399660 540918 399896
rect 541154 399660 541196 399896
rect 540876 399576 541196 399660
rect 540876 399340 540918 399576
rect 541154 399340 541196 399576
rect 540876 399308 541196 399340
rect 539910 398656 540230 398688
rect 539910 398420 539952 398656
rect 540188 398420 540230 398656
rect 539910 398336 540230 398420
rect 539910 398100 539952 398336
rect 540188 398100 540230 398336
rect 539910 398068 540230 398100
rect 541574 373151 541634 409261
rect 542808 399896 543128 399928
rect 542808 399660 542850 399896
rect 543086 399660 543128 399896
rect 542808 399576 543128 399660
rect 542808 399340 542850 399576
rect 543086 399340 543128 399576
rect 542808 399308 543128 399340
rect 541842 398656 542162 398688
rect 541842 398420 541884 398656
rect 542120 398420 542162 398656
rect 541842 398336 542162 398420
rect 541842 398100 541884 398336
rect 542120 398100 542162 398336
rect 541842 398068 542162 398100
rect 543774 398656 544094 398688
rect 543774 398420 543816 398656
rect 544052 398420 544094 398656
rect 543774 398336 544094 398420
rect 543774 398100 543816 398336
rect 544052 398100 544094 398336
rect 543774 398068 544094 398100
rect 544334 373151 544394 409261
rect 547194 404856 547814 440300
rect 547194 404620 547226 404856
rect 547462 404620 547546 404856
rect 547782 404620 547814 404856
rect 547194 404536 547814 404620
rect 547194 404300 547226 404536
rect 547462 404300 547546 404536
rect 547782 404300 547814 404536
rect 544740 399896 545060 399928
rect 544740 399660 544782 399896
rect 545018 399660 545060 399896
rect 544740 399576 545060 399660
rect 544740 399340 544782 399576
rect 545018 399340 545060 399576
rect 544740 399308 545060 399340
rect 546672 399896 546992 399928
rect 546672 399660 546714 399896
rect 546950 399660 546992 399896
rect 546672 399576 546992 399660
rect 546672 399340 546714 399576
rect 546950 399340 546992 399576
rect 546672 399308 546992 399340
rect 545706 398656 546026 398688
rect 545706 398420 545748 398656
rect 545984 398420 546026 398656
rect 545706 398336 546026 398420
rect 545706 398100 545748 398336
rect 545984 398100 546026 398336
rect 545706 398068 546026 398100
rect 541571 373150 541637 373151
rect 541571 373086 541572 373150
rect 541636 373086 541637 373150
rect 541571 373085 541637 373086
rect 544331 373150 544397 373151
rect 544331 373086 544332 373150
rect 544396 373086 544397 373150
rect 544331 373085 544397 373086
rect 513674 371100 513706 371336
rect 513942 371100 514026 371336
rect 514262 371100 514294 371336
rect 513674 371016 514294 371100
rect 513674 370780 513706 371016
rect 513942 370780 514026 371016
rect 514262 370780 514294 371016
rect 513674 335336 514294 370780
rect 540876 363896 541196 363928
rect 540876 363660 540918 363896
rect 541154 363660 541196 363896
rect 540876 363576 541196 363660
rect 540876 363340 540918 363576
rect 541154 363340 541196 363576
rect 540876 363308 541196 363340
rect 539910 362656 540230 362688
rect 539910 362420 539952 362656
rect 540188 362420 540230 362656
rect 539910 362336 540230 362420
rect 539910 362100 539952 362336
rect 540188 362100 540230 362336
rect 539910 362068 540230 362100
rect 541574 339559 541634 373085
rect 542808 363896 543128 363928
rect 542808 363660 542850 363896
rect 543086 363660 543128 363896
rect 542808 363576 543128 363660
rect 542808 363340 542850 363576
rect 543086 363340 543128 363576
rect 542808 363308 543128 363340
rect 541842 362656 542162 362688
rect 541842 362420 541884 362656
rect 542120 362420 542162 362656
rect 541842 362336 542162 362420
rect 541842 362100 541884 362336
rect 542120 362100 542162 362336
rect 541842 362068 542162 362100
rect 543774 362656 544094 362688
rect 543774 362420 543816 362656
rect 544052 362420 544094 362656
rect 543774 362336 544094 362420
rect 543774 362100 543816 362336
rect 544052 362100 544094 362336
rect 543774 362068 544094 362100
rect 544334 339559 544394 373085
rect 547194 368856 547814 404300
rect 547194 368620 547226 368856
rect 547462 368620 547546 368856
rect 547782 368620 547814 368856
rect 547194 368536 547814 368620
rect 547194 368300 547226 368536
rect 547462 368300 547546 368536
rect 547782 368300 547814 368536
rect 544740 363896 545060 363928
rect 544740 363660 544782 363896
rect 545018 363660 545060 363896
rect 544740 363576 545060 363660
rect 544740 363340 544782 363576
rect 545018 363340 545060 363576
rect 544740 363308 545060 363340
rect 546672 363896 546992 363928
rect 546672 363660 546714 363896
rect 546950 363660 546992 363896
rect 546672 363576 546992 363660
rect 546672 363340 546714 363576
rect 546950 363340 546992 363576
rect 546672 363308 546992 363340
rect 545706 362656 546026 362688
rect 545706 362420 545748 362656
rect 545984 362420 546026 362656
rect 545706 362336 546026 362420
rect 545706 362100 545748 362336
rect 545984 362100 546026 362336
rect 545706 362068 546026 362100
rect 541571 339558 541637 339559
rect 541571 339494 541572 339558
rect 541636 339494 541637 339558
rect 541571 339493 541637 339494
rect 544331 339558 544397 339559
rect 544331 339494 544332 339558
rect 544396 339494 544397 339558
rect 544331 339493 544397 339494
rect 513674 335100 513706 335336
rect 513942 335100 514026 335336
rect 514262 335100 514294 335336
rect 513674 335016 514294 335100
rect 513674 334780 513706 335016
rect 513942 334780 514026 335016
rect 514262 334780 514294 335016
rect 513674 299336 514294 334780
rect 540876 327896 541196 327928
rect 540876 327660 540918 327896
rect 541154 327660 541196 327896
rect 540876 327576 541196 327660
rect 540876 327340 540918 327576
rect 541154 327340 541196 327576
rect 540876 327308 541196 327340
rect 539910 326656 540230 326688
rect 539910 326420 539952 326656
rect 540188 326420 540230 326656
rect 539910 326336 540230 326420
rect 539910 326100 539952 326336
rect 540188 326100 540230 326336
rect 539910 326068 540230 326100
rect 541574 303791 541634 339493
rect 542808 327896 543128 327928
rect 542808 327660 542850 327896
rect 543086 327660 543128 327896
rect 542808 327576 543128 327660
rect 542808 327340 542850 327576
rect 543086 327340 543128 327576
rect 542808 327308 543128 327340
rect 541842 326656 542162 326688
rect 541842 326420 541884 326656
rect 542120 326420 542162 326656
rect 541842 326336 542162 326420
rect 541842 326100 541884 326336
rect 542120 326100 542162 326336
rect 541842 326068 542162 326100
rect 543774 326656 544094 326688
rect 543774 326420 543816 326656
rect 544052 326420 544094 326656
rect 543774 326336 544094 326420
rect 543774 326100 543816 326336
rect 544052 326100 544094 326336
rect 543774 326068 544094 326100
rect 544334 303791 544394 339493
rect 547194 332856 547814 368300
rect 547194 332620 547226 332856
rect 547462 332620 547546 332856
rect 547782 332620 547814 332856
rect 547194 332536 547814 332620
rect 547194 332300 547226 332536
rect 547462 332300 547546 332536
rect 547782 332300 547814 332536
rect 544740 327896 545060 327928
rect 544740 327660 544782 327896
rect 545018 327660 545060 327896
rect 544740 327576 545060 327660
rect 544740 327340 544782 327576
rect 545018 327340 545060 327576
rect 544740 327308 545060 327340
rect 546672 327896 546992 327928
rect 546672 327660 546714 327896
rect 546950 327660 546992 327896
rect 546672 327576 546992 327660
rect 546672 327340 546714 327576
rect 546950 327340 546992 327576
rect 546672 327308 546992 327340
rect 545706 326656 546026 326688
rect 545706 326420 545748 326656
rect 545984 326420 546026 326656
rect 545706 326336 546026 326420
rect 545706 326100 545748 326336
rect 545984 326100 546026 326336
rect 545706 326068 546026 326100
rect 541571 303790 541637 303791
rect 541571 303726 541572 303790
rect 541636 303726 541637 303790
rect 541571 303725 541637 303726
rect 544331 303790 544397 303791
rect 544331 303726 544332 303790
rect 544396 303726 544397 303790
rect 544331 303725 544397 303726
rect 513674 299100 513706 299336
rect 513942 299100 514026 299336
rect 514262 299100 514294 299336
rect 513674 299016 514294 299100
rect 513674 298780 513706 299016
rect 513942 298780 514026 299016
rect 514262 298780 514294 299016
rect 513674 263336 514294 298780
rect 547194 296856 547814 332300
rect 547194 296620 547226 296856
rect 547462 296620 547546 296856
rect 547782 296620 547814 296856
rect 547194 296536 547814 296620
rect 547194 296300 547226 296536
rect 547462 296300 547546 296536
rect 547782 296300 547814 296536
rect 540876 291896 541196 291928
rect 540876 291660 540918 291896
rect 541154 291660 541196 291896
rect 540876 291576 541196 291660
rect 540876 291340 540918 291576
rect 541154 291340 541196 291576
rect 540876 291308 541196 291340
rect 542808 291896 543128 291928
rect 542808 291660 542850 291896
rect 543086 291660 543128 291896
rect 542808 291576 543128 291660
rect 542808 291340 542850 291576
rect 543086 291340 543128 291576
rect 542808 291308 543128 291340
rect 544740 291896 545060 291928
rect 544740 291660 544782 291896
rect 545018 291660 545060 291896
rect 544740 291576 545060 291660
rect 544740 291340 544782 291576
rect 545018 291340 545060 291576
rect 544740 291308 545060 291340
rect 546672 291896 546992 291928
rect 546672 291660 546714 291896
rect 546950 291660 546992 291896
rect 546672 291576 546992 291660
rect 546672 291340 546714 291576
rect 546950 291340 546992 291576
rect 546672 291308 546992 291340
rect 539910 290656 540230 290688
rect 539910 290420 539952 290656
rect 540188 290420 540230 290656
rect 539910 290336 540230 290420
rect 539910 290100 539952 290336
rect 540188 290100 540230 290336
rect 539910 290068 540230 290100
rect 541842 290656 542162 290688
rect 541842 290420 541884 290656
rect 542120 290420 542162 290656
rect 541842 290336 542162 290420
rect 541842 290100 541884 290336
rect 542120 290100 542162 290336
rect 541842 290068 542162 290100
rect 543774 290656 544094 290688
rect 543774 290420 543816 290656
rect 544052 290420 544094 290656
rect 543774 290336 544094 290420
rect 543774 290100 543816 290336
rect 544052 290100 544094 290336
rect 543774 290068 544094 290100
rect 545706 290656 546026 290688
rect 545706 290420 545748 290656
rect 545984 290420 546026 290656
rect 545706 290336 546026 290420
rect 545706 290100 545748 290336
rect 545984 290100 546026 290336
rect 545706 290068 546026 290100
rect 513674 263100 513706 263336
rect 513942 263100 514026 263336
rect 514262 263100 514294 263336
rect 513674 263016 514294 263100
rect 513674 262780 513706 263016
rect 513942 262780 514026 263016
rect 514262 262780 514294 263016
rect 513674 227336 514294 262780
rect 513674 227100 513706 227336
rect 513942 227100 514026 227336
rect 514262 227100 514294 227336
rect 513674 227016 514294 227100
rect 513674 226780 513706 227016
rect 513942 226780 514026 227016
rect 514262 226780 514294 227016
rect 513674 191336 514294 226780
rect 513674 191100 513706 191336
rect 513942 191100 514026 191336
rect 514262 191100 514294 191336
rect 513674 191016 514294 191100
rect 513674 190780 513706 191016
rect 513942 190780 514026 191016
rect 514262 190780 514294 191016
rect 513674 155336 514294 190780
rect 513674 155100 513706 155336
rect 513942 155100 514026 155336
rect 514262 155100 514294 155336
rect 513674 155016 514294 155100
rect 513674 154780 513706 155016
rect 513942 154780 514026 155016
rect 514262 154780 514294 155016
rect 513674 119336 514294 154780
rect 513674 119100 513706 119336
rect 513942 119100 514026 119336
rect 514262 119100 514294 119336
rect 513674 119016 514294 119100
rect 513674 118780 513706 119016
rect 513942 118780 514026 119016
rect 514262 118780 514294 119016
rect 513674 83336 514294 118780
rect 513674 83100 513706 83336
rect 513942 83100 514026 83336
rect 514262 83100 514294 83336
rect 513674 83016 514294 83100
rect 513674 82780 513706 83016
rect 513942 82780 514026 83016
rect 514262 82780 514294 83016
rect 513674 47336 514294 82780
rect 513674 47100 513706 47336
rect 513942 47100 514026 47336
rect 514262 47100 514294 47336
rect 513674 47016 514294 47100
rect 513674 46780 513706 47016
rect 513942 46780 514026 47016
rect 514262 46780 514294 47016
rect 513674 11336 514294 46780
rect 513674 11100 513706 11336
rect 513942 11100 514026 11336
rect 514262 11100 514294 11336
rect 513674 11016 514294 11100
rect 513674 10780 513706 11016
rect 513942 10780 514026 11016
rect 514262 10780 514294 11016
rect 513674 -7064 514294 10780
rect 513674 -7300 513706 -7064
rect 513942 -7300 514026 -7064
rect 514262 -7300 514294 -7064
rect 513674 -7384 514294 -7300
rect 513674 -7620 513706 -7384
rect 513942 -7620 514026 -7384
rect 514262 -7620 514294 -7384
rect 513674 -7652 514294 -7620
rect 540994 254656 541614 279790
rect 540994 254420 541026 254656
rect 541262 254420 541346 254656
rect 541582 254420 541614 254656
rect 540994 254336 541614 254420
rect 540994 254100 541026 254336
rect 541262 254100 541346 254336
rect 541582 254100 541614 254336
rect 540994 218656 541614 254100
rect 540994 218420 541026 218656
rect 541262 218420 541346 218656
rect 541582 218420 541614 218656
rect 540994 218336 541614 218420
rect 540994 218100 541026 218336
rect 541262 218100 541346 218336
rect 541582 218100 541614 218336
rect 540994 182656 541614 218100
rect 540994 182420 541026 182656
rect 541262 182420 541346 182656
rect 541582 182420 541614 182656
rect 540994 182336 541614 182420
rect 540994 182100 541026 182336
rect 541262 182100 541346 182336
rect 541582 182100 541614 182336
rect 540994 146656 541614 182100
rect 540994 146420 541026 146656
rect 541262 146420 541346 146656
rect 541582 146420 541614 146656
rect 540994 146336 541614 146420
rect 540994 146100 541026 146336
rect 541262 146100 541346 146336
rect 541582 146100 541614 146336
rect 540994 110656 541614 146100
rect 540994 110420 541026 110656
rect 541262 110420 541346 110656
rect 541582 110420 541614 110656
rect 540994 110336 541614 110420
rect 540994 110100 541026 110336
rect 541262 110100 541346 110336
rect 541582 110100 541614 110336
rect 540994 74656 541614 110100
rect 540994 74420 541026 74656
rect 541262 74420 541346 74656
rect 541582 74420 541614 74656
rect 540994 74336 541614 74420
rect 540994 74100 541026 74336
rect 541262 74100 541346 74336
rect 541582 74100 541614 74336
rect 540994 38656 541614 74100
rect 540994 38420 541026 38656
rect 541262 38420 541346 38656
rect 541582 38420 541614 38656
rect 540994 38336 541614 38420
rect 540994 38100 541026 38336
rect 541262 38100 541346 38336
rect 541582 38100 541614 38336
rect 540994 2656 541614 38100
rect 540994 2420 541026 2656
rect 541262 2420 541346 2656
rect 541582 2420 541614 2656
rect 540994 2336 541614 2420
rect 540994 2100 541026 2336
rect 541262 2100 541346 2336
rect 541582 2100 541614 2336
rect 540994 -344 541614 2100
rect 540994 -580 541026 -344
rect 541262 -580 541346 -344
rect 541582 -580 541614 -344
rect 540994 -664 541614 -580
rect 540994 -900 541026 -664
rect 541262 -900 541346 -664
rect 541582 -900 541614 -664
rect 540994 -7652 541614 -900
rect 542234 255896 542854 279790
rect 542234 255660 542266 255896
rect 542502 255660 542586 255896
rect 542822 255660 542854 255896
rect 542234 255576 542854 255660
rect 542234 255340 542266 255576
rect 542502 255340 542586 255576
rect 542822 255340 542854 255576
rect 542234 219896 542854 255340
rect 542234 219660 542266 219896
rect 542502 219660 542586 219896
rect 542822 219660 542854 219896
rect 542234 219576 542854 219660
rect 542234 219340 542266 219576
rect 542502 219340 542586 219576
rect 542822 219340 542854 219576
rect 542234 183896 542854 219340
rect 542234 183660 542266 183896
rect 542502 183660 542586 183896
rect 542822 183660 542854 183896
rect 542234 183576 542854 183660
rect 542234 183340 542266 183576
rect 542502 183340 542586 183576
rect 542822 183340 542854 183576
rect 542234 147896 542854 183340
rect 542234 147660 542266 147896
rect 542502 147660 542586 147896
rect 542822 147660 542854 147896
rect 542234 147576 542854 147660
rect 542234 147340 542266 147576
rect 542502 147340 542586 147576
rect 542822 147340 542854 147576
rect 542234 111896 542854 147340
rect 542234 111660 542266 111896
rect 542502 111660 542586 111896
rect 542822 111660 542854 111896
rect 542234 111576 542854 111660
rect 542234 111340 542266 111576
rect 542502 111340 542586 111576
rect 542822 111340 542854 111576
rect 542234 75896 542854 111340
rect 542234 75660 542266 75896
rect 542502 75660 542586 75896
rect 542822 75660 542854 75896
rect 542234 75576 542854 75660
rect 542234 75340 542266 75576
rect 542502 75340 542586 75576
rect 542822 75340 542854 75576
rect 542234 39896 542854 75340
rect 542234 39660 542266 39896
rect 542502 39660 542586 39896
rect 542822 39660 542854 39896
rect 542234 39576 542854 39660
rect 542234 39340 542266 39576
rect 542502 39340 542586 39576
rect 542822 39340 542854 39576
rect 542234 3896 542854 39340
rect 542234 3660 542266 3896
rect 542502 3660 542586 3896
rect 542822 3660 542854 3896
rect 542234 3576 542854 3660
rect 542234 3340 542266 3576
rect 542502 3340 542586 3576
rect 542822 3340 542854 3576
rect 542234 -1304 542854 3340
rect 542234 -1540 542266 -1304
rect 542502 -1540 542586 -1304
rect 542822 -1540 542854 -1304
rect 542234 -1624 542854 -1540
rect 542234 -1860 542266 -1624
rect 542502 -1860 542586 -1624
rect 542822 -1860 542854 -1624
rect 542234 -7652 542854 -1860
rect 543474 257136 544094 279790
rect 543474 256900 543506 257136
rect 543742 256900 543826 257136
rect 544062 256900 544094 257136
rect 543474 256816 544094 256900
rect 543474 256580 543506 256816
rect 543742 256580 543826 256816
rect 544062 256580 544094 256816
rect 543474 221136 544094 256580
rect 543474 220900 543506 221136
rect 543742 220900 543826 221136
rect 544062 220900 544094 221136
rect 543474 220816 544094 220900
rect 543474 220580 543506 220816
rect 543742 220580 543826 220816
rect 544062 220580 544094 220816
rect 543474 185136 544094 220580
rect 543474 184900 543506 185136
rect 543742 184900 543826 185136
rect 544062 184900 544094 185136
rect 543474 184816 544094 184900
rect 543474 184580 543506 184816
rect 543742 184580 543826 184816
rect 544062 184580 544094 184816
rect 543474 149136 544094 184580
rect 543474 148900 543506 149136
rect 543742 148900 543826 149136
rect 544062 148900 544094 149136
rect 543474 148816 544094 148900
rect 543474 148580 543506 148816
rect 543742 148580 543826 148816
rect 544062 148580 544094 148816
rect 543474 113136 544094 148580
rect 543474 112900 543506 113136
rect 543742 112900 543826 113136
rect 544062 112900 544094 113136
rect 543474 112816 544094 112900
rect 543474 112580 543506 112816
rect 543742 112580 543826 112816
rect 544062 112580 544094 112816
rect 543474 77136 544094 112580
rect 543474 76900 543506 77136
rect 543742 76900 543826 77136
rect 544062 76900 544094 77136
rect 543474 76816 544094 76900
rect 543474 76580 543506 76816
rect 543742 76580 543826 76816
rect 544062 76580 544094 76816
rect 543474 41136 544094 76580
rect 543474 40900 543506 41136
rect 543742 40900 543826 41136
rect 544062 40900 544094 41136
rect 543474 40816 544094 40900
rect 543474 40580 543506 40816
rect 543742 40580 543826 40816
rect 544062 40580 544094 40816
rect 543474 5136 544094 40580
rect 543474 4900 543506 5136
rect 543742 4900 543826 5136
rect 544062 4900 544094 5136
rect 543474 4816 544094 4900
rect 543474 4580 543506 4816
rect 543742 4580 543826 4816
rect 544062 4580 544094 4816
rect 543474 -2264 544094 4580
rect 543474 -2500 543506 -2264
rect 543742 -2500 543826 -2264
rect 544062 -2500 544094 -2264
rect 543474 -2584 544094 -2500
rect 543474 -2820 543506 -2584
rect 543742 -2820 543826 -2584
rect 544062 -2820 544094 -2584
rect 543474 -7652 544094 -2820
rect 544714 258376 545334 279790
rect 544714 258140 544746 258376
rect 544982 258140 545066 258376
rect 545302 258140 545334 258376
rect 544714 258056 545334 258140
rect 544714 257820 544746 258056
rect 544982 257820 545066 258056
rect 545302 257820 545334 258056
rect 544714 222376 545334 257820
rect 544714 222140 544746 222376
rect 544982 222140 545066 222376
rect 545302 222140 545334 222376
rect 544714 222056 545334 222140
rect 544714 221820 544746 222056
rect 544982 221820 545066 222056
rect 545302 221820 545334 222056
rect 544714 186376 545334 221820
rect 544714 186140 544746 186376
rect 544982 186140 545066 186376
rect 545302 186140 545334 186376
rect 544714 186056 545334 186140
rect 544714 185820 544746 186056
rect 544982 185820 545066 186056
rect 545302 185820 545334 186056
rect 544714 150376 545334 185820
rect 544714 150140 544746 150376
rect 544982 150140 545066 150376
rect 545302 150140 545334 150376
rect 544714 150056 545334 150140
rect 544714 149820 544746 150056
rect 544982 149820 545066 150056
rect 545302 149820 545334 150056
rect 544714 114376 545334 149820
rect 544714 114140 544746 114376
rect 544982 114140 545066 114376
rect 545302 114140 545334 114376
rect 544714 114056 545334 114140
rect 544714 113820 544746 114056
rect 544982 113820 545066 114056
rect 545302 113820 545334 114056
rect 544714 78376 545334 113820
rect 544714 78140 544746 78376
rect 544982 78140 545066 78376
rect 545302 78140 545334 78376
rect 544714 78056 545334 78140
rect 544714 77820 544746 78056
rect 544982 77820 545066 78056
rect 545302 77820 545334 78056
rect 544714 42376 545334 77820
rect 544714 42140 544746 42376
rect 544982 42140 545066 42376
rect 545302 42140 545334 42376
rect 544714 42056 545334 42140
rect 544714 41820 544746 42056
rect 544982 41820 545066 42056
rect 545302 41820 545334 42056
rect 544714 6376 545334 41820
rect 544714 6140 544746 6376
rect 544982 6140 545066 6376
rect 545302 6140 545334 6376
rect 544714 6056 545334 6140
rect 544714 5820 544746 6056
rect 544982 5820 545066 6056
rect 545302 5820 545334 6056
rect 544714 -3224 545334 5820
rect 544714 -3460 544746 -3224
rect 544982 -3460 545066 -3224
rect 545302 -3460 545334 -3224
rect 544714 -3544 545334 -3460
rect 544714 -3780 544746 -3544
rect 544982 -3780 545066 -3544
rect 545302 -3780 545334 -3544
rect 544714 -7652 545334 -3780
rect 545954 259616 546574 279790
rect 545954 259380 545986 259616
rect 546222 259380 546306 259616
rect 546542 259380 546574 259616
rect 545954 259296 546574 259380
rect 545954 259060 545986 259296
rect 546222 259060 546306 259296
rect 546542 259060 546574 259296
rect 545954 223616 546574 259060
rect 545954 223380 545986 223616
rect 546222 223380 546306 223616
rect 546542 223380 546574 223616
rect 545954 223296 546574 223380
rect 545954 223060 545986 223296
rect 546222 223060 546306 223296
rect 546542 223060 546574 223296
rect 545954 187616 546574 223060
rect 545954 187380 545986 187616
rect 546222 187380 546306 187616
rect 546542 187380 546574 187616
rect 545954 187296 546574 187380
rect 545954 187060 545986 187296
rect 546222 187060 546306 187296
rect 546542 187060 546574 187296
rect 545954 151616 546574 187060
rect 545954 151380 545986 151616
rect 546222 151380 546306 151616
rect 546542 151380 546574 151616
rect 545954 151296 546574 151380
rect 545954 151060 545986 151296
rect 546222 151060 546306 151296
rect 546542 151060 546574 151296
rect 545954 115616 546574 151060
rect 545954 115380 545986 115616
rect 546222 115380 546306 115616
rect 546542 115380 546574 115616
rect 545954 115296 546574 115380
rect 545954 115060 545986 115296
rect 546222 115060 546306 115296
rect 546542 115060 546574 115296
rect 545954 79616 546574 115060
rect 545954 79380 545986 79616
rect 546222 79380 546306 79616
rect 546542 79380 546574 79616
rect 545954 79296 546574 79380
rect 545954 79060 545986 79296
rect 546222 79060 546306 79296
rect 546542 79060 546574 79296
rect 545954 43616 546574 79060
rect 545954 43380 545986 43616
rect 546222 43380 546306 43616
rect 546542 43380 546574 43616
rect 545954 43296 546574 43380
rect 545954 43060 545986 43296
rect 546222 43060 546306 43296
rect 546542 43060 546574 43296
rect 545954 7616 546574 43060
rect 545954 7380 545986 7616
rect 546222 7380 546306 7616
rect 546542 7380 546574 7616
rect 545954 7296 546574 7380
rect 545954 7060 545986 7296
rect 546222 7060 546306 7296
rect 546542 7060 546574 7296
rect 545954 -4184 546574 7060
rect 545954 -4420 545986 -4184
rect 546222 -4420 546306 -4184
rect 546542 -4420 546574 -4184
rect 545954 -4504 546574 -4420
rect 545954 -4740 545986 -4504
rect 546222 -4740 546306 -4504
rect 546542 -4740 546574 -4504
rect 545954 -7652 546574 -4740
rect 547194 260856 547814 296300
rect 547194 260620 547226 260856
rect 547462 260620 547546 260856
rect 547782 260620 547814 260856
rect 547194 260536 547814 260620
rect 547194 260300 547226 260536
rect 547462 260300 547546 260536
rect 547782 260300 547814 260536
rect 547194 224856 547814 260300
rect 547194 224620 547226 224856
rect 547462 224620 547546 224856
rect 547782 224620 547814 224856
rect 547194 224536 547814 224620
rect 547194 224300 547226 224536
rect 547462 224300 547546 224536
rect 547782 224300 547814 224536
rect 547194 188856 547814 224300
rect 547194 188620 547226 188856
rect 547462 188620 547546 188856
rect 547782 188620 547814 188856
rect 547194 188536 547814 188620
rect 547194 188300 547226 188536
rect 547462 188300 547546 188536
rect 547782 188300 547814 188536
rect 547194 152856 547814 188300
rect 547194 152620 547226 152856
rect 547462 152620 547546 152856
rect 547782 152620 547814 152856
rect 547194 152536 547814 152620
rect 547194 152300 547226 152536
rect 547462 152300 547546 152536
rect 547782 152300 547814 152536
rect 547194 116856 547814 152300
rect 547194 116620 547226 116856
rect 547462 116620 547546 116856
rect 547782 116620 547814 116856
rect 547194 116536 547814 116620
rect 547194 116300 547226 116536
rect 547462 116300 547546 116536
rect 547782 116300 547814 116536
rect 547194 80856 547814 116300
rect 547194 80620 547226 80856
rect 547462 80620 547546 80856
rect 547782 80620 547814 80856
rect 547194 80536 547814 80620
rect 547194 80300 547226 80536
rect 547462 80300 547546 80536
rect 547782 80300 547814 80536
rect 547194 44856 547814 80300
rect 547194 44620 547226 44856
rect 547462 44620 547546 44856
rect 547782 44620 547814 44856
rect 547194 44536 547814 44620
rect 547194 44300 547226 44536
rect 547462 44300 547546 44536
rect 547782 44300 547814 44536
rect 547194 8856 547814 44300
rect 547194 8620 547226 8856
rect 547462 8620 547546 8856
rect 547782 8620 547814 8856
rect 547194 8536 547814 8620
rect 547194 8300 547226 8536
rect 547462 8300 547546 8536
rect 547782 8300 547814 8536
rect 547194 -5144 547814 8300
rect 547194 -5380 547226 -5144
rect 547462 -5380 547546 -5144
rect 547782 -5380 547814 -5144
rect 547194 -5464 547814 -5380
rect 547194 -5700 547226 -5464
rect 547462 -5700 547546 -5464
rect 547782 -5700 547814 -5464
rect 547194 -7652 547814 -5700
rect 548434 710600 549054 711592
rect 548434 710364 548466 710600
rect 548702 710364 548786 710600
rect 549022 710364 549054 710600
rect 548434 710280 549054 710364
rect 548434 710044 548466 710280
rect 548702 710044 548786 710280
rect 549022 710044 549054 710280
rect 548434 694096 549054 710044
rect 548434 693860 548466 694096
rect 548702 693860 548786 694096
rect 549022 693860 549054 694096
rect 548434 693776 549054 693860
rect 548434 693540 548466 693776
rect 548702 693540 548786 693776
rect 549022 693540 549054 693776
rect 548434 658096 549054 693540
rect 548434 657860 548466 658096
rect 548702 657860 548786 658096
rect 549022 657860 549054 658096
rect 548434 657776 549054 657860
rect 548434 657540 548466 657776
rect 548702 657540 548786 657776
rect 549022 657540 549054 657776
rect 548434 622096 549054 657540
rect 548434 621860 548466 622096
rect 548702 621860 548786 622096
rect 549022 621860 549054 622096
rect 548434 621776 549054 621860
rect 548434 621540 548466 621776
rect 548702 621540 548786 621776
rect 549022 621540 549054 621776
rect 548434 586096 549054 621540
rect 548434 585860 548466 586096
rect 548702 585860 548786 586096
rect 549022 585860 549054 586096
rect 548434 585776 549054 585860
rect 548434 585540 548466 585776
rect 548702 585540 548786 585776
rect 549022 585540 549054 585776
rect 548434 550096 549054 585540
rect 548434 549860 548466 550096
rect 548702 549860 548786 550096
rect 549022 549860 549054 550096
rect 548434 549776 549054 549860
rect 548434 549540 548466 549776
rect 548702 549540 548786 549776
rect 549022 549540 549054 549776
rect 548434 514096 549054 549540
rect 548434 513860 548466 514096
rect 548702 513860 548786 514096
rect 549022 513860 549054 514096
rect 548434 513776 549054 513860
rect 548434 513540 548466 513776
rect 548702 513540 548786 513776
rect 549022 513540 549054 513776
rect 548434 478096 549054 513540
rect 548434 477860 548466 478096
rect 548702 477860 548786 478096
rect 549022 477860 549054 478096
rect 548434 477776 549054 477860
rect 548434 477540 548466 477776
rect 548702 477540 548786 477776
rect 549022 477540 549054 477776
rect 548434 442096 549054 477540
rect 548434 441860 548466 442096
rect 548702 441860 548786 442096
rect 549022 441860 549054 442096
rect 548434 441776 549054 441860
rect 548434 441540 548466 441776
rect 548702 441540 548786 441776
rect 549022 441540 549054 441776
rect 548434 406096 549054 441540
rect 548434 405860 548466 406096
rect 548702 405860 548786 406096
rect 549022 405860 549054 406096
rect 548434 405776 549054 405860
rect 548434 405540 548466 405776
rect 548702 405540 548786 405776
rect 549022 405540 549054 405776
rect 548434 370096 549054 405540
rect 548434 369860 548466 370096
rect 548702 369860 548786 370096
rect 549022 369860 549054 370096
rect 548434 369776 549054 369860
rect 548434 369540 548466 369776
rect 548702 369540 548786 369776
rect 549022 369540 549054 369776
rect 548434 334096 549054 369540
rect 548434 333860 548466 334096
rect 548702 333860 548786 334096
rect 549022 333860 549054 334096
rect 548434 333776 549054 333860
rect 548434 333540 548466 333776
rect 548702 333540 548786 333776
rect 549022 333540 549054 333776
rect 548434 298096 549054 333540
rect 548434 297860 548466 298096
rect 548702 297860 548786 298096
rect 549022 297860 549054 298096
rect 548434 297776 549054 297860
rect 548434 297540 548466 297776
rect 548702 297540 548786 297776
rect 549022 297540 549054 297776
rect 548434 262096 549054 297540
rect 548434 261860 548466 262096
rect 548702 261860 548786 262096
rect 549022 261860 549054 262096
rect 548434 261776 549054 261860
rect 548434 261540 548466 261776
rect 548702 261540 548786 261776
rect 549022 261540 549054 261776
rect 548434 226096 549054 261540
rect 548434 225860 548466 226096
rect 548702 225860 548786 226096
rect 549022 225860 549054 226096
rect 548434 225776 549054 225860
rect 548434 225540 548466 225776
rect 548702 225540 548786 225776
rect 549022 225540 549054 225776
rect 548434 190096 549054 225540
rect 548434 189860 548466 190096
rect 548702 189860 548786 190096
rect 549022 189860 549054 190096
rect 548434 189776 549054 189860
rect 548434 189540 548466 189776
rect 548702 189540 548786 189776
rect 549022 189540 549054 189776
rect 548434 154096 549054 189540
rect 548434 153860 548466 154096
rect 548702 153860 548786 154096
rect 549022 153860 549054 154096
rect 548434 153776 549054 153860
rect 548434 153540 548466 153776
rect 548702 153540 548786 153776
rect 549022 153540 549054 153776
rect 548434 118096 549054 153540
rect 548434 117860 548466 118096
rect 548702 117860 548786 118096
rect 549022 117860 549054 118096
rect 548434 117776 549054 117860
rect 548434 117540 548466 117776
rect 548702 117540 548786 117776
rect 549022 117540 549054 117776
rect 548434 82096 549054 117540
rect 548434 81860 548466 82096
rect 548702 81860 548786 82096
rect 549022 81860 549054 82096
rect 548434 81776 549054 81860
rect 548434 81540 548466 81776
rect 548702 81540 548786 81776
rect 549022 81540 549054 81776
rect 548434 46096 549054 81540
rect 548434 45860 548466 46096
rect 548702 45860 548786 46096
rect 549022 45860 549054 46096
rect 548434 45776 549054 45860
rect 548434 45540 548466 45776
rect 548702 45540 548786 45776
rect 549022 45540 549054 45776
rect 548434 10096 549054 45540
rect 548434 9860 548466 10096
rect 548702 9860 548786 10096
rect 549022 9860 549054 10096
rect 548434 9776 549054 9860
rect 548434 9540 548466 9776
rect 548702 9540 548786 9776
rect 549022 9540 549054 9776
rect 548434 -6104 549054 9540
rect 548434 -6340 548466 -6104
rect 548702 -6340 548786 -6104
rect 549022 -6340 549054 -6104
rect 548434 -6424 549054 -6340
rect 548434 -6660 548466 -6424
rect 548702 -6660 548786 -6424
rect 549022 -6660 549054 -6424
rect 548434 -7652 549054 -6660
rect 549674 711560 550294 711592
rect 549674 711324 549706 711560
rect 549942 711324 550026 711560
rect 550262 711324 550294 711560
rect 549674 711240 550294 711324
rect 549674 711004 549706 711240
rect 549942 711004 550026 711240
rect 550262 711004 550294 711240
rect 549674 695336 550294 711004
rect 549674 695100 549706 695336
rect 549942 695100 550026 695336
rect 550262 695100 550294 695336
rect 549674 695016 550294 695100
rect 549674 694780 549706 695016
rect 549942 694780 550026 695016
rect 550262 694780 550294 695016
rect 549674 659336 550294 694780
rect 549674 659100 549706 659336
rect 549942 659100 550026 659336
rect 550262 659100 550294 659336
rect 549674 659016 550294 659100
rect 549674 658780 549706 659016
rect 549942 658780 550026 659016
rect 550262 658780 550294 659016
rect 549674 623336 550294 658780
rect 549674 623100 549706 623336
rect 549942 623100 550026 623336
rect 550262 623100 550294 623336
rect 549674 623016 550294 623100
rect 549674 622780 549706 623016
rect 549942 622780 550026 623016
rect 550262 622780 550294 623016
rect 549674 587336 550294 622780
rect 549674 587100 549706 587336
rect 549942 587100 550026 587336
rect 550262 587100 550294 587336
rect 549674 587016 550294 587100
rect 549674 586780 549706 587016
rect 549942 586780 550026 587016
rect 550262 586780 550294 587016
rect 549674 551336 550294 586780
rect 549674 551100 549706 551336
rect 549942 551100 550026 551336
rect 550262 551100 550294 551336
rect 549674 551016 550294 551100
rect 549674 550780 549706 551016
rect 549942 550780 550026 551016
rect 550262 550780 550294 551016
rect 549674 515336 550294 550780
rect 549674 515100 549706 515336
rect 549942 515100 550026 515336
rect 550262 515100 550294 515336
rect 549674 515016 550294 515100
rect 549674 514780 549706 515016
rect 549942 514780 550026 515016
rect 550262 514780 550294 515016
rect 549674 479336 550294 514780
rect 549674 479100 549706 479336
rect 549942 479100 550026 479336
rect 550262 479100 550294 479336
rect 549674 479016 550294 479100
rect 549674 478780 549706 479016
rect 549942 478780 550026 479016
rect 550262 478780 550294 479016
rect 549674 443336 550294 478780
rect 549674 443100 549706 443336
rect 549942 443100 550026 443336
rect 550262 443100 550294 443336
rect 549674 443016 550294 443100
rect 549674 442780 549706 443016
rect 549942 442780 550026 443016
rect 550262 442780 550294 443016
rect 549674 407336 550294 442780
rect 549674 407100 549706 407336
rect 549942 407100 550026 407336
rect 550262 407100 550294 407336
rect 549674 407016 550294 407100
rect 549674 406780 549706 407016
rect 549942 406780 550026 407016
rect 550262 406780 550294 407016
rect 549674 371336 550294 406780
rect 549674 371100 549706 371336
rect 549942 371100 550026 371336
rect 550262 371100 550294 371336
rect 549674 371016 550294 371100
rect 549674 370780 549706 371016
rect 549942 370780 550026 371016
rect 550262 370780 550294 371016
rect 549674 335336 550294 370780
rect 549674 335100 549706 335336
rect 549942 335100 550026 335336
rect 550262 335100 550294 335336
rect 549674 335016 550294 335100
rect 549674 334780 549706 335016
rect 549942 334780 550026 335016
rect 550262 334780 550294 335016
rect 549674 299336 550294 334780
rect 549674 299100 549706 299336
rect 549942 299100 550026 299336
rect 550262 299100 550294 299336
rect 549674 299016 550294 299100
rect 549674 298780 549706 299016
rect 549942 298780 550026 299016
rect 550262 298780 550294 299016
rect 549674 263336 550294 298780
rect 549674 263100 549706 263336
rect 549942 263100 550026 263336
rect 550262 263100 550294 263336
rect 549674 263016 550294 263100
rect 549674 262780 549706 263016
rect 549942 262780 550026 263016
rect 550262 262780 550294 263016
rect 549674 227336 550294 262780
rect 549674 227100 549706 227336
rect 549942 227100 550026 227336
rect 550262 227100 550294 227336
rect 549674 227016 550294 227100
rect 549674 226780 549706 227016
rect 549942 226780 550026 227016
rect 550262 226780 550294 227016
rect 549674 191336 550294 226780
rect 549674 191100 549706 191336
rect 549942 191100 550026 191336
rect 550262 191100 550294 191336
rect 549674 191016 550294 191100
rect 549674 190780 549706 191016
rect 549942 190780 550026 191016
rect 550262 190780 550294 191016
rect 549674 155336 550294 190780
rect 549674 155100 549706 155336
rect 549942 155100 550026 155336
rect 550262 155100 550294 155336
rect 549674 155016 550294 155100
rect 549674 154780 549706 155016
rect 549942 154780 550026 155016
rect 550262 154780 550294 155016
rect 549674 119336 550294 154780
rect 549674 119100 549706 119336
rect 549942 119100 550026 119336
rect 550262 119100 550294 119336
rect 549674 119016 550294 119100
rect 549674 118780 549706 119016
rect 549942 118780 550026 119016
rect 550262 118780 550294 119016
rect 549674 83336 550294 118780
rect 549674 83100 549706 83336
rect 549942 83100 550026 83336
rect 550262 83100 550294 83336
rect 549674 83016 550294 83100
rect 549674 82780 549706 83016
rect 549942 82780 550026 83016
rect 550262 82780 550294 83016
rect 549674 47336 550294 82780
rect 549674 47100 549706 47336
rect 549942 47100 550026 47336
rect 550262 47100 550294 47336
rect 549674 47016 550294 47100
rect 549674 46780 549706 47016
rect 549942 46780 550026 47016
rect 550262 46780 550294 47016
rect 549674 11336 550294 46780
rect 549674 11100 549706 11336
rect 549942 11100 550026 11336
rect 550262 11100 550294 11336
rect 549674 11016 550294 11100
rect 549674 10780 549706 11016
rect 549942 10780 550026 11016
rect 550262 10780 550294 11016
rect 549674 -7064 550294 10780
rect 549674 -7300 549706 -7064
rect 549942 -7300 550026 -7064
rect 550262 -7300 550294 -7064
rect 549674 -7384 550294 -7300
rect 549674 -7620 549706 -7384
rect 549942 -7620 550026 -7384
rect 550262 -7620 550294 -7384
rect 549674 -7652 550294 -7620
rect 576994 704840 577614 711592
rect 576994 704604 577026 704840
rect 577262 704604 577346 704840
rect 577582 704604 577614 704840
rect 576994 704520 577614 704604
rect 576994 704284 577026 704520
rect 577262 704284 577346 704520
rect 577582 704284 577614 704520
rect 576994 697910 577614 704284
rect 576994 697846 577032 697910
rect 577096 697846 577112 697910
rect 577176 697846 577192 697910
rect 577256 697846 577272 697910
rect 577336 697846 577352 697910
rect 577416 697846 577432 697910
rect 577496 697846 577512 697910
rect 577576 697846 577614 697910
rect 576994 697830 577614 697846
rect 576994 697766 577032 697830
rect 577096 697766 577112 697830
rect 577176 697766 577192 697830
rect 577256 697766 577272 697830
rect 577336 697766 577352 697830
rect 577416 697766 577432 697830
rect 577496 697766 577512 697830
rect 577576 697766 577614 697830
rect 576994 697750 577614 697766
rect 576994 697686 577032 697750
rect 577096 697686 577112 697750
rect 577176 697686 577192 697750
rect 577256 697686 577272 697750
rect 577336 697686 577352 697750
rect 577416 697686 577432 697750
rect 577496 697686 577512 697750
rect 577576 697686 577614 697750
rect 576994 697670 577614 697686
rect 576994 697606 577032 697670
rect 577096 697606 577112 697670
rect 577176 697606 577192 697670
rect 577256 697606 577272 697670
rect 577336 697606 577352 697670
rect 577416 697606 577432 697670
rect 577496 697606 577512 697670
rect 577576 697606 577614 697670
rect 576994 686656 577614 697606
rect 576994 686420 577026 686656
rect 577262 686420 577346 686656
rect 577582 686420 577614 686656
rect 576994 686336 577614 686420
rect 576994 686100 577026 686336
rect 577262 686100 577346 686336
rect 577582 686100 577614 686336
rect 576994 650656 577614 686100
rect 576994 650420 577026 650656
rect 577262 650420 577346 650656
rect 577582 650420 577614 650656
rect 576994 650336 577614 650420
rect 576994 650100 577026 650336
rect 577262 650100 577346 650336
rect 577582 650100 577614 650336
rect 576994 644734 577614 650100
rect 576994 644670 577032 644734
rect 577096 644670 577112 644734
rect 577176 644670 577192 644734
rect 577256 644670 577272 644734
rect 577336 644670 577352 644734
rect 577416 644670 577432 644734
rect 577496 644670 577512 644734
rect 577576 644670 577614 644734
rect 576994 644654 577614 644670
rect 576994 644590 577032 644654
rect 577096 644590 577112 644654
rect 577176 644590 577192 644654
rect 577256 644590 577272 644654
rect 577336 644590 577352 644654
rect 577416 644590 577432 644654
rect 577496 644590 577512 644654
rect 577576 644590 577614 644654
rect 576994 644574 577614 644590
rect 576994 644510 577032 644574
rect 577096 644510 577112 644574
rect 577176 644510 577192 644574
rect 577256 644510 577272 644574
rect 577336 644510 577352 644574
rect 577416 644510 577432 644574
rect 577496 644510 577512 644574
rect 577576 644510 577614 644574
rect 576994 644494 577614 644510
rect 576994 644430 577032 644494
rect 577096 644430 577112 644494
rect 577176 644430 577192 644494
rect 577256 644430 577272 644494
rect 577336 644430 577352 644494
rect 577416 644430 577432 644494
rect 577496 644430 577512 644494
rect 577576 644430 577614 644494
rect 576994 614656 577614 644430
rect 576994 614420 577026 614656
rect 577262 614420 577346 614656
rect 577582 614420 577614 614656
rect 576994 614336 577614 614420
rect 576994 614100 577026 614336
rect 577262 614100 577346 614336
rect 577582 614100 577614 614336
rect 576994 591694 577614 614100
rect 576994 591630 577032 591694
rect 577096 591630 577112 591694
rect 577176 591630 577192 591694
rect 577256 591630 577272 591694
rect 577336 591630 577352 591694
rect 577416 591630 577432 591694
rect 577496 591630 577512 591694
rect 577576 591630 577614 591694
rect 576994 591614 577614 591630
rect 576994 591550 577032 591614
rect 577096 591550 577112 591614
rect 577176 591550 577192 591614
rect 577256 591550 577272 591614
rect 577336 591550 577352 591614
rect 577416 591550 577432 591614
rect 577496 591550 577512 591614
rect 577576 591550 577614 591614
rect 576994 591534 577614 591550
rect 576994 591470 577032 591534
rect 577096 591470 577112 591534
rect 577176 591470 577192 591534
rect 577256 591470 577272 591534
rect 577336 591470 577352 591534
rect 577416 591470 577432 591534
rect 577496 591470 577512 591534
rect 577576 591470 577614 591534
rect 576994 591454 577614 591470
rect 576994 591390 577032 591454
rect 577096 591390 577112 591454
rect 577176 591390 577192 591454
rect 577256 591390 577272 591454
rect 577336 591390 577352 591454
rect 577416 591390 577432 591454
rect 577496 591390 577512 591454
rect 577576 591390 577614 591454
rect 576994 578656 577614 591390
rect 576994 578420 577026 578656
rect 577262 578420 577346 578656
rect 577582 578420 577614 578656
rect 576994 578336 577614 578420
rect 576994 578100 577026 578336
rect 577262 578100 577346 578336
rect 577582 578100 577614 578336
rect 576994 542656 577614 578100
rect 576994 542420 577026 542656
rect 577262 542420 577346 542656
rect 577582 542420 577614 542656
rect 576994 542336 577614 542420
rect 576994 542100 577026 542336
rect 577262 542100 577346 542336
rect 577582 542100 577614 542336
rect 576994 538518 577614 542100
rect 576994 538454 577032 538518
rect 577096 538454 577112 538518
rect 577176 538454 577192 538518
rect 577256 538454 577272 538518
rect 577336 538454 577352 538518
rect 577416 538454 577432 538518
rect 577496 538454 577512 538518
rect 577576 538454 577614 538518
rect 576994 538438 577614 538454
rect 576994 538374 577032 538438
rect 577096 538374 577112 538438
rect 577176 538374 577192 538438
rect 577256 538374 577272 538438
rect 577336 538374 577352 538438
rect 577416 538374 577432 538438
rect 577496 538374 577512 538438
rect 577576 538374 577614 538438
rect 576994 538358 577614 538374
rect 576994 538294 577032 538358
rect 577096 538294 577112 538358
rect 577176 538294 577192 538358
rect 577256 538294 577272 538358
rect 577336 538294 577352 538358
rect 577416 538294 577432 538358
rect 577496 538294 577512 538358
rect 577576 538294 577614 538358
rect 576994 538278 577614 538294
rect 576994 538214 577032 538278
rect 577096 538214 577112 538278
rect 577176 538214 577192 538278
rect 577256 538214 577272 538278
rect 577336 538214 577352 538278
rect 577416 538214 577432 538278
rect 577496 538214 577512 538278
rect 577576 538214 577614 538278
rect 576994 506656 577614 538214
rect 576994 506420 577026 506656
rect 577262 506420 577346 506656
rect 577582 506420 577614 506656
rect 576994 506336 577614 506420
rect 576994 506100 577026 506336
rect 577262 506100 577346 506336
rect 577582 506100 577614 506336
rect 576994 485342 577614 506100
rect 576994 485278 577032 485342
rect 577096 485278 577112 485342
rect 577176 485278 577192 485342
rect 577256 485278 577272 485342
rect 577336 485278 577352 485342
rect 577416 485278 577432 485342
rect 577496 485278 577512 485342
rect 577576 485278 577614 485342
rect 576994 485262 577614 485278
rect 576994 485198 577032 485262
rect 577096 485198 577112 485262
rect 577176 485198 577192 485262
rect 577256 485198 577272 485262
rect 577336 485198 577352 485262
rect 577416 485198 577432 485262
rect 577496 485198 577512 485262
rect 577576 485198 577614 485262
rect 576994 485182 577614 485198
rect 576994 485118 577032 485182
rect 577096 485118 577112 485182
rect 577176 485118 577192 485182
rect 577256 485118 577272 485182
rect 577336 485118 577352 485182
rect 577416 485118 577432 485182
rect 577496 485118 577512 485182
rect 577576 485118 577614 485182
rect 576994 485102 577614 485118
rect 576994 485038 577032 485102
rect 577096 485038 577112 485102
rect 577176 485038 577192 485102
rect 577256 485038 577272 485102
rect 577336 485038 577352 485102
rect 577416 485038 577432 485102
rect 577496 485038 577512 485102
rect 577576 485038 577614 485102
rect 576994 470656 577614 485038
rect 576994 470420 577026 470656
rect 577262 470420 577346 470656
rect 577582 470420 577614 470656
rect 576994 470336 577614 470420
rect 576994 470100 577026 470336
rect 577262 470100 577346 470336
rect 577582 470100 577614 470336
rect 576994 434656 577614 470100
rect 576994 434420 577026 434656
rect 577262 434420 577346 434656
rect 577582 434420 577614 434656
rect 576994 434336 577614 434420
rect 576994 434100 577026 434336
rect 577262 434100 577346 434336
rect 577582 434100 577614 434336
rect 576994 432302 577614 434100
rect 576994 432238 577032 432302
rect 577096 432238 577112 432302
rect 577176 432238 577192 432302
rect 577256 432238 577272 432302
rect 577336 432238 577352 432302
rect 577416 432238 577432 432302
rect 577496 432238 577512 432302
rect 577576 432238 577614 432302
rect 576994 432222 577614 432238
rect 576994 432158 577032 432222
rect 577096 432158 577112 432222
rect 577176 432158 577192 432222
rect 577256 432158 577272 432222
rect 577336 432158 577352 432222
rect 577416 432158 577432 432222
rect 577496 432158 577512 432222
rect 577576 432158 577614 432222
rect 576994 432142 577614 432158
rect 576994 432078 577032 432142
rect 577096 432078 577112 432142
rect 577176 432078 577192 432142
rect 577256 432078 577272 432142
rect 577336 432078 577352 432142
rect 577416 432078 577432 432142
rect 577496 432078 577512 432142
rect 577576 432078 577614 432142
rect 576994 432062 577614 432078
rect 576994 431998 577032 432062
rect 577096 431998 577112 432062
rect 577176 431998 577192 432062
rect 577256 431998 577272 432062
rect 577336 431998 577352 432062
rect 577416 431998 577432 432062
rect 577496 431998 577512 432062
rect 577576 431998 577614 432062
rect 576994 398656 577614 431998
rect 576994 398420 577026 398656
rect 577262 398420 577346 398656
rect 577582 398420 577614 398656
rect 576994 398336 577614 398420
rect 576994 398100 577026 398336
rect 577262 398100 577346 398336
rect 577582 398100 577614 398336
rect 576994 379126 577614 398100
rect 576994 379062 577032 379126
rect 577096 379062 577112 379126
rect 577176 379062 577192 379126
rect 577256 379062 577272 379126
rect 577336 379062 577352 379126
rect 577416 379062 577432 379126
rect 577496 379062 577512 379126
rect 577576 379062 577614 379126
rect 576994 379046 577614 379062
rect 576994 378982 577032 379046
rect 577096 378982 577112 379046
rect 577176 378982 577192 379046
rect 577256 378982 577272 379046
rect 577336 378982 577352 379046
rect 577416 378982 577432 379046
rect 577496 378982 577512 379046
rect 577576 378982 577614 379046
rect 576994 378966 577614 378982
rect 576994 378902 577032 378966
rect 577096 378902 577112 378966
rect 577176 378902 577192 378966
rect 577256 378902 577272 378966
rect 577336 378902 577352 378966
rect 577416 378902 577432 378966
rect 577496 378902 577512 378966
rect 577576 378902 577614 378966
rect 576994 378886 577614 378902
rect 576994 378822 577032 378886
rect 577096 378822 577112 378886
rect 577176 378822 577192 378886
rect 577256 378822 577272 378886
rect 577336 378822 577352 378886
rect 577416 378822 577432 378886
rect 577496 378822 577512 378886
rect 577576 378822 577614 378886
rect 576994 362656 577614 378822
rect 576994 362420 577026 362656
rect 577262 362420 577346 362656
rect 577582 362420 577614 362656
rect 576994 362336 577614 362420
rect 576994 362100 577026 362336
rect 577262 362100 577346 362336
rect 577582 362100 577614 362336
rect 576994 326656 577614 362100
rect 576994 326420 577026 326656
rect 577262 326420 577346 326656
rect 577582 326420 577614 326656
rect 576994 326336 577614 326420
rect 576994 326100 577026 326336
rect 577262 326100 577346 326336
rect 577582 326100 577614 326336
rect 576994 325950 577614 326100
rect 576994 325886 577032 325950
rect 577096 325886 577112 325950
rect 577176 325886 577192 325950
rect 577256 325886 577272 325950
rect 577336 325886 577352 325950
rect 577416 325886 577432 325950
rect 577496 325886 577512 325950
rect 577576 325886 577614 325950
rect 576994 325870 577614 325886
rect 576994 325806 577032 325870
rect 577096 325806 577112 325870
rect 577176 325806 577192 325870
rect 577256 325806 577272 325870
rect 577336 325806 577352 325870
rect 577416 325806 577432 325870
rect 577496 325806 577512 325870
rect 577576 325806 577614 325870
rect 576994 325790 577614 325806
rect 576994 325726 577032 325790
rect 577096 325726 577112 325790
rect 577176 325726 577192 325790
rect 577256 325726 577272 325790
rect 577336 325726 577352 325790
rect 577416 325726 577432 325790
rect 577496 325726 577512 325790
rect 577576 325726 577614 325790
rect 576994 325710 577614 325726
rect 576994 325646 577032 325710
rect 577096 325646 577112 325710
rect 577176 325646 577192 325710
rect 577256 325646 577272 325710
rect 577336 325646 577352 325710
rect 577416 325646 577432 325710
rect 577496 325646 577512 325710
rect 577576 325646 577614 325710
rect 576994 290656 577614 325646
rect 576994 290420 577026 290656
rect 577262 290420 577346 290656
rect 577582 290420 577614 290656
rect 576994 290336 577614 290420
rect 576994 290100 577026 290336
rect 577262 290100 577346 290336
rect 577582 290100 577614 290336
rect 576994 272910 577614 290100
rect 576994 272846 577032 272910
rect 577096 272846 577112 272910
rect 577176 272846 577192 272910
rect 577256 272846 577272 272910
rect 577336 272846 577352 272910
rect 577416 272846 577432 272910
rect 577496 272846 577512 272910
rect 577576 272846 577614 272910
rect 576994 272830 577614 272846
rect 576994 272766 577032 272830
rect 577096 272766 577112 272830
rect 577176 272766 577192 272830
rect 577256 272766 577272 272830
rect 577336 272766 577352 272830
rect 577416 272766 577432 272830
rect 577496 272766 577512 272830
rect 577576 272766 577614 272830
rect 576994 272750 577614 272766
rect 576994 272686 577032 272750
rect 577096 272686 577112 272750
rect 577176 272686 577192 272750
rect 577256 272686 577272 272750
rect 577336 272686 577352 272750
rect 577416 272686 577432 272750
rect 577496 272686 577512 272750
rect 577576 272686 577614 272750
rect 576994 272670 577614 272686
rect 576994 272606 577032 272670
rect 577096 272606 577112 272670
rect 577176 272606 577192 272670
rect 577256 272606 577272 272670
rect 577336 272606 577352 272670
rect 577416 272606 577432 272670
rect 577496 272606 577512 272670
rect 577576 272606 577614 272670
rect 576994 254656 577614 272606
rect 576994 254420 577026 254656
rect 577262 254420 577346 254656
rect 577582 254420 577614 254656
rect 576994 254336 577614 254420
rect 576994 254100 577026 254336
rect 577262 254100 577346 254336
rect 577582 254100 577614 254336
rect 576994 233063 577614 254100
rect 576994 232999 577032 233063
rect 577096 232999 577112 233063
rect 577176 232999 577192 233063
rect 577256 232999 577272 233063
rect 577336 232999 577352 233063
rect 577416 232999 577432 233063
rect 577496 232999 577512 233063
rect 577576 232999 577614 233063
rect 576994 232983 577614 232999
rect 576994 232919 577032 232983
rect 577096 232919 577112 232983
rect 577176 232919 577192 232983
rect 577256 232919 577272 232983
rect 577336 232919 577352 232983
rect 577416 232919 577432 232983
rect 577496 232919 577512 232983
rect 577576 232919 577614 232983
rect 576994 232903 577614 232919
rect 576994 232839 577032 232903
rect 577096 232839 577112 232903
rect 577176 232839 577192 232903
rect 577256 232839 577272 232903
rect 577336 232839 577352 232903
rect 577416 232839 577432 232903
rect 577496 232839 577512 232903
rect 577576 232839 577614 232903
rect 576994 232823 577614 232839
rect 576994 232759 577032 232823
rect 577096 232759 577112 232823
rect 577176 232759 577192 232823
rect 577256 232759 577272 232823
rect 577336 232759 577352 232823
rect 577416 232759 577432 232823
rect 577496 232759 577512 232823
rect 577576 232759 577614 232823
rect 576994 218656 577614 232759
rect 576994 218420 577026 218656
rect 577262 218420 577346 218656
rect 577582 218420 577614 218656
rect 576994 218336 577614 218420
rect 576994 218100 577026 218336
rect 577262 218100 577346 218336
rect 577582 218100 577614 218336
rect 576994 182656 577614 218100
rect 576994 182420 577026 182656
rect 577262 182420 577346 182656
rect 577582 182420 577614 182656
rect 576994 182336 577614 182420
rect 576994 182100 577026 182336
rect 577262 182100 577346 182336
rect 577582 182100 577614 182336
rect 576994 146656 577614 182100
rect 576994 146420 577026 146656
rect 577262 146420 577346 146656
rect 577582 146420 577614 146656
rect 576994 146336 577614 146420
rect 576994 146100 577026 146336
rect 577262 146100 577346 146336
rect 577582 146100 577614 146336
rect 576994 110656 577614 146100
rect 576994 110420 577026 110656
rect 577262 110420 577346 110656
rect 577582 110420 577614 110656
rect 576994 110336 577614 110420
rect 576994 110100 577026 110336
rect 577262 110100 577346 110336
rect 577582 110100 577614 110336
rect 576994 74656 577614 110100
rect 576994 74420 577026 74656
rect 577262 74420 577346 74656
rect 577582 74420 577614 74656
rect 576994 74336 577614 74420
rect 576994 74100 577026 74336
rect 577262 74100 577346 74336
rect 577582 74100 577614 74336
rect 576994 38656 577614 74100
rect 576994 38420 577026 38656
rect 577262 38420 577346 38656
rect 577582 38420 577614 38656
rect 576994 38336 577614 38420
rect 576994 38100 577026 38336
rect 577262 38100 577346 38336
rect 577582 38100 577614 38336
rect 576994 2656 577614 38100
rect 576994 2420 577026 2656
rect 577262 2420 577346 2656
rect 577582 2420 577614 2656
rect 576994 2336 577614 2420
rect 576994 2100 577026 2336
rect 577262 2100 577346 2336
rect 577582 2100 577614 2336
rect 576994 -344 577614 2100
rect 576994 -580 577026 -344
rect 577262 -580 577346 -344
rect 577582 -580 577614 -344
rect 576994 -664 577614 -580
rect 576994 -900 577026 -664
rect 577262 -900 577346 -664
rect 577582 -900 577614 -664
rect 576994 -7652 577614 -900
rect 578234 705800 578854 711592
rect 578234 705564 578266 705800
rect 578502 705564 578586 705800
rect 578822 705564 578854 705800
rect 578234 705480 578854 705564
rect 578234 705244 578266 705480
rect 578502 705244 578586 705480
rect 578822 705244 578854 705480
rect 578234 697115 578854 705244
rect 578234 697051 578272 697115
rect 578336 697051 578352 697115
rect 578416 697051 578432 697115
rect 578496 697051 578512 697115
rect 578576 697051 578592 697115
rect 578656 697051 578672 697115
rect 578736 697051 578752 697115
rect 578816 697051 578854 697115
rect 578234 697035 578854 697051
rect 578234 696971 578272 697035
rect 578336 696971 578352 697035
rect 578416 696971 578432 697035
rect 578496 696971 578512 697035
rect 578576 696971 578592 697035
rect 578656 696971 578672 697035
rect 578736 696971 578752 697035
rect 578816 696971 578854 697035
rect 578234 696955 578854 696971
rect 578234 696891 578272 696955
rect 578336 696891 578352 696955
rect 578416 696891 578432 696955
rect 578496 696891 578512 696955
rect 578576 696891 578592 696955
rect 578656 696891 578672 696955
rect 578736 696891 578752 696955
rect 578816 696891 578854 696955
rect 578234 696875 578854 696891
rect 578234 696811 578272 696875
rect 578336 696811 578352 696875
rect 578416 696811 578432 696875
rect 578496 696811 578512 696875
rect 578576 696811 578592 696875
rect 578656 696811 578672 696875
rect 578736 696811 578752 696875
rect 578816 696811 578854 696875
rect 578234 687896 578854 696811
rect 578234 687660 578266 687896
rect 578502 687660 578586 687896
rect 578822 687660 578854 687896
rect 578234 687576 578854 687660
rect 578234 687340 578266 687576
rect 578502 687340 578586 687576
rect 578822 687340 578854 687576
rect 578234 651896 578854 687340
rect 578234 651660 578266 651896
rect 578502 651660 578586 651896
rect 578822 651660 578854 651896
rect 578234 651576 578854 651660
rect 578234 651340 578266 651576
rect 578502 651340 578586 651576
rect 578822 651340 578854 651576
rect 578234 643939 578854 651340
rect 578234 643875 578272 643939
rect 578336 643875 578352 643939
rect 578416 643875 578432 643939
rect 578496 643875 578512 643939
rect 578576 643875 578592 643939
rect 578656 643875 578672 643939
rect 578736 643875 578752 643939
rect 578816 643875 578854 643939
rect 578234 643859 578854 643875
rect 578234 643795 578272 643859
rect 578336 643795 578352 643859
rect 578416 643795 578432 643859
rect 578496 643795 578512 643859
rect 578576 643795 578592 643859
rect 578656 643795 578672 643859
rect 578736 643795 578752 643859
rect 578816 643795 578854 643859
rect 578234 643779 578854 643795
rect 578234 643715 578272 643779
rect 578336 643715 578352 643779
rect 578416 643715 578432 643779
rect 578496 643715 578512 643779
rect 578576 643715 578592 643779
rect 578656 643715 578672 643779
rect 578736 643715 578752 643779
rect 578816 643715 578854 643779
rect 578234 643699 578854 643715
rect 578234 643635 578272 643699
rect 578336 643635 578352 643699
rect 578416 643635 578432 643699
rect 578496 643635 578512 643699
rect 578576 643635 578592 643699
rect 578656 643635 578672 643699
rect 578736 643635 578752 643699
rect 578816 643635 578854 643699
rect 578234 615896 578854 643635
rect 578234 615660 578266 615896
rect 578502 615660 578586 615896
rect 578822 615660 578854 615896
rect 578234 615576 578854 615660
rect 578234 615340 578266 615576
rect 578502 615340 578586 615576
rect 578822 615340 578854 615576
rect 578234 590899 578854 615340
rect 578234 590835 578272 590899
rect 578336 590835 578352 590899
rect 578416 590835 578432 590899
rect 578496 590835 578512 590899
rect 578576 590835 578592 590899
rect 578656 590835 578672 590899
rect 578736 590835 578752 590899
rect 578816 590835 578854 590899
rect 578234 590819 578854 590835
rect 578234 590755 578272 590819
rect 578336 590755 578352 590819
rect 578416 590755 578432 590819
rect 578496 590755 578512 590819
rect 578576 590755 578592 590819
rect 578656 590755 578672 590819
rect 578736 590755 578752 590819
rect 578816 590755 578854 590819
rect 578234 590739 578854 590755
rect 578234 590675 578272 590739
rect 578336 590675 578352 590739
rect 578416 590675 578432 590739
rect 578496 590675 578512 590739
rect 578576 590675 578592 590739
rect 578656 590675 578672 590739
rect 578736 590675 578752 590739
rect 578816 590675 578854 590739
rect 578234 590659 578854 590675
rect 578234 590595 578272 590659
rect 578336 590595 578352 590659
rect 578416 590595 578432 590659
rect 578496 590595 578512 590659
rect 578576 590595 578592 590659
rect 578656 590595 578672 590659
rect 578736 590595 578752 590659
rect 578816 590595 578854 590659
rect 578234 579896 578854 590595
rect 578234 579660 578266 579896
rect 578502 579660 578586 579896
rect 578822 579660 578854 579896
rect 578234 579576 578854 579660
rect 578234 579340 578266 579576
rect 578502 579340 578586 579576
rect 578822 579340 578854 579576
rect 578234 543896 578854 579340
rect 578234 543660 578266 543896
rect 578502 543660 578586 543896
rect 578822 543660 578854 543896
rect 578234 543576 578854 543660
rect 578234 543340 578266 543576
rect 578502 543340 578586 543576
rect 578822 543340 578854 543576
rect 578234 537723 578854 543340
rect 578234 537659 578272 537723
rect 578336 537659 578352 537723
rect 578416 537659 578432 537723
rect 578496 537659 578512 537723
rect 578576 537659 578592 537723
rect 578656 537659 578672 537723
rect 578736 537659 578752 537723
rect 578816 537659 578854 537723
rect 578234 537643 578854 537659
rect 578234 537579 578272 537643
rect 578336 537579 578352 537643
rect 578416 537579 578432 537643
rect 578496 537579 578512 537643
rect 578576 537579 578592 537643
rect 578656 537579 578672 537643
rect 578736 537579 578752 537643
rect 578816 537579 578854 537643
rect 578234 537563 578854 537579
rect 578234 537499 578272 537563
rect 578336 537499 578352 537563
rect 578416 537499 578432 537563
rect 578496 537499 578512 537563
rect 578576 537499 578592 537563
rect 578656 537499 578672 537563
rect 578736 537499 578752 537563
rect 578816 537499 578854 537563
rect 578234 537483 578854 537499
rect 578234 537419 578272 537483
rect 578336 537419 578352 537483
rect 578416 537419 578432 537483
rect 578496 537419 578512 537483
rect 578576 537419 578592 537483
rect 578656 537419 578672 537483
rect 578736 537419 578752 537483
rect 578816 537419 578854 537483
rect 578234 507896 578854 537419
rect 578234 507660 578266 507896
rect 578502 507660 578586 507896
rect 578822 507660 578854 507896
rect 578234 507576 578854 507660
rect 578234 507340 578266 507576
rect 578502 507340 578586 507576
rect 578822 507340 578854 507576
rect 578234 484547 578854 507340
rect 578234 484483 578272 484547
rect 578336 484483 578352 484547
rect 578416 484483 578432 484547
rect 578496 484483 578512 484547
rect 578576 484483 578592 484547
rect 578656 484483 578672 484547
rect 578736 484483 578752 484547
rect 578816 484483 578854 484547
rect 578234 484467 578854 484483
rect 578234 484403 578272 484467
rect 578336 484403 578352 484467
rect 578416 484403 578432 484467
rect 578496 484403 578512 484467
rect 578576 484403 578592 484467
rect 578656 484403 578672 484467
rect 578736 484403 578752 484467
rect 578816 484403 578854 484467
rect 578234 484387 578854 484403
rect 578234 484323 578272 484387
rect 578336 484323 578352 484387
rect 578416 484323 578432 484387
rect 578496 484323 578512 484387
rect 578576 484323 578592 484387
rect 578656 484323 578672 484387
rect 578736 484323 578752 484387
rect 578816 484323 578854 484387
rect 578234 484307 578854 484323
rect 578234 484243 578272 484307
rect 578336 484243 578352 484307
rect 578416 484243 578432 484307
rect 578496 484243 578512 484307
rect 578576 484243 578592 484307
rect 578656 484243 578672 484307
rect 578736 484243 578752 484307
rect 578816 484243 578854 484307
rect 578234 471896 578854 484243
rect 578234 471660 578266 471896
rect 578502 471660 578586 471896
rect 578822 471660 578854 471896
rect 578234 471576 578854 471660
rect 578234 471340 578266 471576
rect 578502 471340 578586 471576
rect 578822 471340 578854 471576
rect 578234 435896 578854 471340
rect 578234 435660 578266 435896
rect 578502 435660 578586 435896
rect 578822 435660 578854 435896
rect 578234 435576 578854 435660
rect 578234 435340 578266 435576
rect 578502 435340 578586 435576
rect 578822 435340 578854 435576
rect 578234 431507 578854 435340
rect 578234 431443 578272 431507
rect 578336 431443 578352 431507
rect 578416 431443 578432 431507
rect 578496 431443 578512 431507
rect 578576 431443 578592 431507
rect 578656 431443 578672 431507
rect 578736 431443 578752 431507
rect 578816 431443 578854 431507
rect 578234 431427 578854 431443
rect 578234 431363 578272 431427
rect 578336 431363 578352 431427
rect 578416 431363 578432 431427
rect 578496 431363 578512 431427
rect 578576 431363 578592 431427
rect 578656 431363 578672 431427
rect 578736 431363 578752 431427
rect 578816 431363 578854 431427
rect 578234 431347 578854 431363
rect 578234 431283 578272 431347
rect 578336 431283 578352 431347
rect 578416 431283 578432 431347
rect 578496 431283 578512 431347
rect 578576 431283 578592 431347
rect 578656 431283 578672 431347
rect 578736 431283 578752 431347
rect 578816 431283 578854 431347
rect 578234 431267 578854 431283
rect 578234 431203 578272 431267
rect 578336 431203 578352 431267
rect 578416 431203 578432 431267
rect 578496 431203 578512 431267
rect 578576 431203 578592 431267
rect 578656 431203 578672 431267
rect 578736 431203 578752 431267
rect 578816 431203 578854 431267
rect 578234 399896 578854 431203
rect 578234 399660 578266 399896
rect 578502 399660 578586 399896
rect 578822 399660 578854 399896
rect 578234 399576 578854 399660
rect 578234 399340 578266 399576
rect 578502 399340 578586 399576
rect 578822 399340 578854 399576
rect 578234 378331 578854 399340
rect 578234 378267 578272 378331
rect 578336 378267 578352 378331
rect 578416 378267 578432 378331
rect 578496 378267 578512 378331
rect 578576 378267 578592 378331
rect 578656 378267 578672 378331
rect 578736 378267 578752 378331
rect 578816 378267 578854 378331
rect 578234 378251 578854 378267
rect 578234 378187 578272 378251
rect 578336 378187 578352 378251
rect 578416 378187 578432 378251
rect 578496 378187 578512 378251
rect 578576 378187 578592 378251
rect 578656 378187 578672 378251
rect 578736 378187 578752 378251
rect 578816 378187 578854 378251
rect 578234 378171 578854 378187
rect 578234 378107 578272 378171
rect 578336 378107 578352 378171
rect 578416 378107 578432 378171
rect 578496 378107 578512 378171
rect 578576 378107 578592 378171
rect 578656 378107 578672 378171
rect 578736 378107 578752 378171
rect 578816 378107 578854 378171
rect 578234 378091 578854 378107
rect 578234 378027 578272 378091
rect 578336 378027 578352 378091
rect 578416 378027 578432 378091
rect 578496 378027 578512 378091
rect 578576 378027 578592 378091
rect 578656 378027 578672 378091
rect 578736 378027 578752 378091
rect 578816 378027 578854 378091
rect 578234 363896 578854 378027
rect 578234 363660 578266 363896
rect 578502 363660 578586 363896
rect 578822 363660 578854 363896
rect 578234 363576 578854 363660
rect 578234 363340 578266 363576
rect 578502 363340 578586 363576
rect 578822 363340 578854 363576
rect 578234 327896 578854 363340
rect 578234 327660 578266 327896
rect 578502 327660 578586 327896
rect 578822 327660 578854 327896
rect 578234 327576 578854 327660
rect 578234 327340 578266 327576
rect 578502 327340 578586 327576
rect 578822 327340 578854 327576
rect 578234 325155 578854 327340
rect 578234 325091 578272 325155
rect 578336 325091 578352 325155
rect 578416 325091 578432 325155
rect 578496 325091 578512 325155
rect 578576 325091 578592 325155
rect 578656 325091 578672 325155
rect 578736 325091 578752 325155
rect 578816 325091 578854 325155
rect 578234 325075 578854 325091
rect 578234 325011 578272 325075
rect 578336 325011 578352 325075
rect 578416 325011 578432 325075
rect 578496 325011 578512 325075
rect 578576 325011 578592 325075
rect 578656 325011 578672 325075
rect 578736 325011 578752 325075
rect 578816 325011 578854 325075
rect 578234 324995 578854 325011
rect 578234 324931 578272 324995
rect 578336 324931 578352 324995
rect 578416 324931 578432 324995
rect 578496 324931 578512 324995
rect 578576 324931 578592 324995
rect 578656 324931 578672 324995
rect 578736 324931 578752 324995
rect 578816 324931 578854 324995
rect 578234 324915 578854 324931
rect 578234 324851 578272 324915
rect 578336 324851 578352 324915
rect 578416 324851 578432 324915
rect 578496 324851 578512 324915
rect 578576 324851 578592 324915
rect 578656 324851 578672 324915
rect 578736 324851 578752 324915
rect 578816 324851 578854 324915
rect 578234 291896 578854 324851
rect 578234 291660 578266 291896
rect 578502 291660 578586 291896
rect 578822 291660 578854 291896
rect 578234 291576 578854 291660
rect 578234 291340 578266 291576
rect 578502 291340 578586 291576
rect 578822 291340 578854 291576
rect 578234 272115 578854 291340
rect 578234 272051 578272 272115
rect 578336 272051 578352 272115
rect 578416 272051 578432 272115
rect 578496 272051 578512 272115
rect 578576 272051 578592 272115
rect 578656 272051 578672 272115
rect 578736 272051 578752 272115
rect 578816 272051 578854 272115
rect 578234 272035 578854 272051
rect 578234 271971 578272 272035
rect 578336 271971 578352 272035
rect 578416 271971 578432 272035
rect 578496 271971 578512 272035
rect 578576 271971 578592 272035
rect 578656 271971 578672 272035
rect 578736 271971 578752 272035
rect 578816 271971 578854 272035
rect 578234 271955 578854 271971
rect 578234 271891 578272 271955
rect 578336 271891 578352 271955
rect 578416 271891 578432 271955
rect 578496 271891 578512 271955
rect 578576 271891 578592 271955
rect 578656 271891 578672 271955
rect 578736 271891 578752 271955
rect 578816 271891 578854 271955
rect 578234 271875 578854 271891
rect 578234 271811 578272 271875
rect 578336 271811 578352 271875
rect 578416 271811 578432 271875
rect 578496 271811 578512 271875
rect 578576 271811 578592 271875
rect 578656 271811 578672 271875
rect 578736 271811 578752 271875
rect 578816 271811 578854 271875
rect 578234 255896 578854 271811
rect 578234 255660 578266 255896
rect 578502 255660 578586 255896
rect 578822 255660 578854 255896
rect 578234 255576 578854 255660
rect 578234 255340 578266 255576
rect 578502 255340 578586 255576
rect 578822 255340 578854 255576
rect 578234 232268 578854 255340
rect 578234 232204 578272 232268
rect 578336 232204 578352 232268
rect 578416 232204 578432 232268
rect 578496 232204 578512 232268
rect 578576 232204 578592 232268
rect 578656 232204 578672 232268
rect 578736 232204 578752 232268
rect 578816 232204 578854 232268
rect 578234 232188 578854 232204
rect 578234 232124 578272 232188
rect 578336 232124 578352 232188
rect 578416 232124 578432 232188
rect 578496 232124 578512 232188
rect 578576 232124 578592 232188
rect 578656 232124 578672 232188
rect 578736 232124 578752 232188
rect 578816 232124 578854 232188
rect 578234 232108 578854 232124
rect 578234 232044 578272 232108
rect 578336 232044 578352 232108
rect 578416 232044 578432 232108
rect 578496 232044 578512 232108
rect 578576 232044 578592 232108
rect 578656 232044 578672 232108
rect 578736 232044 578752 232108
rect 578816 232044 578854 232108
rect 578234 232028 578854 232044
rect 578234 231964 578272 232028
rect 578336 231964 578352 232028
rect 578416 231964 578432 232028
rect 578496 231964 578512 232028
rect 578576 231964 578592 232028
rect 578656 231964 578672 232028
rect 578736 231964 578752 232028
rect 578816 231964 578854 232028
rect 578234 219896 578854 231964
rect 578234 219660 578266 219896
rect 578502 219660 578586 219896
rect 578822 219660 578854 219896
rect 578234 219576 578854 219660
rect 578234 219340 578266 219576
rect 578502 219340 578586 219576
rect 578822 219340 578854 219576
rect 578234 183896 578854 219340
rect 578234 183660 578266 183896
rect 578502 183660 578586 183896
rect 578822 183660 578854 183896
rect 578234 183576 578854 183660
rect 578234 183340 578266 183576
rect 578502 183340 578586 183576
rect 578822 183340 578854 183576
rect 578234 147896 578854 183340
rect 578234 147660 578266 147896
rect 578502 147660 578586 147896
rect 578822 147660 578854 147896
rect 578234 147576 578854 147660
rect 578234 147340 578266 147576
rect 578502 147340 578586 147576
rect 578822 147340 578854 147576
rect 578234 111896 578854 147340
rect 578234 111660 578266 111896
rect 578502 111660 578586 111896
rect 578822 111660 578854 111896
rect 578234 111576 578854 111660
rect 578234 111340 578266 111576
rect 578502 111340 578586 111576
rect 578822 111340 578854 111576
rect 578234 75896 578854 111340
rect 578234 75660 578266 75896
rect 578502 75660 578586 75896
rect 578822 75660 578854 75896
rect 578234 75576 578854 75660
rect 578234 75340 578266 75576
rect 578502 75340 578586 75576
rect 578822 75340 578854 75576
rect 578234 39896 578854 75340
rect 578234 39660 578266 39896
rect 578502 39660 578586 39896
rect 578822 39660 578854 39896
rect 578234 39576 578854 39660
rect 578234 39340 578266 39576
rect 578502 39340 578586 39576
rect 578822 39340 578854 39576
rect 578234 3896 578854 39340
rect 578234 3660 578266 3896
rect 578502 3660 578586 3896
rect 578822 3660 578854 3896
rect 578234 3576 578854 3660
rect 578234 3340 578266 3576
rect 578502 3340 578586 3576
rect 578822 3340 578854 3576
rect 578234 -1304 578854 3340
rect 578234 -1540 578266 -1304
rect 578502 -1540 578586 -1304
rect 578822 -1540 578854 -1304
rect 578234 -1624 578854 -1540
rect 578234 -1860 578266 -1624
rect 578502 -1860 578586 -1624
rect 578822 -1860 578854 -1624
rect 578234 -7652 578854 -1860
rect 579474 706760 580094 711592
rect 579474 706524 579506 706760
rect 579742 706524 579826 706760
rect 580062 706524 580094 706760
rect 579474 706440 580094 706524
rect 579474 706204 579506 706440
rect 579742 706204 579826 706440
rect 580062 706204 580094 706440
rect 579474 689136 580094 706204
rect 579474 688900 579506 689136
rect 579742 688900 579826 689136
rect 580062 688900 580094 689136
rect 579474 688816 580094 688900
rect 579474 688580 579506 688816
rect 579742 688580 579826 688816
rect 580062 688580 580094 688816
rect 579474 653136 580094 688580
rect 579474 652900 579506 653136
rect 579742 652900 579826 653136
rect 580062 652900 580094 653136
rect 579474 652816 580094 652900
rect 579474 652580 579506 652816
rect 579742 652580 579826 652816
rect 580062 652580 580094 652816
rect 579474 617136 580094 652580
rect 579474 616900 579506 617136
rect 579742 616900 579826 617136
rect 580062 616900 580094 617136
rect 579474 616816 580094 616900
rect 579474 616580 579506 616816
rect 579742 616580 579826 616816
rect 580062 616580 580094 616816
rect 579474 581136 580094 616580
rect 579474 580900 579506 581136
rect 579742 580900 579826 581136
rect 580062 580900 580094 581136
rect 579474 580816 580094 580900
rect 579474 580580 579506 580816
rect 579742 580580 579826 580816
rect 580062 580580 580094 580816
rect 579474 545136 580094 580580
rect 579474 544900 579506 545136
rect 579742 544900 579826 545136
rect 580062 544900 580094 545136
rect 579474 544816 580094 544900
rect 579474 544580 579506 544816
rect 579742 544580 579826 544816
rect 580062 544580 580094 544816
rect 579474 509136 580094 544580
rect 579474 508900 579506 509136
rect 579742 508900 579826 509136
rect 580062 508900 580094 509136
rect 579474 508816 580094 508900
rect 579474 508580 579506 508816
rect 579742 508580 579826 508816
rect 580062 508580 580094 508816
rect 579474 473136 580094 508580
rect 579474 472900 579506 473136
rect 579742 472900 579826 473136
rect 580062 472900 580094 473136
rect 579474 472816 580094 472900
rect 579474 472580 579506 472816
rect 579742 472580 579826 472816
rect 580062 472580 580094 472816
rect 579474 437136 580094 472580
rect 579474 436900 579506 437136
rect 579742 436900 579826 437136
rect 580062 436900 580094 437136
rect 579474 436816 580094 436900
rect 579474 436580 579506 436816
rect 579742 436580 579826 436816
rect 580062 436580 580094 436816
rect 579474 401136 580094 436580
rect 579474 400900 579506 401136
rect 579742 400900 579826 401136
rect 580062 400900 580094 401136
rect 579474 400816 580094 400900
rect 579474 400580 579506 400816
rect 579742 400580 579826 400816
rect 580062 400580 580094 400816
rect 579474 365136 580094 400580
rect 579474 364900 579506 365136
rect 579742 364900 579826 365136
rect 580062 364900 580094 365136
rect 579474 364816 580094 364900
rect 579474 364580 579506 364816
rect 579742 364580 579826 364816
rect 580062 364580 580094 364816
rect 579474 329136 580094 364580
rect 579474 328900 579506 329136
rect 579742 328900 579826 329136
rect 580062 328900 580094 329136
rect 579474 328816 580094 328900
rect 579474 328580 579506 328816
rect 579742 328580 579826 328816
rect 580062 328580 580094 328816
rect 579474 293136 580094 328580
rect 579474 292900 579506 293136
rect 579742 292900 579826 293136
rect 580062 292900 580094 293136
rect 579474 292816 580094 292900
rect 579474 292580 579506 292816
rect 579742 292580 579826 292816
rect 580062 292580 580094 292816
rect 579474 257136 580094 292580
rect 579474 256900 579506 257136
rect 579742 256900 579826 257136
rect 580062 256900 580094 257136
rect 579474 256816 580094 256900
rect 579474 256580 579506 256816
rect 579742 256580 579826 256816
rect 580062 256580 580094 256816
rect 579474 221136 580094 256580
rect 579474 220900 579506 221136
rect 579742 220900 579826 221136
rect 580062 220900 580094 221136
rect 579474 220816 580094 220900
rect 579474 220580 579506 220816
rect 579742 220580 579826 220816
rect 580062 220580 580094 220816
rect 579474 185136 580094 220580
rect 579474 184900 579506 185136
rect 579742 184900 579826 185136
rect 580062 184900 580094 185136
rect 579474 184816 580094 184900
rect 579474 184580 579506 184816
rect 579742 184580 579826 184816
rect 580062 184580 580094 184816
rect 579474 149136 580094 184580
rect 579474 148900 579506 149136
rect 579742 148900 579826 149136
rect 580062 148900 580094 149136
rect 579474 148816 580094 148900
rect 579474 148580 579506 148816
rect 579742 148580 579826 148816
rect 580062 148580 580094 148816
rect 579474 113136 580094 148580
rect 579474 112900 579506 113136
rect 579742 112900 579826 113136
rect 580062 112900 580094 113136
rect 579474 112816 580094 112900
rect 579474 112580 579506 112816
rect 579742 112580 579826 112816
rect 580062 112580 580094 112816
rect 579474 77136 580094 112580
rect 579474 76900 579506 77136
rect 579742 76900 579826 77136
rect 580062 76900 580094 77136
rect 579474 76816 580094 76900
rect 579474 76580 579506 76816
rect 579742 76580 579826 76816
rect 580062 76580 580094 76816
rect 579474 41136 580094 76580
rect 579474 40900 579506 41136
rect 579742 40900 579826 41136
rect 580062 40900 580094 41136
rect 579474 40816 580094 40900
rect 579474 40580 579506 40816
rect 579742 40580 579826 40816
rect 580062 40580 580094 40816
rect 579474 5136 580094 40580
rect 579474 4900 579506 5136
rect 579742 4900 579826 5136
rect 580062 4900 580094 5136
rect 579474 4816 580094 4900
rect 579474 4580 579506 4816
rect 579742 4580 579826 4816
rect 580062 4580 580094 4816
rect 579474 -2264 580094 4580
rect 579474 -2500 579506 -2264
rect 579742 -2500 579826 -2264
rect 580062 -2500 580094 -2264
rect 579474 -2584 580094 -2500
rect 579474 -2820 579506 -2584
rect 579742 -2820 579826 -2584
rect 580062 -2820 580094 -2584
rect 579474 -7652 580094 -2820
rect 580714 707720 581334 711592
rect 580714 707484 580746 707720
rect 580982 707484 581066 707720
rect 581302 707484 581334 707720
rect 580714 707400 581334 707484
rect 580714 707164 580746 707400
rect 580982 707164 581066 707400
rect 581302 707164 581334 707400
rect 580714 690376 581334 707164
rect 580714 690140 580746 690376
rect 580982 690140 581066 690376
rect 581302 690140 581334 690376
rect 580714 690056 581334 690140
rect 580714 689820 580746 690056
rect 580982 689820 581066 690056
rect 581302 689820 581334 690056
rect 580714 654376 581334 689820
rect 580714 654140 580746 654376
rect 580982 654140 581066 654376
rect 581302 654140 581334 654376
rect 580714 654056 581334 654140
rect 580714 653820 580746 654056
rect 580982 653820 581066 654056
rect 581302 653820 581334 654056
rect 580714 618376 581334 653820
rect 580714 618140 580746 618376
rect 580982 618140 581066 618376
rect 581302 618140 581334 618376
rect 580714 618056 581334 618140
rect 580714 617820 580746 618056
rect 580982 617820 581066 618056
rect 581302 617820 581334 618056
rect 580714 582376 581334 617820
rect 580714 582140 580746 582376
rect 580982 582140 581066 582376
rect 581302 582140 581334 582376
rect 580714 582056 581334 582140
rect 580714 581820 580746 582056
rect 580982 581820 581066 582056
rect 581302 581820 581334 582056
rect 580714 546376 581334 581820
rect 580714 546140 580746 546376
rect 580982 546140 581066 546376
rect 581302 546140 581334 546376
rect 580714 546056 581334 546140
rect 580714 545820 580746 546056
rect 580982 545820 581066 546056
rect 581302 545820 581334 546056
rect 580714 510376 581334 545820
rect 580714 510140 580746 510376
rect 580982 510140 581066 510376
rect 581302 510140 581334 510376
rect 580714 510056 581334 510140
rect 580714 509820 580746 510056
rect 580982 509820 581066 510056
rect 581302 509820 581334 510056
rect 580714 474376 581334 509820
rect 580714 474140 580746 474376
rect 580982 474140 581066 474376
rect 581302 474140 581334 474376
rect 580714 474056 581334 474140
rect 580714 473820 580746 474056
rect 580982 473820 581066 474056
rect 581302 473820 581334 474056
rect 580714 438376 581334 473820
rect 580714 438140 580746 438376
rect 580982 438140 581066 438376
rect 581302 438140 581334 438376
rect 580714 438056 581334 438140
rect 580714 437820 580746 438056
rect 580982 437820 581066 438056
rect 581302 437820 581334 438056
rect 580714 402376 581334 437820
rect 580714 402140 580746 402376
rect 580982 402140 581066 402376
rect 581302 402140 581334 402376
rect 580714 402056 581334 402140
rect 580714 401820 580746 402056
rect 580982 401820 581066 402056
rect 581302 401820 581334 402056
rect 580714 366376 581334 401820
rect 580714 366140 580746 366376
rect 580982 366140 581066 366376
rect 581302 366140 581334 366376
rect 580714 366056 581334 366140
rect 580714 365820 580746 366056
rect 580982 365820 581066 366056
rect 581302 365820 581334 366056
rect 580714 330376 581334 365820
rect 580714 330140 580746 330376
rect 580982 330140 581066 330376
rect 581302 330140 581334 330376
rect 580714 330056 581334 330140
rect 580714 329820 580746 330056
rect 580982 329820 581066 330056
rect 581302 329820 581334 330056
rect 580714 294376 581334 329820
rect 580714 294140 580746 294376
rect 580982 294140 581066 294376
rect 581302 294140 581334 294376
rect 580714 294056 581334 294140
rect 580714 293820 580746 294056
rect 580982 293820 581066 294056
rect 581302 293820 581334 294056
rect 580714 258376 581334 293820
rect 580714 258140 580746 258376
rect 580982 258140 581066 258376
rect 581302 258140 581334 258376
rect 580714 258056 581334 258140
rect 580714 257820 580746 258056
rect 580982 257820 581066 258056
rect 581302 257820 581334 258056
rect 580714 222376 581334 257820
rect 580714 222140 580746 222376
rect 580982 222140 581066 222376
rect 581302 222140 581334 222376
rect 580714 222056 581334 222140
rect 580714 221820 580746 222056
rect 580982 221820 581066 222056
rect 581302 221820 581334 222056
rect 580714 186376 581334 221820
rect 580714 186140 580746 186376
rect 580982 186140 581066 186376
rect 581302 186140 581334 186376
rect 580714 186056 581334 186140
rect 580714 185820 580746 186056
rect 580982 185820 581066 186056
rect 581302 185820 581334 186056
rect 580714 150376 581334 185820
rect 580714 150140 580746 150376
rect 580982 150140 581066 150376
rect 581302 150140 581334 150376
rect 580714 150056 581334 150140
rect 580714 149820 580746 150056
rect 580982 149820 581066 150056
rect 581302 149820 581334 150056
rect 580714 114376 581334 149820
rect 580714 114140 580746 114376
rect 580982 114140 581066 114376
rect 581302 114140 581334 114376
rect 580714 114056 581334 114140
rect 580714 113820 580746 114056
rect 580982 113820 581066 114056
rect 581302 113820 581334 114056
rect 580714 78376 581334 113820
rect 580714 78140 580746 78376
rect 580982 78140 581066 78376
rect 581302 78140 581334 78376
rect 580714 78056 581334 78140
rect 580714 77820 580746 78056
rect 580982 77820 581066 78056
rect 581302 77820 581334 78056
rect 580714 42376 581334 77820
rect 580714 42140 580746 42376
rect 580982 42140 581066 42376
rect 581302 42140 581334 42376
rect 580714 42056 581334 42140
rect 580714 41820 580746 42056
rect 580982 41820 581066 42056
rect 581302 41820 581334 42056
rect 580714 6376 581334 41820
rect 580714 6140 580746 6376
rect 580982 6140 581066 6376
rect 581302 6140 581334 6376
rect 580714 6056 581334 6140
rect 580714 5820 580746 6056
rect 580982 5820 581066 6056
rect 581302 5820 581334 6056
rect 580714 -3224 581334 5820
rect 580714 -3460 580746 -3224
rect 580982 -3460 581066 -3224
rect 581302 -3460 581334 -3224
rect 580714 -3544 581334 -3460
rect 580714 -3780 580746 -3544
rect 580982 -3780 581066 -3544
rect 581302 -3780 581334 -3544
rect 580714 -7652 581334 -3780
rect 581954 708680 582574 711592
rect 592030 711560 592650 711592
rect 592030 711324 592062 711560
rect 592298 711324 592382 711560
rect 592618 711324 592650 711560
rect 592030 711240 592650 711324
rect 592030 711004 592062 711240
rect 592298 711004 592382 711240
rect 592618 711004 592650 711240
rect 591070 710600 591690 710632
rect 591070 710364 591102 710600
rect 591338 710364 591422 710600
rect 591658 710364 591690 710600
rect 591070 710280 591690 710364
rect 591070 710044 591102 710280
rect 591338 710044 591422 710280
rect 591658 710044 591690 710280
rect 590110 709640 590730 709672
rect 590110 709404 590142 709640
rect 590378 709404 590462 709640
rect 590698 709404 590730 709640
rect 590110 709320 590730 709404
rect 590110 709084 590142 709320
rect 590378 709084 590462 709320
rect 590698 709084 590730 709320
rect 581954 708444 581986 708680
rect 582222 708444 582306 708680
rect 582542 708444 582574 708680
rect 581954 708360 582574 708444
rect 581954 708124 581986 708360
rect 582222 708124 582306 708360
rect 582542 708124 582574 708360
rect 581954 691616 582574 708124
rect 589150 708680 589770 708712
rect 589150 708444 589182 708680
rect 589418 708444 589502 708680
rect 589738 708444 589770 708680
rect 589150 708360 589770 708444
rect 589150 708124 589182 708360
rect 589418 708124 589502 708360
rect 589738 708124 589770 708360
rect 588190 707720 588810 707752
rect 588190 707484 588222 707720
rect 588458 707484 588542 707720
rect 588778 707484 588810 707720
rect 588190 707400 588810 707484
rect 588190 707164 588222 707400
rect 588458 707164 588542 707400
rect 588778 707164 588810 707400
rect 587230 706760 587850 706792
rect 587230 706524 587262 706760
rect 587498 706524 587582 706760
rect 587818 706524 587850 706760
rect 587230 706440 587850 706524
rect 587230 706204 587262 706440
rect 587498 706204 587582 706440
rect 587818 706204 587850 706440
rect 586270 705800 586890 705832
rect 586270 705564 586302 705800
rect 586538 705564 586622 705800
rect 586858 705564 586890 705800
rect 586270 705480 586890 705564
rect 586270 705244 586302 705480
rect 586538 705244 586622 705480
rect 586858 705244 586890 705480
rect 581954 691380 581986 691616
rect 582222 691380 582306 691616
rect 582542 691380 582574 691616
rect 581954 691296 582574 691380
rect 581954 691060 581986 691296
rect 582222 691060 582306 691296
rect 582542 691060 582574 691296
rect 581954 655616 582574 691060
rect 581954 655380 581986 655616
rect 582222 655380 582306 655616
rect 582542 655380 582574 655616
rect 581954 655296 582574 655380
rect 581954 655060 581986 655296
rect 582222 655060 582306 655296
rect 582542 655060 582574 655296
rect 581954 619616 582574 655060
rect 581954 619380 581986 619616
rect 582222 619380 582306 619616
rect 582542 619380 582574 619616
rect 581954 619296 582574 619380
rect 581954 619060 581986 619296
rect 582222 619060 582306 619296
rect 582542 619060 582574 619296
rect 581954 583616 582574 619060
rect 581954 583380 581986 583616
rect 582222 583380 582306 583616
rect 582542 583380 582574 583616
rect 581954 583296 582574 583380
rect 581954 583060 581986 583296
rect 582222 583060 582306 583296
rect 582542 583060 582574 583296
rect 581954 547616 582574 583060
rect 581954 547380 581986 547616
rect 582222 547380 582306 547616
rect 582542 547380 582574 547616
rect 581954 547296 582574 547380
rect 581954 547060 581986 547296
rect 582222 547060 582306 547296
rect 582542 547060 582574 547296
rect 581954 511616 582574 547060
rect 581954 511380 581986 511616
rect 582222 511380 582306 511616
rect 582542 511380 582574 511616
rect 581954 511296 582574 511380
rect 581954 511060 581986 511296
rect 582222 511060 582306 511296
rect 582542 511060 582574 511296
rect 581954 475616 582574 511060
rect 581954 475380 581986 475616
rect 582222 475380 582306 475616
rect 582542 475380 582574 475616
rect 581954 475296 582574 475380
rect 581954 475060 581986 475296
rect 582222 475060 582306 475296
rect 582542 475060 582574 475296
rect 581954 439616 582574 475060
rect 581954 439380 581986 439616
rect 582222 439380 582306 439616
rect 582542 439380 582574 439616
rect 581954 439296 582574 439380
rect 581954 439060 581986 439296
rect 582222 439060 582306 439296
rect 582542 439060 582574 439296
rect 581954 403616 582574 439060
rect 581954 403380 581986 403616
rect 582222 403380 582306 403616
rect 582542 403380 582574 403616
rect 581954 403296 582574 403380
rect 581954 403060 581986 403296
rect 582222 403060 582306 403296
rect 582542 403060 582574 403296
rect 581954 367616 582574 403060
rect 581954 367380 581986 367616
rect 582222 367380 582306 367616
rect 582542 367380 582574 367616
rect 581954 367296 582574 367380
rect 581954 367060 581986 367296
rect 582222 367060 582306 367296
rect 582542 367060 582574 367296
rect 581954 331616 582574 367060
rect 581954 331380 581986 331616
rect 582222 331380 582306 331616
rect 582542 331380 582574 331616
rect 581954 331296 582574 331380
rect 581954 331060 581986 331296
rect 582222 331060 582306 331296
rect 582542 331060 582574 331296
rect 581954 295616 582574 331060
rect 581954 295380 581986 295616
rect 582222 295380 582306 295616
rect 582542 295380 582574 295616
rect 581954 295296 582574 295380
rect 581954 295060 581986 295296
rect 582222 295060 582306 295296
rect 582542 295060 582574 295296
rect 581954 259616 582574 295060
rect 581954 259380 581986 259616
rect 582222 259380 582306 259616
rect 582542 259380 582574 259616
rect 581954 259296 582574 259380
rect 581954 259060 581986 259296
rect 582222 259060 582306 259296
rect 582542 259060 582574 259296
rect 581954 223616 582574 259060
rect 581954 223380 581986 223616
rect 582222 223380 582306 223616
rect 582542 223380 582574 223616
rect 581954 223296 582574 223380
rect 581954 223060 581986 223296
rect 582222 223060 582306 223296
rect 582542 223060 582574 223296
rect 581954 187616 582574 223060
rect 581954 187380 581986 187616
rect 582222 187380 582306 187616
rect 582542 187380 582574 187616
rect 581954 187296 582574 187380
rect 581954 187060 581986 187296
rect 582222 187060 582306 187296
rect 582542 187060 582574 187296
rect 581954 151616 582574 187060
rect 581954 151380 581986 151616
rect 582222 151380 582306 151616
rect 582542 151380 582574 151616
rect 581954 151296 582574 151380
rect 581954 151060 581986 151296
rect 582222 151060 582306 151296
rect 582542 151060 582574 151296
rect 581954 115616 582574 151060
rect 581954 115380 581986 115616
rect 582222 115380 582306 115616
rect 582542 115380 582574 115616
rect 581954 115296 582574 115380
rect 581954 115060 581986 115296
rect 582222 115060 582306 115296
rect 582542 115060 582574 115296
rect 581954 79616 582574 115060
rect 581954 79380 581986 79616
rect 582222 79380 582306 79616
rect 582542 79380 582574 79616
rect 581954 79296 582574 79380
rect 581954 79060 581986 79296
rect 582222 79060 582306 79296
rect 582542 79060 582574 79296
rect 581954 43616 582574 79060
rect 581954 43380 581986 43616
rect 582222 43380 582306 43616
rect 582542 43380 582574 43616
rect 581954 43296 582574 43380
rect 581954 43060 581986 43296
rect 582222 43060 582306 43296
rect 582542 43060 582574 43296
rect 581954 7616 582574 43060
rect 581954 7380 581986 7616
rect 582222 7380 582306 7616
rect 582542 7380 582574 7616
rect 581954 7296 582574 7380
rect 581954 7060 581986 7296
rect 582222 7060 582306 7296
rect 582542 7060 582574 7296
rect 581954 -4184 582574 7060
rect 585310 704840 585930 704872
rect 585310 704604 585342 704840
rect 585578 704604 585662 704840
rect 585898 704604 585930 704840
rect 585310 704520 585930 704604
rect 585310 704284 585342 704520
rect 585578 704284 585662 704520
rect 585898 704284 585930 704520
rect 585310 686656 585930 704284
rect 585310 686420 585342 686656
rect 585578 686420 585662 686656
rect 585898 686420 585930 686656
rect 585310 686336 585930 686420
rect 585310 686100 585342 686336
rect 585578 686100 585662 686336
rect 585898 686100 585930 686336
rect 585310 650656 585930 686100
rect 585310 650420 585342 650656
rect 585578 650420 585662 650656
rect 585898 650420 585930 650656
rect 585310 650336 585930 650420
rect 585310 650100 585342 650336
rect 585578 650100 585662 650336
rect 585898 650100 585930 650336
rect 585310 614656 585930 650100
rect 585310 614420 585342 614656
rect 585578 614420 585662 614656
rect 585898 614420 585930 614656
rect 585310 614336 585930 614420
rect 585310 614100 585342 614336
rect 585578 614100 585662 614336
rect 585898 614100 585930 614336
rect 585310 578656 585930 614100
rect 585310 578420 585342 578656
rect 585578 578420 585662 578656
rect 585898 578420 585930 578656
rect 585310 578336 585930 578420
rect 585310 578100 585342 578336
rect 585578 578100 585662 578336
rect 585898 578100 585930 578336
rect 585310 542656 585930 578100
rect 585310 542420 585342 542656
rect 585578 542420 585662 542656
rect 585898 542420 585930 542656
rect 585310 542336 585930 542420
rect 585310 542100 585342 542336
rect 585578 542100 585662 542336
rect 585898 542100 585930 542336
rect 585310 506656 585930 542100
rect 585310 506420 585342 506656
rect 585578 506420 585662 506656
rect 585898 506420 585930 506656
rect 585310 506336 585930 506420
rect 585310 506100 585342 506336
rect 585578 506100 585662 506336
rect 585898 506100 585930 506336
rect 585310 470656 585930 506100
rect 585310 470420 585342 470656
rect 585578 470420 585662 470656
rect 585898 470420 585930 470656
rect 585310 470336 585930 470420
rect 585310 470100 585342 470336
rect 585578 470100 585662 470336
rect 585898 470100 585930 470336
rect 585310 434656 585930 470100
rect 585310 434420 585342 434656
rect 585578 434420 585662 434656
rect 585898 434420 585930 434656
rect 585310 434336 585930 434420
rect 585310 434100 585342 434336
rect 585578 434100 585662 434336
rect 585898 434100 585930 434336
rect 585310 398656 585930 434100
rect 585310 398420 585342 398656
rect 585578 398420 585662 398656
rect 585898 398420 585930 398656
rect 585310 398336 585930 398420
rect 585310 398100 585342 398336
rect 585578 398100 585662 398336
rect 585898 398100 585930 398336
rect 585310 362656 585930 398100
rect 585310 362420 585342 362656
rect 585578 362420 585662 362656
rect 585898 362420 585930 362656
rect 585310 362336 585930 362420
rect 585310 362100 585342 362336
rect 585578 362100 585662 362336
rect 585898 362100 585930 362336
rect 585310 326656 585930 362100
rect 585310 326420 585342 326656
rect 585578 326420 585662 326656
rect 585898 326420 585930 326656
rect 585310 326336 585930 326420
rect 585310 326100 585342 326336
rect 585578 326100 585662 326336
rect 585898 326100 585930 326336
rect 585310 290656 585930 326100
rect 585310 290420 585342 290656
rect 585578 290420 585662 290656
rect 585898 290420 585930 290656
rect 585310 290336 585930 290420
rect 585310 290100 585342 290336
rect 585578 290100 585662 290336
rect 585898 290100 585930 290336
rect 585310 254656 585930 290100
rect 585310 254420 585342 254656
rect 585578 254420 585662 254656
rect 585898 254420 585930 254656
rect 585310 254336 585930 254420
rect 585310 254100 585342 254336
rect 585578 254100 585662 254336
rect 585898 254100 585930 254336
rect 585310 218656 585930 254100
rect 585310 218420 585342 218656
rect 585578 218420 585662 218656
rect 585898 218420 585930 218656
rect 585310 218336 585930 218420
rect 585310 218100 585342 218336
rect 585578 218100 585662 218336
rect 585898 218100 585930 218336
rect 585310 182656 585930 218100
rect 585310 182420 585342 182656
rect 585578 182420 585662 182656
rect 585898 182420 585930 182656
rect 585310 182336 585930 182420
rect 585310 182100 585342 182336
rect 585578 182100 585662 182336
rect 585898 182100 585930 182336
rect 585310 146656 585930 182100
rect 585310 146420 585342 146656
rect 585578 146420 585662 146656
rect 585898 146420 585930 146656
rect 585310 146336 585930 146420
rect 585310 146100 585342 146336
rect 585578 146100 585662 146336
rect 585898 146100 585930 146336
rect 585310 110656 585930 146100
rect 585310 110420 585342 110656
rect 585578 110420 585662 110656
rect 585898 110420 585930 110656
rect 585310 110336 585930 110420
rect 585310 110100 585342 110336
rect 585578 110100 585662 110336
rect 585898 110100 585930 110336
rect 585310 74656 585930 110100
rect 585310 74420 585342 74656
rect 585578 74420 585662 74656
rect 585898 74420 585930 74656
rect 585310 74336 585930 74420
rect 585310 74100 585342 74336
rect 585578 74100 585662 74336
rect 585898 74100 585930 74336
rect 585310 38656 585930 74100
rect 585310 38420 585342 38656
rect 585578 38420 585662 38656
rect 585898 38420 585930 38656
rect 585310 38336 585930 38420
rect 585310 38100 585342 38336
rect 585578 38100 585662 38336
rect 585898 38100 585930 38336
rect 585310 2656 585930 38100
rect 585310 2420 585342 2656
rect 585578 2420 585662 2656
rect 585898 2420 585930 2656
rect 585310 2336 585930 2420
rect 585310 2100 585342 2336
rect 585578 2100 585662 2336
rect 585898 2100 585930 2336
rect 585310 -344 585930 2100
rect 585310 -580 585342 -344
rect 585578 -580 585662 -344
rect 585898 -580 585930 -344
rect 585310 -664 585930 -580
rect 585310 -900 585342 -664
rect 585578 -900 585662 -664
rect 585898 -900 585930 -664
rect 585310 -932 585930 -900
rect 586270 687896 586890 705244
rect 586270 687660 586302 687896
rect 586538 687660 586622 687896
rect 586858 687660 586890 687896
rect 586270 687576 586890 687660
rect 586270 687340 586302 687576
rect 586538 687340 586622 687576
rect 586858 687340 586890 687576
rect 586270 651896 586890 687340
rect 586270 651660 586302 651896
rect 586538 651660 586622 651896
rect 586858 651660 586890 651896
rect 586270 651576 586890 651660
rect 586270 651340 586302 651576
rect 586538 651340 586622 651576
rect 586858 651340 586890 651576
rect 586270 615896 586890 651340
rect 586270 615660 586302 615896
rect 586538 615660 586622 615896
rect 586858 615660 586890 615896
rect 586270 615576 586890 615660
rect 586270 615340 586302 615576
rect 586538 615340 586622 615576
rect 586858 615340 586890 615576
rect 586270 579896 586890 615340
rect 586270 579660 586302 579896
rect 586538 579660 586622 579896
rect 586858 579660 586890 579896
rect 586270 579576 586890 579660
rect 586270 579340 586302 579576
rect 586538 579340 586622 579576
rect 586858 579340 586890 579576
rect 586270 543896 586890 579340
rect 586270 543660 586302 543896
rect 586538 543660 586622 543896
rect 586858 543660 586890 543896
rect 586270 543576 586890 543660
rect 586270 543340 586302 543576
rect 586538 543340 586622 543576
rect 586858 543340 586890 543576
rect 586270 507896 586890 543340
rect 586270 507660 586302 507896
rect 586538 507660 586622 507896
rect 586858 507660 586890 507896
rect 586270 507576 586890 507660
rect 586270 507340 586302 507576
rect 586538 507340 586622 507576
rect 586858 507340 586890 507576
rect 586270 471896 586890 507340
rect 586270 471660 586302 471896
rect 586538 471660 586622 471896
rect 586858 471660 586890 471896
rect 586270 471576 586890 471660
rect 586270 471340 586302 471576
rect 586538 471340 586622 471576
rect 586858 471340 586890 471576
rect 586270 435896 586890 471340
rect 586270 435660 586302 435896
rect 586538 435660 586622 435896
rect 586858 435660 586890 435896
rect 586270 435576 586890 435660
rect 586270 435340 586302 435576
rect 586538 435340 586622 435576
rect 586858 435340 586890 435576
rect 586270 399896 586890 435340
rect 586270 399660 586302 399896
rect 586538 399660 586622 399896
rect 586858 399660 586890 399896
rect 586270 399576 586890 399660
rect 586270 399340 586302 399576
rect 586538 399340 586622 399576
rect 586858 399340 586890 399576
rect 586270 363896 586890 399340
rect 586270 363660 586302 363896
rect 586538 363660 586622 363896
rect 586858 363660 586890 363896
rect 586270 363576 586890 363660
rect 586270 363340 586302 363576
rect 586538 363340 586622 363576
rect 586858 363340 586890 363576
rect 586270 327896 586890 363340
rect 586270 327660 586302 327896
rect 586538 327660 586622 327896
rect 586858 327660 586890 327896
rect 586270 327576 586890 327660
rect 586270 327340 586302 327576
rect 586538 327340 586622 327576
rect 586858 327340 586890 327576
rect 586270 291896 586890 327340
rect 586270 291660 586302 291896
rect 586538 291660 586622 291896
rect 586858 291660 586890 291896
rect 586270 291576 586890 291660
rect 586270 291340 586302 291576
rect 586538 291340 586622 291576
rect 586858 291340 586890 291576
rect 586270 255896 586890 291340
rect 586270 255660 586302 255896
rect 586538 255660 586622 255896
rect 586858 255660 586890 255896
rect 586270 255576 586890 255660
rect 586270 255340 586302 255576
rect 586538 255340 586622 255576
rect 586858 255340 586890 255576
rect 586270 219896 586890 255340
rect 586270 219660 586302 219896
rect 586538 219660 586622 219896
rect 586858 219660 586890 219896
rect 586270 219576 586890 219660
rect 586270 219340 586302 219576
rect 586538 219340 586622 219576
rect 586858 219340 586890 219576
rect 586270 183896 586890 219340
rect 586270 183660 586302 183896
rect 586538 183660 586622 183896
rect 586858 183660 586890 183896
rect 586270 183576 586890 183660
rect 586270 183340 586302 183576
rect 586538 183340 586622 183576
rect 586858 183340 586890 183576
rect 586270 147896 586890 183340
rect 586270 147660 586302 147896
rect 586538 147660 586622 147896
rect 586858 147660 586890 147896
rect 586270 147576 586890 147660
rect 586270 147340 586302 147576
rect 586538 147340 586622 147576
rect 586858 147340 586890 147576
rect 586270 111896 586890 147340
rect 586270 111660 586302 111896
rect 586538 111660 586622 111896
rect 586858 111660 586890 111896
rect 586270 111576 586890 111660
rect 586270 111340 586302 111576
rect 586538 111340 586622 111576
rect 586858 111340 586890 111576
rect 586270 75896 586890 111340
rect 586270 75660 586302 75896
rect 586538 75660 586622 75896
rect 586858 75660 586890 75896
rect 586270 75576 586890 75660
rect 586270 75340 586302 75576
rect 586538 75340 586622 75576
rect 586858 75340 586890 75576
rect 586270 39896 586890 75340
rect 586270 39660 586302 39896
rect 586538 39660 586622 39896
rect 586858 39660 586890 39896
rect 586270 39576 586890 39660
rect 586270 39340 586302 39576
rect 586538 39340 586622 39576
rect 586858 39340 586890 39576
rect 586270 3896 586890 39340
rect 586270 3660 586302 3896
rect 586538 3660 586622 3896
rect 586858 3660 586890 3896
rect 586270 3576 586890 3660
rect 586270 3340 586302 3576
rect 586538 3340 586622 3576
rect 586858 3340 586890 3576
rect 586270 -1304 586890 3340
rect 586270 -1540 586302 -1304
rect 586538 -1540 586622 -1304
rect 586858 -1540 586890 -1304
rect 586270 -1624 586890 -1540
rect 586270 -1860 586302 -1624
rect 586538 -1860 586622 -1624
rect 586858 -1860 586890 -1624
rect 586270 -1892 586890 -1860
rect 587230 689136 587850 706204
rect 587230 688900 587262 689136
rect 587498 688900 587582 689136
rect 587818 688900 587850 689136
rect 587230 688816 587850 688900
rect 587230 688580 587262 688816
rect 587498 688580 587582 688816
rect 587818 688580 587850 688816
rect 587230 653136 587850 688580
rect 587230 652900 587262 653136
rect 587498 652900 587582 653136
rect 587818 652900 587850 653136
rect 587230 652816 587850 652900
rect 587230 652580 587262 652816
rect 587498 652580 587582 652816
rect 587818 652580 587850 652816
rect 587230 617136 587850 652580
rect 587230 616900 587262 617136
rect 587498 616900 587582 617136
rect 587818 616900 587850 617136
rect 587230 616816 587850 616900
rect 587230 616580 587262 616816
rect 587498 616580 587582 616816
rect 587818 616580 587850 616816
rect 587230 581136 587850 616580
rect 587230 580900 587262 581136
rect 587498 580900 587582 581136
rect 587818 580900 587850 581136
rect 587230 580816 587850 580900
rect 587230 580580 587262 580816
rect 587498 580580 587582 580816
rect 587818 580580 587850 580816
rect 587230 545136 587850 580580
rect 587230 544900 587262 545136
rect 587498 544900 587582 545136
rect 587818 544900 587850 545136
rect 587230 544816 587850 544900
rect 587230 544580 587262 544816
rect 587498 544580 587582 544816
rect 587818 544580 587850 544816
rect 587230 509136 587850 544580
rect 587230 508900 587262 509136
rect 587498 508900 587582 509136
rect 587818 508900 587850 509136
rect 587230 508816 587850 508900
rect 587230 508580 587262 508816
rect 587498 508580 587582 508816
rect 587818 508580 587850 508816
rect 587230 473136 587850 508580
rect 587230 472900 587262 473136
rect 587498 472900 587582 473136
rect 587818 472900 587850 473136
rect 587230 472816 587850 472900
rect 587230 472580 587262 472816
rect 587498 472580 587582 472816
rect 587818 472580 587850 472816
rect 587230 437136 587850 472580
rect 587230 436900 587262 437136
rect 587498 436900 587582 437136
rect 587818 436900 587850 437136
rect 587230 436816 587850 436900
rect 587230 436580 587262 436816
rect 587498 436580 587582 436816
rect 587818 436580 587850 436816
rect 587230 401136 587850 436580
rect 587230 400900 587262 401136
rect 587498 400900 587582 401136
rect 587818 400900 587850 401136
rect 587230 400816 587850 400900
rect 587230 400580 587262 400816
rect 587498 400580 587582 400816
rect 587818 400580 587850 400816
rect 587230 365136 587850 400580
rect 587230 364900 587262 365136
rect 587498 364900 587582 365136
rect 587818 364900 587850 365136
rect 587230 364816 587850 364900
rect 587230 364580 587262 364816
rect 587498 364580 587582 364816
rect 587818 364580 587850 364816
rect 587230 329136 587850 364580
rect 587230 328900 587262 329136
rect 587498 328900 587582 329136
rect 587818 328900 587850 329136
rect 587230 328816 587850 328900
rect 587230 328580 587262 328816
rect 587498 328580 587582 328816
rect 587818 328580 587850 328816
rect 587230 293136 587850 328580
rect 587230 292900 587262 293136
rect 587498 292900 587582 293136
rect 587818 292900 587850 293136
rect 587230 292816 587850 292900
rect 587230 292580 587262 292816
rect 587498 292580 587582 292816
rect 587818 292580 587850 292816
rect 587230 257136 587850 292580
rect 587230 256900 587262 257136
rect 587498 256900 587582 257136
rect 587818 256900 587850 257136
rect 587230 256816 587850 256900
rect 587230 256580 587262 256816
rect 587498 256580 587582 256816
rect 587818 256580 587850 256816
rect 587230 221136 587850 256580
rect 587230 220900 587262 221136
rect 587498 220900 587582 221136
rect 587818 220900 587850 221136
rect 587230 220816 587850 220900
rect 587230 220580 587262 220816
rect 587498 220580 587582 220816
rect 587818 220580 587850 220816
rect 587230 185136 587850 220580
rect 587230 184900 587262 185136
rect 587498 184900 587582 185136
rect 587818 184900 587850 185136
rect 587230 184816 587850 184900
rect 587230 184580 587262 184816
rect 587498 184580 587582 184816
rect 587818 184580 587850 184816
rect 587230 149136 587850 184580
rect 587230 148900 587262 149136
rect 587498 148900 587582 149136
rect 587818 148900 587850 149136
rect 587230 148816 587850 148900
rect 587230 148580 587262 148816
rect 587498 148580 587582 148816
rect 587818 148580 587850 148816
rect 587230 113136 587850 148580
rect 587230 112900 587262 113136
rect 587498 112900 587582 113136
rect 587818 112900 587850 113136
rect 587230 112816 587850 112900
rect 587230 112580 587262 112816
rect 587498 112580 587582 112816
rect 587818 112580 587850 112816
rect 587230 77136 587850 112580
rect 587230 76900 587262 77136
rect 587498 76900 587582 77136
rect 587818 76900 587850 77136
rect 587230 76816 587850 76900
rect 587230 76580 587262 76816
rect 587498 76580 587582 76816
rect 587818 76580 587850 76816
rect 587230 41136 587850 76580
rect 587230 40900 587262 41136
rect 587498 40900 587582 41136
rect 587818 40900 587850 41136
rect 587230 40816 587850 40900
rect 587230 40580 587262 40816
rect 587498 40580 587582 40816
rect 587818 40580 587850 40816
rect 587230 5136 587850 40580
rect 587230 4900 587262 5136
rect 587498 4900 587582 5136
rect 587818 4900 587850 5136
rect 587230 4816 587850 4900
rect 587230 4580 587262 4816
rect 587498 4580 587582 4816
rect 587818 4580 587850 4816
rect 587230 -2264 587850 4580
rect 587230 -2500 587262 -2264
rect 587498 -2500 587582 -2264
rect 587818 -2500 587850 -2264
rect 587230 -2584 587850 -2500
rect 587230 -2820 587262 -2584
rect 587498 -2820 587582 -2584
rect 587818 -2820 587850 -2584
rect 587230 -2852 587850 -2820
rect 588190 690376 588810 707164
rect 588190 690140 588222 690376
rect 588458 690140 588542 690376
rect 588778 690140 588810 690376
rect 588190 690056 588810 690140
rect 588190 689820 588222 690056
rect 588458 689820 588542 690056
rect 588778 689820 588810 690056
rect 588190 654376 588810 689820
rect 588190 654140 588222 654376
rect 588458 654140 588542 654376
rect 588778 654140 588810 654376
rect 588190 654056 588810 654140
rect 588190 653820 588222 654056
rect 588458 653820 588542 654056
rect 588778 653820 588810 654056
rect 588190 618376 588810 653820
rect 588190 618140 588222 618376
rect 588458 618140 588542 618376
rect 588778 618140 588810 618376
rect 588190 618056 588810 618140
rect 588190 617820 588222 618056
rect 588458 617820 588542 618056
rect 588778 617820 588810 618056
rect 588190 582376 588810 617820
rect 588190 582140 588222 582376
rect 588458 582140 588542 582376
rect 588778 582140 588810 582376
rect 588190 582056 588810 582140
rect 588190 581820 588222 582056
rect 588458 581820 588542 582056
rect 588778 581820 588810 582056
rect 588190 546376 588810 581820
rect 588190 546140 588222 546376
rect 588458 546140 588542 546376
rect 588778 546140 588810 546376
rect 588190 546056 588810 546140
rect 588190 545820 588222 546056
rect 588458 545820 588542 546056
rect 588778 545820 588810 546056
rect 588190 510376 588810 545820
rect 588190 510140 588222 510376
rect 588458 510140 588542 510376
rect 588778 510140 588810 510376
rect 588190 510056 588810 510140
rect 588190 509820 588222 510056
rect 588458 509820 588542 510056
rect 588778 509820 588810 510056
rect 588190 474376 588810 509820
rect 588190 474140 588222 474376
rect 588458 474140 588542 474376
rect 588778 474140 588810 474376
rect 588190 474056 588810 474140
rect 588190 473820 588222 474056
rect 588458 473820 588542 474056
rect 588778 473820 588810 474056
rect 588190 438376 588810 473820
rect 588190 438140 588222 438376
rect 588458 438140 588542 438376
rect 588778 438140 588810 438376
rect 588190 438056 588810 438140
rect 588190 437820 588222 438056
rect 588458 437820 588542 438056
rect 588778 437820 588810 438056
rect 588190 402376 588810 437820
rect 588190 402140 588222 402376
rect 588458 402140 588542 402376
rect 588778 402140 588810 402376
rect 588190 402056 588810 402140
rect 588190 401820 588222 402056
rect 588458 401820 588542 402056
rect 588778 401820 588810 402056
rect 588190 366376 588810 401820
rect 588190 366140 588222 366376
rect 588458 366140 588542 366376
rect 588778 366140 588810 366376
rect 588190 366056 588810 366140
rect 588190 365820 588222 366056
rect 588458 365820 588542 366056
rect 588778 365820 588810 366056
rect 588190 330376 588810 365820
rect 588190 330140 588222 330376
rect 588458 330140 588542 330376
rect 588778 330140 588810 330376
rect 588190 330056 588810 330140
rect 588190 329820 588222 330056
rect 588458 329820 588542 330056
rect 588778 329820 588810 330056
rect 588190 294376 588810 329820
rect 588190 294140 588222 294376
rect 588458 294140 588542 294376
rect 588778 294140 588810 294376
rect 588190 294056 588810 294140
rect 588190 293820 588222 294056
rect 588458 293820 588542 294056
rect 588778 293820 588810 294056
rect 588190 258376 588810 293820
rect 588190 258140 588222 258376
rect 588458 258140 588542 258376
rect 588778 258140 588810 258376
rect 588190 258056 588810 258140
rect 588190 257820 588222 258056
rect 588458 257820 588542 258056
rect 588778 257820 588810 258056
rect 588190 222376 588810 257820
rect 588190 222140 588222 222376
rect 588458 222140 588542 222376
rect 588778 222140 588810 222376
rect 588190 222056 588810 222140
rect 588190 221820 588222 222056
rect 588458 221820 588542 222056
rect 588778 221820 588810 222056
rect 588190 186376 588810 221820
rect 588190 186140 588222 186376
rect 588458 186140 588542 186376
rect 588778 186140 588810 186376
rect 588190 186056 588810 186140
rect 588190 185820 588222 186056
rect 588458 185820 588542 186056
rect 588778 185820 588810 186056
rect 588190 150376 588810 185820
rect 588190 150140 588222 150376
rect 588458 150140 588542 150376
rect 588778 150140 588810 150376
rect 588190 150056 588810 150140
rect 588190 149820 588222 150056
rect 588458 149820 588542 150056
rect 588778 149820 588810 150056
rect 588190 114376 588810 149820
rect 588190 114140 588222 114376
rect 588458 114140 588542 114376
rect 588778 114140 588810 114376
rect 588190 114056 588810 114140
rect 588190 113820 588222 114056
rect 588458 113820 588542 114056
rect 588778 113820 588810 114056
rect 588190 78376 588810 113820
rect 588190 78140 588222 78376
rect 588458 78140 588542 78376
rect 588778 78140 588810 78376
rect 588190 78056 588810 78140
rect 588190 77820 588222 78056
rect 588458 77820 588542 78056
rect 588778 77820 588810 78056
rect 588190 42376 588810 77820
rect 588190 42140 588222 42376
rect 588458 42140 588542 42376
rect 588778 42140 588810 42376
rect 588190 42056 588810 42140
rect 588190 41820 588222 42056
rect 588458 41820 588542 42056
rect 588778 41820 588810 42056
rect 588190 6376 588810 41820
rect 588190 6140 588222 6376
rect 588458 6140 588542 6376
rect 588778 6140 588810 6376
rect 588190 6056 588810 6140
rect 588190 5820 588222 6056
rect 588458 5820 588542 6056
rect 588778 5820 588810 6056
rect 588190 -3224 588810 5820
rect 588190 -3460 588222 -3224
rect 588458 -3460 588542 -3224
rect 588778 -3460 588810 -3224
rect 588190 -3544 588810 -3460
rect 588190 -3780 588222 -3544
rect 588458 -3780 588542 -3544
rect 588778 -3780 588810 -3544
rect 588190 -3812 588810 -3780
rect 589150 691616 589770 708124
rect 589150 691380 589182 691616
rect 589418 691380 589502 691616
rect 589738 691380 589770 691616
rect 589150 691296 589770 691380
rect 589150 691060 589182 691296
rect 589418 691060 589502 691296
rect 589738 691060 589770 691296
rect 589150 655616 589770 691060
rect 589150 655380 589182 655616
rect 589418 655380 589502 655616
rect 589738 655380 589770 655616
rect 589150 655296 589770 655380
rect 589150 655060 589182 655296
rect 589418 655060 589502 655296
rect 589738 655060 589770 655296
rect 589150 619616 589770 655060
rect 589150 619380 589182 619616
rect 589418 619380 589502 619616
rect 589738 619380 589770 619616
rect 589150 619296 589770 619380
rect 589150 619060 589182 619296
rect 589418 619060 589502 619296
rect 589738 619060 589770 619296
rect 589150 583616 589770 619060
rect 589150 583380 589182 583616
rect 589418 583380 589502 583616
rect 589738 583380 589770 583616
rect 589150 583296 589770 583380
rect 589150 583060 589182 583296
rect 589418 583060 589502 583296
rect 589738 583060 589770 583296
rect 589150 547616 589770 583060
rect 589150 547380 589182 547616
rect 589418 547380 589502 547616
rect 589738 547380 589770 547616
rect 589150 547296 589770 547380
rect 589150 547060 589182 547296
rect 589418 547060 589502 547296
rect 589738 547060 589770 547296
rect 589150 511616 589770 547060
rect 589150 511380 589182 511616
rect 589418 511380 589502 511616
rect 589738 511380 589770 511616
rect 589150 511296 589770 511380
rect 589150 511060 589182 511296
rect 589418 511060 589502 511296
rect 589738 511060 589770 511296
rect 589150 475616 589770 511060
rect 589150 475380 589182 475616
rect 589418 475380 589502 475616
rect 589738 475380 589770 475616
rect 589150 475296 589770 475380
rect 589150 475060 589182 475296
rect 589418 475060 589502 475296
rect 589738 475060 589770 475296
rect 589150 439616 589770 475060
rect 589150 439380 589182 439616
rect 589418 439380 589502 439616
rect 589738 439380 589770 439616
rect 589150 439296 589770 439380
rect 589150 439060 589182 439296
rect 589418 439060 589502 439296
rect 589738 439060 589770 439296
rect 589150 403616 589770 439060
rect 589150 403380 589182 403616
rect 589418 403380 589502 403616
rect 589738 403380 589770 403616
rect 589150 403296 589770 403380
rect 589150 403060 589182 403296
rect 589418 403060 589502 403296
rect 589738 403060 589770 403296
rect 589150 367616 589770 403060
rect 589150 367380 589182 367616
rect 589418 367380 589502 367616
rect 589738 367380 589770 367616
rect 589150 367296 589770 367380
rect 589150 367060 589182 367296
rect 589418 367060 589502 367296
rect 589738 367060 589770 367296
rect 589150 331616 589770 367060
rect 589150 331380 589182 331616
rect 589418 331380 589502 331616
rect 589738 331380 589770 331616
rect 589150 331296 589770 331380
rect 589150 331060 589182 331296
rect 589418 331060 589502 331296
rect 589738 331060 589770 331296
rect 589150 295616 589770 331060
rect 589150 295380 589182 295616
rect 589418 295380 589502 295616
rect 589738 295380 589770 295616
rect 589150 295296 589770 295380
rect 589150 295060 589182 295296
rect 589418 295060 589502 295296
rect 589738 295060 589770 295296
rect 589150 259616 589770 295060
rect 589150 259380 589182 259616
rect 589418 259380 589502 259616
rect 589738 259380 589770 259616
rect 589150 259296 589770 259380
rect 589150 259060 589182 259296
rect 589418 259060 589502 259296
rect 589738 259060 589770 259296
rect 589150 223616 589770 259060
rect 589150 223380 589182 223616
rect 589418 223380 589502 223616
rect 589738 223380 589770 223616
rect 589150 223296 589770 223380
rect 589150 223060 589182 223296
rect 589418 223060 589502 223296
rect 589738 223060 589770 223296
rect 589150 187616 589770 223060
rect 589150 187380 589182 187616
rect 589418 187380 589502 187616
rect 589738 187380 589770 187616
rect 589150 187296 589770 187380
rect 589150 187060 589182 187296
rect 589418 187060 589502 187296
rect 589738 187060 589770 187296
rect 589150 151616 589770 187060
rect 589150 151380 589182 151616
rect 589418 151380 589502 151616
rect 589738 151380 589770 151616
rect 589150 151296 589770 151380
rect 589150 151060 589182 151296
rect 589418 151060 589502 151296
rect 589738 151060 589770 151296
rect 589150 115616 589770 151060
rect 589150 115380 589182 115616
rect 589418 115380 589502 115616
rect 589738 115380 589770 115616
rect 589150 115296 589770 115380
rect 589150 115060 589182 115296
rect 589418 115060 589502 115296
rect 589738 115060 589770 115296
rect 589150 79616 589770 115060
rect 589150 79380 589182 79616
rect 589418 79380 589502 79616
rect 589738 79380 589770 79616
rect 589150 79296 589770 79380
rect 589150 79060 589182 79296
rect 589418 79060 589502 79296
rect 589738 79060 589770 79296
rect 589150 43616 589770 79060
rect 589150 43380 589182 43616
rect 589418 43380 589502 43616
rect 589738 43380 589770 43616
rect 589150 43296 589770 43380
rect 589150 43060 589182 43296
rect 589418 43060 589502 43296
rect 589738 43060 589770 43296
rect 589150 7616 589770 43060
rect 589150 7380 589182 7616
rect 589418 7380 589502 7616
rect 589738 7380 589770 7616
rect 589150 7296 589770 7380
rect 589150 7060 589182 7296
rect 589418 7060 589502 7296
rect 589738 7060 589770 7296
rect 581954 -4420 581986 -4184
rect 582222 -4420 582306 -4184
rect 582542 -4420 582574 -4184
rect 581954 -4504 582574 -4420
rect 581954 -4740 581986 -4504
rect 582222 -4740 582306 -4504
rect 582542 -4740 582574 -4504
rect 581954 -7652 582574 -4740
rect 589150 -4184 589770 7060
rect 589150 -4420 589182 -4184
rect 589418 -4420 589502 -4184
rect 589738 -4420 589770 -4184
rect 589150 -4504 589770 -4420
rect 589150 -4740 589182 -4504
rect 589418 -4740 589502 -4504
rect 589738 -4740 589770 -4504
rect 589150 -4772 589770 -4740
rect 590110 692856 590730 709084
rect 590110 692620 590142 692856
rect 590378 692620 590462 692856
rect 590698 692620 590730 692856
rect 590110 692536 590730 692620
rect 590110 692300 590142 692536
rect 590378 692300 590462 692536
rect 590698 692300 590730 692536
rect 590110 656856 590730 692300
rect 590110 656620 590142 656856
rect 590378 656620 590462 656856
rect 590698 656620 590730 656856
rect 590110 656536 590730 656620
rect 590110 656300 590142 656536
rect 590378 656300 590462 656536
rect 590698 656300 590730 656536
rect 590110 620856 590730 656300
rect 590110 620620 590142 620856
rect 590378 620620 590462 620856
rect 590698 620620 590730 620856
rect 590110 620536 590730 620620
rect 590110 620300 590142 620536
rect 590378 620300 590462 620536
rect 590698 620300 590730 620536
rect 590110 584856 590730 620300
rect 590110 584620 590142 584856
rect 590378 584620 590462 584856
rect 590698 584620 590730 584856
rect 590110 584536 590730 584620
rect 590110 584300 590142 584536
rect 590378 584300 590462 584536
rect 590698 584300 590730 584536
rect 590110 548856 590730 584300
rect 590110 548620 590142 548856
rect 590378 548620 590462 548856
rect 590698 548620 590730 548856
rect 590110 548536 590730 548620
rect 590110 548300 590142 548536
rect 590378 548300 590462 548536
rect 590698 548300 590730 548536
rect 590110 512856 590730 548300
rect 590110 512620 590142 512856
rect 590378 512620 590462 512856
rect 590698 512620 590730 512856
rect 590110 512536 590730 512620
rect 590110 512300 590142 512536
rect 590378 512300 590462 512536
rect 590698 512300 590730 512536
rect 590110 476856 590730 512300
rect 590110 476620 590142 476856
rect 590378 476620 590462 476856
rect 590698 476620 590730 476856
rect 590110 476536 590730 476620
rect 590110 476300 590142 476536
rect 590378 476300 590462 476536
rect 590698 476300 590730 476536
rect 590110 440856 590730 476300
rect 590110 440620 590142 440856
rect 590378 440620 590462 440856
rect 590698 440620 590730 440856
rect 590110 440536 590730 440620
rect 590110 440300 590142 440536
rect 590378 440300 590462 440536
rect 590698 440300 590730 440536
rect 590110 404856 590730 440300
rect 590110 404620 590142 404856
rect 590378 404620 590462 404856
rect 590698 404620 590730 404856
rect 590110 404536 590730 404620
rect 590110 404300 590142 404536
rect 590378 404300 590462 404536
rect 590698 404300 590730 404536
rect 590110 368856 590730 404300
rect 590110 368620 590142 368856
rect 590378 368620 590462 368856
rect 590698 368620 590730 368856
rect 590110 368536 590730 368620
rect 590110 368300 590142 368536
rect 590378 368300 590462 368536
rect 590698 368300 590730 368536
rect 590110 332856 590730 368300
rect 590110 332620 590142 332856
rect 590378 332620 590462 332856
rect 590698 332620 590730 332856
rect 590110 332536 590730 332620
rect 590110 332300 590142 332536
rect 590378 332300 590462 332536
rect 590698 332300 590730 332536
rect 590110 296856 590730 332300
rect 590110 296620 590142 296856
rect 590378 296620 590462 296856
rect 590698 296620 590730 296856
rect 590110 296536 590730 296620
rect 590110 296300 590142 296536
rect 590378 296300 590462 296536
rect 590698 296300 590730 296536
rect 590110 260856 590730 296300
rect 590110 260620 590142 260856
rect 590378 260620 590462 260856
rect 590698 260620 590730 260856
rect 590110 260536 590730 260620
rect 590110 260300 590142 260536
rect 590378 260300 590462 260536
rect 590698 260300 590730 260536
rect 590110 224856 590730 260300
rect 590110 224620 590142 224856
rect 590378 224620 590462 224856
rect 590698 224620 590730 224856
rect 590110 224536 590730 224620
rect 590110 224300 590142 224536
rect 590378 224300 590462 224536
rect 590698 224300 590730 224536
rect 590110 188856 590730 224300
rect 590110 188620 590142 188856
rect 590378 188620 590462 188856
rect 590698 188620 590730 188856
rect 590110 188536 590730 188620
rect 590110 188300 590142 188536
rect 590378 188300 590462 188536
rect 590698 188300 590730 188536
rect 590110 152856 590730 188300
rect 590110 152620 590142 152856
rect 590378 152620 590462 152856
rect 590698 152620 590730 152856
rect 590110 152536 590730 152620
rect 590110 152300 590142 152536
rect 590378 152300 590462 152536
rect 590698 152300 590730 152536
rect 590110 116856 590730 152300
rect 590110 116620 590142 116856
rect 590378 116620 590462 116856
rect 590698 116620 590730 116856
rect 590110 116536 590730 116620
rect 590110 116300 590142 116536
rect 590378 116300 590462 116536
rect 590698 116300 590730 116536
rect 590110 80856 590730 116300
rect 590110 80620 590142 80856
rect 590378 80620 590462 80856
rect 590698 80620 590730 80856
rect 590110 80536 590730 80620
rect 590110 80300 590142 80536
rect 590378 80300 590462 80536
rect 590698 80300 590730 80536
rect 590110 44856 590730 80300
rect 590110 44620 590142 44856
rect 590378 44620 590462 44856
rect 590698 44620 590730 44856
rect 590110 44536 590730 44620
rect 590110 44300 590142 44536
rect 590378 44300 590462 44536
rect 590698 44300 590730 44536
rect 590110 8856 590730 44300
rect 590110 8620 590142 8856
rect 590378 8620 590462 8856
rect 590698 8620 590730 8856
rect 590110 8536 590730 8620
rect 590110 8300 590142 8536
rect 590378 8300 590462 8536
rect 590698 8300 590730 8536
rect 590110 -5144 590730 8300
rect 590110 -5380 590142 -5144
rect 590378 -5380 590462 -5144
rect 590698 -5380 590730 -5144
rect 590110 -5464 590730 -5380
rect 590110 -5700 590142 -5464
rect 590378 -5700 590462 -5464
rect 590698 -5700 590730 -5464
rect 590110 -5732 590730 -5700
rect 591070 694096 591690 710044
rect 591070 693860 591102 694096
rect 591338 693860 591422 694096
rect 591658 693860 591690 694096
rect 591070 693776 591690 693860
rect 591070 693540 591102 693776
rect 591338 693540 591422 693776
rect 591658 693540 591690 693776
rect 591070 658096 591690 693540
rect 591070 657860 591102 658096
rect 591338 657860 591422 658096
rect 591658 657860 591690 658096
rect 591070 657776 591690 657860
rect 591070 657540 591102 657776
rect 591338 657540 591422 657776
rect 591658 657540 591690 657776
rect 591070 622096 591690 657540
rect 591070 621860 591102 622096
rect 591338 621860 591422 622096
rect 591658 621860 591690 622096
rect 591070 621776 591690 621860
rect 591070 621540 591102 621776
rect 591338 621540 591422 621776
rect 591658 621540 591690 621776
rect 591070 586096 591690 621540
rect 591070 585860 591102 586096
rect 591338 585860 591422 586096
rect 591658 585860 591690 586096
rect 591070 585776 591690 585860
rect 591070 585540 591102 585776
rect 591338 585540 591422 585776
rect 591658 585540 591690 585776
rect 591070 550096 591690 585540
rect 591070 549860 591102 550096
rect 591338 549860 591422 550096
rect 591658 549860 591690 550096
rect 591070 549776 591690 549860
rect 591070 549540 591102 549776
rect 591338 549540 591422 549776
rect 591658 549540 591690 549776
rect 591070 514096 591690 549540
rect 591070 513860 591102 514096
rect 591338 513860 591422 514096
rect 591658 513860 591690 514096
rect 591070 513776 591690 513860
rect 591070 513540 591102 513776
rect 591338 513540 591422 513776
rect 591658 513540 591690 513776
rect 591070 478096 591690 513540
rect 591070 477860 591102 478096
rect 591338 477860 591422 478096
rect 591658 477860 591690 478096
rect 591070 477776 591690 477860
rect 591070 477540 591102 477776
rect 591338 477540 591422 477776
rect 591658 477540 591690 477776
rect 591070 442096 591690 477540
rect 591070 441860 591102 442096
rect 591338 441860 591422 442096
rect 591658 441860 591690 442096
rect 591070 441776 591690 441860
rect 591070 441540 591102 441776
rect 591338 441540 591422 441776
rect 591658 441540 591690 441776
rect 591070 406096 591690 441540
rect 591070 405860 591102 406096
rect 591338 405860 591422 406096
rect 591658 405860 591690 406096
rect 591070 405776 591690 405860
rect 591070 405540 591102 405776
rect 591338 405540 591422 405776
rect 591658 405540 591690 405776
rect 591070 370096 591690 405540
rect 591070 369860 591102 370096
rect 591338 369860 591422 370096
rect 591658 369860 591690 370096
rect 591070 369776 591690 369860
rect 591070 369540 591102 369776
rect 591338 369540 591422 369776
rect 591658 369540 591690 369776
rect 591070 334096 591690 369540
rect 591070 333860 591102 334096
rect 591338 333860 591422 334096
rect 591658 333860 591690 334096
rect 591070 333776 591690 333860
rect 591070 333540 591102 333776
rect 591338 333540 591422 333776
rect 591658 333540 591690 333776
rect 591070 298096 591690 333540
rect 591070 297860 591102 298096
rect 591338 297860 591422 298096
rect 591658 297860 591690 298096
rect 591070 297776 591690 297860
rect 591070 297540 591102 297776
rect 591338 297540 591422 297776
rect 591658 297540 591690 297776
rect 591070 262096 591690 297540
rect 591070 261860 591102 262096
rect 591338 261860 591422 262096
rect 591658 261860 591690 262096
rect 591070 261776 591690 261860
rect 591070 261540 591102 261776
rect 591338 261540 591422 261776
rect 591658 261540 591690 261776
rect 591070 226096 591690 261540
rect 591070 225860 591102 226096
rect 591338 225860 591422 226096
rect 591658 225860 591690 226096
rect 591070 225776 591690 225860
rect 591070 225540 591102 225776
rect 591338 225540 591422 225776
rect 591658 225540 591690 225776
rect 591070 190096 591690 225540
rect 591070 189860 591102 190096
rect 591338 189860 591422 190096
rect 591658 189860 591690 190096
rect 591070 189776 591690 189860
rect 591070 189540 591102 189776
rect 591338 189540 591422 189776
rect 591658 189540 591690 189776
rect 591070 154096 591690 189540
rect 591070 153860 591102 154096
rect 591338 153860 591422 154096
rect 591658 153860 591690 154096
rect 591070 153776 591690 153860
rect 591070 153540 591102 153776
rect 591338 153540 591422 153776
rect 591658 153540 591690 153776
rect 591070 118096 591690 153540
rect 591070 117860 591102 118096
rect 591338 117860 591422 118096
rect 591658 117860 591690 118096
rect 591070 117776 591690 117860
rect 591070 117540 591102 117776
rect 591338 117540 591422 117776
rect 591658 117540 591690 117776
rect 591070 82096 591690 117540
rect 591070 81860 591102 82096
rect 591338 81860 591422 82096
rect 591658 81860 591690 82096
rect 591070 81776 591690 81860
rect 591070 81540 591102 81776
rect 591338 81540 591422 81776
rect 591658 81540 591690 81776
rect 591070 46096 591690 81540
rect 591070 45860 591102 46096
rect 591338 45860 591422 46096
rect 591658 45860 591690 46096
rect 591070 45776 591690 45860
rect 591070 45540 591102 45776
rect 591338 45540 591422 45776
rect 591658 45540 591690 45776
rect 591070 10096 591690 45540
rect 591070 9860 591102 10096
rect 591338 9860 591422 10096
rect 591658 9860 591690 10096
rect 591070 9776 591690 9860
rect 591070 9540 591102 9776
rect 591338 9540 591422 9776
rect 591658 9540 591690 9776
rect 591070 -6104 591690 9540
rect 591070 -6340 591102 -6104
rect 591338 -6340 591422 -6104
rect 591658 -6340 591690 -6104
rect 591070 -6424 591690 -6340
rect 591070 -6660 591102 -6424
rect 591338 -6660 591422 -6424
rect 591658 -6660 591690 -6424
rect 591070 -6692 591690 -6660
rect 592030 695336 592650 711004
rect 592030 695100 592062 695336
rect 592298 695100 592382 695336
rect 592618 695100 592650 695336
rect 592030 695016 592650 695100
rect 592030 694780 592062 695016
rect 592298 694780 592382 695016
rect 592618 694780 592650 695016
rect 592030 659336 592650 694780
rect 592030 659100 592062 659336
rect 592298 659100 592382 659336
rect 592618 659100 592650 659336
rect 592030 659016 592650 659100
rect 592030 658780 592062 659016
rect 592298 658780 592382 659016
rect 592618 658780 592650 659016
rect 592030 623336 592650 658780
rect 592030 623100 592062 623336
rect 592298 623100 592382 623336
rect 592618 623100 592650 623336
rect 592030 623016 592650 623100
rect 592030 622780 592062 623016
rect 592298 622780 592382 623016
rect 592618 622780 592650 623016
rect 592030 587336 592650 622780
rect 592030 587100 592062 587336
rect 592298 587100 592382 587336
rect 592618 587100 592650 587336
rect 592030 587016 592650 587100
rect 592030 586780 592062 587016
rect 592298 586780 592382 587016
rect 592618 586780 592650 587016
rect 592030 551336 592650 586780
rect 592030 551100 592062 551336
rect 592298 551100 592382 551336
rect 592618 551100 592650 551336
rect 592030 551016 592650 551100
rect 592030 550780 592062 551016
rect 592298 550780 592382 551016
rect 592618 550780 592650 551016
rect 592030 515336 592650 550780
rect 592030 515100 592062 515336
rect 592298 515100 592382 515336
rect 592618 515100 592650 515336
rect 592030 515016 592650 515100
rect 592030 514780 592062 515016
rect 592298 514780 592382 515016
rect 592618 514780 592650 515016
rect 592030 479336 592650 514780
rect 592030 479100 592062 479336
rect 592298 479100 592382 479336
rect 592618 479100 592650 479336
rect 592030 479016 592650 479100
rect 592030 478780 592062 479016
rect 592298 478780 592382 479016
rect 592618 478780 592650 479016
rect 592030 443336 592650 478780
rect 592030 443100 592062 443336
rect 592298 443100 592382 443336
rect 592618 443100 592650 443336
rect 592030 443016 592650 443100
rect 592030 442780 592062 443016
rect 592298 442780 592382 443016
rect 592618 442780 592650 443016
rect 592030 407336 592650 442780
rect 592030 407100 592062 407336
rect 592298 407100 592382 407336
rect 592618 407100 592650 407336
rect 592030 407016 592650 407100
rect 592030 406780 592062 407016
rect 592298 406780 592382 407016
rect 592618 406780 592650 407016
rect 592030 371336 592650 406780
rect 592030 371100 592062 371336
rect 592298 371100 592382 371336
rect 592618 371100 592650 371336
rect 592030 371016 592650 371100
rect 592030 370780 592062 371016
rect 592298 370780 592382 371016
rect 592618 370780 592650 371016
rect 592030 335336 592650 370780
rect 592030 335100 592062 335336
rect 592298 335100 592382 335336
rect 592618 335100 592650 335336
rect 592030 335016 592650 335100
rect 592030 334780 592062 335016
rect 592298 334780 592382 335016
rect 592618 334780 592650 335016
rect 592030 299336 592650 334780
rect 592030 299100 592062 299336
rect 592298 299100 592382 299336
rect 592618 299100 592650 299336
rect 592030 299016 592650 299100
rect 592030 298780 592062 299016
rect 592298 298780 592382 299016
rect 592618 298780 592650 299016
rect 592030 263336 592650 298780
rect 592030 263100 592062 263336
rect 592298 263100 592382 263336
rect 592618 263100 592650 263336
rect 592030 263016 592650 263100
rect 592030 262780 592062 263016
rect 592298 262780 592382 263016
rect 592618 262780 592650 263016
rect 592030 227336 592650 262780
rect 592030 227100 592062 227336
rect 592298 227100 592382 227336
rect 592618 227100 592650 227336
rect 592030 227016 592650 227100
rect 592030 226780 592062 227016
rect 592298 226780 592382 227016
rect 592618 226780 592650 227016
rect 592030 191336 592650 226780
rect 592030 191100 592062 191336
rect 592298 191100 592382 191336
rect 592618 191100 592650 191336
rect 592030 191016 592650 191100
rect 592030 190780 592062 191016
rect 592298 190780 592382 191016
rect 592618 190780 592650 191016
rect 592030 155336 592650 190780
rect 592030 155100 592062 155336
rect 592298 155100 592382 155336
rect 592618 155100 592650 155336
rect 592030 155016 592650 155100
rect 592030 154780 592062 155016
rect 592298 154780 592382 155016
rect 592618 154780 592650 155016
rect 592030 119336 592650 154780
rect 592030 119100 592062 119336
rect 592298 119100 592382 119336
rect 592618 119100 592650 119336
rect 592030 119016 592650 119100
rect 592030 118780 592062 119016
rect 592298 118780 592382 119016
rect 592618 118780 592650 119016
rect 592030 83336 592650 118780
rect 592030 83100 592062 83336
rect 592298 83100 592382 83336
rect 592618 83100 592650 83336
rect 592030 83016 592650 83100
rect 592030 82780 592062 83016
rect 592298 82780 592382 83016
rect 592618 82780 592650 83016
rect 592030 47336 592650 82780
rect 592030 47100 592062 47336
rect 592298 47100 592382 47336
rect 592618 47100 592650 47336
rect 592030 47016 592650 47100
rect 592030 46780 592062 47016
rect 592298 46780 592382 47016
rect 592618 46780 592650 47016
rect 592030 11336 592650 46780
rect 592030 11100 592062 11336
rect 592298 11100 592382 11336
rect 592618 11100 592650 11336
rect 592030 11016 592650 11100
rect 592030 10780 592062 11016
rect 592298 10780 592382 11016
rect 592618 10780 592650 11016
rect 592030 -7064 592650 10780
rect 592030 -7300 592062 -7064
rect 592298 -7300 592382 -7064
rect 592618 -7300 592650 -7064
rect 592030 -7384 592650 -7300
rect 592030 -7620 592062 -7384
rect 592298 -7620 592382 -7384
rect 592618 -7620 592650 -7384
rect 592030 -7652 592650 -7620
<< via4 >>
rect -8694 711324 -8458 711560
rect -8374 711324 -8138 711560
rect -8694 711004 -8458 711240
rect -8374 711004 -8138 711240
rect -8694 695100 -8458 695336
rect -8374 695100 -8138 695336
rect -8694 694780 -8458 695016
rect -8374 694780 -8138 695016
rect -8694 659100 -8458 659336
rect -8374 659100 -8138 659336
rect -8694 658780 -8458 659016
rect -8374 658780 -8138 659016
rect -8694 623100 -8458 623336
rect -8374 623100 -8138 623336
rect -8694 622780 -8458 623016
rect -8374 622780 -8138 623016
rect -8694 587100 -8458 587336
rect -8374 587100 -8138 587336
rect -8694 586780 -8458 587016
rect -8374 586780 -8138 587016
rect -8694 551100 -8458 551336
rect -8374 551100 -8138 551336
rect -8694 550780 -8458 551016
rect -8374 550780 -8138 551016
rect -8694 515100 -8458 515336
rect -8374 515100 -8138 515336
rect -8694 514780 -8458 515016
rect -8374 514780 -8138 515016
rect -8694 479100 -8458 479336
rect -8374 479100 -8138 479336
rect -8694 478780 -8458 479016
rect -8374 478780 -8138 479016
rect -8694 443100 -8458 443336
rect -8374 443100 -8138 443336
rect -8694 442780 -8458 443016
rect -8374 442780 -8138 443016
rect -8694 407100 -8458 407336
rect -8374 407100 -8138 407336
rect -8694 406780 -8458 407016
rect -8374 406780 -8138 407016
rect -8694 371100 -8458 371336
rect -8374 371100 -8138 371336
rect -8694 370780 -8458 371016
rect -8374 370780 -8138 371016
rect -8694 335100 -8458 335336
rect -8374 335100 -8138 335336
rect -8694 334780 -8458 335016
rect -8374 334780 -8138 335016
rect -8694 299100 -8458 299336
rect -8374 299100 -8138 299336
rect -8694 298780 -8458 299016
rect -8374 298780 -8138 299016
rect -8694 263100 -8458 263336
rect -8374 263100 -8138 263336
rect -8694 262780 -8458 263016
rect -8374 262780 -8138 263016
rect -8694 227100 -8458 227336
rect -8374 227100 -8138 227336
rect -8694 226780 -8458 227016
rect -8374 226780 -8138 227016
rect -8694 191100 -8458 191336
rect -8374 191100 -8138 191336
rect -8694 190780 -8458 191016
rect -8374 190780 -8138 191016
rect -8694 155100 -8458 155336
rect -8374 155100 -8138 155336
rect -8694 154780 -8458 155016
rect -8374 154780 -8138 155016
rect -8694 119100 -8458 119336
rect -8374 119100 -8138 119336
rect -8694 118780 -8458 119016
rect -8374 118780 -8138 119016
rect -8694 83100 -8458 83336
rect -8374 83100 -8138 83336
rect -8694 82780 -8458 83016
rect -8374 82780 -8138 83016
rect -8694 47100 -8458 47336
rect -8374 47100 -8138 47336
rect -8694 46780 -8458 47016
rect -8374 46780 -8138 47016
rect -8694 11100 -8458 11336
rect -8374 11100 -8138 11336
rect -8694 10780 -8458 11016
rect -8374 10780 -8138 11016
rect -7734 710364 -7498 710600
rect -7414 710364 -7178 710600
rect -7734 710044 -7498 710280
rect -7414 710044 -7178 710280
rect -7734 693860 -7498 694096
rect -7414 693860 -7178 694096
rect -7734 693540 -7498 693776
rect -7414 693540 -7178 693776
rect -7734 657860 -7498 658096
rect -7414 657860 -7178 658096
rect -7734 657540 -7498 657776
rect -7414 657540 -7178 657776
rect -7734 621860 -7498 622096
rect -7414 621860 -7178 622096
rect -7734 621540 -7498 621776
rect -7414 621540 -7178 621776
rect -7734 585860 -7498 586096
rect -7414 585860 -7178 586096
rect -7734 585540 -7498 585776
rect -7414 585540 -7178 585776
rect -7734 549860 -7498 550096
rect -7414 549860 -7178 550096
rect -7734 549540 -7498 549776
rect -7414 549540 -7178 549776
rect -7734 513860 -7498 514096
rect -7414 513860 -7178 514096
rect -7734 513540 -7498 513776
rect -7414 513540 -7178 513776
rect -7734 477860 -7498 478096
rect -7414 477860 -7178 478096
rect -7734 477540 -7498 477776
rect -7414 477540 -7178 477776
rect -7734 441860 -7498 442096
rect -7414 441860 -7178 442096
rect -7734 441540 -7498 441776
rect -7414 441540 -7178 441776
rect -7734 405860 -7498 406096
rect -7414 405860 -7178 406096
rect -7734 405540 -7498 405776
rect -7414 405540 -7178 405776
rect -7734 369860 -7498 370096
rect -7414 369860 -7178 370096
rect -7734 369540 -7498 369776
rect -7414 369540 -7178 369776
rect -7734 333860 -7498 334096
rect -7414 333860 -7178 334096
rect -7734 333540 -7498 333776
rect -7414 333540 -7178 333776
rect -7734 297860 -7498 298096
rect -7414 297860 -7178 298096
rect -7734 297540 -7498 297776
rect -7414 297540 -7178 297776
rect -7734 261860 -7498 262096
rect -7414 261860 -7178 262096
rect -7734 261540 -7498 261776
rect -7414 261540 -7178 261776
rect -7734 225860 -7498 226096
rect -7414 225860 -7178 226096
rect -7734 225540 -7498 225776
rect -7414 225540 -7178 225776
rect -7734 189860 -7498 190096
rect -7414 189860 -7178 190096
rect -7734 189540 -7498 189776
rect -7414 189540 -7178 189776
rect -7734 153860 -7498 154096
rect -7414 153860 -7178 154096
rect -7734 153540 -7498 153776
rect -7414 153540 -7178 153776
rect -7734 117860 -7498 118096
rect -7414 117860 -7178 118096
rect -7734 117540 -7498 117776
rect -7414 117540 -7178 117776
rect -7734 81860 -7498 82096
rect -7414 81860 -7178 82096
rect -7734 81540 -7498 81776
rect -7414 81540 -7178 81776
rect -7734 45860 -7498 46096
rect -7414 45860 -7178 46096
rect -7734 45540 -7498 45776
rect -7414 45540 -7178 45776
rect -7734 9860 -7498 10096
rect -7414 9860 -7178 10096
rect -7734 9540 -7498 9776
rect -7414 9540 -7178 9776
rect -6774 709404 -6538 709640
rect -6454 709404 -6218 709640
rect -6774 709084 -6538 709320
rect -6454 709084 -6218 709320
rect -6774 692620 -6538 692856
rect -6454 692620 -6218 692856
rect -6774 692300 -6538 692536
rect -6454 692300 -6218 692536
rect -6774 656620 -6538 656856
rect -6454 656620 -6218 656856
rect -6774 656300 -6538 656536
rect -6454 656300 -6218 656536
rect -6774 620620 -6538 620856
rect -6454 620620 -6218 620856
rect -6774 620300 -6538 620536
rect -6454 620300 -6218 620536
rect -6774 584620 -6538 584856
rect -6454 584620 -6218 584856
rect -6774 584300 -6538 584536
rect -6454 584300 -6218 584536
rect -6774 548620 -6538 548856
rect -6454 548620 -6218 548856
rect -6774 548300 -6538 548536
rect -6454 548300 -6218 548536
rect -6774 512620 -6538 512856
rect -6454 512620 -6218 512856
rect -6774 512300 -6538 512536
rect -6454 512300 -6218 512536
rect -6774 476620 -6538 476856
rect -6454 476620 -6218 476856
rect -6774 476300 -6538 476536
rect -6454 476300 -6218 476536
rect -6774 440620 -6538 440856
rect -6454 440620 -6218 440856
rect -6774 440300 -6538 440536
rect -6454 440300 -6218 440536
rect -6774 404620 -6538 404856
rect -6454 404620 -6218 404856
rect -6774 404300 -6538 404536
rect -6454 404300 -6218 404536
rect -6774 368620 -6538 368856
rect -6454 368620 -6218 368856
rect -6774 368300 -6538 368536
rect -6454 368300 -6218 368536
rect -6774 332620 -6538 332856
rect -6454 332620 -6218 332856
rect -6774 332300 -6538 332536
rect -6454 332300 -6218 332536
rect -6774 296620 -6538 296856
rect -6454 296620 -6218 296856
rect -6774 296300 -6538 296536
rect -6454 296300 -6218 296536
rect -6774 260620 -6538 260856
rect -6454 260620 -6218 260856
rect -6774 260300 -6538 260536
rect -6454 260300 -6218 260536
rect -6774 224620 -6538 224856
rect -6454 224620 -6218 224856
rect -6774 224300 -6538 224536
rect -6454 224300 -6218 224536
rect -6774 188620 -6538 188856
rect -6454 188620 -6218 188856
rect -6774 188300 -6538 188536
rect -6454 188300 -6218 188536
rect -6774 152620 -6538 152856
rect -6454 152620 -6218 152856
rect -6774 152300 -6538 152536
rect -6454 152300 -6218 152536
rect -6774 116620 -6538 116856
rect -6454 116620 -6218 116856
rect -6774 116300 -6538 116536
rect -6454 116300 -6218 116536
rect -6774 80620 -6538 80856
rect -6454 80620 -6218 80856
rect -6774 80300 -6538 80536
rect -6454 80300 -6218 80536
rect -6774 44620 -6538 44856
rect -6454 44620 -6218 44856
rect -6774 44300 -6538 44536
rect -6454 44300 -6218 44536
rect -6774 8620 -6538 8856
rect -6454 8620 -6218 8856
rect -6774 8300 -6538 8536
rect -6454 8300 -6218 8536
rect -5814 708444 -5578 708680
rect -5494 708444 -5258 708680
rect -5814 708124 -5578 708360
rect -5494 708124 -5258 708360
rect -5814 691380 -5578 691616
rect -5494 691380 -5258 691616
rect -5814 691060 -5578 691296
rect -5494 691060 -5258 691296
rect -5814 655380 -5578 655616
rect -5494 655380 -5258 655616
rect -5814 655060 -5578 655296
rect -5494 655060 -5258 655296
rect -5814 619380 -5578 619616
rect -5494 619380 -5258 619616
rect -5814 619060 -5578 619296
rect -5494 619060 -5258 619296
rect -5814 583380 -5578 583616
rect -5494 583380 -5258 583616
rect -5814 583060 -5578 583296
rect -5494 583060 -5258 583296
rect -5814 547380 -5578 547616
rect -5494 547380 -5258 547616
rect -5814 547060 -5578 547296
rect -5494 547060 -5258 547296
rect -5814 511380 -5578 511616
rect -5494 511380 -5258 511616
rect -5814 511060 -5578 511296
rect -5494 511060 -5258 511296
rect -5814 475380 -5578 475616
rect -5494 475380 -5258 475616
rect -5814 475060 -5578 475296
rect -5494 475060 -5258 475296
rect -5814 439380 -5578 439616
rect -5494 439380 -5258 439616
rect -5814 439060 -5578 439296
rect -5494 439060 -5258 439296
rect -5814 403380 -5578 403616
rect -5494 403380 -5258 403616
rect -5814 403060 -5578 403296
rect -5494 403060 -5258 403296
rect -5814 367380 -5578 367616
rect -5494 367380 -5258 367616
rect -5814 367060 -5578 367296
rect -5494 367060 -5258 367296
rect -5814 331380 -5578 331616
rect -5494 331380 -5258 331616
rect -5814 331060 -5578 331296
rect -5494 331060 -5258 331296
rect -5814 295380 -5578 295616
rect -5494 295380 -5258 295616
rect -5814 295060 -5578 295296
rect -5494 295060 -5258 295296
rect -5814 259380 -5578 259616
rect -5494 259380 -5258 259616
rect -5814 259060 -5578 259296
rect -5494 259060 -5258 259296
rect -5814 223380 -5578 223616
rect -5494 223380 -5258 223616
rect -5814 223060 -5578 223296
rect -5494 223060 -5258 223296
rect -5814 187380 -5578 187616
rect -5494 187380 -5258 187616
rect -5814 187060 -5578 187296
rect -5494 187060 -5258 187296
rect -5814 151380 -5578 151616
rect -5494 151380 -5258 151616
rect -5814 151060 -5578 151296
rect -5494 151060 -5258 151296
rect -5814 115380 -5578 115616
rect -5494 115380 -5258 115616
rect -5814 115060 -5578 115296
rect -5494 115060 -5258 115296
rect -5814 79380 -5578 79616
rect -5494 79380 -5258 79616
rect -5814 79060 -5578 79296
rect -5494 79060 -5258 79296
rect -5814 43380 -5578 43616
rect -5494 43380 -5258 43616
rect -5814 43060 -5578 43296
rect -5494 43060 -5258 43296
rect -5814 7380 -5578 7616
rect -5494 7380 -5258 7616
rect -5814 7060 -5578 7296
rect -5494 7060 -5258 7296
rect -4854 707484 -4618 707720
rect -4534 707484 -4298 707720
rect -4854 707164 -4618 707400
rect -4534 707164 -4298 707400
rect -4854 690140 -4618 690376
rect -4534 690140 -4298 690376
rect -4854 689820 -4618 690056
rect -4534 689820 -4298 690056
rect -4854 654140 -4618 654376
rect -4534 654140 -4298 654376
rect -4854 653820 -4618 654056
rect -4534 653820 -4298 654056
rect -4854 618140 -4618 618376
rect -4534 618140 -4298 618376
rect -4854 617820 -4618 618056
rect -4534 617820 -4298 618056
rect -4854 582140 -4618 582376
rect -4534 582140 -4298 582376
rect -4854 581820 -4618 582056
rect -4534 581820 -4298 582056
rect -4854 546140 -4618 546376
rect -4534 546140 -4298 546376
rect -4854 545820 -4618 546056
rect -4534 545820 -4298 546056
rect -4854 510140 -4618 510376
rect -4534 510140 -4298 510376
rect -4854 509820 -4618 510056
rect -4534 509820 -4298 510056
rect -4854 474140 -4618 474376
rect -4534 474140 -4298 474376
rect -4854 473820 -4618 474056
rect -4534 473820 -4298 474056
rect -4854 438140 -4618 438376
rect -4534 438140 -4298 438376
rect -4854 437820 -4618 438056
rect -4534 437820 -4298 438056
rect -4854 402140 -4618 402376
rect -4534 402140 -4298 402376
rect -4854 401820 -4618 402056
rect -4534 401820 -4298 402056
rect -4854 366140 -4618 366376
rect -4534 366140 -4298 366376
rect -4854 365820 -4618 366056
rect -4534 365820 -4298 366056
rect -4854 330140 -4618 330376
rect -4534 330140 -4298 330376
rect -4854 329820 -4618 330056
rect -4534 329820 -4298 330056
rect -4854 294140 -4618 294376
rect -4534 294140 -4298 294376
rect -4854 293820 -4618 294056
rect -4534 293820 -4298 294056
rect -4854 258140 -4618 258376
rect -4534 258140 -4298 258376
rect -4854 257820 -4618 258056
rect -4534 257820 -4298 258056
rect -4854 222140 -4618 222376
rect -4534 222140 -4298 222376
rect -4854 221820 -4618 222056
rect -4534 221820 -4298 222056
rect -4854 186140 -4618 186376
rect -4534 186140 -4298 186376
rect -4854 185820 -4618 186056
rect -4534 185820 -4298 186056
rect -4854 150140 -4618 150376
rect -4534 150140 -4298 150376
rect -4854 149820 -4618 150056
rect -4534 149820 -4298 150056
rect -4854 114140 -4618 114376
rect -4534 114140 -4298 114376
rect -4854 113820 -4618 114056
rect -4534 113820 -4298 114056
rect -4854 78140 -4618 78376
rect -4534 78140 -4298 78376
rect -4854 77820 -4618 78056
rect -4534 77820 -4298 78056
rect -4854 42140 -4618 42376
rect -4534 42140 -4298 42376
rect -4854 41820 -4618 42056
rect -4534 41820 -4298 42056
rect -4854 6140 -4618 6376
rect -4534 6140 -4298 6376
rect -4854 5820 -4618 6056
rect -4534 5820 -4298 6056
rect -3894 706524 -3658 706760
rect -3574 706524 -3338 706760
rect -3894 706204 -3658 706440
rect -3574 706204 -3338 706440
rect -3894 688900 -3658 689136
rect -3574 688900 -3338 689136
rect -3894 688580 -3658 688816
rect -3574 688580 -3338 688816
rect -3894 652900 -3658 653136
rect -3574 652900 -3338 653136
rect -3894 652580 -3658 652816
rect -3574 652580 -3338 652816
rect -3894 616900 -3658 617136
rect -3574 616900 -3338 617136
rect -3894 616580 -3658 616816
rect -3574 616580 -3338 616816
rect -3894 580900 -3658 581136
rect -3574 580900 -3338 581136
rect -3894 580580 -3658 580816
rect -3574 580580 -3338 580816
rect -3894 544900 -3658 545136
rect -3574 544900 -3338 545136
rect -3894 544580 -3658 544816
rect -3574 544580 -3338 544816
rect -3894 508900 -3658 509136
rect -3574 508900 -3338 509136
rect -3894 508580 -3658 508816
rect -3574 508580 -3338 508816
rect -3894 472900 -3658 473136
rect -3574 472900 -3338 473136
rect -3894 472580 -3658 472816
rect -3574 472580 -3338 472816
rect -3894 436900 -3658 437136
rect -3574 436900 -3338 437136
rect -3894 436580 -3658 436816
rect -3574 436580 -3338 436816
rect -3894 400900 -3658 401136
rect -3574 400900 -3338 401136
rect -3894 400580 -3658 400816
rect -3574 400580 -3338 400816
rect -3894 364900 -3658 365136
rect -3574 364900 -3338 365136
rect -3894 364580 -3658 364816
rect -3574 364580 -3338 364816
rect -3894 328900 -3658 329136
rect -3574 328900 -3338 329136
rect -3894 328580 -3658 328816
rect -3574 328580 -3338 328816
rect -3894 292900 -3658 293136
rect -3574 292900 -3338 293136
rect -3894 292580 -3658 292816
rect -3574 292580 -3338 292816
rect -3894 256900 -3658 257136
rect -3574 256900 -3338 257136
rect -3894 256580 -3658 256816
rect -3574 256580 -3338 256816
rect -3894 220900 -3658 221136
rect -3574 220900 -3338 221136
rect -3894 220580 -3658 220816
rect -3574 220580 -3338 220816
rect -3894 184900 -3658 185136
rect -3574 184900 -3338 185136
rect -3894 184580 -3658 184816
rect -3574 184580 -3338 184816
rect -3894 148900 -3658 149136
rect -3574 148900 -3338 149136
rect -3894 148580 -3658 148816
rect -3574 148580 -3338 148816
rect -3894 112900 -3658 113136
rect -3574 112900 -3338 113136
rect -3894 112580 -3658 112816
rect -3574 112580 -3338 112816
rect -3894 76900 -3658 77136
rect -3574 76900 -3338 77136
rect -3894 76580 -3658 76816
rect -3574 76580 -3338 76816
rect -3894 40900 -3658 41136
rect -3574 40900 -3338 41136
rect -3894 40580 -3658 40816
rect -3574 40580 -3338 40816
rect -3894 4900 -3658 5136
rect -3574 4900 -3338 5136
rect -3894 4580 -3658 4816
rect -3574 4580 -3338 4816
rect -2934 705564 -2698 705800
rect -2614 705564 -2378 705800
rect -2934 705244 -2698 705480
rect -2614 705244 -2378 705480
rect -2934 687660 -2698 687896
rect -2614 687660 -2378 687896
rect -2934 687340 -2698 687576
rect -2614 687340 -2378 687576
rect -2934 651660 -2698 651896
rect -2614 651660 -2378 651896
rect -2934 651340 -2698 651576
rect -2614 651340 -2378 651576
rect -2934 615660 -2698 615896
rect -2614 615660 -2378 615896
rect -2934 615340 -2698 615576
rect -2614 615340 -2378 615576
rect -2934 579660 -2698 579896
rect -2614 579660 -2378 579896
rect -2934 579340 -2698 579576
rect -2614 579340 -2378 579576
rect -2934 543660 -2698 543896
rect -2614 543660 -2378 543896
rect -2934 543340 -2698 543576
rect -2614 543340 -2378 543576
rect -2934 507660 -2698 507896
rect -2614 507660 -2378 507896
rect -2934 507340 -2698 507576
rect -2614 507340 -2378 507576
rect -2934 471660 -2698 471896
rect -2614 471660 -2378 471896
rect -2934 471340 -2698 471576
rect -2614 471340 -2378 471576
rect -2934 435660 -2698 435896
rect -2614 435660 -2378 435896
rect -2934 435340 -2698 435576
rect -2614 435340 -2378 435576
rect -2934 399660 -2698 399896
rect -2614 399660 -2378 399896
rect -2934 399340 -2698 399576
rect -2614 399340 -2378 399576
rect -2934 363660 -2698 363896
rect -2614 363660 -2378 363896
rect -2934 363340 -2698 363576
rect -2614 363340 -2378 363576
rect -2934 327660 -2698 327896
rect -2614 327660 -2378 327896
rect -2934 327340 -2698 327576
rect -2614 327340 -2378 327576
rect -2934 291660 -2698 291896
rect -2614 291660 -2378 291896
rect -2934 291340 -2698 291576
rect -2614 291340 -2378 291576
rect -2934 255660 -2698 255896
rect -2614 255660 -2378 255896
rect -2934 255340 -2698 255576
rect -2614 255340 -2378 255576
rect -2934 219660 -2698 219896
rect -2614 219660 -2378 219896
rect -2934 219340 -2698 219576
rect -2614 219340 -2378 219576
rect -2934 183660 -2698 183896
rect -2614 183660 -2378 183896
rect -2934 183340 -2698 183576
rect -2614 183340 -2378 183576
rect -2934 147660 -2698 147896
rect -2614 147660 -2378 147896
rect -2934 147340 -2698 147576
rect -2614 147340 -2378 147576
rect -2934 111660 -2698 111896
rect -2614 111660 -2378 111896
rect -2934 111340 -2698 111576
rect -2614 111340 -2378 111576
rect -2934 75660 -2698 75896
rect -2614 75660 -2378 75896
rect -2934 75340 -2698 75576
rect -2614 75340 -2378 75576
rect -2934 39660 -2698 39896
rect -2614 39660 -2378 39896
rect -2934 39340 -2698 39576
rect -2614 39340 -2378 39576
rect -2934 3660 -2698 3896
rect -2614 3660 -2378 3896
rect -2934 3340 -2698 3576
rect -2614 3340 -2378 3576
rect -1974 704604 -1738 704840
rect -1654 704604 -1418 704840
rect -1974 704284 -1738 704520
rect -1654 704284 -1418 704520
rect -1974 686420 -1738 686656
rect -1654 686420 -1418 686656
rect -1974 686100 -1738 686336
rect -1654 686100 -1418 686336
rect -1974 650420 -1738 650656
rect -1654 650420 -1418 650656
rect -1974 650100 -1738 650336
rect -1654 650100 -1418 650336
rect -1974 614420 -1738 614656
rect -1654 614420 -1418 614656
rect -1974 614100 -1738 614336
rect -1654 614100 -1418 614336
rect -1974 578420 -1738 578656
rect -1654 578420 -1418 578656
rect -1974 578100 -1738 578336
rect -1654 578100 -1418 578336
rect -1974 542420 -1738 542656
rect -1654 542420 -1418 542656
rect -1974 542100 -1738 542336
rect -1654 542100 -1418 542336
rect -1974 506420 -1738 506656
rect -1654 506420 -1418 506656
rect -1974 506100 -1738 506336
rect -1654 506100 -1418 506336
rect -1974 470420 -1738 470656
rect -1654 470420 -1418 470656
rect -1974 470100 -1738 470336
rect -1654 470100 -1418 470336
rect -1974 434420 -1738 434656
rect -1654 434420 -1418 434656
rect -1974 434100 -1738 434336
rect -1654 434100 -1418 434336
rect -1974 398420 -1738 398656
rect -1654 398420 -1418 398656
rect -1974 398100 -1738 398336
rect -1654 398100 -1418 398336
rect -1974 362420 -1738 362656
rect -1654 362420 -1418 362656
rect -1974 362100 -1738 362336
rect -1654 362100 -1418 362336
rect -1974 326420 -1738 326656
rect -1654 326420 -1418 326656
rect -1974 326100 -1738 326336
rect -1654 326100 -1418 326336
rect -1974 290420 -1738 290656
rect -1654 290420 -1418 290656
rect -1974 290100 -1738 290336
rect -1654 290100 -1418 290336
rect -1974 254420 -1738 254656
rect -1654 254420 -1418 254656
rect -1974 254100 -1738 254336
rect -1654 254100 -1418 254336
rect -1974 218420 -1738 218656
rect -1654 218420 -1418 218656
rect -1974 218100 -1738 218336
rect -1654 218100 -1418 218336
rect -1974 182420 -1738 182656
rect -1654 182420 -1418 182656
rect -1974 182100 -1738 182336
rect -1654 182100 -1418 182336
rect -1974 146420 -1738 146656
rect -1654 146420 -1418 146656
rect -1974 146100 -1738 146336
rect -1654 146100 -1418 146336
rect -1974 110420 -1738 110656
rect -1654 110420 -1418 110656
rect -1974 110100 -1738 110336
rect -1654 110100 -1418 110336
rect -1974 74420 -1738 74656
rect -1654 74420 -1418 74656
rect -1974 74100 -1738 74336
rect -1654 74100 -1418 74336
rect -1974 38420 -1738 38656
rect -1654 38420 -1418 38656
rect -1974 38100 -1738 38336
rect -1654 38100 -1418 38336
rect -1974 2420 -1738 2656
rect -1654 2420 -1418 2656
rect -1974 2100 -1738 2336
rect -1654 2100 -1418 2336
rect -1974 -580 -1738 -344
rect -1654 -580 -1418 -344
rect -1974 -900 -1738 -664
rect -1654 -900 -1418 -664
rect 1026 704604 1262 704840
rect 1346 704604 1582 704840
rect 1026 704284 1262 704520
rect 1346 704284 1582 704520
rect 1026 686420 1262 686656
rect 1346 686420 1582 686656
rect 1026 686100 1262 686336
rect 1346 686100 1582 686336
rect 1026 650420 1262 650656
rect 1346 650420 1582 650656
rect 1026 650100 1262 650336
rect 1346 650100 1582 650336
rect 1026 614420 1262 614656
rect 1346 614420 1582 614656
rect 1026 614100 1262 614336
rect 1346 614100 1582 614336
rect 1026 578420 1262 578656
rect 1346 578420 1582 578656
rect 1026 578100 1262 578336
rect 1346 578100 1582 578336
rect 1026 542420 1262 542656
rect 1346 542420 1582 542656
rect 1026 542100 1262 542336
rect 1346 542100 1582 542336
rect 1026 506420 1262 506656
rect 1346 506420 1582 506656
rect 1026 506100 1262 506336
rect 1346 506100 1582 506336
rect 1026 470420 1262 470656
rect 1346 470420 1582 470656
rect 1026 470100 1262 470336
rect 1346 470100 1582 470336
rect 1026 434420 1262 434656
rect 1346 434420 1582 434656
rect 1026 434100 1262 434336
rect 1346 434100 1582 434336
rect 1026 398420 1262 398656
rect 1346 398420 1582 398656
rect 1026 398100 1262 398336
rect 1346 398100 1582 398336
rect 1026 362420 1262 362656
rect 1346 362420 1582 362656
rect 1026 362100 1262 362336
rect 1346 362100 1582 362336
rect 1026 326420 1262 326656
rect 1346 326420 1582 326656
rect 1026 326100 1262 326336
rect 1346 326100 1582 326336
rect 1026 290420 1262 290656
rect 1346 290420 1582 290656
rect 1026 290100 1262 290336
rect 1346 290100 1582 290336
rect 1026 254420 1262 254656
rect 1346 254420 1582 254656
rect 1026 254100 1262 254336
rect 1346 254100 1582 254336
rect 1026 218420 1262 218656
rect 1346 218420 1582 218656
rect 1026 218100 1262 218336
rect 1346 218100 1582 218336
rect 1026 182420 1262 182656
rect 1346 182420 1582 182656
rect 1026 182100 1262 182336
rect 1346 182100 1582 182336
rect 1026 146420 1262 146656
rect 1346 146420 1582 146656
rect 1026 146100 1262 146336
rect 1346 146100 1582 146336
rect 1026 110420 1262 110656
rect 1346 110420 1582 110656
rect 1026 110100 1262 110336
rect 1346 110100 1582 110336
rect 1026 74420 1262 74656
rect 1346 74420 1582 74656
rect 1026 74100 1262 74336
rect 1346 74100 1582 74336
rect 1026 38420 1262 38656
rect 1346 38420 1582 38656
rect 1026 38100 1262 38336
rect 1346 38100 1582 38336
rect 1026 2420 1262 2656
rect 1346 2420 1582 2656
rect 1026 2100 1262 2336
rect 1346 2100 1582 2336
rect 1026 -580 1262 -344
rect 1346 -580 1582 -344
rect 1026 -900 1262 -664
rect 1346 -900 1582 -664
rect -2934 -1540 -2698 -1304
rect -2614 -1540 -2378 -1304
rect -2934 -1860 -2698 -1624
rect -2614 -1860 -2378 -1624
rect -3894 -2500 -3658 -2264
rect -3574 -2500 -3338 -2264
rect -3894 -2820 -3658 -2584
rect -3574 -2820 -3338 -2584
rect -4854 -3460 -4618 -3224
rect -4534 -3460 -4298 -3224
rect -4854 -3780 -4618 -3544
rect -4534 -3780 -4298 -3544
rect -5814 -4420 -5578 -4184
rect -5494 -4420 -5258 -4184
rect -5814 -4740 -5578 -4504
rect -5494 -4740 -5258 -4504
rect -6774 -5380 -6538 -5144
rect -6454 -5380 -6218 -5144
rect -6774 -5700 -6538 -5464
rect -6454 -5700 -6218 -5464
rect -7734 -6340 -7498 -6104
rect -7414 -6340 -7178 -6104
rect -7734 -6660 -7498 -6424
rect -7414 -6660 -7178 -6424
rect -8694 -7300 -8458 -7064
rect -8374 -7300 -8138 -7064
rect -8694 -7620 -8458 -7384
rect -8374 -7620 -8138 -7384
rect 2266 705564 2502 705800
rect 2586 705564 2822 705800
rect 2266 705244 2502 705480
rect 2586 705244 2822 705480
rect 2266 687660 2502 687896
rect 2586 687660 2822 687896
rect 2266 687340 2502 687576
rect 2586 687340 2822 687576
rect 2266 651660 2502 651896
rect 2586 651660 2822 651896
rect 2266 651340 2502 651576
rect 2586 651340 2822 651576
rect 2266 615660 2502 615896
rect 2586 615660 2822 615896
rect 2266 615340 2502 615576
rect 2586 615340 2822 615576
rect 2266 579660 2502 579896
rect 2586 579660 2822 579896
rect 2266 579340 2502 579576
rect 2586 579340 2822 579576
rect 2266 543660 2502 543896
rect 2586 543660 2822 543896
rect 2266 543340 2502 543576
rect 2586 543340 2822 543576
rect 2266 507660 2502 507896
rect 2586 507660 2822 507896
rect 2266 507340 2502 507576
rect 2586 507340 2822 507576
rect 2266 471660 2502 471896
rect 2586 471660 2822 471896
rect 2266 471340 2502 471576
rect 2586 471340 2822 471576
rect 2266 435660 2502 435896
rect 2586 435660 2822 435896
rect 2266 435340 2502 435576
rect 2586 435340 2822 435576
rect 2266 399660 2502 399896
rect 2586 399660 2822 399896
rect 2266 399340 2502 399576
rect 2586 399340 2822 399576
rect 2266 363660 2502 363896
rect 2586 363660 2822 363896
rect 2266 363340 2502 363576
rect 2586 363340 2822 363576
rect 2266 327660 2502 327896
rect 2586 327660 2822 327896
rect 2266 327340 2502 327576
rect 2586 327340 2822 327576
rect 2266 291660 2502 291896
rect 2586 291660 2822 291896
rect 2266 291340 2502 291576
rect 2586 291340 2822 291576
rect 2266 255660 2502 255896
rect 2586 255660 2822 255896
rect 2266 255340 2502 255576
rect 2586 255340 2822 255576
rect 2266 219660 2502 219896
rect 2586 219660 2822 219896
rect 2266 219340 2502 219576
rect 2586 219340 2822 219576
rect 2266 183660 2502 183896
rect 2586 183660 2822 183896
rect 2266 183340 2502 183576
rect 2586 183340 2822 183576
rect 2266 147660 2502 147896
rect 2586 147660 2822 147896
rect 2266 147340 2502 147576
rect 2586 147340 2822 147576
rect 2266 111660 2502 111896
rect 2586 111660 2822 111896
rect 2266 111340 2502 111576
rect 2586 111340 2822 111576
rect 2266 75660 2502 75896
rect 2586 75660 2822 75896
rect 2266 75340 2502 75576
rect 2586 75340 2822 75576
rect 2266 39660 2502 39896
rect 2586 39660 2822 39896
rect 2266 39340 2502 39576
rect 2586 39340 2822 39576
rect 2266 3660 2502 3896
rect 2586 3660 2822 3896
rect 2266 3340 2502 3576
rect 2586 3340 2822 3576
rect 2266 -1540 2502 -1304
rect 2586 -1540 2822 -1304
rect 2266 -1860 2502 -1624
rect 2586 -1860 2822 -1624
rect 3506 706524 3742 706760
rect 3826 706524 4062 706760
rect 3506 706204 3742 706440
rect 3826 706204 4062 706440
rect 3506 688900 3742 689136
rect 3826 688900 4062 689136
rect 3506 688580 3742 688816
rect 3826 688580 4062 688816
rect 3506 652900 3742 653136
rect 3826 652900 4062 653136
rect 3506 652580 3742 652816
rect 3826 652580 4062 652816
rect 3506 616900 3742 617136
rect 3826 616900 4062 617136
rect 3506 616580 3742 616816
rect 3826 616580 4062 616816
rect 3506 580900 3742 581136
rect 3826 580900 4062 581136
rect 3506 580580 3742 580816
rect 3826 580580 4062 580816
rect 3506 544900 3742 545136
rect 3826 544900 4062 545136
rect 3506 544580 3742 544816
rect 3826 544580 4062 544816
rect 3506 508900 3742 509136
rect 3826 508900 4062 509136
rect 3506 508580 3742 508816
rect 3826 508580 4062 508816
rect 3506 472900 3742 473136
rect 3826 472900 4062 473136
rect 3506 472580 3742 472816
rect 3826 472580 4062 472816
rect 3506 436900 3742 437136
rect 3826 436900 4062 437136
rect 3506 436580 3742 436816
rect 3826 436580 4062 436816
rect 3506 400900 3742 401136
rect 3826 400900 4062 401136
rect 3506 400580 3742 400816
rect 3826 400580 4062 400816
rect 3506 364900 3742 365136
rect 3826 364900 4062 365136
rect 3506 364580 3742 364816
rect 3826 364580 4062 364816
rect 3506 328900 3742 329136
rect 3826 328900 4062 329136
rect 3506 328580 3742 328816
rect 3826 328580 4062 328816
rect 3506 292900 3742 293136
rect 3826 292900 4062 293136
rect 3506 292580 3742 292816
rect 3826 292580 4062 292816
rect 3506 256900 3742 257136
rect 3826 256900 4062 257136
rect 3506 256580 3742 256816
rect 3826 256580 4062 256816
rect 3506 220900 3742 221136
rect 3826 220900 4062 221136
rect 3506 220580 3742 220816
rect 3826 220580 4062 220816
rect 3506 184900 3742 185136
rect 3826 184900 4062 185136
rect 3506 184580 3742 184816
rect 3826 184580 4062 184816
rect 3506 148900 3742 149136
rect 3826 148900 4062 149136
rect 3506 148580 3742 148816
rect 3826 148580 4062 148816
rect 3506 112900 3742 113136
rect 3826 112900 4062 113136
rect 3506 112580 3742 112816
rect 3826 112580 4062 112816
rect 3506 76900 3742 77136
rect 3826 76900 4062 77136
rect 3506 76580 3742 76816
rect 3826 76580 4062 76816
rect 3506 40900 3742 41136
rect 3826 40900 4062 41136
rect 3506 40580 3742 40816
rect 3826 40580 4062 40816
rect 3506 4900 3742 5136
rect 3826 4900 4062 5136
rect 3506 4580 3742 4816
rect 3826 4580 4062 4816
rect 3506 -2500 3742 -2264
rect 3826 -2500 4062 -2264
rect 3506 -2820 3742 -2584
rect 3826 -2820 4062 -2584
rect 4746 707484 4982 707720
rect 5066 707484 5302 707720
rect 4746 707164 4982 707400
rect 5066 707164 5302 707400
rect 4746 690140 4982 690376
rect 5066 690140 5302 690376
rect 4746 689820 4982 690056
rect 5066 689820 5302 690056
rect 4746 654140 4982 654376
rect 5066 654140 5302 654376
rect 4746 653820 4982 654056
rect 5066 653820 5302 654056
rect 4746 618140 4982 618376
rect 5066 618140 5302 618376
rect 4746 617820 4982 618056
rect 5066 617820 5302 618056
rect 4746 582140 4982 582376
rect 5066 582140 5302 582376
rect 4746 581820 4982 582056
rect 5066 581820 5302 582056
rect 4746 546140 4982 546376
rect 5066 546140 5302 546376
rect 4746 545820 4982 546056
rect 5066 545820 5302 546056
rect 4746 510140 4982 510376
rect 5066 510140 5302 510376
rect 4746 509820 4982 510056
rect 5066 509820 5302 510056
rect 4746 474140 4982 474376
rect 5066 474140 5302 474376
rect 4746 473820 4982 474056
rect 5066 473820 5302 474056
rect 4746 438140 4982 438376
rect 5066 438140 5302 438376
rect 4746 437820 4982 438056
rect 5066 437820 5302 438056
rect 4746 402140 4982 402376
rect 5066 402140 5302 402376
rect 4746 401820 4982 402056
rect 5066 401820 5302 402056
rect 4746 366140 4982 366376
rect 5066 366140 5302 366376
rect 4746 365820 4982 366056
rect 5066 365820 5302 366056
rect 4746 330140 4982 330376
rect 5066 330140 5302 330376
rect 4746 329820 4982 330056
rect 5066 329820 5302 330056
rect 4746 294140 4982 294376
rect 5066 294140 5302 294376
rect 4746 293820 4982 294056
rect 5066 293820 5302 294056
rect 4746 258140 4982 258376
rect 5066 258140 5302 258376
rect 4746 257820 4982 258056
rect 5066 257820 5302 258056
rect 4746 222140 4982 222376
rect 5066 222140 5302 222376
rect 4746 221820 4982 222056
rect 5066 221820 5302 222056
rect 4746 186140 4982 186376
rect 5066 186140 5302 186376
rect 4746 185820 4982 186056
rect 5066 185820 5302 186056
rect 4746 150140 4982 150376
rect 5066 150140 5302 150376
rect 4746 149820 4982 150056
rect 5066 149820 5302 150056
rect 4746 114140 4982 114376
rect 5066 114140 5302 114376
rect 4746 113820 4982 114056
rect 5066 113820 5302 114056
rect 4746 78140 4982 78376
rect 5066 78140 5302 78376
rect 4746 77820 4982 78056
rect 5066 77820 5302 78056
rect 4746 42140 4982 42376
rect 5066 42140 5302 42376
rect 4746 41820 4982 42056
rect 5066 41820 5302 42056
rect 4746 6140 4982 6376
rect 5066 6140 5302 6376
rect 4746 5820 4982 6056
rect 5066 5820 5302 6056
rect 4746 -3460 4982 -3224
rect 5066 -3460 5302 -3224
rect 4746 -3780 4982 -3544
rect 5066 -3780 5302 -3544
rect 5986 708444 6222 708680
rect 6306 708444 6542 708680
rect 5986 708124 6222 708360
rect 6306 708124 6542 708360
rect 5986 691380 6222 691616
rect 6306 691380 6542 691616
rect 5986 691060 6222 691296
rect 6306 691060 6542 691296
rect 5986 655380 6222 655616
rect 6306 655380 6542 655616
rect 5986 655060 6222 655296
rect 6306 655060 6542 655296
rect 5986 619380 6222 619616
rect 6306 619380 6542 619616
rect 5986 619060 6222 619296
rect 6306 619060 6542 619296
rect 5986 583380 6222 583616
rect 6306 583380 6542 583616
rect 5986 583060 6222 583296
rect 6306 583060 6542 583296
rect 5986 547380 6222 547616
rect 6306 547380 6542 547616
rect 5986 547060 6222 547296
rect 6306 547060 6542 547296
rect 5986 511380 6222 511616
rect 6306 511380 6542 511616
rect 5986 511060 6222 511296
rect 6306 511060 6542 511296
rect 5986 475380 6222 475616
rect 6306 475380 6542 475616
rect 5986 475060 6222 475296
rect 6306 475060 6542 475296
rect 5986 439380 6222 439616
rect 6306 439380 6542 439616
rect 5986 439060 6222 439296
rect 6306 439060 6542 439296
rect 5986 403380 6222 403616
rect 6306 403380 6542 403616
rect 5986 403060 6222 403296
rect 6306 403060 6542 403296
rect 5986 367380 6222 367616
rect 6306 367380 6542 367616
rect 5986 367060 6222 367296
rect 6306 367060 6542 367296
rect 5986 331380 6222 331616
rect 6306 331380 6542 331616
rect 5986 331060 6222 331296
rect 6306 331060 6542 331296
rect 5986 295380 6222 295616
rect 6306 295380 6542 295616
rect 5986 295060 6222 295296
rect 6306 295060 6542 295296
rect 5986 259380 6222 259616
rect 6306 259380 6542 259616
rect 5986 259060 6222 259296
rect 6306 259060 6542 259296
rect 5986 223380 6222 223616
rect 6306 223380 6542 223616
rect 5986 223060 6222 223296
rect 6306 223060 6542 223296
rect 5986 187380 6222 187616
rect 6306 187380 6542 187616
rect 5986 187060 6222 187296
rect 6306 187060 6542 187296
rect 5986 151380 6222 151616
rect 6306 151380 6542 151616
rect 5986 151060 6222 151296
rect 6306 151060 6542 151296
rect 5986 115380 6222 115616
rect 6306 115380 6542 115616
rect 5986 115060 6222 115296
rect 6306 115060 6542 115296
rect 5986 79380 6222 79616
rect 6306 79380 6542 79616
rect 5986 79060 6222 79296
rect 6306 79060 6542 79296
rect 5986 43380 6222 43616
rect 6306 43380 6542 43616
rect 5986 43060 6222 43296
rect 6306 43060 6542 43296
rect 5986 7380 6222 7616
rect 6306 7380 6542 7616
rect 5986 7060 6222 7296
rect 6306 7060 6542 7296
rect 5986 -4420 6222 -4184
rect 6306 -4420 6542 -4184
rect 5986 -4740 6222 -4504
rect 6306 -4740 6542 -4504
rect 7226 709404 7462 709640
rect 7546 709404 7782 709640
rect 7226 709084 7462 709320
rect 7546 709084 7782 709320
rect 7226 692620 7462 692856
rect 7546 692620 7782 692856
rect 7226 692300 7462 692536
rect 7546 692300 7782 692536
rect 7226 656620 7462 656856
rect 7546 656620 7782 656856
rect 7226 656300 7462 656536
rect 7546 656300 7782 656536
rect 7226 620620 7462 620856
rect 7546 620620 7782 620856
rect 7226 620300 7462 620536
rect 7546 620300 7782 620536
rect 7226 584620 7462 584856
rect 7546 584620 7782 584856
rect 7226 584300 7462 584536
rect 7546 584300 7782 584536
rect 7226 548620 7462 548856
rect 7546 548620 7782 548856
rect 7226 548300 7462 548536
rect 7546 548300 7782 548536
rect 7226 512620 7462 512856
rect 7546 512620 7782 512856
rect 7226 512300 7462 512536
rect 7546 512300 7782 512536
rect 7226 476620 7462 476856
rect 7546 476620 7782 476856
rect 7226 476300 7462 476536
rect 7546 476300 7782 476536
rect 7226 440620 7462 440856
rect 7546 440620 7782 440856
rect 7226 440300 7462 440536
rect 7546 440300 7782 440536
rect 7226 404620 7462 404856
rect 7546 404620 7782 404856
rect 7226 404300 7462 404536
rect 7546 404300 7782 404536
rect 7226 368620 7462 368856
rect 7546 368620 7782 368856
rect 7226 368300 7462 368536
rect 7546 368300 7782 368536
rect 7226 332620 7462 332856
rect 7546 332620 7782 332856
rect 7226 332300 7462 332536
rect 7546 332300 7782 332536
rect 7226 296620 7462 296856
rect 7546 296620 7782 296856
rect 7226 296300 7462 296536
rect 7546 296300 7782 296536
rect 7226 260620 7462 260856
rect 7546 260620 7782 260856
rect 7226 260300 7462 260536
rect 7546 260300 7782 260536
rect 7226 224620 7462 224856
rect 7546 224620 7782 224856
rect 7226 224300 7462 224536
rect 7546 224300 7782 224536
rect 7226 188620 7462 188856
rect 7546 188620 7782 188856
rect 7226 188300 7462 188536
rect 7546 188300 7782 188536
rect 7226 152620 7462 152856
rect 7546 152620 7782 152856
rect 7226 152300 7462 152536
rect 7546 152300 7782 152536
rect 7226 116620 7462 116856
rect 7546 116620 7782 116856
rect 7226 116300 7462 116536
rect 7546 116300 7782 116536
rect 7226 80620 7462 80856
rect 7546 80620 7782 80856
rect 7226 80300 7462 80536
rect 7546 80300 7782 80536
rect 7226 44620 7462 44856
rect 7546 44620 7782 44856
rect 7226 44300 7462 44536
rect 7546 44300 7782 44536
rect 7226 8620 7462 8856
rect 7546 8620 7782 8856
rect 7226 8300 7462 8536
rect 7546 8300 7782 8536
rect 7226 -5380 7462 -5144
rect 7546 -5380 7782 -5144
rect 7226 -5700 7462 -5464
rect 7546 -5700 7782 -5464
rect 8466 710364 8702 710600
rect 8786 710364 9022 710600
rect 8466 710044 8702 710280
rect 8786 710044 9022 710280
rect 8466 693860 8702 694096
rect 8786 693860 9022 694096
rect 8466 693540 8702 693776
rect 8786 693540 9022 693776
rect 8466 657860 8702 658096
rect 8786 657860 9022 658096
rect 8466 657540 8702 657776
rect 8786 657540 9022 657776
rect 8466 621860 8702 622096
rect 8786 621860 9022 622096
rect 8466 621540 8702 621776
rect 8786 621540 9022 621776
rect 8466 585860 8702 586096
rect 8786 585860 9022 586096
rect 8466 585540 8702 585776
rect 8786 585540 9022 585776
rect 8466 549860 8702 550096
rect 8786 549860 9022 550096
rect 8466 549540 8702 549776
rect 8786 549540 9022 549776
rect 8466 513860 8702 514096
rect 8786 513860 9022 514096
rect 8466 513540 8702 513776
rect 8786 513540 9022 513776
rect 8466 477860 8702 478096
rect 8786 477860 9022 478096
rect 8466 477540 8702 477776
rect 8786 477540 9022 477776
rect 8466 441860 8702 442096
rect 8786 441860 9022 442096
rect 8466 441540 8702 441776
rect 8786 441540 9022 441776
rect 8466 405860 8702 406096
rect 8786 405860 9022 406096
rect 8466 405540 8702 405776
rect 8786 405540 9022 405776
rect 8466 369860 8702 370096
rect 8786 369860 9022 370096
rect 8466 369540 8702 369776
rect 8786 369540 9022 369776
rect 8466 333860 8702 334096
rect 8786 333860 9022 334096
rect 8466 333540 8702 333776
rect 8786 333540 9022 333776
rect 8466 297860 8702 298096
rect 8786 297860 9022 298096
rect 8466 297540 8702 297776
rect 8786 297540 9022 297776
rect 8466 261860 8702 262096
rect 8786 261860 9022 262096
rect 8466 261540 8702 261776
rect 8786 261540 9022 261776
rect 8466 225860 8702 226096
rect 8786 225860 9022 226096
rect 8466 225540 8702 225776
rect 8786 225540 9022 225776
rect 8466 189860 8702 190096
rect 8786 189860 9022 190096
rect 8466 189540 8702 189776
rect 8786 189540 9022 189776
rect 8466 153860 8702 154096
rect 8786 153860 9022 154096
rect 8466 153540 8702 153776
rect 8786 153540 9022 153776
rect 8466 117860 8702 118096
rect 8786 117860 9022 118096
rect 8466 117540 8702 117776
rect 8786 117540 9022 117776
rect 8466 81860 8702 82096
rect 8786 81860 9022 82096
rect 8466 81540 8702 81776
rect 8786 81540 9022 81776
rect 8466 45860 8702 46096
rect 8786 45860 9022 46096
rect 8466 45540 8702 45776
rect 8786 45540 9022 45776
rect 8466 9860 8702 10096
rect 8786 9860 9022 10096
rect 8466 9540 8702 9776
rect 8786 9540 9022 9776
rect 8466 -6340 8702 -6104
rect 8786 -6340 9022 -6104
rect 8466 -6660 8702 -6424
rect 8786 -6660 9022 -6424
rect 9706 711324 9942 711560
rect 10026 711324 10262 711560
rect 9706 711004 9942 711240
rect 10026 711004 10262 711240
rect 9706 695100 9942 695336
rect 10026 695100 10262 695336
rect 9706 694780 9942 695016
rect 10026 694780 10262 695016
rect 9706 659100 9942 659336
rect 10026 659100 10262 659336
rect 9706 658780 9942 659016
rect 10026 658780 10262 659016
rect 9706 623100 9942 623336
rect 10026 623100 10262 623336
rect 9706 622780 9942 623016
rect 10026 622780 10262 623016
rect 9706 587100 9942 587336
rect 10026 587100 10262 587336
rect 9706 586780 9942 587016
rect 10026 586780 10262 587016
rect 9706 551100 9942 551336
rect 10026 551100 10262 551336
rect 9706 550780 9942 551016
rect 10026 550780 10262 551016
rect 9706 515100 9942 515336
rect 10026 515100 10262 515336
rect 9706 514780 9942 515016
rect 10026 514780 10262 515016
rect 9706 479100 9942 479336
rect 10026 479100 10262 479336
rect 9706 478780 9942 479016
rect 10026 478780 10262 479016
rect 9706 443100 9942 443336
rect 10026 443100 10262 443336
rect 9706 442780 9942 443016
rect 10026 442780 10262 443016
rect 9706 407100 9942 407336
rect 10026 407100 10262 407336
rect 9706 406780 9942 407016
rect 10026 406780 10262 407016
rect 9706 371100 9942 371336
rect 10026 371100 10262 371336
rect 9706 370780 9942 371016
rect 10026 370780 10262 371016
rect 9706 335100 9942 335336
rect 10026 335100 10262 335336
rect 9706 334780 9942 335016
rect 10026 334780 10262 335016
rect 9706 299100 9942 299336
rect 10026 299100 10262 299336
rect 9706 298780 9942 299016
rect 10026 298780 10262 299016
rect 9706 263100 9942 263336
rect 10026 263100 10262 263336
rect 9706 262780 9942 263016
rect 10026 262780 10262 263016
rect 9706 227100 9942 227336
rect 10026 227100 10262 227336
rect 9706 226780 9942 227016
rect 10026 226780 10262 227016
rect 9706 191100 9942 191336
rect 10026 191100 10262 191336
rect 9706 190780 9942 191016
rect 10026 190780 10262 191016
rect 9706 155100 9942 155336
rect 10026 155100 10262 155336
rect 9706 154780 9942 155016
rect 10026 154780 10262 155016
rect 9706 119100 9942 119336
rect 10026 119100 10262 119336
rect 9706 118780 9942 119016
rect 10026 118780 10262 119016
rect 9706 83100 9942 83336
rect 10026 83100 10262 83336
rect 9706 82780 9942 83016
rect 10026 82780 10262 83016
rect 9706 47100 9942 47336
rect 10026 47100 10262 47336
rect 9706 46780 9942 47016
rect 10026 46780 10262 47016
rect 9706 11100 9942 11336
rect 10026 11100 10262 11336
rect 9706 10780 9942 11016
rect 10026 10780 10262 11016
rect 9706 -7300 9942 -7064
rect 10026 -7300 10262 -7064
rect 9706 -7620 9942 -7384
rect 10026 -7620 10262 -7384
rect 37026 704604 37262 704840
rect 37346 704604 37582 704840
rect 37026 704284 37262 704520
rect 37346 704284 37582 704520
rect 37026 686420 37262 686656
rect 37346 686420 37582 686656
rect 37026 686100 37262 686336
rect 37346 686100 37582 686336
rect 37026 650420 37262 650656
rect 37346 650420 37582 650656
rect 37026 650100 37262 650336
rect 37346 650100 37582 650336
rect 37026 614420 37262 614656
rect 37346 614420 37582 614656
rect 37026 614100 37262 614336
rect 37346 614100 37582 614336
rect 37026 578420 37262 578656
rect 37346 578420 37582 578656
rect 37026 578100 37262 578336
rect 37346 578100 37582 578336
rect 37026 542420 37262 542656
rect 37346 542420 37582 542656
rect 37026 542100 37262 542336
rect 37346 542100 37582 542336
rect 37026 506420 37262 506656
rect 37346 506420 37582 506656
rect 37026 506100 37262 506336
rect 37346 506100 37582 506336
rect 37026 470420 37262 470656
rect 37346 470420 37582 470656
rect 37026 470100 37262 470336
rect 37346 470100 37582 470336
rect 37026 434420 37262 434656
rect 37346 434420 37582 434656
rect 37026 434100 37262 434336
rect 37346 434100 37582 434336
rect 37026 398420 37262 398656
rect 37346 398420 37582 398656
rect 37026 398100 37262 398336
rect 37346 398100 37582 398336
rect 37026 362420 37262 362656
rect 37346 362420 37582 362656
rect 37026 362100 37262 362336
rect 37346 362100 37582 362336
rect 37026 326420 37262 326656
rect 37346 326420 37582 326656
rect 37026 326100 37262 326336
rect 37346 326100 37582 326336
rect 37026 290420 37262 290656
rect 37346 290420 37582 290656
rect 37026 290100 37262 290336
rect 37346 290100 37582 290336
rect 37026 254420 37262 254656
rect 37346 254420 37582 254656
rect 37026 254100 37262 254336
rect 37346 254100 37582 254336
rect 37026 218420 37262 218656
rect 37346 218420 37582 218656
rect 37026 218100 37262 218336
rect 37346 218100 37582 218336
rect 37026 182420 37262 182656
rect 37346 182420 37582 182656
rect 37026 182100 37262 182336
rect 37346 182100 37582 182336
rect 37026 146420 37262 146656
rect 37346 146420 37582 146656
rect 37026 146100 37262 146336
rect 37346 146100 37582 146336
rect 37026 110420 37262 110656
rect 37346 110420 37582 110656
rect 37026 110100 37262 110336
rect 37346 110100 37582 110336
rect 37026 74420 37262 74656
rect 37346 74420 37582 74656
rect 37026 74100 37262 74336
rect 37346 74100 37582 74336
rect 37026 38420 37262 38656
rect 37346 38420 37582 38656
rect 37026 38100 37262 38336
rect 37346 38100 37582 38336
rect 37026 2420 37262 2656
rect 37346 2420 37582 2656
rect 37026 2100 37262 2336
rect 37346 2100 37582 2336
rect 37026 -580 37262 -344
rect 37346 -580 37582 -344
rect 37026 -900 37262 -664
rect 37346 -900 37582 -664
rect 38266 705564 38502 705800
rect 38586 705564 38822 705800
rect 38266 705244 38502 705480
rect 38586 705244 38822 705480
rect 38266 687660 38502 687896
rect 38586 687660 38822 687896
rect 38266 687340 38502 687576
rect 38586 687340 38822 687576
rect 38266 651660 38502 651896
rect 38586 651660 38822 651896
rect 38266 651340 38502 651576
rect 38586 651340 38822 651576
rect 38266 615660 38502 615896
rect 38586 615660 38822 615896
rect 38266 615340 38502 615576
rect 38586 615340 38822 615576
rect 38266 579660 38502 579896
rect 38586 579660 38822 579896
rect 38266 579340 38502 579576
rect 38586 579340 38822 579576
rect 38266 543660 38502 543896
rect 38586 543660 38822 543896
rect 38266 543340 38502 543576
rect 38586 543340 38822 543576
rect 38266 507660 38502 507896
rect 38586 507660 38822 507896
rect 38266 507340 38502 507576
rect 38586 507340 38822 507576
rect 38266 471660 38502 471896
rect 38586 471660 38822 471896
rect 38266 471340 38502 471576
rect 38586 471340 38822 471576
rect 38266 435660 38502 435896
rect 38586 435660 38822 435896
rect 38266 435340 38502 435576
rect 38586 435340 38822 435576
rect 38266 399660 38502 399896
rect 38586 399660 38822 399896
rect 38266 399340 38502 399576
rect 38586 399340 38822 399576
rect 38266 363660 38502 363896
rect 38586 363660 38822 363896
rect 38266 363340 38502 363576
rect 38586 363340 38822 363576
rect 38266 327660 38502 327896
rect 38586 327660 38822 327896
rect 38266 327340 38502 327576
rect 38586 327340 38822 327576
rect 38266 291660 38502 291896
rect 38586 291660 38822 291896
rect 38266 291340 38502 291576
rect 38586 291340 38822 291576
rect 38266 255660 38502 255896
rect 38586 255660 38822 255896
rect 38266 255340 38502 255576
rect 38586 255340 38822 255576
rect 38266 219660 38502 219896
rect 38586 219660 38822 219896
rect 38266 219340 38502 219576
rect 38586 219340 38822 219576
rect 38266 183660 38502 183896
rect 38586 183660 38822 183896
rect 38266 183340 38502 183576
rect 38586 183340 38822 183576
rect 38266 147660 38502 147896
rect 38586 147660 38822 147896
rect 38266 147340 38502 147576
rect 38586 147340 38822 147576
rect 38266 111660 38502 111896
rect 38586 111660 38822 111896
rect 38266 111340 38502 111576
rect 38586 111340 38822 111576
rect 38266 75660 38502 75896
rect 38586 75660 38822 75896
rect 38266 75340 38502 75576
rect 38586 75340 38822 75576
rect 38266 39660 38502 39896
rect 38586 39660 38822 39896
rect 38266 39340 38502 39576
rect 38586 39340 38822 39576
rect 38266 3660 38502 3896
rect 38586 3660 38822 3896
rect 38266 3340 38502 3576
rect 38586 3340 38822 3576
rect 38266 -1540 38502 -1304
rect 38586 -1540 38822 -1304
rect 38266 -1860 38502 -1624
rect 38586 -1860 38822 -1624
rect 39506 706524 39742 706760
rect 39826 706524 40062 706760
rect 39506 706204 39742 706440
rect 39826 706204 40062 706440
rect 39506 688900 39742 689136
rect 39826 688900 40062 689136
rect 39506 688580 39742 688816
rect 39826 688580 40062 688816
rect 39506 652900 39742 653136
rect 39826 652900 40062 653136
rect 39506 652580 39742 652816
rect 39826 652580 40062 652816
rect 39506 616900 39742 617136
rect 39826 616900 40062 617136
rect 39506 616580 39742 616816
rect 39826 616580 40062 616816
rect 39506 580900 39742 581136
rect 39826 580900 40062 581136
rect 39506 580580 39742 580816
rect 39826 580580 40062 580816
rect 39506 544900 39742 545136
rect 39826 544900 40062 545136
rect 39506 544580 39742 544816
rect 39826 544580 40062 544816
rect 39506 508900 39742 509136
rect 39826 508900 40062 509136
rect 39506 508580 39742 508816
rect 39826 508580 40062 508816
rect 39506 472900 39742 473136
rect 39826 472900 40062 473136
rect 39506 472580 39742 472816
rect 39826 472580 40062 472816
rect 39506 436900 39742 437136
rect 39826 436900 40062 437136
rect 39506 436580 39742 436816
rect 39826 436580 40062 436816
rect 39506 400900 39742 401136
rect 39826 400900 40062 401136
rect 39506 400580 39742 400816
rect 39826 400580 40062 400816
rect 39506 364900 39742 365136
rect 39826 364900 40062 365136
rect 39506 364580 39742 364816
rect 39826 364580 40062 364816
rect 39506 328900 39742 329136
rect 39826 328900 40062 329136
rect 39506 328580 39742 328816
rect 39826 328580 40062 328816
rect 39506 292900 39742 293136
rect 39826 292900 40062 293136
rect 39506 292580 39742 292816
rect 39826 292580 40062 292816
rect 39506 256900 39742 257136
rect 39826 256900 40062 257136
rect 39506 256580 39742 256816
rect 39826 256580 40062 256816
rect 39506 220900 39742 221136
rect 39826 220900 40062 221136
rect 39506 220580 39742 220816
rect 39826 220580 40062 220816
rect 39506 184900 39742 185136
rect 39826 184900 40062 185136
rect 39506 184580 39742 184816
rect 39826 184580 40062 184816
rect 39506 148900 39742 149136
rect 39826 148900 40062 149136
rect 39506 148580 39742 148816
rect 39826 148580 40062 148816
rect 39506 112900 39742 113136
rect 39826 112900 40062 113136
rect 39506 112580 39742 112816
rect 39826 112580 40062 112816
rect 39506 76900 39742 77136
rect 39826 76900 40062 77136
rect 39506 76580 39742 76816
rect 39826 76580 40062 76816
rect 39506 40900 39742 41136
rect 39826 40900 40062 41136
rect 39506 40580 39742 40816
rect 39826 40580 40062 40816
rect 39506 4900 39742 5136
rect 39826 4900 40062 5136
rect 39506 4580 39742 4816
rect 39826 4580 40062 4816
rect 39506 -2500 39742 -2264
rect 39826 -2500 40062 -2264
rect 39506 -2820 39742 -2584
rect 39826 -2820 40062 -2584
rect 40746 707484 40982 707720
rect 41066 707484 41302 707720
rect 40746 707164 40982 707400
rect 41066 707164 41302 707400
rect 40746 690140 40982 690376
rect 41066 690140 41302 690376
rect 40746 689820 40982 690056
rect 41066 689820 41302 690056
rect 40746 654140 40982 654376
rect 41066 654140 41302 654376
rect 40746 653820 40982 654056
rect 41066 653820 41302 654056
rect 40746 618140 40982 618376
rect 41066 618140 41302 618376
rect 40746 617820 40982 618056
rect 41066 617820 41302 618056
rect 40746 582140 40982 582376
rect 41066 582140 41302 582376
rect 40746 581820 40982 582056
rect 41066 581820 41302 582056
rect 40746 546140 40982 546376
rect 41066 546140 41302 546376
rect 40746 545820 40982 546056
rect 41066 545820 41302 546056
rect 40746 510140 40982 510376
rect 41066 510140 41302 510376
rect 40746 509820 40982 510056
rect 41066 509820 41302 510056
rect 40746 474140 40982 474376
rect 41066 474140 41302 474376
rect 40746 473820 40982 474056
rect 41066 473820 41302 474056
rect 40746 438140 40982 438376
rect 41066 438140 41302 438376
rect 40746 437820 40982 438056
rect 41066 437820 41302 438056
rect 40746 402140 40982 402376
rect 41066 402140 41302 402376
rect 40746 401820 40982 402056
rect 41066 401820 41302 402056
rect 40746 366140 40982 366376
rect 41066 366140 41302 366376
rect 40746 365820 40982 366056
rect 41066 365820 41302 366056
rect 40746 330140 40982 330376
rect 41066 330140 41302 330376
rect 40746 329820 40982 330056
rect 41066 329820 41302 330056
rect 40746 294140 40982 294376
rect 41066 294140 41302 294376
rect 40746 293820 40982 294056
rect 41066 293820 41302 294056
rect 40746 258140 40982 258376
rect 41066 258140 41302 258376
rect 40746 257820 40982 258056
rect 41066 257820 41302 258056
rect 40746 222140 40982 222376
rect 41066 222140 41302 222376
rect 40746 221820 40982 222056
rect 41066 221820 41302 222056
rect 40746 186140 40982 186376
rect 41066 186140 41302 186376
rect 40746 185820 40982 186056
rect 41066 185820 41302 186056
rect 40746 150140 40982 150376
rect 41066 150140 41302 150376
rect 40746 149820 40982 150056
rect 41066 149820 41302 150056
rect 40746 114140 40982 114376
rect 41066 114140 41302 114376
rect 40746 113820 40982 114056
rect 41066 113820 41302 114056
rect 40746 78140 40982 78376
rect 41066 78140 41302 78376
rect 40746 77820 40982 78056
rect 41066 77820 41302 78056
rect 40746 42140 40982 42376
rect 41066 42140 41302 42376
rect 40746 41820 40982 42056
rect 41066 41820 41302 42056
rect 40746 6140 40982 6376
rect 41066 6140 41302 6376
rect 40746 5820 40982 6056
rect 41066 5820 41302 6056
rect 40746 -3460 40982 -3224
rect 41066 -3460 41302 -3224
rect 40746 -3780 40982 -3544
rect 41066 -3780 41302 -3544
rect 41986 708444 42222 708680
rect 42306 708444 42542 708680
rect 41986 708124 42222 708360
rect 42306 708124 42542 708360
rect 41986 691380 42222 691616
rect 42306 691380 42542 691616
rect 41986 691060 42222 691296
rect 42306 691060 42542 691296
rect 41986 655380 42222 655616
rect 42306 655380 42542 655616
rect 41986 655060 42222 655296
rect 42306 655060 42542 655296
rect 41986 619380 42222 619616
rect 42306 619380 42542 619616
rect 41986 619060 42222 619296
rect 42306 619060 42542 619296
rect 41986 583380 42222 583616
rect 42306 583380 42542 583616
rect 41986 583060 42222 583296
rect 42306 583060 42542 583296
rect 41986 547380 42222 547616
rect 42306 547380 42542 547616
rect 41986 547060 42222 547296
rect 42306 547060 42542 547296
rect 41986 511380 42222 511616
rect 42306 511380 42542 511616
rect 41986 511060 42222 511296
rect 42306 511060 42542 511296
rect 41986 475380 42222 475616
rect 42306 475380 42542 475616
rect 41986 475060 42222 475296
rect 42306 475060 42542 475296
rect 41986 439380 42222 439616
rect 42306 439380 42542 439616
rect 41986 439060 42222 439296
rect 42306 439060 42542 439296
rect 41986 403380 42222 403616
rect 42306 403380 42542 403616
rect 41986 403060 42222 403296
rect 42306 403060 42542 403296
rect 41986 367380 42222 367616
rect 42306 367380 42542 367616
rect 41986 367060 42222 367296
rect 42306 367060 42542 367296
rect 41986 331380 42222 331616
rect 42306 331380 42542 331616
rect 41986 331060 42222 331296
rect 42306 331060 42542 331296
rect 41986 295380 42222 295616
rect 42306 295380 42542 295616
rect 41986 295060 42222 295296
rect 42306 295060 42542 295296
rect 41986 259380 42222 259616
rect 42306 259380 42542 259616
rect 41986 259060 42222 259296
rect 42306 259060 42542 259296
rect 41986 223380 42222 223616
rect 42306 223380 42542 223616
rect 41986 223060 42222 223296
rect 42306 223060 42542 223296
rect 41986 187380 42222 187616
rect 42306 187380 42542 187616
rect 41986 187060 42222 187296
rect 42306 187060 42542 187296
rect 41986 151380 42222 151616
rect 42306 151380 42542 151616
rect 41986 151060 42222 151296
rect 42306 151060 42542 151296
rect 41986 115380 42222 115616
rect 42306 115380 42542 115616
rect 41986 115060 42222 115296
rect 42306 115060 42542 115296
rect 41986 79380 42222 79616
rect 42306 79380 42542 79616
rect 41986 79060 42222 79296
rect 42306 79060 42542 79296
rect 41986 43380 42222 43616
rect 42306 43380 42542 43616
rect 41986 43060 42222 43296
rect 42306 43060 42542 43296
rect 41986 7380 42222 7616
rect 42306 7380 42542 7616
rect 41986 7060 42222 7296
rect 42306 7060 42542 7296
rect 41986 -4420 42222 -4184
rect 42306 -4420 42542 -4184
rect 41986 -4740 42222 -4504
rect 42306 -4740 42542 -4504
rect 43226 709404 43462 709640
rect 43546 709404 43782 709640
rect 43226 709084 43462 709320
rect 43546 709084 43782 709320
rect 43226 692620 43462 692856
rect 43546 692620 43782 692856
rect 43226 692300 43462 692536
rect 43546 692300 43782 692536
rect 43226 656620 43462 656856
rect 43546 656620 43782 656856
rect 43226 656300 43462 656536
rect 43546 656300 43782 656536
rect 43226 620620 43462 620856
rect 43546 620620 43782 620856
rect 43226 620300 43462 620536
rect 43546 620300 43782 620536
rect 43226 584620 43462 584856
rect 43546 584620 43782 584856
rect 43226 584300 43462 584536
rect 43546 584300 43782 584536
rect 43226 548620 43462 548856
rect 43546 548620 43782 548856
rect 43226 548300 43462 548536
rect 43546 548300 43782 548536
rect 43226 512620 43462 512856
rect 43546 512620 43782 512856
rect 43226 512300 43462 512536
rect 43546 512300 43782 512536
rect 43226 476620 43462 476856
rect 43546 476620 43782 476856
rect 43226 476300 43462 476536
rect 43546 476300 43782 476536
rect 43226 440620 43462 440856
rect 43546 440620 43782 440856
rect 43226 440300 43462 440536
rect 43546 440300 43782 440536
rect 43226 404620 43462 404856
rect 43546 404620 43782 404856
rect 43226 404300 43462 404536
rect 43546 404300 43782 404536
rect 43226 368620 43462 368856
rect 43546 368620 43782 368856
rect 43226 368300 43462 368536
rect 43546 368300 43782 368536
rect 43226 332620 43462 332856
rect 43546 332620 43782 332856
rect 43226 332300 43462 332536
rect 43546 332300 43782 332536
rect 43226 296620 43462 296856
rect 43546 296620 43782 296856
rect 43226 296300 43462 296536
rect 43546 296300 43782 296536
rect 43226 260620 43462 260856
rect 43546 260620 43782 260856
rect 43226 260300 43462 260536
rect 43546 260300 43782 260536
rect 43226 224620 43462 224856
rect 43546 224620 43782 224856
rect 43226 224300 43462 224536
rect 43546 224300 43782 224536
rect 43226 188620 43462 188856
rect 43546 188620 43782 188856
rect 43226 188300 43462 188536
rect 43546 188300 43782 188536
rect 43226 152620 43462 152856
rect 43546 152620 43782 152856
rect 43226 152300 43462 152536
rect 43546 152300 43782 152536
rect 43226 116620 43462 116856
rect 43546 116620 43782 116856
rect 43226 116300 43462 116536
rect 43546 116300 43782 116536
rect 43226 80620 43462 80856
rect 43546 80620 43782 80856
rect 43226 80300 43462 80536
rect 43546 80300 43782 80536
rect 43226 44620 43462 44856
rect 43546 44620 43782 44856
rect 43226 44300 43462 44536
rect 43546 44300 43782 44536
rect 43226 8620 43462 8856
rect 43546 8620 43782 8856
rect 43226 8300 43462 8536
rect 43546 8300 43782 8536
rect 43226 -5380 43462 -5144
rect 43546 -5380 43782 -5144
rect 43226 -5700 43462 -5464
rect 43546 -5700 43782 -5464
rect 44466 710364 44702 710600
rect 44786 710364 45022 710600
rect 44466 710044 44702 710280
rect 44786 710044 45022 710280
rect 44466 693860 44702 694096
rect 44786 693860 45022 694096
rect 44466 693540 44702 693776
rect 44786 693540 45022 693776
rect 44466 657860 44702 658096
rect 44786 657860 45022 658096
rect 44466 657540 44702 657776
rect 44786 657540 45022 657776
rect 44466 621860 44702 622096
rect 44786 621860 45022 622096
rect 44466 621540 44702 621776
rect 44786 621540 45022 621776
rect 44466 585860 44702 586096
rect 44786 585860 45022 586096
rect 44466 585540 44702 585776
rect 44786 585540 45022 585776
rect 44466 549860 44702 550096
rect 44786 549860 45022 550096
rect 44466 549540 44702 549776
rect 44786 549540 45022 549776
rect 44466 513860 44702 514096
rect 44786 513860 45022 514096
rect 44466 513540 44702 513776
rect 44786 513540 45022 513776
rect 44466 477860 44702 478096
rect 44786 477860 45022 478096
rect 44466 477540 44702 477776
rect 44786 477540 45022 477776
rect 44466 441860 44702 442096
rect 44786 441860 45022 442096
rect 44466 441540 44702 441776
rect 44786 441540 45022 441776
rect 44466 405860 44702 406096
rect 44786 405860 45022 406096
rect 44466 405540 44702 405776
rect 44786 405540 45022 405776
rect 44466 369860 44702 370096
rect 44786 369860 45022 370096
rect 44466 369540 44702 369776
rect 44786 369540 45022 369776
rect 44466 333860 44702 334096
rect 44786 333860 45022 334096
rect 44466 333540 44702 333776
rect 44786 333540 45022 333776
rect 44466 297860 44702 298096
rect 44786 297860 45022 298096
rect 44466 297540 44702 297776
rect 44786 297540 45022 297776
rect 44466 261860 44702 262096
rect 44786 261860 45022 262096
rect 44466 261540 44702 261776
rect 44786 261540 45022 261776
rect 44466 225860 44702 226096
rect 44786 225860 45022 226096
rect 44466 225540 44702 225776
rect 44786 225540 45022 225776
rect 44466 189860 44702 190096
rect 44786 189860 45022 190096
rect 44466 189540 44702 189776
rect 44786 189540 45022 189776
rect 44466 153860 44702 154096
rect 44786 153860 45022 154096
rect 44466 153540 44702 153776
rect 44786 153540 45022 153776
rect 44466 117860 44702 118096
rect 44786 117860 45022 118096
rect 44466 117540 44702 117776
rect 44786 117540 45022 117776
rect 44466 81860 44702 82096
rect 44786 81860 45022 82096
rect 44466 81540 44702 81776
rect 44786 81540 45022 81776
rect 44466 45860 44702 46096
rect 44786 45860 45022 46096
rect 44466 45540 44702 45776
rect 44786 45540 45022 45776
rect 44466 9860 44702 10096
rect 44786 9860 45022 10096
rect 44466 9540 44702 9776
rect 44786 9540 45022 9776
rect 44466 -6340 44702 -6104
rect 44786 -6340 45022 -6104
rect 44466 -6660 44702 -6424
rect 44786 -6660 45022 -6424
rect 45706 711324 45942 711560
rect 46026 711324 46262 711560
rect 45706 711004 45942 711240
rect 46026 711004 46262 711240
rect 45706 695100 45942 695336
rect 46026 695100 46262 695336
rect 45706 694780 45942 695016
rect 46026 694780 46262 695016
rect 45706 659100 45942 659336
rect 46026 659100 46262 659336
rect 45706 658780 45942 659016
rect 46026 658780 46262 659016
rect 45706 623100 45942 623336
rect 46026 623100 46262 623336
rect 45706 622780 45942 623016
rect 46026 622780 46262 623016
rect 45706 587100 45942 587336
rect 46026 587100 46262 587336
rect 45706 586780 45942 587016
rect 46026 586780 46262 587016
rect 45706 551100 45942 551336
rect 46026 551100 46262 551336
rect 45706 550780 45942 551016
rect 46026 550780 46262 551016
rect 45706 515100 45942 515336
rect 46026 515100 46262 515336
rect 45706 514780 45942 515016
rect 46026 514780 46262 515016
rect 45706 479100 45942 479336
rect 46026 479100 46262 479336
rect 45706 478780 45942 479016
rect 46026 478780 46262 479016
rect 45706 443100 45942 443336
rect 46026 443100 46262 443336
rect 45706 442780 45942 443016
rect 46026 442780 46262 443016
rect 45706 407100 45942 407336
rect 46026 407100 46262 407336
rect 45706 406780 45942 407016
rect 46026 406780 46262 407016
rect 45706 371100 45942 371336
rect 46026 371100 46262 371336
rect 45706 370780 45942 371016
rect 46026 370780 46262 371016
rect 45706 335100 45942 335336
rect 46026 335100 46262 335336
rect 45706 334780 45942 335016
rect 46026 334780 46262 335016
rect 45706 299100 45942 299336
rect 46026 299100 46262 299336
rect 45706 298780 45942 299016
rect 46026 298780 46262 299016
rect 45706 263100 45942 263336
rect 46026 263100 46262 263336
rect 45706 262780 45942 263016
rect 46026 262780 46262 263016
rect 45706 227100 45942 227336
rect 46026 227100 46262 227336
rect 45706 226780 45942 227016
rect 46026 226780 46262 227016
rect 45706 191100 45942 191336
rect 46026 191100 46262 191336
rect 45706 190780 45942 191016
rect 46026 190780 46262 191016
rect 45706 155100 45942 155336
rect 46026 155100 46262 155336
rect 45706 154780 45942 155016
rect 46026 154780 46262 155016
rect 45706 119100 45942 119336
rect 46026 119100 46262 119336
rect 45706 118780 45942 119016
rect 46026 118780 46262 119016
rect 45706 83100 45942 83336
rect 46026 83100 46262 83336
rect 45706 82780 45942 83016
rect 46026 82780 46262 83016
rect 45706 47100 45942 47336
rect 46026 47100 46262 47336
rect 45706 46780 45942 47016
rect 46026 46780 46262 47016
rect 45706 11100 45942 11336
rect 46026 11100 46262 11336
rect 45706 10780 45942 11016
rect 46026 10780 46262 11016
rect 45706 -7300 45942 -7064
rect 46026 -7300 46262 -7064
rect 45706 -7620 45942 -7384
rect 46026 -7620 46262 -7384
rect 73026 704604 73262 704840
rect 73346 704604 73582 704840
rect 73026 704284 73262 704520
rect 73346 704284 73582 704520
rect 73026 686420 73262 686656
rect 73346 686420 73582 686656
rect 73026 686100 73262 686336
rect 73346 686100 73582 686336
rect 73026 650420 73262 650656
rect 73346 650420 73582 650656
rect 73026 650100 73262 650336
rect 73346 650100 73582 650336
rect 73026 614420 73262 614656
rect 73346 614420 73582 614656
rect 73026 614100 73262 614336
rect 73346 614100 73582 614336
rect 73026 578420 73262 578656
rect 73346 578420 73582 578656
rect 73026 578100 73262 578336
rect 73346 578100 73582 578336
rect 73026 542420 73262 542656
rect 73346 542420 73582 542656
rect 73026 542100 73262 542336
rect 73346 542100 73582 542336
rect 73026 506420 73262 506656
rect 73346 506420 73582 506656
rect 73026 506100 73262 506336
rect 73346 506100 73582 506336
rect 73026 470420 73262 470656
rect 73346 470420 73582 470656
rect 73026 470100 73262 470336
rect 73346 470100 73582 470336
rect 73026 434420 73262 434656
rect 73346 434420 73582 434656
rect 73026 434100 73262 434336
rect 73346 434100 73582 434336
rect 73026 398420 73262 398656
rect 73346 398420 73582 398656
rect 73026 398100 73262 398336
rect 73346 398100 73582 398336
rect 73026 362420 73262 362656
rect 73346 362420 73582 362656
rect 73026 362100 73262 362336
rect 73346 362100 73582 362336
rect 73026 326420 73262 326656
rect 73346 326420 73582 326656
rect 73026 326100 73262 326336
rect 73346 326100 73582 326336
rect 73026 290420 73262 290656
rect 73346 290420 73582 290656
rect 73026 290100 73262 290336
rect 73346 290100 73582 290336
rect 73026 254420 73262 254656
rect 73346 254420 73582 254656
rect 73026 254100 73262 254336
rect 73346 254100 73582 254336
rect 73026 218420 73262 218656
rect 73346 218420 73582 218656
rect 73026 218100 73262 218336
rect 73346 218100 73582 218336
rect 73026 182420 73262 182656
rect 73346 182420 73582 182656
rect 73026 182100 73262 182336
rect 73346 182100 73582 182336
rect 73026 146420 73262 146656
rect 73346 146420 73582 146656
rect 73026 146100 73262 146336
rect 73346 146100 73582 146336
rect 73026 110420 73262 110656
rect 73346 110420 73582 110656
rect 73026 110100 73262 110336
rect 73346 110100 73582 110336
rect 73026 74420 73262 74656
rect 73346 74420 73582 74656
rect 73026 74100 73262 74336
rect 73346 74100 73582 74336
rect 73026 38420 73262 38656
rect 73346 38420 73582 38656
rect 73026 38100 73262 38336
rect 73346 38100 73582 38336
rect 73026 2420 73262 2656
rect 73346 2420 73582 2656
rect 73026 2100 73262 2336
rect 73346 2100 73582 2336
rect 73026 -580 73262 -344
rect 73346 -580 73582 -344
rect 73026 -900 73262 -664
rect 73346 -900 73582 -664
rect 74266 705564 74502 705800
rect 74586 705564 74822 705800
rect 74266 705244 74502 705480
rect 74586 705244 74822 705480
rect 74266 687660 74502 687896
rect 74586 687660 74822 687896
rect 74266 687340 74502 687576
rect 74586 687340 74822 687576
rect 74266 651660 74502 651896
rect 74586 651660 74822 651896
rect 74266 651340 74502 651576
rect 74586 651340 74822 651576
rect 74266 615660 74502 615896
rect 74586 615660 74822 615896
rect 74266 615340 74502 615576
rect 74586 615340 74822 615576
rect 74266 579660 74502 579896
rect 74586 579660 74822 579896
rect 74266 579340 74502 579576
rect 74586 579340 74822 579576
rect 74266 543660 74502 543896
rect 74586 543660 74822 543896
rect 74266 543340 74502 543576
rect 74586 543340 74822 543576
rect 74266 507660 74502 507896
rect 74586 507660 74822 507896
rect 74266 507340 74502 507576
rect 74586 507340 74822 507576
rect 74266 471660 74502 471896
rect 74586 471660 74822 471896
rect 74266 471340 74502 471576
rect 74586 471340 74822 471576
rect 74266 435660 74502 435896
rect 74586 435660 74822 435896
rect 74266 435340 74502 435576
rect 74586 435340 74822 435576
rect 74266 399660 74502 399896
rect 74586 399660 74822 399896
rect 74266 399340 74502 399576
rect 74586 399340 74822 399576
rect 74266 363660 74502 363896
rect 74586 363660 74822 363896
rect 74266 363340 74502 363576
rect 74586 363340 74822 363576
rect 74266 327660 74502 327896
rect 74586 327660 74822 327896
rect 74266 327340 74502 327576
rect 74586 327340 74822 327576
rect 74266 291660 74502 291896
rect 74586 291660 74822 291896
rect 74266 291340 74502 291576
rect 74586 291340 74822 291576
rect 74266 255660 74502 255896
rect 74586 255660 74822 255896
rect 74266 255340 74502 255576
rect 74586 255340 74822 255576
rect 74266 219660 74502 219896
rect 74586 219660 74822 219896
rect 74266 219340 74502 219576
rect 74586 219340 74822 219576
rect 74266 183660 74502 183896
rect 74586 183660 74822 183896
rect 74266 183340 74502 183576
rect 74586 183340 74822 183576
rect 74266 147660 74502 147896
rect 74586 147660 74822 147896
rect 74266 147340 74502 147576
rect 74586 147340 74822 147576
rect 74266 111660 74502 111896
rect 74586 111660 74822 111896
rect 74266 111340 74502 111576
rect 74586 111340 74822 111576
rect 74266 75660 74502 75896
rect 74586 75660 74822 75896
rect 74266 75340 74502 75576
rect 74586 75340 74822 75576
rect 74266 39660 74502 39896
rect 74586 39660 74822 39896
rect 74266 39340 74502 39576
rect 74586 39340 74822 39576
rect 74266 3660 74502 3896
rect 74586 3660 74822 3896
rect 74266 3340 74502 3576
rect 74586 3340 74822 3576
rect 74266 -1540 74502 -1304
rect 74586 -1540 74822 -1304
rect 74266 -1860 74502 -1624
rect 74586 -1860 74822 -1624
rect 75506 706524 75742 706760
rect 75826 706524 76062 706760
rect 75506 706204 75742 706440
rect 75826 706204 76062 706440
rect 75506 688900 75742 689136
rect 75826 688900 76062 689136
rect 75506 688580 75742 688816
rect 75826 688580 76062 688816
rect 75506 652900 75742 653136
rect 75826 652900 76062 653136
rect 75506 652580 75742 652816
rect 75826 652580 76062 652816
rect 75506 616900 75742 617136
rect 75826 616900 76062 617136
rect 75506 616580 75742 616816
rect 75826 616580 76062 616816
rect 75506 580900 75742 581136
rect 75826 580900 76062 581136
rect 75506 580580 75742 580816
rect 75826 580580 76062 580816
rect 75506 544900 75742 545136
rect 75826 544900 76062 545136
rect 75506 544580 75742 544816
rect 75826 544580 76062 544816
rect 75506 508900 75742 509136
rect 75826 508900 76062 509136
rect 75506 508580 75742 508816
rect 75826 508580 76062 508816
rect 75506 472900 75742 473136
rect 75826 472900 76062 473136
rect 75506 472580 75742 472816
rect 75826 472580 76062 472816
rect 75506 436900 75742 437136
rect 75826 436900 76062 437136
rect 75506 436580 75742 436816
rect 75826 436580 76062 436816
rect 75506 400900 75742 401136
rect 75826 400900 76062 401136
rect 75506 400580 75742 400816
rect 75826 400580 76062 400816
rect 75506 364900 75742 365136
rect 75826 364900 76062 365136
rect 75506 364580 75742 364816
rect 75826 364580 76062 364816
rect 75506 328900 75742 329136
rect 75826 328900 76062 329136
rect 75506 328580 75742 328816
rect 75826 328580 76062 328816
rect 75506 292900 75742 293136
rect 75826 292900 76062 293136
rect 75506 292580 75742 292816
rect 75826 292580 76062 292816
rect 75506 256900 75742 257136
rect 75826 256900 76062 257136
rect 75506 256580 75742 256816
rect 75826 256580 76062 256816
rect 75506 220900 75742 221136
rect 75826 220900 76062 221136
rect 75506 220580 75742 220816
rect 75826 220580 76062 220816
rect 75506 184900 75742 185136
rect 75826 184900 76062 185136
rect 75506 184580 75742 184816
rect 75826 184580 76062 184816
rect 75506 148900 75742 149136
rect 75826 148900 76062 149136
rect 75506 148580 75742 148816
rect 75826 148580 76062 148816
rect 75506 112900 75742 113136
rect 75826 112900 76062 113136
rect 75506 112580 75742 112816
rect 75826 112580 76062 112816
rect 75506 76900 75742 77136
rect 75826 76900 76062 77136
rect 75506 76580 75742 76816
rect 75826 76580 76062 76816
rect 75506 40900 75742 41136
rect 75826 40900 76062 41136
rect 75506 40580 75742 40816
rect 75826 40580 76062 40816
rect 75506 4900 75742 5136
rect 75826 4900 76062 5136
rect 75506 4580 75742 4816
rect 75826 4580 76062 4816
rect 75506 -2500 75742 -2264
rect 75826 -2500 76062 -2264
rect 75506 -2820 75742 -2584
rect 75826 -2820 76062 -2584
rect 76746 707484 76982 707720
rect 77066 707484 77302 707720
rect 76746 707164 76982 707400
rect 77066 707164 77302 707400
rect 76746 690140 76982 690376
rect 77066 690140 77302 690376
rect 76746 689820 76982 690056
rect 77066 689820 77302 690056
rect 76746 654140 76982 654376
rect 77066 654140 77302 654376
rect 76746 653820 76982 654056
rect 77066 653820 77302 654056
rect 76746 618140 76982 618376
rect 77066 618140 77302 618376
rect 76746 617820 76982 618056
rect 77066 617820 77302 618056
rect 76746 582140 76982 582376
rect 77066 582140 77302 582376
rect 76746 581820 76982 582056
rect 77066 581820 77302 582056
rect 76746 546140 76982 546376
rect 77066 546140 77302 546376
rect 76746 545820 76982 546056
rect 77066 545820 77302 546056
rect 76746 510140 76982 510376
rect 77066 510140 77302 510376
rect 76746 509820 76982 510056
rect 77066 509820 77302 510056
rect 76746 474140 76982 474376
rect 77066 474140 77302 474376
rect 76746 473820 76982 474056
rect 77066 473820 77302 474056
rect 76746 438140 76982 438376
rect 77066 438140 77302 438376
rect 76746 437820 76982 438056
rect 77066 437820 77302 438056
rect 76746 402140 76982 402376
rect 77066 402140 77302 402376
rect 76746 401820 76982 402056
rect 77066 401820 77302 402056
rect 76746 366140 76982 366376
rect 77066 366140 77302 366376
rect 76746 365820 76982 366056
rect 77066 365820 77302 366056
rect 76746 330140 76982 330376
rect 77066 330140 77302 330376
rect 76746 329820 76982 330056
rect 77066 329820 77302 330056
rect 76746 294140 76982 294376
rect 77066 294140 77302 294376
rect 76746 293820 76982 294056
rect 77066 293820 77302 294056
rect 76746 258140 76982 258376
rect 77066 258140 77302 258376
rect 76746 257820 76982 258056
rect 77066 257820 77302 258056
rect 76746 222140 76982 222376
rect 77066 222140 77302 222376
rect 76746 221820 76982 222056
rect 77066 221820 77302 222056
rect 76746 186140 76982 186376
rect 77066 186140 77302 186376
rect 76746 185820 76982 186056
rect 77066 185820 77302 186056
rect 76746 150140 76982 150376
rect 77066 150140 77302 150376
rect 76746 149820 76982 150056
rect 77066 149820 77302 150056
rect 76746 114140 76982 114376
rect 77066 114140 77302 114376
rect 76746 113820 76982 114056
rect 77066 113820 77302 114056
rect 76746 78140 76982 78376
rect 77066 78140 77302 78376
rect 76746 77820 76982 78056
rect 77066 77820 77302 78056
rect 76746 42140 76982 42376
rect 77066 42140 77302 42376
rect 76746 41820 76982 42056
rect 77066 41820 77302 42056
rect 76746 6140 76982 6376
rect 77066 6140 77302 6376
rect 76746 5820 76982 6056
rect 77066 5820 77302 6056
rect 76746 -3460 76982 -3224
rect 77066 -3460 77302 -3224
rect 76746 -3780 76982 -3544
rect 77066 -3780 77302 -3544
rect 77986 708444 78222 708680
rect 78306 708444 78542 708680
rect 77986 708124 78222 708360
rect 78306 708124 78542 708360
rect 77986 691380 78222 691616
rect 78306 691380 78542 691616
rect 77986 691060 78222 691296
rect 78306 691060 78542 691296
rect 77986 655380 78222 655616
rect 78306 655380 78542 655616
rect 77986 655060 78222 655296
rect 78306 655060 78542 655296
rect 77986 619380 78222 619616
rect 78306 619380 78542 619616
rect 77986 619060 78222 619296
rect 78306 619060 78542 619296
rect 77986 583380 78222 583616
rect 78306 583380 78542 583616
rect 77986 583060 78222 583296
rect 78306 583060 78542 583296
rect 77986 547380 78222 547616
rect 78306 547380 78542 547616
rect 77986 547060 78222 547296
rect 78306 547060 78542 547296
rect 77986 511380 78222 511616
rect 78306 511380 78542 511616
rect 77986 511060 78222 511296
rect 78306 511060 78542 511296
rect 77986 475380 78222 475616
rect 78306 475380 78542 475616
rect 77986 475060 78222 475296
rect 78306 475060 78542 475296
rect 77986 439380 78222 439616
rect 78306 439380 78542 439616
rect 77986 439060 78222 439296
rect 78306 439060 78542 439296
rect 77986 403380 78222 403616
rect 78306 403380 78542 403616
rect 77986 403060 78222 403296
rect 78306 403060 78542 403296
rect 77986 367380 78222 367616
rect 78306 367380 78542 367616
rect 77986 367060 78222 367296
rect 78306 367060 78542 367296
rect 77986 331380 78222 331616
rect 78306 331380 78542 331616
rect 77986 331060 78222 331296
rect 78306 331060 78542 331296
rect 77986 295380 78222 295616
rect 78306 295380 78542 295616
rect 77986 295060 78222 295296
rect 78306 295060 78542 295296
rect 77986 259380 78222 259616
rect 78306 259380 78542 259616
rect 77986 259060 78222 259296
rect 78306 259060 78542 259296
rect 77986 223380 78222 223616
rect 78306 223380 78542 223616
rect 77986 223060 78222 223296
rect 78306 223060 78542 223296
rect 77986 187380 78222 187616
rect 78306 187380 78542 187616
rect 77986 187060 78222 187296
rect 78306 187060 78542 187296
rect 77986 151380 78222 151616
rect 78306 151380 78542 151616
rect 77986 151060 78222 151296
rect 78306 151060 78542 151296
rect 77986 115380 78222 115616
rect 78306 115380 78542 115616
rect 77986 115060 78222 115296
rect 78306 115060 78542 115296
rect 77986 79380 78222 79616
rect 78306 79380 78542 79616
rect 77986 79060 78222 79296
rect 78306 79060 78542 79296
rect 77986 43380 78222 43616
rect 78306 43380 78542 43616
rect 77986 43060 78222 43296
rect 78306 43060 78542 43296
rect 77986 7380 78222 7616
rect 78306 7380 78542 7616
rect 77986 7060 78222 7296
rect 78306 7060 78542 7296
rect 77986 -4420 78222 -4184
rect 78306 -4420 78542 -4184
rect 77986 -4740 78222 -4504
rect 78306 -4740 78542 -4504
rect 79226 709404 79462 709640
rect 79546 709404 79782 709640
rect 79226 709084 79462 709320
rect 79546 709084 79782 709320
rect 79226 692620 79462 692856
rect 79546 692620 79782 692856
rect 79226 692300 79462 692536
rect 79546 692300 79782 692536
rect 79226 656620 79462 656856
rect 79546 656620 79782 656856
rect 79226 656300 79462 656536
rect 79546 656300 79782 656536
rect 79226 620620 79462 620856
rect 79546 620620 79782 620856
rect 79226 620300 79462 620536
rect 79546 620300 79782 620536
rect 79226 584620 79462 584856
rect 79546 584620 79782 584856
rect 79226 584300 79462 584536
rect 79546 584300 79782 584536
rect 79226 548620 79462 548856
rect 79546 548620 79782 548856
rect 79226 548300 79462 548536
rect 79546 548300 79782 548536
rect 79226 512620 79462 512856
rect 79546 512620 79782 512856
rect 79226 512300 79462 512536
rect 79546 512300 79782 512536
rect 79226 476620 79462 476856
rect 79546 476620 79782 476856
rect 79226 476300 79462 476536
rect 79546 476300 79782 476536
rect 79226 440620 79462 440856
rect 79546 440620 79782 440856
rect 79226 440300 79462 440536
rect 79546 440300 79782 440536
rect 79226 404620 79462 404856
rect 79546 404620 79782 404856
rect 79226 404300 79462 404536
rect 79546 404300 79782 404536
rect 79226 368620 79462 368856
rect 79546 368620 79782 368856
rect 79226 368300 79462 368536
rect 79546 368300 79782 368536
rect 79226 332620 79462 332856
rect 79546 332620 79782 332856
rect 79226 332300 79462 332536
rect 79546 332300 79782 332536
rect 79226 296620 79462 296856
rect 79546 296620 79782 296856
rect 79226 296300 79462 296536
rect 79546 296300 79782 296536
rect 79226 260620 79462 260856
rect 79546 260620 79782 260856
rect 79226 260300 79462 260536
rect 79546 260300 79782 260536
rect 79226 224620 79462 224856
rect 79546 224620 79782 224856
rect 79226 224300 79462 224536
rect 79546 224300 79782 224536
rect 79226 188620 79462 188856
rect 79546 188620 79782 188856
rect 79226 188300 79462 188536
rect 79546 188300 79782 188536
rect 79226 152620 79462 152856
rect 79546 152620 79782 152856
rect 79226 152300 79462 152536
rect 79546 152300 79782 152536
rect 79226 116620 79462 116856
rect 79546 116620 79782 116856
rect 79226 116300 79462 116536
rect 79546 116300 79782 116536
rect 79226 80620 79462 80856
rect 79546 80620 79782 80856
rect 79226 80300 79462 80536
rect 79546 80300 79782 80536
rect 79226 44620 79462 44856
rect 79546 44620 79782 44856
rect 79226 44300 79462 44536
rect 79546 44300 79782 44536
rect 79226 8620 79462 8856
rect 79546 8620 79782 8856
rect 79226 8300 79462 8536
rect 79546 8300 79782 8536
rect 79226 -5380 79462 -5144
rect 79546 -5380 79782 -5144
rect 79226 -5700 79462 -5464
rect 79546 -5700 79782 -5464
rect 80466 710364 80702 710600
rect 80786 710364 81022 710600
rect 80466 710044 80702 710280
rect 80786 710044 81022 710280
rect 80466 693860 80702 694096
rect 80786 693860 81022 694096
rect 80466 693540 80702 693776
rect 80786 693540 81022 693776
rect 80466 657860 80702 658096
rect 80786 657860 81022 658096
rect 80466 657540 80702 657776
rect 80786 657540 81022 657776
rect 80466 621860 80702 622096
rect 80786 621860 81022 622096
rect 80466 621540 80702 621776
rect 80786 621540 81022 621776
rect 80466 585860 80702 586096
rect 80786 585860 81022 586096
rect 80466 585540 80702 585776
rect 80786 585540 81022 585776
rect 80466 549860 80702 550096
rect 80786 549860 81022 550096
rect 80466 549540 80702 549776
rect 80786 549540 81022 549776
rect 80466 513860 80702 514096
rect 80786 513860 81022 514096
rect 80466 513540 80702 513776
rect 80786 513540 81022 513776
rect 80466 477860 80702 478096
rect 80786 477860 81022 478096
rect 80466 477540 80702 477776
rect 80786 477540 81022 477776
rect 80466 441860 80702 442096
rect 80786 441860 81022 442096
rect 80466 441540 80702 441776
rect 80786 441540 81022 441776
rect 80466 405860 80702 406096
rect 80786 405860 81022 406096
rect 80466 405540 80702 405776
rect 80786 405540 81022 405776
rect 80466 369860 80702 370096
rect 80786 369860 81022 370096
rect 80466 369540 80702 369776
rect 80786 369540 81022 369776
rect 80466 333860 80702 334096
rect 80786 333860 81022 334096
rect 80466 333540 80702 333776
rect 80786 333540 81022 333776
rect 80466 297860 80702 298096
rect 80786 297860 81022 298096
rect 80466 297540 80702 297776
rect 80786 297540 81022 297776
rect 80466 261860 80702 262096
rect 80786 261860 81022 262096
rect 80466 261540 80702 261776
rect 80786 261540 81022 261776
rect 80466 225860 80702 226096
rect 80786 225860 81022 226096
rect 80466 225540 80702 225776
rect 80786 225540 81022 225776
rect 80466 189860 80702 190096
rect 80786 189860 81022 190096
rect 80466 189540 80702 189776
rect 80786 189540 81022 189776
rect 80466 153860 80702 154096
rect 80786 153860 81022 154096
rect 80466 153540 80702 153776
rect 80786 153540 81022 153776
rect 80466 117860 80702 118096
rect 80786 117860 81022 118096
rect 80466 117540 80702 117776
rect 80786 117540 81022 117776
rect 80466 81860 80702 82096
rect 80786 81860 81022 82096
rect 80466 81540 80702 81776
rect 80786 81540 81022 81776
rect 80466 45860 80702 46096
rect 80786 45860 81022 46096
rect 80466 45540 80702 45776
rect 80786 45540 81022 45776
rect 80466 9860 80702 10096
rect 80786 9860 81022 10096
rect 80466 9540 80702 9776
rect 80786 9540 81022 9776
rect 80466 -6340 80702 -6104
rect 80786 -6340 81022 -6104
rect 80466 -6660 80702 -6424
rect 80786 -6660 81022 -6424
rect 81706 711324 81942 711560
rect 82026 711324 82262 711560
rect 81706 711004 81942 711240
rect 82026 711004 82262 711240
rect 81706 695100 81942 695336
rect 82026 695100 82262 695336
rect 81706 694780 81942 695016
rect 82026 694780 82262 695016
rect 81706 659100 81942 659336
rect 82026 659100 82262 659336
rect 81706 658780 81942 659016
rect 82026 658780 82262 659016
rect 81706 623100 81942 623336
rect 82026 623100 82262 623336
rect 81706 622780 81942 623016
rect 82026 622780 82262 623016
rect 81706 587100 81942 587336
rect 82026 587100 82262 587336
rect 81706 586780 81942 587016
rect 82026 586780 82262 587016
rect 81706 551100 81942 551336
rect 82026 551100 82262 551336
rect 81706 550780 81942 551016
rect 82026 550780 82262 551016
rect 81706 515100 81942 515336
rect 82026 515100 82262 515336
rect 81706 514780 81942 515016
rect 82026 514780 82262 515016
rect 81706 479100 81942 479336
rect 82026 479100 82262 479336
rect 81706 478780 81942 479016
rect 82026 478780 82262 479016
rect 81706 443100 81942 443336
rect 82026 443100 82262 443336
rect 81706 442780 81942 443016
rect 82026 442780 82262 443016
rect 81706 407100 81942 407336
rect 82026 407100 82262 407336
rect 81706 406780 81942 407016
rect 82026 406780 82262 407016
rect 81706 371100 81942 371336
rect 82026 371100 82262 371336
rect 81706 370780 81942 371016
rect 82026 370780 82262 371016
rect 81706 335100 81942 335336
rect 82026 335100 82262 335336
rect 81706 334780 81942 335016
rect 82026 334780 82262 335016
rect 81706 299100 81942 299336
rect 82026 299100 82262 299336
rect 81706 298780 81942 299016
rect 82026 298780 82262 299016
rect 81706 263100 81942 263336
rect 82026 263100 82262 263336
rect 81706 262780 81942 263016
rect 82026 262780 82262 263016
rect 81706 227100 81942 227336
rect 82026 227100 82262 227336
rect 81706 226780 81942 227016
rect 82026 226780 82262 227016
rect 81706 191100 81942 191336
rect 82026 191100 82262 191336
rect 81706 190780 81942 191016
rect 82026 190780 82262 191016
rect 81706 155100 81942 155336
rect 82026 155100 82262 155336
rect 81706 154780 81942 155016
rect 82026 154780 82262 155016
rect 81706 119100 81942 119336
rect 82026 119100 82262 119336
rect 81706 118780 81942 119016
rect 82026 118780 82262 119016
rect 81706 83100 81942 83336
rect 82026 83100 82262 83336
rect 81706 82780 81942 83016
rect 82026 82780 82262 83016
rect 81706 47100 81942 47336
rect 82026 47100 82262 47336
rect 81706 46780 81942 47016
rect 82026 46780 82262 47016
rect 81706 11100 81942 11336
rect 82026 11100 82262 11336
rect 81706 10780 81942 11016
rect 82026 10780 82262 11016
rect 81706 -7300 81942 -7064
rect 82026 -7300 82262 -7064
rect 81706 -7620 81942 -7384
rect 82026 -7620 82262 -7384
rect 109026 704604 109262 704840
rect 109346 704604 109582 704840
rect 109026 704284 109262 704520
rect 109346 704284 109582 704520
rect 109026 686420 109262 686656
rect 109346 686420 109582 686656
rect 109026 686100 109262 686336
rect 109346 686100 109582 686336
rect 109026 650420 109262 650656
rect 109346 650420 109582 650656
rect 109026 650100 109262 650336
rect 109346 650100 109582 650336
rect 109026 614420 109262 614656
rect 109346 614420 109582 614656
rect 109026 614100 109262 614336
rect 109346 614100 109582 614336
rect 109026 578420 109262 578656
rect 109346 578420 109582 578656
rect 109026 578100 109262 578336
rect 109346 578100 109582 578336
rect 109026 542420 109262 542656
rect 109346 542420 109582 542656
rect 109026 542100 109262 542336
rect 109346 542100 109582 542336
rect 109026 506420 109262 506656
rect 109346 506420 109582 506656
rect 109026 506100 109262 506336
rect 109346 506100 109582 506336
rect 109026 470420 109262 470656
rect 109346 470420 109582 470656
rect 109026 470100 109262 470336
rect 109346 470100 109582 470336
rect 109026 434420 109262 434656
rect 109346 434420 109582 434656
rect 109026 434100 109262 434336
rect 109346 434100 109582 434336
rect 109026 398420 109262 398656
rect 109346 398420 109582 398656
rect 109026 398100 109262 398336
rect 109346 398100 109582 398336
rect 109026 362420 109262 362656
rect 109346 362420 109582 362656
rect 109026 362100 109262 362336
rect 109346 362100 109582 362336
rect 109026 326420 109262 326656
rect 109346 326420 109582 326656
rect 109026 326100 109262 326336
rect 109346 326100 109582 326336
rect 109026 290420 109262 290656
rect 109346 290420 109582 290656
rect 109026 290100 109262 290336
rect 109346 290100 109582 290336
rect 109026 254420 109262 254656
rect 109346 254420 109582 254656
rect 109026 254100 109262 254336
rect 109346 254100 109582 254336
rect 109026 218420 109262 218656
rect 109346 218420 109582 218656
rect 109026 218100 109262 218336
rect 109346 218100 109582 218336
rect 109026 182420 109262 182656
rect 109346 182420 109582 182656
rect 109026 182100 109262 182336
rect 109346 182100 109582 182336
rect 109026 146420 109262 146656
rect 109346 146420 109582 146656
rect 109026 146100 109262 146336
rect 109346 146100 109582 146336
rect 109026 110420 109262 110656
rect 109346 110420 109582 110656
rect 109026 110100 109262 110336
rect 109346 110100 109582 110336
rect 109026 74420 109262 74656
rect 109346 74420 109582 74656
rect 109026 74100 109262 74336
rect 109346 74100 109582 74336
rect 109026 38420 109262 38656
rect 109346 38420 109582 38656
rect 109026 38100 109262 38336
rect 109346 38100 109582 38336
rect 109026 2420 109262 2656
rect 109346 2420 109582 2656
rect 109026 2100 109262 2336
rect 109346 2100 109582 2336
rect 109026 -580 109262 -344
rect 109346 -580 109582 -344
rect 109026 -900 109262 -664
rect 109346 -900 109582 -664
rect 110266 705564 110502 705800
rect 110586 705564 110822 705800
rect 110266 705244 110502 705480
rect 110586 705244 110822 705480
rect 110266 687660 110502 687896
rect 110586 687660 110822 687896
rect 110266 687340 110502 687576
rect 110586 687340 110822 687576
rect 110266 651660 110502 651896
rect 110586 651660 110822 651896
rect 110266 651340 110502 651576
rect 110586 651340 110822 651576
rect 110266 615660 110502 615896
rect 110586 615660 110822 615896
rect 110266 615340 110502 615576
rect 110586 615340 110822 615576
rect 110266 579660 110502 579896
rect 110586 579660 110822 579896
rect 110266 579340 110502 579576
rect 110586 579340 110822 579576
rect 110266 543660 110502 543896
rect 110586 543660 110822 543896
rect 110266 543340 110502 543576
rect 110586 543340 110822 543576
rect 110266 507660 110502 507896
rect 110586 507660 110822 507896
rect 110266 507340 110502 507576
rect 110586 507340 110822 507576
rect 110266 471660 110502 471896
rect 110586 471660 110822 471896
rect 110266 471340 110502 471576
rect 110586 471340 110822 471576
rect 110266 435660 110502 435896
rect 110586 435660 110822 435896
rect 110266 435340 110502 435576
rect 110586 435340 110822 435576
rect 110266 399660 110502 399896
rect 110586 399660 110822 399896
rect 110266 399340 110502 399576
rect 110586 399340 110822 399576
rect 110266 363660 110502 363896
rect 110586 363660 110822 363896
rect 110266 363340 110502 363576
rect 110586 363340 110822 363576
rect 110266 327660 110502 327896
rect 110586 327660 110822 327896
rect 110266 327340 110502 327576
rect 110586 327340 110822 327576
rect 110266 291660 110502 291896
rect 110586 291660 110822 291896
rect 110266 291340 110502 291576
rect 110586 291340 110822 291576
rect 110266 255660 110502 255896
rect 110586 255660 110822 255896
rect 110266 255340 110502 255576
rect 110586 255340 110822 255576
rect 110266 219660 110502 219896
rect 110586 219660 110822 219896
rect 110266 219340 110502 219576
rect 110586 219340 110822 219576
rect 110266 183660 110502 183896
rect 110586 183660 110822 183896
rect 110266 183340 110502 183576
rect 110586 183340 110822 183576
rect 110266 147660 110502 147896
rect 110586 147660 110822 147896
rect 110266 147340 110502 147576
rect 110586 147340 110822 147576
rect 110266 111660 110502 111896
rect 110586 111660 110822 111896
rect 110266 111340 110502 111576
rect 110586 111340 110822 111576
rect 110266 75660 110502 75896
rect 110586 75660 110822 75896
rect 110266 75340 110502 75576
rect 110586 75340 110822 75576
rect 110266 39660 110502 39896
rect 110586 39660 110822 39896
rect 110266 39340 110502 39576
rect 110586 39340 110822 39576
rect 110266 3660 110502 3896
rect 110586 3660 110822 3896
rect 110266 3340 110502 3576
rect 110586 3340 110822 3576
rect 110266 -1540 110502 -1304
rect 110586 -1540 110822 -1304
rect 110266 -1860 110502 -1624
rect 110586 -1860 110822 -1624
rect 111506 706524 111742 706760
rect 111826 706524 112062 706760
rect 111506 706204 111742 706440
rect 111826 706204 112062 706440
rect 111506 688900 111742 689136
rect 111826 688900 112062 689136
rect 111506 688580 111742 688816
rect 111826 688580 112062 688816
rect 111506 652900 111742 653136
rect 111826 652900 112062 653136
rect 111506 652580 111742 652816
rect 111826 652580 112062 652816
rect 111506 616900 111742 617136
rect 111826 616900 112062 617136
rect 111506 616580 111742 616816
rect 111826 616580 112062 616816
rect 111506 580900 111742 581136
rect 111826 580900 112062 581136
rect 111506 580580 111742 580816
rect 111826 580580 112062 580816
rect 111506 544900 111742 545136
rect 111826 544900 112062 545136
rect 111506 544580 111742 544816
rect 111826 544580 112062 544816
rect 111506 508900 111742 509136
rect 111826 508900 112062 509136
rect 111506 508580 111742 508816
rect 111826 508580 112062 508816
rect 111506 472900 111742 473136
rect 111826 472900 112062 473136
rect 111506 472580 111742 472816
rect 111826 472580 112062 472816
rect 111506 436900 111742 437136
rect 111826 436900 112062 437136
rect 111506 436580 111742 436816
rect 111826 436580 112062 436816
rect 111506 400900 111742 401136
rect 111826 400900 112062 401136
rect 111506 400580 111742 400816
rect 111826 400580 112062 400816
rect 111506 364900 111742 365136
rect 111826 364900 112062 365136
rect 111506 364580 111742 364816
rect 111826 364580 112062 364816
rect 111506 328900 111742 329136
rect 111826 328900 112062 329136
rect 111506 328580 111742 328816
rect 111826 328580 112062 328816
rect 111506 292900 111742 293136
rect 111826 292900 112062 293136
rect 111506 292580 111742 292816
rect 111826 292580 112062 292816
rect 111506 256900 111742 257136
rect 111826 256900 112062 257136
rect 111506 256580 111742 256816
rect 111826 256580 112062 256816
rect 111506 220900 111742 221136
rect 111826 220900 112062 221136
rect 111506 220580 111742 220816
rect 111826 220580 112062 220816
rect 111506 184900 111742 185136
rect 111826 184900 112062 185136
rect 111506 184580 111742 184816
rect 111826 184580 112062 184816
rect 111506 148900 111742 149136
rect 111826 148900 112062 149136
rect 111506 148580 111742 148816
rect 111826 148580 112062 148816
rect 111506 112900 111742 113136
rect 111826 112900 112062 113136
rect 111506 112580 111742 112816
rect 111826 112580 112062 112816
rect 111506 76900 111742 77136
rect 111826 76900 112062 77136
rect 111506 76580 111742 76816
rect 111826 76580 112062 76816
rect 111506 40900 111742 41136
rect 111826 40900 112062 41136
rect 111506 40580 111742 40816
rect 111826 40580 112062 40816
rect 111506 4900 111742 5136
rect 111826 4900 112062 5136
rect 111506 4580 111742 4816
rect 111826 4580 112062 4816
rect 111506 -2500 111742 -2264
rect 111826 -2500 112062 -2264
rect 111506 -2820 111742 -2584
rect 111826 -2820 112062 -2584
rect 112746 707484 112982 707720
rect 113066 707484 113302 707720
rect 112746 707164 112982 707400
rect 113066 707164 113302 707400
rect 112746 690140 112982 690376
rect 113066 690140 113302 690376
rect 112746 689820 112982 690056
rect 113066 689820 113302 690056
rect 112746 654140 112982 654376
rect 113066 654140 113302 654376
rect 112746 653820 112982 654056
rect 113066 653820 113302 654056
rect 112746 618140 112982 618376
rect 113066 618140 113302 618376
rect 112746 617820 112982 618056
rect 113066 617820 113302 618056
rect 112746 582140 112982 582376
rect 113066 582140 113302 582376
rect 112746 581820 112982 582056
rect 113066 581820 113302 582056
rect 112746 546140 112982 546376
rect 113066 546140 113302 546376
rect 112746 545820 112982 546056
rect 113066 545820 113302 546056
rect 112746 510140 112982 510376
rect 113066 510140 113302 510376
rect 112746 509820 112982 510056
rect 113066 509820 113302 510056
rect 112746 474140 112982 474376
rect 113066 474140 113302 474376
rect 112746 473820 112982 474056
rect 113066 473820 113302 474056
rect 112746 438140 112982 438376
rect 113066 438140 113302 438376
rect 112746 437820 112982 438056
rect 113066 437820 113302 438056
rect 112746 402140 112982 402376
rect 113066 402140 113302 402376
rect 112746 401820 112982 402056
rect 113066 401820 113302 402056
rect 112746 366140 112982 366376
rect 113066 366140 113302 366376
rect 112746 365820 112982 366056
rect 113066 365820 113302 366056
rect 112746 330140 112982 330376
rect 113066 330140 113302 330376
rect 112746 329820 112982 330056
rect 113066 329820 113302 330056
rect 112746 294140 112982 294376
rect 113066 294140 113302 294376
rect 112746 293820 112982 294056
rect 113066 293820 113302 294056
rect 112746 258140 112982 258376
rect 113066 258140 113302 258376
rect 112746 257820 112982 258056
rect 113066 257820 113302 258056
rect 112746 222140 112982 222376
rect 113066 222140 113302 222376
rect 112746 221820 112982 222056
rect 113066 221820 113302 222056
rect 112746 186140 112982 186376
rect 113066 186140 113302 186376
rect 112746 185820 112982 186056
rect 113066 185820 113302 186056
rect 112746 150140 112982 150376
rect 113066 150140 113302 150376
rect 112746 149820 112982 150056
rect 113066 149820 113302 150056
rect 112746 114140 112982 114376
rect 113066 114140 113302 114376
rect 112746 113820 112982 114056
rect 113066 113820 113302 114056
rect 112746 78140 112982 78376
rect 113066 78140 113302 78376
rect 112746 77820 112982 78056
rect 113066 77820 113302 78056
rect 112746 42140 112982 42376
rect 113066 42140 113302 42376
rect 112746 41820 112982 42056
rect 113066 41820 113302 42056
rect 112746 6140 112982 6376
rect 113066 6140 113302 6376
rect 112746 5820 112982 6056
rect 113066 5820 113302 6056
rect 112746 -3460 112982 -3224
rect 113066 -3460 113302 -3224
rect 112746 -3780 112982 -3544
rect 113066 -3780 113302 -3544
rect 113986 708444 114222 708680
rect 114306 708444 114542 708680
rect 113986 708124 114222 708360
rect 114306 708124 114542 708360
rect 113986 691380 114222 691616
rect 114306 691380 114542 691616
rect 113986 691060 114222 691296
rect 114306 691060 114542 691296
rect 113986 655380 114222 655616
rect 114306 655380 114542 655616
rect 113986 655060 114222 655296
rect 114306 655060 114542 655296
rect 113986 619380 114222 619616
rect 114306 619380 114542 619616
rect 113986 619060 114222 619296
rect 114306 619060 114542 619296
rect 113986 583380 114222 583616
rect 114306 583380 114542 583616
rect 113986 583060 114222 583296
rect 114306 583060 114542 583296
rect 113986 547380 114222 547616
rect 114306 547380 114542 547616
rect 113986 547060 114222 547296
rect 114306 547060 114542 547296
rect 113986 511380 114222 511616
rect 114306 511380 114542 511616
rect 113986 511060 114222 511296
rect 114306 511060 114542 511296
rect 113986 475380 114222 475616
rect 114306 475380 114542 475616
rect 113986 475060 114222 475296
rect 114306 475060 114542 475296
rect 113986 439380 114222 439616
rect 114306 439380 114542 439616
rect 113986 439060 114222 439296
rect 114306 439060 114542 439296
rect 113986 403380 114222 403616
rect 114306 403380 114542 403616
rect 113986 403060 114222 403296
rect 114306 403060 114542 403296
rect 113986 367380 114222 367616
rect 114306 367380 114542 367616
rect 113986 367060 114222 367296
rect 114306 367060 114542 367296
rect 113986 331380 114222 331616
rect 114306 331380 114542 331616
rect 113986 331060 114222 331296
rect 114306 331060 114542 331296
rect 113986 295380 114222 295616
rect 114306 295380 114542 295616
rect 113986 295060 114222 295296
rect 114306 295060 114542 295296
rect 113986 259380 114222 259616
rect 114306 259380 114542 259616
rect 113986 259060 114222 259296
rect 114306 259060 114542 259296
rect 113986 223380 114222 223616
rect 114306 223380 114542 223616
rect 113986 223060 114222 223296
rect 114306 223060 114542 223296
rect 113986 187380 114222 187616
rect 114306 187380 114542 187616
rect 113986 187060 114222 187296
rect 114306 187060 114542 187296
rect 113986 151380 114222 151616
rect 114306 151380 114542 151616
rect 113986 151060 114222 151296
rect 114306 151060 114542 151296
rect 113986 115380 114222 115616
rect 114306 115380 114542 115616
rect 113986 115060 114222 115296
rect 114306 115060 114542 115296
rect 113986 79380 114222 79616
rect 114306 79380 114542 79616
rect 113986 79060 114222 79296
rect 114306 79060 114542 79296
rect 113986 43380 114222 43616
rect 114306 43380 114542 43616
rect 113986 43060 114222 43296
rect 114306 43060 114542 43296
rect 113986 7380 114222 7616
rect 114306 7380 114542 7616
rect 113986 7060 114222 7296
rect 114306 7060 114542 7296
rect 113986 -4420 114222 -4184
rect 114306 -4420 114542 -4184
rect 113986 -4740 114222 -4504
rect 114306 -4740 114542 -4504
rect 115226 709404 115462 709640
rect 115546 709404 115782 709640
rect 115226 709084 115462 709320
rect 115546 709084 115782 709320
rect 115226 692620 115462 692856
rect 115546 692620 115782 692856
rect 115226 692300 115462 692536
rect 115546 692300 115782 692536
rect 115226 656620 115462 656856
rect 115546 656620 115782 656856
rect 115226 656300 115462 656536
rect 115546 656300 115782 656536
rect 115226 620620 115462 620856
rect 115546 620620 115782 620856
rect 115226 620300 115462 620536
rect 115546 620300 115782 620536
rect 115226 584620 115462 584856
rect 115546 584620 115782 584856
rect 115226 584300 115462 584536
rect 115546 584300 115782 584536
rect 115226 548620 115462 548856
rect 115546 548620 115782 548856
rect 115226 548300 115462 548536
rect 115546 548300 115782 548536
rect 115226 512620 115462 512856
rect 115546 512620 115782 512856
rect 115226 512300 115462 512536
rect 115546 512300 115782 512536
rect 115226 476620 115462 476856
rect 115546 476620 115782 476856
rect 115226 476300 115462 476536
rect 115546 476300 115782 476536
rect 115226 440620 115462 440856
rect 115546 440620 115782 440856
rect 115226 440300 115462 440536
rect 115546 440300 115782 440536
rect 115226 404620 115462 404856
rect 115546 404620 115782 404856
rect 115226 404300 115462 404536
rect 115546 404300 115782 404536
rect 115226 368620 115462 368856
rect 115546 368620 115782 368856
rect 115226 368300 115462 368536
rect 115546 368300 115782 368536
rect 115226 332620 115462 332856
rect 115546 332620 115782 332856
rect 115226 332300 115462 332536
rect 115546 332300 115782 332536
rect 115226 296620 115462 296856
rect 115546 296620 115782 296856
rect 115226 296300 115462 296536
rect 115546 296300 115782 296536
rect 115226 260620 115462 260856
rect 115546 260620 115782 260856
rect 115226 260300 115462 260536
rect 115546 260300 115782 260536
rect 115226 224620 115462 224856
rect 115546 224620 115782 224856
rect 115226 224300 115462 224536
rect 115546 224300 115782 224536
rect 115226 188620 115462 188856
rect 115546 188620 115782 188856
rect 115226 188300 115462 188536
rect 115546 188300 115782 188536
rect 115226 152620 115462 152856
rect 115546 152620 115782 152856
rect 115226 152300 115462 152536
rect 115546 152300 115782 152536
rect 115226 116620 115462 116856
rect 115546 116620 115782 116856
rect 115226 116300 115462 116536
rect 115546 116300 115782 116536
rect 115226 80620 115462 80856
rect 115546 80620 115782 80856
rect 115226 80300 115462 80536
rect 115546 80300 115782 80536
rect 115226 44620 115462 44856
rect 115546 44620 115782 44856
rect 115226 44300 115462 44536
rect 115546 44300 115782 44536
rect 115226 8620 115462 8856
rect 115546 8620 115782 8856
rect 115226 8300 115462 8536
rect 115546 8300 115782 8536
rect 115226 -5380 115462 -5144
rect 115546 -5380 115782 -5144
rect 115226 -5700 115462 -5464
rect 115546 -5700 115782 -5464
rect 116466 710364 116702 710600
rect 116786 710364 117022 710600
rect 116466 710044 116702 710280
rect 116786 710044 117022 710280
rect 116466 693860 116702 694096
rect 116786 693860 117022 694096
rect 116466 693540 116702 693776
rect 116786 693540 117022 693776
rect 116466 657860 116702 658096
rect 116786 657860 117022 658096
rect 116466 657540 116702 657776
rect 116786 657540 117022 657776
rect 116466 621860 116702 622096
rect 116786 621860 117022 622096
rect 116466 621540 116702 621776
rect 116786 621540 117022 621776
rect 116466 585860 116702 586096
rect 116786 585860 117022 586096
rect 116466 585540 116702 585776
rect 116786 585540 117022 585776
rect 116466 549860 116702 550096
rect 116786 549860 117022 550096
rect 116466 549540 116702 549776
rect 116786 549540 117022 549776
rect 116466 513860 116702 514096
rect 116786 513860 117022 514096
rect 116466 513540 116702 513776
rect 116786 513540 117022 513776
rect 116466 477860 116702 478096
rect 116786 477860 117022 478096
rect 116466 477540 116702 477776
rect 116786 477540 117022 477776
rect 116466 441860 116702 442096
rect 116786 441860 117022 442096
rect 116466 441540 116702 441776
rect 116786 441540 117022 441776
rect 116466 405860 116702 406096
rect 116786 405860 117022 406096
rect 116466 405540 116702 405776
rect 116786 405540 117022 405776
rect 116466 369860 116702 370096
rect 116786 369860 117022 370096
rect 116466 369540 116702 369776
rect 116786 369540 117022 369776
rect 116466 333860 116702 334096
rect 116786 333860 117022 334096
rect 116466 333540 116702 333776
rect 116786 333540 117022 333776
rect 116466 297860 116702 298096
rect 116786 297860 117022 298096
rect 116466 297540 116702 297776
rect 116786 297540 117022 297776
rect 116466 261860 116702 262096
rect 116786 261860 117022 262096
rect 116466 261540 116702 261776
rect 116786 261540 117022 261776
rect 116466 225860 116702 226096
rect 116786 225860 117022 226096
rect 116466 225540 116702 225776
rect 116786 225540 117022 225776
rect 116466 189860 116702 190096
rect 116786 189860 117022 190096
rect 116466 189540 116702 189776
rect 116786 189540 117022 189776
rect 116466 153860 116702 154096
rect 116786 153860 117022 154096
rect 116466 153540 116702 153776
rect 116786 153540 117022 153776
rect 116466 117860 116702 118096
rect 116786 117860 117022 118096
rect 116466 117540 116702 117776
rect 116786 117540 117022 117776
rect 116466 81860 116702 82096
rect 116786 81860 117022 82096
rect 116466 81540 116702 81776
rect 116786 81540 117022 81776
rect 116466 45860 116702 46096
rect 116786 45860 117022 46096
rect 116466 45540 116702 45776
rect 116786 45540 117022 45776
rect 116466 9860 116702 10096
rect 116786 9860 117022 10096
rect 116466 9540 116702 9776
rect 116786 9540 117022 9776
rect 116466 -6340 116702 -6104
rect 116786 -6340 117022 -6104
rect 116466 -6660 116702 -6424
rect 116786 -6660 117022 -6424
rect 117706 711324 117942 711560
rect 118026 711324 118262 711560
rect 117706 711004 117942 711240
rect 118026 711004 118262 711240
rect 117706 695100 117942 695336
rect 118026 695100 118262 695336
rect 117706 694780 117942 695016
rect 118026 694780 118262 695016
rect 117706 659100 117942 659336
rect 118026 659100 118262 659336
rect 117706 658780 117942 659016
rect 118026 658780 118262 659016
rect 117706 623100 117942 623336
rect 118026 623100 118262 623336
rect 117706 622780 117942 623016
rect 118026 622780 118262 623016
rect 117706 587100 117942 587336
rect 118026 587100 118262 587336
rect 117706 586780 117942 587016
rect 118026 586780 118262 587016
rect 117706 551100 117942 551336
rect 118026 551100 118262 551336
rect 117706 550780 117942 551016
rect 118026 550780 118262 551016
rect 117706 515100 117942 515336
rect 118026 515100 118262 515336
rect 117706 514780 117942 515016
rect 118026 514780 118262 515016
rect 117706 479100 117942 479336
rect 118026 479100 118262 479336
rect 117706 478780 117942 479016
rect 118026 478780 118262 479016
rect 117706 443100 117942 443336
rect 118026 443100 118262 443336
rect 117706 442780 117942 443016
rect 118026 442780 118262 443016
rect 117706 407100 117942 407336
rect 118026 407100 118262 407336
rect 117706 406780 117942 407016
rect 118026 406780 118262 407016
rect 117706 371100 117942 371336
rect 118026 371100 118262 371336
rect 117706 370780 117942 371016
rect 118026 370780 118262 371016
rect 117706 335100 117942 335336
rect 118026 335100 118262 335336
rect 117706 334780 117942 335016
rect 118026 334780 118262 335016
rect 117706 299100 117942 299336
rect 118026 299100 118262 299336
rect 117706 298780 117942 299016
rect 118026 298780 118262 299016
rect 117706 263100 117942 263336
rect 118026 263100 118262 263336
rect 117706 262780 117942 263016
rect 118026 262780 118262 263016
rect 117706 227100 117942 227336
rect 118026 227100 118262 227336
rect 117706 226780 117942 227016
rect 118026 226780 118262 227016
rect 117706 191100 117942 191336
rect 118026 191100 118262 191336
rect 117706 190780 117942 191016
rect 118026 190780 118262 191016
rect 117706 155100 117942 155336
rect 118026 155100 118262 155336
rect 117706 154780 117942 155016
rect 118026 154780 118262 155016
rect 117706 119100 117942 119336
rect 118026 119100 118262 119336
rect 117706 118780 117942 119016
rect 118026 118780 118262 119016
rect 117706 83100 117942 83336
rect 118026 83100 118262 83336
rect 117706 82780 117942 83016
rect 118026 82780 118262 83016
rect 117706 47100 117942 47336
rect 118026 47100 118262 47336
rect 117706 46780 117942 47016
rect 118026 46780 118262 47016
rect 117706 11100 117942 11336
rect 118026 11100 118262 11336
rect 117706 10780 117942 11016
rect 118026 10780 118262 11016
rect 117706 -7300 117942 -7064
rect 118026 -7300 118262 -7064
rect 117706 -7620 117942 -7384
rect 118026 -7620 118262 -7384
rect 145026 704604 145262 704840
rect 145346 704604 145582 704840
rect 145026 704284 145262 704520
rect 145346 704284 145582 704520
rect 145026 686420 145262 686656
rect 145346 686420 145582 686656
rect 145026 686100 145262 686336
rect 145346 686100 145582 686336
rect 145026 650420 145262 650656
rect 145346 650420 145582 650656
rect 145026 650100 145262 650336
rect 145346 650100 145582 650336
rect 145026 614420 145262 614656
rect 145346 614420 145582 614656
rect 145026 614100 145262 614336
rect 145346 614100 145582 614336
rect 145026 578420 145262 578656
rect 145346 578420 145582 578656
rect 145026 578100 145262 578336
rect 145346 578100 145582 578336
rect 145026 542420 145262 542656
rect 145346 542420 145582 542656
rect 145026 542100 145262 542336
rect 145346 542100 145582 542336
rect 145026 506420 145262 506656
rect 145346 506420 145582 506656
rect 145026 506100 145262 506336
rect 145346 506100 145582 506336
rect 145026 470420 145262 470656
rect 145346 470420 145582 470656
rect 145026 470100 145262 470336
rect 145346 470100 145582 470336
rect 145026 434420 145262 434656
rect 145346 434420 145582 434656
rect 145026 434100 145262 434336
rect 145346 434100 145582 434336
rect 145026 398420 145262 398656
rect 145346 398420 145582 398656
rect 145026 398100 145262 398336
rect 145346 398100 145582 398336
rect 145026 362420 145262 362656
rect 145346 362420 145582 362656
rect 145026 362100 145262 362336
rect 145346 362100 145582 362336
rect 145026 326420 145262 326656
rect 145346 326420 145582 326656
rect 145026 326100 145262 326336
rect 145346 326100 145582 326336
rect 145026 290420 145262 290656
rect 145346 290420 145582 290656
rect 145026 290100 145262 290336
rect 145346 290100 145582 290336
rect 145026 254420 145262 254656
rect 145346 254420 145582 254656
rect 145026 254100 145262 254336
rect 145346 254100 145582 254336
rect 145026 218420 145262 218656
rect 145346 218420 145582 218656
rect 145026 218100 145262 218336
rect 145346 218100 145582 218336
rect 145026 182420 145262 182656
rect 145346 182420 145582 182656
rect 145026 182100 145262 182336
rect 145346 182100 145582 182336
rect 145026 146420 145262 146656
rect 145346 146420 145582 146656
rect 145026 146100 145262 146336
rect 145346 146100 145582 146336
rect 145026 110420 145262 110656
rect 145346 110420 145582 110656
rect 145026 110100 145262 110336
rect 145346 110100 145582 110336
rect 145026 74420 145262 74656
rect 145346 74420 145582 74656
rect 145026 74100 145262 74336
rect 145346 74100 145582 74336
rect 145026 38420 145262 38656
rect 145346 38420 145582 38656
rect 145026 38100 145262 38336
rect 145346 38100 145582 38336
rect 145026 2420 145262 2656
rect 145346 2420 145582 2656
rect 145026 2100 145262 2336
rect 145346 2100 145582 2336
rect 145026 -580 145262 -344
rect 145346 -580 145582 -344
rect 145026 -900 145262 -664
rect 145346 -900 145582 -664
rect 146266 705564 146502 705800
rect 146586 705564 146822 705800
rect 146266 705244 146502 705480
rect 146586 705244 146822 705480
rect 146266 687660 146502 687896
rect 146586 687660 146822 687896
rect 146266 687340 146502 687576
rect 146586 687340 146822 687576
rect 146266 651660 146502 651896
rect 146586 651660 146822 651896
rect 146266 651340 146502 651576
rect 146586 651340 146822 651576
rect 146266 615660 146502 615896
rect 146586 615660 146822 615896
rect 146266 615340 146502 615576
rect 146586 615340 146822 615576
rect 146266 579660 146502 579896
rect 146586 579660 146822 579896
rect 146266 579340 146502 579576
rect 146586 579340 146822 579576
rect 146266 543660 146502 543896
rect 146586 543660 146822 543896
rect 146266 543340 146502 543576
rect 146586 543340 146822 543576
rect 146266 507660 146502 507896
rect 146586 507660 146822 507896
rect 146266 507340 146502 507576
rect 146586 507340 146822 507576
rect 146266 471660 146502 471896
rect 146586 471660 146822 471896
rect 146266 471340 146502 471576
rect 146586 471340 146822 471576
rect 146266 435660 146502 435896
rect 146586 435660 146822 435896
rect 146266 435340 146502 435576
rect 146586 435340 146822 435576
rect 146266 399660 146502 399896
rect 146586 399660 146822 399896
rect 146266 399340 146502 399576
rect 146586 399340 146822 399576
rect 146266 363660 146502 363896
rect 146586 363660 146822 363896
rect 146266 363340 146502 363576
rect 146586 363340 146822 363576
rect 146266 327660 146502 327896
rect 146586 327660 146822 327896
rect 146266 327340 146502 327576
rect 146586 327340 146822 327576
rect 146266 291660 146502 291896
rect 146586 291660 146822 291896
rect 146266 291340 146502 291576
rect 146586 291340 146822 291576
rect 146266 255660 146502 255896
rect 146586 255660 146822 255896
rect 146266 255340 146502 255576
rect 146586 255340 146822 255576
rect 146266 219660 146502 219896
rect 146586 219660 146822 219896
rect 146266 219340 146502 219576
rect 146586 219340 146822 219576
rect 146266 183660 146502 183896
rect 146586 183660 146822 183896
rect 146266 183340 146502 183576
rect 146586 183340 146822 183576
rect 146266 147660 146502 147896
rect 146586 147660 146822 147896
rect 146266 147340 146502 147576
rect 146586 147340 146822 147576
rect 146266 111660 146502 111896
rect 146586 111660 146822 111896
rect 146266 111340 146502 111576
rect 146586 111340 146822 111576
rect 146266 75660 146502 75896
rect 146586 75660 146822 75896
rect 146266 75340 146502 75576
rect 146586 75340 146822 75576
rect 146266 39660 146502 39896
rect 146586 39660 146822 39896
rect 146266 39340 146502 39576
rect 146586 39340 146822 39576
rect 146266 3660 146502 3896
rect 146586 3660 146822 3896
rect 146266 3340 146502 3576
rect 146586 3340 146822 3576
rect 146266 -1540 146502 -1304
rect 146586 -1540 146822 -1304
rect 146266 -1860 146502 -1624
rect 146586 -1860 146822 -1624
rect 147506 706524 147742 706760
rect 147826 706524 148062 706760
rect 147506 706204 147742 706440
rect 147826 706204 148062 706440
rect 147506 688900 147742 689136
rect 147826 688900 148062 689136
rect 147506 688580 147742 688816
rect 147826 688580 148062 688816
rect 147506 652900 147742 653136
rect 147826 652900 148062 653136
rect 147506 652580 147742 652816
rect 147826 652580 148062 652816
rect 147506 616900 147742 617136
rect 147826 616900 148062 617136
rect 147506 616580 147742 616816
rect 147826 616580 148062 616816
rect 147506 580900 147742 581136
rect 147826 580900 148062 581136
rect 147506 580580 147742 580816
rect 147826 580580 148062 580816
rect 147506 544900 147742 545136
rect 147826 544900 148062 545136
rect 147506 544580 147742 544816
rect 147826 544580 148062 544816
rect 147506 508900 147742 509136
rect 147826 508900 148062 509136
rect 147506 508580 147742 508816
rect 147826 508580 148062 508816
rect 147506 472900 147742 473136
rect 147826 472900 148062 473136
rect 147506 472580 147742 472816
rect 147826 472580 148062 472816
rect 147506 436900 147742 437136
rect 147826 436900 148062 437136
rect 147506 436580 147742 436816
rect 147826 436580 148062 436816
rect 147506 400900 147742 401136
rect 147826 400900 148062 401136
rect 147506 400580 147742 400816
rect 147826 400580 148062 400816
rect 147506 364900 147742 365136
rect 147826 364900 148062 365136
rect 147506 364580 147742 364816
rect 147826 364580 148062 364816
rect 147506 328900 147742 329136
rect 147826 328900 148062 329136
rect 147506 328580 147742 328816
rect 147826 328580 148062 328816
rect 147506 292900 147742 293136
rect 147826 292900 148062 293136
rect 147506 292580 147742 292816
rect 147826 292580 148062 292816
rect 147506 256900 147742 257136
rect 147826 256900 148062 257136
rect 147506 256580 147742 256816
rect 147826 256580 148062 256816
rect 147506 220900 147742 221136
rect 147826 220900 148062 221136
rect 147506 220580 147742 220816
rect 147826 220580 148062 220816
rect 147506 184900 147742 185136
rect 147826 184900 148062 185136
rect 147506 184580 147742 184816
rect 147826 184580 148062 184816
rect 147506 148900 147742 149136
rect 147826 148900 148062 149136
rect 147506 148580 147742 148816
rect 147826 148580 148062 148816
rect 147506 112900 147742 113136
rect 147826 112900 148062 113136
rect 147506 112580 147742 112816
rect 147826 112580 148062 112816
rect 147506 76900 147742 77136
rect 147826 76900 148062 77136
rect 147506 76580 147742 76816
rect 147826 76580 148062 76816
rect 147506 40900 147742 41136
rect 147826 40900 148062 41136
rect 147506 40580 147742 40816
rect 147826 40580 148062 40816
rect 147506 4900 147742 5136
rect 147826 4900 148062 5136
rect 147506 4580 147742 4816
rect 147826 4580 148062 4816
rect 147506 -2500 147742 -2264
rect 147826 -2500 148062 -2264
rect 147506 -2820 147742 -2584
rect 147826 -2820 148062 -2584
rect 148746 707484 148982 707720
rect 149066 707484 149302 707720
rect 148746 707164 148982 707400
rect 149066 707164 149302 707400
rect 148746 690140 148982 690376
rect 149066 690140 149302 690376
rect 148746 689820 148982 690056
rect 149066 689820 149302 690056
rect 148746 654140 148982 654376
rect 149066 654140 149302 654376
rect 148746 653820 148982 654056
rect 149066 653820 149302 654056
rect 148746 618140 148982 618376
rect 149066 618140 149302 618376
rect 148746 617820 148982 618056
rect 149066 617820 149302 618056
rect 148746 582140 148982 582376
rect 149066 582140 149302 582376
rect 148746 581820 148982 582056
rect 149066 581820 149302 582056
rect 148746 546140 148982 546376
rect 149066 546140 149302 546376
rect 148746 545820 148982 546056
rect 149066 545820 149302 546056
rect 148746 510140 148982 510376
rect 149066 510140 149302 510376
rect 148746 509820 148982 510056
rect 149066 509820 149302 510056
rect 148746 474140 148982 474376
rect 149066 474140 149302 474376
rect 148746 473820 148982 474056
rect 149066 473820 149302 474056
rect 148746 438140 148982 438376
rect 149066 438140 149302 438376
rect 148746 437820 148982 438056
rect 149066 437820 149302 438056
rect 148746 402140 148982 402376
rect 149066 402140 149302 402376
rect 148746 401820 148982 402056
rect 149066 401820 149302 402056
rect 148746 366140 148982 366376
rect 149066 366140 149302 366376
rect 148746 365820 148982 366056
rect 149066 365820 149302 366056
rect 148746 330140 148982 330376
rect 149066 330140 149302 330376
rect 148746 329820 148982 330056
rect 149066 329820 149302 330056
rect 148746 294140 148982 294376
rect 149066 294140 149302 294376
rect 148746 293820 148982 294056
rect 149066 293820 149302 294056
rect 148746 258140 148982 258376
rect 149066 258140 149302 258376
rect 148746 257820 148982 258056
rect 149066 257820 149302 258056
rect 148746 222140 148982 222376
rect 149066 222140 149302 222376
rect 148746 221820 148982 222056
rect 149066 221820 149302 222056
rect 148746 186140 148982 186376
rect 149066 186140 149302 186376
rect 148746 185820 148982 186056
rect 149066 185820 149302 186056
rect 148746 150140 148982 150376
rect 149066 150140 149302 150376
rect 148746 149820 148982 150056
rect 149066 149820 149302 150056
rect 148746 114140 148982 114376
rect 149066 114140 149302 114376
rect 148746 113820 148982 114056
rect 149066 113820 149302 114056
rect 148746 78140 148982 78376
rect 149066 78140 149302 78376
rect 148746 77820 148982 78056
rect 149066 77820 149302 78056
rect 148746 42140 148982 42376
rect 149066 42140 149302 42376
rect 148746 41820 148982 42056
rect 149066 41820 149302 42056
rect 148746 6140 148982 6376
rect 149066 6140 149302 6376
rect 148746 5820 148982 6056
rect 149066 5820 149302 6056
rect 148746 -3460 148982 -3224
rect 149066 -3460 149302 -3224
rect 148746 -3780 148982 -3544
rect 149066 -3780 149302 -3544
rect 149986 708444 150222 708680
rect 150306 708444 150542 708680
rect 149986 708124 150222 708360
rect 150306 708124 150542 708360
rect 149986 691380 150222 691616
rect 150306 691380 150542 691616
rect 149986 691060 150222 691296
rect 150306 691060 150542 691296
rect 149986 655380 150222 655616
rect 150306 655380 150542 655616
rect 149986 655060 150222 655296
rect 150306 655060 150542 655296
rect 149986 619380 150222 619616
rect 150306 619380 150542 619616
rect 149986 619060 150222 619296
rect 150306 619060 150542 619296
rect 149986 583380 150222 583616
rect 150306 583380 150542 583616
rect 149986 583060 150222 583296
rect 150306 583060 150542 583296
rect 149986 547380 150222 547616
rect 150306 547380 150542 547616
rect 149986 547060 150222 547296
rect 150306 547060 150542 547296
rect 149986 511380 150222 511616
rect 150306 511380 150542 511616
rect 149986 511060 150222 511296
rect 150306 511060 150542 511296
rect 149986 475380 150222 475616
rect 150306 475380 150542 475616
rect 149986 475060 150222 475296
rect 150306 475060 150542 475296
rect 149986 439380 150222 439616
rect 150306 439380 150542 439616
rect 149986 439060 150222 439296
rect 150306 439060 150542 439296
rect 149986 403380 150222 403616
rect 150306 403380 150542 403616
rect 149986 403060 150222 403296
rect 150306 403060 150542 403296
rect 149986 367380 150222 367616
rect 150306 367380 150542 367616
rect 149986 367060 150222 367296
rect 150306 367060 150542 367296
rect 149986 331380 150222 331616
rect 150306 331380 150542 331616
rect 149986 331060 150222 331296
rect 150306 331060 150542 331296
rect 149986 295380 150222 295616
rect 150306 295380 150542 295616
rect 149986 295060 150222 295296
rect 150306 295060 150542 295296
rect 149986 259380 150222 259616
rect 150306 259380 150542 259616
rect 149986 259060 150222 259296
rect 150306 259060 150542 259296
rect 149986 223380 150222 223616
rect 150306 223380 150542 223616
rect 149986 223060 150222 223296
rect 150306 223060 150542 223296
rect 149986 187380 150222 187616
rect 150306 187380 150542 187616
rect 149986 187060 150222 187296
rect 150306 187060 150542 187296
rect 149986 151380 150222 151616
rect 150306 151380 150542 151616
rect 149986 151060 150222 151296
rect 150306 151060 150542 151296
rect 149986 115380 150222 115616
rect 150306 115380 150542 115616
rect 149986 115060 150222 115296
rect 150306 115060 150542 115296
rect 149986 79380 150222 79616
rect 150306 79380 150542 79616
rect 149986 79060 150222 79296
rect 150306 79060 150542 79296
rect 149986 43380 150222 43616
rect 150306 43380 150542 43616
rect 149986 43060 150222 43296
rect 150306 43060 150542 43296
rect 149986 7380 150222 7616
rect 150306 7380 150542 7616
rect 149986 7060 150222 7296
rect 150306 7060 150542 7296
rect 149986 -4420 150222 -4184
rect 150306 -4420 150542 -4184
rect 149986 -4740 150222 -4504
rect 150306 -4740 150542 -4504
rect 151226 709404 151462 709640
rect 151546 709404 151782 709640
rect 151226 709084 151462 709320
rect 151546 709084 151782 709320
rect 151226 692620 151462 692856
rect 151546 692620 151782 692856
rect 151226 692300 151462 692536
rect 151546 692300 151782 692536
rect 151226 656620 151462 656856
rect 151546 656620 151782 656856
rect 151226 656300 151462 656536
rect 151546 656300 151782 656536
rect 151226 620620 151462 620856
rect 151546 620620 151782 620856
rect 151226 620300 151462 620536
rect 151546 620300 151782 620536
rect 151226 584620 151462 584856
rect 151546 584620 151782 584856
rect 151226 584300 151462 584536
rect 151546 584300 151782 584536
rect 151226 548620 151462 548856
rect 151546 548620 151782 548856
rect 151226 548300 151462 548536
rect 151546 548300 151782 548536
rect 151226 512620 151462 512856
rect 151546 512620 151782 512856
rect 151226 512300 151462 512536
rect 151546 512300 151782 512536
rect 151226 476620 151462 476856
rect 151546 476620 151782 476856
rect 151226 476300 151462 476536
rect 151546 476300 151782 476536
rect 151226 440620 151462 440856
rect 151546 440620 151782 440856
rect 151226 440300 151462 440536
rect 151546 440300 151782 440536
rect 151226 404620 151462 404856
rect 151546 404620 151782 404856
rect 151226 404300 151462 404536
rect 151546 404300 151782 404536
rect 151226 368620 151462 368856
rect 151546 368620 151782 368856
rect 151226 368300 151462 368536
rect 151546 368300 151782 368536
rect 151226 332620 151462 332856
rect 151546 332620 151782 332856
rect 151226 332300 151462 332536
rect 151546 332300 151782 332536
rect 151226 296620 151462 296856
rect 151546 296620 151782 296856
rect 151226 296300 151462 296536
rect 151546 296300 151782 296536
rect 151226 260620 151462 260856
rect 151546 260620 151782 260856
rect 151226 260300 151462 260536
rect 151546 260300 151782 260536
rect 151226 224620 151462 224856
rect 151546 224620 151782 224856
rect 151226 224300 151462 224536
rect 151546 224300 151782 224536
rect 151226 188620 151462 188856
rect 151546 188620 151782 188856
rect 151226 188300 151462 188536
rect 151546 188300 151782 188536
rect 151226 152620 151462 152856
rect 151546 152620 151782 152856
rect 151226 152300 151462 152536
rect 151546 152300 151782 152536
rect 151226 116620 151462 116856
rect 151546 116620 151782 116856
rect 151226 116300 151462 116536
rect 151546 116300 151782 116536
rect 151226 80620 151462 80856
rect 151546 80620 151782 80856
rect 151226 80300 151462 80536
rect 151546 80300 151782 80536
rect 151226 44620 151462 44856
rect 151546 44620 151782 44856
rect 151226 44300 151462 44536
rect 151546 44300 151782 44536
rect 151226 8620 151462 8856
rect 151546 8620 151782 8856
rect 151226 8300 151462 8536
rect 151546 8300 151782 8536
rect 151226 -5380 151462 -5144
rect 151546 -5380 151782 -5144
rect 151226 -5700 151462 -5464
rect 151546 -5700 151782 -5464
rect 152466 710364 152702 710600
rect 152786 710364 153022 710600
rect 152466 710044 152702 710280
rect 152786 710044 153022 710280
rect 152466 693860 152702 694096
rect 152786 693860 153022 694096
rect 152466 693540 152702 693776
rect 152786 693540 153022 693776
rect 152466 657860 152702 658096
rect 152786 657860 153022 658096
rect 152466 657540 152702 657776
rect 152786 657540 153022 657776
rect 152466 621860 152702 622096
rect 152786 621860 153022 622096
rect 152466 621540 152702 621776
rect 152786 621540 153022 621776
rect 152466 585860 152702 586096
rect 152786 585860 153022 586096
rect 152466 585540 152702 585776
rect 152786 585540 153022 585776
rect 152466 549860 152702 550096
rect 152786 549860 153022 550096
rect 152466 549540 152702 549776
rect 152786 549540 153022 549776
rect 152466 513860 152702 514096
rect 152786 513860 153022 514096
rect 152466 513540 152702 513776
rect 152786 513540 153022 513776
rect 152466 477860 152702 478096
rect 152786 477860 153022 478096
rect 152466 477540 152702 477776
rect 152786 477540 153022 477776
rect 152466 441860 152702 442096
rect 152786 441860 153022 442096
rect 152466 441540 152702 441776
rect 152786 441540 153022 441776
rect 152466 405860 152702 406096
rect 152786 405860 153022 406096
rect 152466 405540 152702 405776
rect 152786 405540 153022 405776
rect 152466 369860 152702 370096
rect 152786 369860 153022 370096
rect 152466 369540 152702 369776
rect 152786 369540 153022 369776
rect 152466 333860 152702 334096
rect 152786 333860 153022 334096
rect 152466 333540 152702 333776
rect 152786 333540 153022 333776
rect 152466 297860 152702 298096
rect 152786 297860 153022 298096
rect 152466 297540 152702 297776
rect 152786 297540 153022 297776
rect 152466 261860 152702 262096
rect 152786 261860 153022 262096
rect 152466 261540 152702 261776
rect 152786 261540 153022 261776
rect 152466 225860 152702 226096
rect 152786 225860 153022 226096
rect 152466 225540 152702 225776
rect 152786 225540 153022 225776
rect 152466 189860 152702 190096
rect 152786 189860 153022 190096
rect 152466 189540 152702 189776
rect 152786 189540 153022 189776
rect 152466 153860 152702 154096
rect 152786 153860 153022 154096
rect 152466 153540 152702 153776
rect 152786 153540 153022 153776
rect 152466 117860 152702 118096
rect 152786 117860 153022 118096
rect 152466 117540 152702 117776
rect 152786 117540 153022 117776
rect 152466 81860 152702 82096
rect 152786 81860 153022 82096
rect 152466 81540 152702 81776
rect 152786 81540 153022 81776
rect 152466 45860 152702 46096
rect 152786 45860 153022 46096
rect 152466 45540 152702 45776
rect 152786 45540 153022 45776
rect 152466 9860 152702 10096
rect 152786 9860 153022 10096
rect 152466 9540 152702 9776
rect 152786 9540 153022 9776
rect 152466 -6340 152702 -6104
rect 152786 -6340 153022 -6104
rect 152466 -6660 152702 -6424
rect 152786 -6660 153022 -6424
rect 153706 711324 153942 711560
rect 154026 711324 154262 711560
rect 153706 711004 153942 711240
rect 154026 711004 154262 711240
rect 153706 695100 153942 695336
rect 154026 695100 154262 695336
rect 153706 694780 153942 695016
rect 154026 694780 154262 695016
rect 153706 659100 153942 659336
rect 154026 659100 154262 659336
rect 153706 658780 153942 659016
rect 154026 658780 154262 659016
rect 153706 623100 153942 623336
rect 154026 623100 154262 623336
rect 153706 622780 153942 623016
rect 154026 622780 154262 623016
rect 153706 587100 153942 587336
rect 154026 587100 154262 587336
rect 153706 586780 153942 587016
rect 154026 586780 154262 587016
rect 153706 551100 153942 551336
rect 154026 551100 154262 551336
rect 153706 550780 153942 551016
rect 154026 550780 154262 551016
rect 153706 515100 153942 515336
rect 154026 515100 154262 515336
rect 153706 514780 153942 515016
rect 154026 514780 154262 515016
rect 153706 479100 153942 479336
rect 154026 479100 154262 479336
rect 153706 478780 153942 479016
rect 154026 478780 154262 479016
rect 153706 443100 153942 443336
rect 154026 443100 154262 443336
rect 153706 442780 153942 443016
rect 154026 442780 154262 443016
rect 153706 407100 153942 407336
rect 154026 407100 154262 407336
rect 153706 406780 153942 407016
rect 154026 406780 154262 407016
rect 153706 371100 153942 371336
rect 154026 371100 154262 371336
rect 153706 370780 153942 371016
rect 154026 370780 154262 371016
rect 153706 335100 153942 335336
rect 154026 335100 154262 335336
rect 153706 334780 153942 335016
rect 154026 334780 154262 335016
rect 153706 299100 153942 299336
rect 154026 299100 154262 299336
rect 153706 298780 153942 299016
rect 154026 298780 154262 299016
rect 153706 263100 153942 263336
rect 154026 263100 154262 263336
rect 153706 262780 153942 263016
rect 154026 262780 154262 263016
rect 153706 227100 153942 227336
rect 154026 227100 154262 227336
rect 153706 226780 153942 227016
rect 154026 226780 154262 227016
rect 153706 191100 153942 191336
rect 154026 191100 154262 191336
rect 153706 190780 153942 191016
rect 154026 190780 154262 191016
rect 153706 155100 153942 155336
rect 154026 155100 154262 155336
rect 153706 154780 153942 155016
rect 154026 154780 154262 155016
rect 153706 119100 153942 119336
rect 154026 119100 154262 119336
rect 153706 118780 153942 119016
rect 154026 118780 154262 119016
rect 153706 83100 153942 83336
rect 154026 83100 154262 83336
rect 153706 82780 153942 83016
rect 154026 82780 154262 83016
rect 153706 47100 153942 47336
rect 154026 47100 154262 47336
rect 153706 46780 153942 47016
rect 154026 46780 154262 47016
rect 153706 11100 153942 11336
rect 154026 11100 154262 11336
rect 153706 10780 153942 11016
rect 154026 10780 154262 11016
rect 153706 -7300 153942 -7064
rect 154026 -7300 154262 -7064
rect 153706 -7620 153942 -7384
rect 154026 -7620 154262 -7384
rect 181026 704604 181262 704840
rect 181346 704604 181582 704840
rect 181026 704284 181262 704520
rect 181346 704284 181582 704520
rect 181026 686420 181262 686656
rect 181346 686420 181582 686656
rect 181026 686100 181262 686336
rect 181346 686100 181582 686336
rect 181026 650420 181262 650656
rect 181346 650420 181582 650656
rect 181026 650100 181262 650336
rect 181346 650100 181582 650336
rect 181026 614420 181262 614656
rect 181346 614420 181582 614656
rect 181026 614100 181262 614336
rect 181346 614100 181582 614336
rect 181026 578420 181262 578656
rect 181346 578420 181582 578656
rect 181026 578100 181262 578336
rect 181346 578100 181582 578336
rect 181026 542420 181262 542656
rect 181346 542420 181582 542656
rect 181026 542100 181262 542336
rect 181346 542100 181582 542336
rect 181026 506420 181262 506656
rect 181346 506420 181582 506656
rect 181026 506100 181262 506336
rect 181346 506100 181582 506336
rect 181026 470420 181262 470656
rect 181346 470420 181582 470656
rect 181026 470100 181262 470336
rect 181346 470100 181582 470336
rect 181026 434420 181262 434656
rect 181346 434420 181582 434656
rect 181026 434100 181262 434336
rect 181346 434100 181582 434336
rect 181026 398420 181262 398656
rect 181346 398420 181582 398656
rect 181026 398100 181262 398336
rect 181346 398100 181582 398336
rect 181026 362420 181262 362656
rect 181346 362420 181582 362656
rect 181026 362100 181262 362336
rect 181346 362100 181582 362336
rect 181026 326420 181262 326656
rect 181346 326420 181582 326656
rect 181026 326100 181262 326336
rect 181346 326100 181582 326336
rect 181026 290420 181262 290656
rect 181346 290420 181582 290656
rect 181026 290100 181262 290336
rect 181346 290100 181582 290336
rect 181026 254420 181262 254656
rect 181346 254420 181582 254656
rect 181026 254100 181262 254336
rect 181346 254100 181582 254336
rect 181026 218420 181262 218656
rect 181346 218420 181582 218656
rect 181026 218100 181262 218336
rect 181346 218100 181582 218336
rect 181026 182420 181262 182656
rect 181346 182420 181582 182656
rect 181026 182100 181262 182336
rect 181346 182100 181582 182336
rect 181026 146420 181262 146656
rect 181346 146420 181582 146656
rect 181026 146100 181262 146336
rect 181346 146100 181582 146336
rect 181026 110420 181262 110656
rect 181346 110420 181582 110656
rect 181026 110100 181262 110336
rect 181346 110100 181582 110336
rect 181026 74420 181262 74656
rect 181346 74420 181582 74656
rect 181026 74100 181262 74336
rect 181346 74100 181582 74336
rect 181026 38420 181262 38656
rect 181346 38420 181582 38656
rect 181026 38100 181262 38336
rect 181346 38100 181582 38336
rect 181026 2420 181262 2656
rect 181346 2420 181582 2656
rect 181026 2100 181262 2336
rect 181346 2100 181582 2336
rect 181026 -580 181262 -344
rect 181346 -580 181582 -344
rect 181026 -900 181262 -664
rect 181346 -900 181582 -664
rect 182266 705564 182502 705800
rect 182586 705564 182822 705800
rect 182266 705244 182502 705480
rect 182586 705244 182822 705480
rect 182266 687660 182502 687896
rect 182586 687660 182822 687896
rect 182266 687340 182502 687576
rect 182586 687340 182822 687576
rect 182266 651660 182502 651896
rect 182586 651660 182822 651896
rect 182266 651340 182502 651576
rect 182586 651340 182822 651576
rect 182266 615660 182502 615896
rect 182586 615660 182822 615896
rect 182266 615340 182502 615576
rect 182586 615340 182822 615576
rect 182266 579660 182502 579896
rect 182586 579660 182822 579896
rect 182266 579340 182502 579576
rect 182586 579340 182822 579576
rect 182266 543660 182502 543896
rect 182586 543660 182822 543896
rect 182266 543340 182502 543576
rect 182586 543340 182822 543576
rect 182266 507660 182502 507896
rect 182586 507660 182822 507896
rect 182266 507340 182502 507576
rect 182586 507340 182822 507576
rect 182266 471660 182502 471896
rect 182586 471660 182822 471896
rect 182266 471340 182502 471576
rect 182586 471340 182822 471576
rect 182266 435660 182502 435896
rect 182586 435660 182822 435896
rect 182266 435340 182502 435576
rect 182586 435340 182822 435576
rect 182266 399660 182502 399896
rect 182586 399660 182822 399896
rect 182266 399340 182502 399576
rect 182586 399340 182822 399576
rect 182266 363660 182502 363896
rect 182586 363660 182822 363896
rect 182266 363340 182502 363576
rect 182586 363340 182822 363576
rect 182266 327660 182502 327896
rect 182586 327660 182822 327896
rect 182266 327340 182502 327576
rect 182586 327340 182822 327576
rect 182266 291660 182502 291896
rect 182586 291660 182822 291896
rect 182266 291340 182502 291576
rect 182586 291340 182822 291576
rect 182266 255660 182502 255896
rect 182586 255660 182822 255896
rect 182266 255340 182502 255576
rect 182586 255340 182822 255576
rect 182266 219660 182502 219896
rect 182586 219660 182822 219896
rect 182266 219340 182502 219576
rect 182586 219340 182822 219576
rect 182266 183660 182502 183896
rect 182586 183660 182822 183896
rect 182266 183340 182502 183576
rect 182586 183340 182822 183576
rect 182266 147660 182502 147896
rect 182586 147660 182822 147896
rect 182266 147340 182502 147576
rect 182586 147340 182822 147576
rect 182266 111660 182502 111896
rect 182586 111660 182822 111896
rect 182266 111340 182502 111576
rect 182586 111340 182822 111576
rect 182266 75660 182502 75896
rect 182586 75660 182822 75896
rect 182266 75340 182502 75576
rect 182586 75340 182822 75576
rect 182266 39660 182502 39896
rect 182586 39660 182822 39896
rect 182266 39340 182502 39576
rect 182586 39340 182822 39576
rect 182266 3660 182502 3896
rect 182586 3660 182822 3896
rect 182266 3340 182502 3576
rect 182586 3340 182822 3576
rect 182266 -1540 182502 -1304
rect 182586 -1540 182822 -1304
rect 182266 -1860 182502 -1624
rect 182586 -1860 182822 -1624
rect 183506 706524 183742 706760
rect 183826 706524 184062 706760
rect 183506 706204 183742 706440
rect 183826 706204 184062 706440
rect 183506 688900 183742 689136
rect 183826 688900 184062 689136
rect 183506 688580 183742 688816
rect 183826 688580 184062 688816
rect 183506 652900 183742 653136
rect 183826 652900 184062 653136
rect 183506 652580 183742 652816
rect 183826 652580 184062 652816
rect 183506 616900 183742 617136
rect 183826 616900 184062 617136
rect 183506 616580 183742 616816
rect 183826 616580 184062 616816
rect 183506 580900 183742 581136
rect 183826 580900 184062 581136
rect 183506 580580 183742 580816
rect 183826 580580 184062 580816
rect 183506 544900 183742 545136
rect 183826 544900 184062 545136
rect 183506 544580 183742 544816
rect 183826 544580 184062 544816
rect 183506 508900 183742 509136
rect 183826 508900 184062 509136
rect 183506 508580 183742 508816
rect 183826 508580 184062 508816
rect 183506 472900 183742 473136
rect 183826 472900 184062 473136
rect 183506 472580 183742 472816
rect 183826 472580 184062 472816
rect 183506 436900 183742 437136
rect 183826 436900 184062 437136
rect 183506 436580 183742 436816
rect 183826 436580 184062 436816
rect 183506 400900 183742 401136
rect 183826 400900 184062 401136
rect 183506 400580 183742 400816
rect 183826 400580 184062 400816
rect 183506 364900 183742 365136
rect 183826 364900 184062 365136
rect 183506 364580 183742 364816
rect 183826 364580 184062 364816
rect 183506 328900 183742 329136
rect 183826 328900 184062 329136
rect 183506 328580 183742 328816
rect 183826 328580 184062 328816
rect 183506 292900 183742 293136
rect 183826 292900 184062 293136
rect 183506 292580 183742 292816
rect 183826 292580 184062 292816
rect 183506 256900 183742 257136
rect 183826 256900 184062 257136
rect 183506 256580 183742 256816
rect 183826 256580 184062 256816
rect 183506 220900 183742 221136
rect 183826 220900 184062 221136
rect 183506 220580 183742 220816
rect 183826 220580 184062 220816
rect 183506 184900 183742 185136
rect 183826 184900 184062 185136
rect 183506 184580 183742 184816
rect 183826 184580 184062 184816
rect 183506 148900 183742 149136
rect 183826 148900 184062 149136
rect 183506 148580 183742 148816
rect 183826 148580 184062 148816
rect 183506 112900 183742 113136
rect 183826 112900 184062 113136
rect 183506 112580 183742 112816
rect 183826 112580 184062 112816
rect 183506 76900 183742 77136
rect 183826 76900 184062 77136
rect 183506 76580 183742 76816
rect 183826 76580 184062 76816
rect 183506 40900 183742 41136
rect 183826 40900 184062 41136
rect 183506 40580 183742 40816
rect 183826 40580 184062 40816
rect 183506 4900 183742 5136
rect 183826 4900 184062 5136
rect 183506 4580 183742 4816
rect 183826 4580 184062 4816
rect 183506 -2500 183742 -2264
rect 183826 -2500 184062 -2264
rect 183506 -2820 183742 -2584
rect 183826 -2820 184062 -2584
rect 184746 707484 184982 707720
rect 185066 707484 185302 707720
rect 184746 707164 184982 707400
rect 185066 707164 185302 707400
rect 184746 690140 184982 690376
rect 185066 690140 185302 690376
rect 184746 689820 184982 690056
rect 185066 689820 185302 690056
rect 184746 654140 184982 654376
rect 185066 654140 185302 654376
rect 184746 653820 184982 654056
rect 185066 653820 185302 654056
rect 184746 618140 184982 618376
rect 185066 618140 185302 618376
rect 184746 617820 184982 618056
rect 185066 617820 185302 618056
rect 184746 582140 184982 582376
rect 185066 582140 185302 582376
rect 184746 581820 184982 582056
rect 185066 581820 185302 582056
rect 184746 546140 184982 546376
rect 185066 546140 185302 546376
rect 184746 545820 184982 546056
rect 185066 545820 185302 546056
rect 184746 510140 184982 510376
rect 185066 510140 185302 510376
rect 184746 509820 184982 510056
rect 185066 509820 185302 510056
rect 184746 474140 184982 474376
rect 185066 474140 185302 474376
rect 184746 473820 184982 474056
rect 185066 473820 185302 474056
rect 184746 438140 184982 438376
rect 185066 438140 185302 438376
rect 184746 437820 184982 438056
rect 185066 437820 185302 438056
rect 184746 402140 184982 402376
rect 185066 402140 185302 402376
rect 184746 401820 184982 402056
rect 185066 401820 185302 402056
rect 184746 366140 184982 366376
rect 185066 366140 185302 366376
rect 184746 365820 184982 366056
rect 185066 365820 185302 366056
rect 184746 330140 184982 330376
rect 185066 330140 185302 330376
rect 184746 329820 184982 330056
rect 185066 329820 185302 330056
rect 184746 294140 184982 294376
rect 185066 294140 185302 294376
rect 184746 293820 184982 294056
rect 185066 293820 185302 294056
rect 184746 258140 184982 258376
rect 185066 258140 185302 258376
rect 184746 257820 184982 258056
rect 185066 257820 185302 258056
rect 184746 222140 184982 222376
rect 185066 222140 185302 222376
rect 184746 221820 184982 222056
rect 185066 221820 185302 222056
rect 184746 186140 184982 186376
rect 185066 186140 185302 186376
rect 184746 185820 184982 186056
rect 185066 185820 185302 186056
rect 184746 150140 184982 150376
rect 185066 150140 185302 150376
rect 184746 149820 184982 150056
rect 185066 149820 185302 150056
rect 184746 114140 184982 114376
rect 185066 114140 185302 114376
rect 184746 113820 184982 114056
rect 185066 113820 185302 114056
rect 184746 78140 184982 78376
rect 185066 78140 185302 78376
rect 184746 77820 184982 78056
rect 185066 77820 185302 78056
rect 184746 42140 184982 42376
rect 185066 42140 185302 42376
rect 184746 41820 184982 42056
rect 185066 41820 185302 42056
rect 184746 6140 184982 6376
rect 185066 6140 185302 6376
rect 184746 5820 184982 6056
rect 185066 5820 185302 6056
rect 184746 -3460 184982 -3224
rect 185066 -3460 185302 -3224
rect 184746 -3780 184982 -3544
rect 185066 -3780 185302 -3544
rect 185986 708444 186222 708680
rect 186306 708444 186542 708680
rect 185986 708124 186222 708360
rect 186306 708124 186542 708360
rect 185986 691380 186222 691616
rect 186306 691380 186542 691616
rect 185986 691060 186222 691296
rect 186306 691060 186542 691296
rect 185986 655380 186222 655616
rect 186306 655380 186542 655616
rect 185986 655060 186222 655296
rect 186306 655060 186542 655296
rect 185986 619380 186222 619616
rect 186306 619380 186542 619616
rect 185986 619060 186222 619296
rect 186306 619060 186542 619296
rect 185986 583380 186222 583616
rect 186306 583380 186542 583616
rect 185986 583060 186222 583296
rect 186306 583060 186542 583296
rect 185986 547380 186222 547616
rect 186306 547380 186542 547616
rect 185986 547060 186222 547296
rect 186306 547060 186542 547296
rect 185986 511380 186222 511616
rect 186306 511380 186542 511616
rect 185986 511060 186222 511296
rect 186306 511060 186542 511296
rect 185986 475380 186222 475616
rect 186306 475380 186542 475616
rect 185986 475060 186222 475296
rect 186306 475060 186542 475296
rect 185986 439380 186222 439616
rect 186306 439380 186542 439616
rect 185986 439060 186222 439296
rect 186306 439060 186542 439296
rect 185986 403380 186222 403616
rect 186306 403380 186542 403616
rect 185986 403060 186222 403296
rect 186306 403060 186542 403296
rect 185986 367380 186222 367616
rect 186306 367380 186542 367616
rect 185986 367060 186222 367296
rect 186306 367060 186542 367296
rect 185986 331380 186222 331616
rect 186306 331380 186542 331616
rect 185986 331060 186222 331296
rect 186306 331060 186542 331296
rect 185986 295380 186222 295616
rect 186306 295380 186542 295616
rect 185986 295060 186222 295296
rect 186306 295060 186542 295296
rect 185986 259380 186222 259616
rect 186306 259380 186542 259616
rect 185986 259060 186222 259296
rect 186306 259060 186542 259296
rect 185986 223380 186222 223616
rect 186306 223380 186542 223616
rect 185986 223060 186222 223296
rect 186306 223060 186542 223296
rect 185986 187380 186222 187616
rect 186306 187380 186542 187616
rect 185986 187060 186222 187296
rect 186306 187060 186542 187296
rect 185986 151380 186222 151616
rect 186306 151380 186542 151616
rect 185986 151060 186222 151296
rect 186306 151060 186542 151296
rect 185986 115380 186222 115616
rect 186306 115380 186542 115616
rect 185986 115060 186222 115296
rect 186306 115060 186542 115296
rect 185986 79380 186222 79616
rect 186306 79380 186542 79616
rect 185986 79060 186222 79296
rect 186306 79060 186542 79296
rect 185986 43380 186222 43616
rect 186306 43380 186542 43616
rect 185986 43060 186222 43296
rect 186306 43060 186542 43296
rect 185986 7380 186222 7616
rect 186306 7380 186542 7616
rect 185986 7060 186222 7296
rect 186306 7060 186542 7296
rect 185986 -4420 186222 -4184
rect 186306 -4420 186542 -4184
rect 185986 -4740 186222 -4504
rect 186306 -4740 186542 -4504
rect 187226 709404 187462 709640
rect 187546 709404 187782 709640
rect 187226 709084 187462 709320
rect 187546 709084 187782 709320
rect 187226 692620 187462 692856
rect 187546 692620 187782 692856
rect 187226 692300 187462 692536
rect 187546 692300 187782 692536
rect 187226 656620 187462 656856
rect 187546 656620 187782 656856
rect 187226 656300 187462 656536
rect 187546 656300 187782 656536
rect 187226 620620 187462 620856
rect 187546 620620 187782 620856
rect 187226 620300 187462 620536
rect 187546 620300 187782 620536
rect 187226 584620 187462 584856
rect 187546 584620 187782 584856
rect 187226 584300 187462 584536
rect 187546 584300 187782 584536
rect 187226 548620 187462 548856
rect 187546 548620 187782 548856
rect 187226 548300 187462 548536
rect 187546 548300 187782 548536
rect 187226 512620 187462 512856
rect 187546 512620 187782 512856
rect 187226 512300 187462 512536
rect 187546 512300 187782 512536
rect 187226 476620 187462 476856
rect 187546 476620 187782 476856
rect 187226 476300 187462 476536
rect 187546 476300 187782 476536
rect 187226 440620 187462 440856
rect 187546 440620 187782 440856
rect 187226 440300 187462 440536
rect 187546 440300 187782 440536
rect 187226 404620 187462 404856
rect 187546 404620 187782 404856
rect 187226 404300 187462 404536
rect 187546 404300 187782 404536
rect 187226 368620 187462 368856
rect 187546 368620 187782 368856
rect 187226 368300 187462 368536
rect 187546 368300 187782 368536
rect 187226 332620 187462 332856
rect 187546 332620 187782 332856
rect 187226 332300 187462 332536
rect 187546 332300 187782 332536
rect 187226 296620 187462 296856
rect 187546 296620 187782 296856
rect 187226 296300 187462 296536
rect 187546 296300 187782 296536
rect 187226 260620 187462 260856
rect 187546 260620 187782 260856
rect 187226 260300 187462 260536
rect 187546 260300 187782 260536
rect 187226 224620 187462 224856
rect 187546 224620 187782 224856
rect 187226 224300 187462 224536
rect 187546 224300 187782 224536
rect 187226 188620 187462 188856
rect 187546 188620 187782 188856
rect 187226 188300 187462 188536
rect 187546 188300 187782 188536
rect 187226 152620 187462 152856
rect 187546 152620 187782 152856
rect 187226 152300 187462 152536
rect 187546 152300 187782 152536
rect 187226 116620 187462 116856
rect 187546 116620 187782 116856
rect 187226 116300 187462 116536
rect 187546 116300 187782 116536
rect 187226 80620 187462 80856
rect 187546 80620 187782 80856
rect 187226 80300 187462 80536
rect 187546 80300 187782 80536
rect 187226 44620 187462 44856
rect 187546 44620 187782 44856
rect 187226 44300 187462 44536
rect 187546 44300 187782 44536
rect 187226 8620 187462 8856
rect 187546 8620 187782 8856
rect 187226 8300 187462 8536
rect 187546 8300 187782 8536
rect 187226 -5380 187462 -5144
rect 187546 -5380 187782 -5144
rect 187226 -5700 187462 -5464
rect 187546 -5700 187782 -5464
rect 188466 710364 188702 710600
rect 188786 710364 189022 710600
rect 188466 710044 188702 710280
rect 188786 710044 189022 710280
rect 188466 693860 188702 694096
rect 188786 693860 189022 694096
rect 188466 693540 188702 693776
rect 188786 693540 189022 693776
rect 188466 657860 188702 658096
rect 188786 657860 189022 658096
rect 188466 657540 188702 657776
rect 188786 657540 189022 657776
rect 188466 621860 188702 622096
rect 188786 621860 189022 622096
rect 188466 621540 188702 621776
rect 188786 621540 189022 621776
rect 188466 585860 188702 586096
rect 188786 585860 189022 586096
rect 188466 585540 188702 585776
rect 188786 585540 189022 585776
rect 188466 549860 188702 550096
rect 188786 549860 189022 550096
rect 188466 549540 188702 549776
rect 188786 549540 189022 549776
rect 188466 513860 188702 514096
rect 188786 513860 189022 514096
rect 188466 513540 188702 513776
rect 188786 513540 189022 513776
rect 188466 477860 188702 478096
rect 188786 477860 189022 478096
rect 188466 477540 188702 477776
rect 188786 477540 189022 477776
rect 188466 441860 188702 442096
rect 188786 441860 189022 442096
rect 188466 441540 188702 441776
rect 188786 441540 189022 441776
rect 188466 405860 188702 406096
rect 188786 405860 189022 406096
rect 188466 405540 188702 405776
rect 188786 405540 189022 405776
rect 188466 369860 188702 370096
rect 188786 369860 189022 370096
rect 188466 369540 188702 369776
rect 188786 369540 189022 369776
rect 188466 333860 188702 334096
rect 188786 333860 189022 334096
rect 188466 333540 188702 333776
rect 188786 333540 189022 333776
rect 188466 297860 188702 298096
rect 188786 297860 189022 298096
rect 188466 297540 188702 297776
rect 188786 297540 189022 297776
rect 188466 261860 188702 262096
rect 188786 261860 189022 262096
rect 188466 261540 188702 261776
rect 188786 261540 189022 261776
rect 188466 225860 188702 226096
rect 188786 225860 189022 226096
rect 188466 225540 188702 225776
rect 188786 225540 189022 225776
rect 188466 189860 188702 190096
rect 188786 189860 189022 190096
rect 188466 189540 188702 189776
rect 188786 189540 189022 189776
rect 188466 153860 188702 154096
rect 188786 153860 189022 154096
rect 188466 153540 188702 153776
rect 188786 153540 189022 153776
rect 188466 117860 188702 118096
rect 188786 117860 189022 118096
rect 188466 117540 188702 117776
rect 188786 117540 189022 117776
rect 188466 81860 188702 82096
rect 188786 81860 189022 82096
rect 188466 81540 188702 81776
rect 188786 81540 189022 81776
rect 188466 45860 188702 46096
rect 188786 45860 189022 46096
rect 188466 45540 188702 45776
rect 188786 45540 189022 45776
rect 188466 9860 188702 10096
rect 188786 9860 189022 10096
rect 188466 9540 188702 9776
rect 188786 9540 189022 9776
rect 188466 -6340 188702 -6104
rect 188786 -6340 189022 -6104
rect 188466 -6660 188702 -6424
rect 188786 -6660 189022 -6424
rect 189706 711324 189942 711560
rect 190026 711324 190262 711560
rect 189706 711004 189942 711240
rect 190026 711004 190262 711240
rect 189706 695100 189942 695336
rect 190026 695100 190262 695336
rect 189706 694780 189942 695016
rect 190026 694780 190262 695016
rect 189706 659100 189942 659336
rect 190026 659100 190262 659336
rect 189706 658780 189942 659016
rect 190026 658780 190262 659016
rect 189706 623100 189942 623336
rect 190026 623100 190262 623336
rect 189706 622780 189942 623016
rect 190026 622780 190262 623016
rect 189706 587100 189942 587336
rect 190026 587100 190262 587336
rect 189706 586780 189942 587016
rect 190026 586780 190262 587016
rect 189706 551100 189942 551336
rect 190026 551100 190262 551336
rect 189706 550780 189942 551016
rect 190026 550780 190262 551016
rect 189706 515100 189942 515336
rect 190026 515100 190262 515336
rect 189706 514780 189942 515016
rect 190026 514780 190262 515016
rect 189706 479100 189942 479336
rect 190026 479100 190262 479336
rect 189706 478780 189942 479016
rect 190026 478780 190262 479016
rect 189706 443100 189942 443336
rect 190026 443100 190262 443336
rect 189706 442780 189942 443016
rect 190026 442780 190262 443016
rect 189706 407100 189942 407336
rect 190026 407100 190262 407336
rect 189706 406780 189942 407016
rect 190026 406780 190262 407016
rect 189706 371100 189942 371336
rect 190026 371100 190262 371336
rect 189706 370780 189942 371016
rect 190026 370780 190262 371016
rect 189706 335100 189942 335336
rect 190026 335100 190262 335336
rect 189706 334780 189942 335016
rect 190026 334780 190262 335016
rect 189706 299100 189942 299336
rect 190026 299100 190262 299336
rect 189706 298780 189942 299016
rect 190026 298780 190262 299016
rect 189706 263100 189942 263336
rect 190026 263100 190262 263336
rect 189706 262780 189942 263016
rect 190026 262780 190262 263016
rect 189706 227100 189942 227336
rect 190026 227100 190262 227336
rect 189706 226780 189942 227016
rect 190026 226780 190262 227016
rect 189706 191100 189942 191336
rect 190026 191100 190262 191336
rect 189706 190780 189942 191016
rect 190026 190780 190262 191016
rect 189706 155100 189942 155336
rect 190026 155100 190262 155336
rect 189706 154780 189942 155016
rect 190026 154780 190262 155016
rect 189706 119100 189942 119336
rect 190026 119100 190262 119336
rect 189706 118780 189942 119016
rect 190026 118780 190262 119016
rect 189706 83100 189942 83336
rect 190026 83100 190262 83336
rect 189706 82780 189942 83016
rect 190026 82780 190262 83016
rect 189706 47100 189942 47336
rect 190026 47100 190262 47336
rect 189706 46780 189942 47016
rect 190026 46780 190262 47016
rect 189706 11100 189942 11336
rect 190026 11100 190262 11336
rect 189706 10780 189942 11016
rect 190026 10780 190262 11016
rect 189706 -7300 189942 -7064
rect 190026 -7300 190262 -7064
rect 189706 -7620 189942 -7384
rect 190026 -7620 190262 -7384
rect 217026 704604 217262 704840
rect 217346 704604 217582 704840
rect 217026 704284 217262 704520
rect 217346 704284 217582 704520
rect 217026 686420 217262 686656
rect 217346 686420 217582 686656
rect 217026 686100 217262 686336
rect 217346 686100 217582 686336
rect 217026 650420 217262 650656
rect 217346 650420 217582 650656
rect 217026 650100 217262 650336
rect 217346 650100 217582 650336
rect 217026 614420 217262 614656
rect 217346 614420 217582 614656
rect 217026 614100 217262 614336
rect 217346 614100 217582 614336
rect 217026 578420 217262 578656
rect 217346 578420 217582 578656
rect 217026 578100 217262 578336
rect 217346 578100 217582 578336
rect 217026 542420 217262 542656
rect 217346 542420 217582 542656
rect 217026 542100 217262 542336
rect 217346 542100 217582 542336
rect 217026 506420 217262 506656
rect 217346 506420 217582 506656
rect 217026 506100 217262 506336
rect 217346 506100 217582 506336
rect 217026 470420 217262 470656
rect 217346 470420 217582 470656
rect 217026 470100 217262 470336
rect 217346 470100 217582 470336
rect 217026 434420 217262 434656
rect 217346 434420 217582 434656
rect 217026 434100 217262 434336
rect 217346 434100 217582 434336
rect 217026 398420 217262 398656
rect 217346 398420 217582 398656
rect 217026 398100 217262 398336
rect 217346 398100 217582 398336
rect 217026 362420 217262 362656
rect 217346 362420 217582 362656
rect 217026 362100 217262 362336
rect 217346 362100 217582 362336
rect 217026 326420 217262 326656
rect 217346 326420 217582 326656
rect 217026 326100 217262 326336
rect 217346 326100 217582 326336
rect 217026 290420 217262 290656
rect 217346 290420 217582 290656
rect 217026 290100 217262 290336
rect 217346 290100 217582 290336
rect 217026 254420 217262 254656
rect 217346 254420 217582 254656
rect 217026 254100 217262 254336
rect 217346 254100 217582 254336
rect 217026 218420 217262 218656
rect 217346 218420 217582 218656
rect 217026 218100 217262 218336
rect 217346 218100 217582 218336
rect 217026 182420 217262 182656
rect 217346 182420 217582 182656
rect 217026 182100 217262 182336
rect 217346 182100 217582 182336
rect 217026 146420 217262 146656
rect 217346 146420 217582 146656
rect 217026 146100 217262 146336
rect 217346 146100 217582 146336
rect 217026 110420 217262 110656
rect 217346 110420 217582 110656
rect 217026 110100 217262 110336
rect 217346 110100 217582 110336
rect 217026 74420 217262 74656
rect 217346 74420 217582 74656
rect 217026 74100 217262 74336
rect 217346 74100 217582 74336
rect 217026 38420 217262 38656
rect 217346 38420 217582 38656
rect 217026 38100 217262 38336
rect 217346 38100 217582 38336
rect 217026 2420 217262 2656
rect 217346 2420 217582 2656
rect 217026 2100 217262 2336
rect 217346 2100 217582 2336
rect 217026 -580 217262 -344
rect 217346 -580 217582 -344
rect 217026 -900 217262 -664
rect 217346 -900 217582 -664
rect 218266 705564 218502 705800
rect 218586 705564 218822 705800
rect 218266 705244 218502 705480
rect 218586 705244 218822 705480
rect 218266 687660 218502 687896
rect 218586 687660 218822 687896
rect 218266 687340 218502 687576
rect 218586 687340 218822 687576
rect 218266 651660 218502 651896
rect 218586 651660 218822 651896
rect 218266 651340 218502 651576
rect 218586 651340 218822 651576
rect 218266 615660 218502 615896
rect 218586 615660 218822 615896
rect 218266 615340 218502 615576
rect 218586 615340 218822 615576
rect 218266 579660 218502 579896
rect 218586 579660 218822 579896
rect 218266 579340 218502 579576
rect 218586 579340 218822 579576
rect 218266 543660 218502 543896
rect 218586 543660 218822 543896
rect 218266 543340 218502 543576
rect 218586 543340 218822 543576
rect 218266 507660 218502 507896
rect 218586 507660 218822 507896
rect 218266 507340 218502 507576
rect 218586 507340 218822 507576
rect 218266 471660 218502 471896
rect 218586 471660 218822 471896
rect 218266 471340 218502 471576
rect 218586 471340 218822 471576
rect 218266 435660 218502 435896
rect 218586 435660 218822 435896
rect 218266 435340 218502 435576
rect 218586 435340 218822 435576
rect 218266 399660 218502 399896
rect 218586 399660 218822 399896
rect 218266 399340 218502 399576
rect 218586 399340 218822 399576
rect 218266 363660 218502 363896
rect 218586 363660 218822 363896
rect 218266 363340 218502 363576
rect 218586 363340 218822 363576
rect 218266 327660 218502 327896
rect 218586 327660 218822 327896
rect 218266 327340 218502 327576
rect 218586 327340 218822 327576
rect 218266 291660 218502 291896
rect 218586 291660 218822 291896
rect 218266 291340 218502 291576
rect 218586 291340 218822 291576
rect 218266 255660 218502 255896
rect 218586 255660 218822 255896
rect 218266 255340 218502 255576
rect 218586 255340 218822 255576
rect 218266 219660 218502 219896
rect 218586 219660 218822 219896
rect 218266 219340 218502 219576
rect 218586 219340 218822 219576
rect 218266 183660 218502 183896
rect 218586 183660 218822 183896
rect 218266 183340 218502 183576
rect 218586 183340 218822 183576
rect 218266 147660 218502 147896
rect 218586 147660 218822 147896
rect 218266 147340 218502 147576
rect 218586 147340 218822 147576
rect 218266 111660 218502 111896
rect 218586 111660 218822 111896
rect 218266 111340 218502 111576
rect 218586 111340 218822 111576
rect 218266 75660 218502 75896
rect 218586 75660 218822 75896
rect 218266 75340 218502 75576
rect 218586 75340 218822 75576
rect 218266 39660 218502 39896
rect 218586 39660 218822 39896
rect 218266 39340 218502 39576
rect 218586 39340 218822 39576
rect 218266 3660 218502 3896
rect 218586 3660 218822 3896
rect 218266 3340 218502 3576
rect 218586 3340 218822 3576
rect 218266 -1540 218502 -1304
rect 218586 -1540 218822 -1304
rect 218266 -1860 218502 -1624
rect 218586 -1860 218822 -1624
rect 219506 706524 219742 706760
rect 219826 706524 220062 706760
rect 219506 706204 219742 706440
rect 219826 706204 220062 706440
rect 219506 688900 219742 689136
rect 219826 688900 220062 689136
rect 219506 688580 219742 688816
rect 219826 688580 220062 688816
rect 219506 652900 219742 653136
rect 219826 652900 220062 653136
rect 219506 652580 219742 652816
rect 219826 652580 220062 652816
rect 219506 616900 219742 617136
rect 219826 616900 220062 617136
rect 219506 616580 219742 616816
rect 219826 616580 220062 616816
rect 219506 580900 219742 581136
rect 219826 580900 220062 581136
rect 219506 580580 219742 580816
rect 219826 580580 220062 580816
rect 219506 544900 219742 545136
rect 219826 544900 220062 545136
rect 219506 544580 219742 544816
rect 219826 544580 220062 544816
rect 219506 508900 219742 509136
rect 219826 508900 220062 509136
rect 219506 508580 219742 508816
rect 219826 508580 220062 508816
rect 219506 472900 219742 473136
rect 219826 472900 220062 473136
rect 219506 472580 219742 472816
rect 219826 472580 220062 472816
rect 219506 436900 219742 437136
rect 219826 436900 220062 437136
rect 219506 436580 219742 436816
rect 219826 436580 220062 436816
rect 219506 400900 219742 401136
rect 219826 400900 220062 401136
rect 219506 400580 219742 400816
rect 219826 400580 220062 400816
rect 219506 364900 219742 365136
rect 219826 364900 220062 365136
rect 219506 364580 219742 364816
rect 219826 364580 220062 364816
rect 219506 328900 219742 329136
rect 219826 328900 220062 329136
rect 219506 328580 219742 328816
rect 219826 328580 220062 328816
rect 219506 292900 219742 293136
rect 219826 292900 220062 293136
rect 219506 292580 219742 292816
rect 219826 292580 220062 292816
rect 219506 256900 219742 257136
rect 219826 256900 220062 257136
rect 219506 256580 219742 256816
rect 219826 256580 220062 256816
rect 219506 220900 219742 221136
rect 219826 220900 220062 221136
rect 219506 220580 219742 220816
rect 219826 220580 220062 220816
rect 219506 184900 219742 185136
rect 219826 184900 220062 185136
rect 219506 184580 219742 184816
rect 219826 184580 220062 184816
rect 219506 148900 219742 149136
rect 219826 148900 220062 149136
rect 219506 148580 219742 148816
rect 219826 148580 220062 148816
rect 219506 112900 219742 113136
rect 219826 112900 220062 113136
rect 219506 112580 219742 112816
rect 219826 112580 220062 112816
rect 219506 76900 219742 77136
rect 219826 76900 220062 77136
rect 219506 76580 219742 76816
rect 219826 76580 220062 76816
rect 219506 40900 219742 41136
rect 219826 40900 220062 41136
rect 219506 40580 219742 40816
rect 219826 40580 220062 40816
rect 219506 4900 219742 5136
rect 219826 4900 220062 5136
rect 219506 4580 219742 4816
rect 219826 4580 220062 4816
rect 219506 -2500 219742 -2264
rect 219826 -2500 220062 -2264
rect 219506 -2820 219742 -2584
rect 219826 -2820 220062 -2584
rect 220746 707484 220982 707720
rect 221066 707484 221302 707720
rect 220746 707164 220982 707400
rect 221066 707164 221302 707400
rect 220746 690140 220982 690376
rect 221066 690140 221302 690376
rect 220746 689820 220982 690056
rect 221066 689820 221302 690056
rect 220746 654140 220982 654376
rect 221066 654140 221302 654376
rect 220746 653820 220982 654056
rect 221066 653820 221302 654056
rect 220746 618140 220982 618376
rect 221066 618140 221302 618376
rect 220746 617820 220982 618056
rect 221066 617820 221302 618056
rect 220746 582140 220982 582376
rect 221066 582140 221302 582376
rect 220746 581820 220982 582056
rect 221066 581820 221302 582056
rect 220746 546140 220982 546376
rect 221066 546140 221302 546376
rect 220746 545820 220982 546056
rect 221066 545820 221302 546056
rect 220746 510140 220982 510376
rect 221066 510140 221302 510376
rect 220746 509820 220982 510056
rect 221066 509820 221302 510056
rect 220746 474140 220982 474376
rect 221066 474140 221302 474376
rect 220746 473820 220982 474056
rect 221066 473820 221302 474056
rect 220746 438140 220982 438376
rect 221066 438140 221302 438376
rect 220746 437820 220982 438056
rect 221066 437820 221302 438056
rect 220746 402140 220982 402376
rect 221066 402140 221302 402376
rect 220746 401820 220982 402056
rect 221066 401820 221302 402056
rect 220746 366140 220982 366376
rect 221066 366140 221302 366376
rect 220746 365820 220982 366056
rect 221066 365820 221302 366056
rect 220746 330140 220982 330376
rect 221066 330140 221302 330376
rect 220746 329820 220982 330056
rect 221066 329820 221302 330056
rect 220746 294140 220982 294376
rect 221066 294140 221302 294376
rect 220746 293820 220982 294056
rect 221066 293820 221302 294056
rect 220746 258140 220982 258376
rect 221066 258140 221302 258376
rect 220746 257820 220982 258056
rect 221066 257820 221302 258056
rect 220746 222140 220982 222376
rect 221066 222140 221302 222376
rect 220746 221820 220982 222056
rect 221066 221820 221302 222056
rect 220746 186140 220982 186376
rect 221066 186140 221302 186376
rect 220746 185820 220982 186056
rect 221066 185820 221302 186056
rect 220746 150140 220982 150376
rect 221066 150140 221302 150376
rect 220746 149820 220982 150056
rect 221066 149820 221302 150056
rect 220746 114140 220982 114376
rect 221066 114140 221302 114376
rect 220746 113820 220982 114056
rect 221066 113820 221302 114056
rect 220746 78140 220982 78376
rect 221066 78140 221302 78376
rect 220746 77820 220982 78056
rect 221066 77820 221302 78056
rect 220746 42140 220982 42376
rect 221066 42140 221302 42376
rect 220746 41820 220982 42056
rect 221066 41820 221302 42056
rect 220746 6140 220982 6376
rect 221066 6140 221302 6376
rect 220746 5820 220982 6056
rect 221066 5820 221302 6056
rect 220746 -3460 220982 -3224
rect 221066 -3460 221302 -3224
rect 220746 -3780 220982 -3544
rect 221066 -3780 221302 -3544
rect 221986 708444 222222 708680
rect 222306 708444 222542 708680
rect 221986 708124 222222 708360
rect 222306 708124 222542 708360
rect 221986 691380 222222 691616
rect 222306 691380 222542 691616
rect 221986 691060 222222 691296
rect 222306 691060 222542 691296
rect 221986 655380 222222 655616
rect 222306 655380 222542 655616
rect 221986 655060 222222 655296
rect 222306 655060 222542 655296
rect 221986 619380 222222 619616
rect 222306 619380 222542 619616
rect 221986 619060 222222 619296
rect 222306 619060 222542 619296
rect 221986 583380 222222 583616
rect 222306 583380 222542 583616
rect 221986 583060 222222 583296
rect 222306 583060 222542 583296
rect 221986 547380 222222 547616
rect 222306 547380 222542 547616
rect 221986 547060 222222 547296
rect 222306 547060 222542 547296
rect 221986 511380 222222 511616
rect 222306 511380 222542 511616
rect 221986 511060 222222 511296
rect 222306 511060 222542 511296
rect 221986 475380 222222 475616
rect 222306 475380 222542 475616
rect 221986 475060 222222 475296
rect 222306 475060 222542 475296
rect 221986 439380 222222 439616
rect 222306 439380 222542 439616
rect 221986 439060 222222 439296
rect 222306 439060 222542 439296
rect 221986 403380 222222 403616
rect 222306 403380 222542 403616
rect 221986 403060 222222 403296
rect 222306 403060 222542 403296
rect 221986 367380 222222 367616
rect 222306 367380 222542 367616
rect 221986 367060 222222 367296
rect 222306 367060 222542 367296
rect 221986 331380 222222 331616
rect 222306 331380 222542 331616
rect 221986 331060 222222 331296
rect 222306 331060 222542 331296
rect 221986 295380 222222 295616
rect 222306 295380 222542 295616
rect 221986 295060 222222 295296
rect 222306 295060 222542 295296
rect 221986 259380 222222 259616
rect 222306 259380 222542 259616
rect 221986 259060 222222 259296
rect 222306 259060 222542 259296
rect 221986 223380 222222 223616
rect 222306 223380 222542 223616
rect 221986 223060 222222 223296
rect 222306 223060 222542 223296
rect 221986 187380 222222 187616
rect 222306 187380 222542 187616
rect 221986 187060 222222 187296
rect 222306 187060 222542 187296
rect 221986 151380 222222 151616
rect 222306 151380 222542 151616
rect 221986 151060 222222 151296
rect 222306 151060 222542 151296
rect 221986 115380 222222 115616
rect 222306 115380 222542 115616
rect 221986 115060 222222 115296
rect 222306 115060 222542 115296
rect 221986 79380 222222 79616
rect 222306 79380 222542 79616
rect 221986 79060 222222 79296
rect 222306 79060 222542 79296
rect 221986 43380 222222 43616
rect 222306 43380 222542 43616
rect 221986 43060 222222 43296
rect 222306 43060 222542 43296
rect 221986 7380 222222 7616
rect 222306 7380 222542 7616
rect 221986 7060 222222 7296
rect 222306 7060 222542 7296
rect 221986 -4420 222222 -4184
rect 222306 -4420 222542 -4184
rect 221986 -4740 222222 -4504
rect 222306 -4740 222542 -4504
rect 223226 709404 223462 709640
rect 223546 709404 223782 709640
rect 223226 709084 223462 709320
rect 223546 709084 223782 709320
rect 223226 692620 223462 692856
rect 223546 692620 223782 692856
rect 223226 692300 223462 692536
rect 223546 692300 223782 692536
rect 223226 656620 223462 656856
rect 223546 656620 223782 656856
rect 223226 656300 223462 656536
rect 223546 656300 223782 656536
rect 223226 620620 223462 620856
rect 223546 620620 223782 620856
rect 223226 620300 223462 620536
rect 223546 620300 223782 620536
rect 223226 584620 223462 584856
rect 223546 584620 223782 584856
rect 223226 584300 223462 584536
rect 223546 584300 223782 584536
rect 223226 548620 223462 548856
rect 223546 548620 223782 548856
rect 223226 548300 223462 548536
rect 223546 548300 223782 548536
rect 223226 512620 223462 512856
rect 223546 512620 223782 512856
rect 223226 512300 223462 512536
rect 223546 512300 223782 512536
rect 223226 476620 223462 476856
rect 223546 476620 223782 476856
rect 223226 476300 223462 476536
rect 223546 476300 223782 476536
rect 223226 440620 223462 440856
rect 223546 440620 223782 440856
rect 223226 440300 223462 440536
rect 223546 440300 223782 440536
rect 223226 404620 223462 404856
rect 223546 404620 223782 404856
rect 223226 404300 223462 404536
rect 223546 404300 223782 404536
rect 223226 368620 223462 368856
rect 223546 368620 223782 368856
rect 223226 368300 223462 368536
rect 223546 368300 223782 368536
rect 223226 332620 223462 332856
rect 223546 332620 223782 332856
rect 223226 332300 223462 332536
rect 223546 332300 223782 332536
rect 223226 296620 223462 296856
rect 223546 296620 223782 296856
rect 223226 296300 223462 296536
rect 223546 296300 223782 296536
rect 223226 260620 223462 260856
rect 223546 260620 223782 260856
rect 223226 260300 223462 260536
rect 223546 260300 223782 260536
rect 223226 224620 223462 224856
rect 223546 224620 223782 224856
rect 223226 224300 223462 224536
rect 223546 224300 223782 224536
rect 223226 188620 223462 188856
rect 223546 188620 223782 188856
rect 223226 188300 223462 188536
rect 223546 188300 223782 188536
rect 223226 152620 223462 152856
rect 223546 152620 223782 152856
rect 223226 152300 223462 152536
rect 223546 152300 223782 152536
rect 223226 116620 223462 116856
rect 223546 116620 223782 116856
rect 223226 116300 223462 116536
rect 223546 116300 223782 116536
rect 223226 80620 223462 80856
rect 223546 80620 223782 80856
rect 223226 80300 223462 80536
rect 223546 80300 223782 80536
rect 223226 44620 223462 44856
rect 223546 44620 223782 44856
rect 223226 44300 223462 44536
rect 223546 44300 223782 44536
rect 223226 8620 223462 8856
rect 223546 8620 223782 8856
rect 223226 8300 223462 8536
rect 223546 8300 223782 8536
rect 223226 -5380 223462 -5144
rect 223546 -5380 223782 -5144
rect 223226 -5700 223462 -5464
rect 223546 -5700 223782 -5464
rect 224466 710364 224702 710600
rect 224786 710364 225022 710600
rect 224466 710044 224702 710280
rect 224786 710044 225022 710280
rect 224466 693860 224702 694096
rect 224786 693860 225022 694096
rect 224466 693540 224702 693776
rect 224786 693540 225022 693776
rect 224466 657860 224702 658096
rect 224786 657860 225022 658096
rect 224466 657540 224702 657776
rect 224786 657540 225022 657776
rect 224466 621860 224702 622096
rect 224786 621860 225022 622096
rect 224466 621540 224702 621776
rect 224786 621540 225022 621776
rect 224466 585860 224702 586096
rect 224786 585860 225022 586096
rect 224466 585540 224702 585776
rect 224786 585540 225022 585776
rect 224466 549860 224702 550096
rect 224786 549860 225022 550096
rect 224466 549540 224702 549776
rect 224786 549540 225022 549776
rect 224466 513860 224702 514096
rect 224786 513860 225022 514096
rect 224466 513540 224702 513776
rect 224786 513540 225022 513776
rect 224466 477860 224702 478096
rect 224786 477860 225022 478096
rect 224466 477540 224702 477776
rect 224786 477540 225022 477776
rect 224466 441860 224702 442096
rect 224786 441860 225022 442096
rect 224466 441540 224702 441776
rect 224786 441540 225022 441776
rect 224466 405860 224702 406096
rect 224786 405860 225022 406096
rect 224466 405540 224702 405776
rect 224786 405540 225022 405776
rect 224466 369860 224702 370096
rect 224786 369860 225022 370096
rect 224466 369540 224702 369776
rect 224786 369540 225022 369776
rect 224466 333860 224702 334096
rect 224786 333860 225022 334096
rect 224466 333540 224702 333776
rect 224786 333540 225022 333776
rect 224466 297860 224702 298096
rect 224786 297860 225022 298096
rect 224466 297540 224702 297776
rect 224786 297540 225022 297776
rect 224466 261860 224702 262096
rect 224786 261860 225022 262096
rect 224466 261540 224702 261776
rect 224786 261540 225022 261776
rect 224466 225860 224702 226096
rect 224786 225860 225022 226096
rect 224466 225540 224702 225776
rect 224786 225540 225022 225776
rect 224466 189860 224702 190096
rect 224786 189860 225022 190096
rect 224466 189540 224702 189776
rect 224786 189540 225022 189776
rect 224466 153860 224702 154096
rect 224786 153860 225022 154096
rect 224466 153540 224702 153776
rect 224786 153540 225022 153776
rect 224466 117860 224702 118096
rect 224786 117860 225022 118096
rect 224466 117540 224702 117776
rect 224786 117540 225022 117776
rect 224466 81860 224702 82096
rect 224786 81860 225022 82096
rect 224466 81540 224702 81776
rect 224786 81540 225022 81776
rect 224466 45860 224702 46096
rect 224786 45860 225022 46096
rect 224466 45540 224702 45776
rect 224786 45540 225022 45776
rect 224466 9860 224702 10096
rect 224786 9860 225022 10096
rect 224466 9540 224702 9776
rect 224786 9540 225022 9776
rect 224466 -6340 224702 -6104
rect 224786 -6340 225022 -6104
rect 224466 -6660 224702 -6424
rect 224786 -6660 225022 -6424
rect 225706 711324 225942 711560
rect 226026 711324 226262 711560
rect 225706 711004 225942 711240
rect 226026 711004 226262 711240
rect 225706 695100 225942 695336
rect 226026 695100 226262 695336
rect 225706 694780 225942 695016
rect 226026 694780 226262 695016
rect 225706 659100 225942 659336
rect 226026 659100 226262 659336
rect 225706 658780 225942 659016
rect 226026 658780 226262 659016
rect 225706 623100 225942 623336
rect 226026 623100 226262 623336
rect 225706 622780 225942 623016
rect 226026 622780 226262 623016
rect 225706 587100 225942 587336
rect 226026 587100 226262 587336
rect 225706 586780 225942 587016
rect 226026 586780 226262 587016
rect 225706 551100 225942 551336
rect 226026 551100 226262 551336
rect 225706 550780 225942 551016
rect 226026 550780 226262 551016
rect 225706 515100 225942 515336
rect 226026 515100 226262 515336
rect 225706 514780 225942 515016
rect 226026 514780 226262 515016
rect 225706 479100 225942 479336
rect 226026 479100 226262 479336
rect 225706 478780 225942 479016
rect 226026 478780 226262 479016
rect 225706 443100 225942 443336
rect 226026 443100 226262 443336
rect 225706 442780 225942 443016
rect 226026 442780 226262 443016
rect 225706 407100 225942 407336
rect 226026 407100 226262 407336
rect 225706 406780 225942 407016
rect 226026 406780 226262 407016
rect 225706 371100 225942 371336
rect 226026 371100 226262 371336
rect 225706 370780 225942 371016
rect 226026 370780 226262 371016
rect 225706 335100 225942 335336
rect 226026 335100 226262 335336
rect 225706 334780 225942 335016
rect 226026 334780 226262 335016
rect 225706 299100 225942 299336
rect 226026 299100 226262 299336
rect 225706 298780 225942 299016
rect 226026 298780 226262 299016
rect 225706 263100 225942 263336
rect 226026 263100 226262 263336
rect 225706 262780 225942 263016
rect 226026 262780 226262 263016
rect 225706 227100 225942 227336
rect 226026 227100 226262 227336
rect 225706 226780 225942 227016
rect 226026 226780 226262 227016
rect 225706 191100 225942 191336
rect 226026 191100 226262 191336
rect 225706 190780 225942 191016
rect 226026 190780 226262 191016
rect 225706 155100 225942 155336
rect 226026 155100 226262 155336
rect 225706 154780 225942 155016
rect 226026 154780 226262 155016
rect 225706 119100 225942 119336
rect 226026 119100 226262 119336
rect 225706 118780 225942 119016
rect 226026 118780 226262 119016
rect 225706 83100 225942 83336
rect 226026 83100 226262 83336
rect 225706 82780 225942 83016
rect 226026 82780 226262 83016
rect 225706 47100 225942 47336
rect 226026 47100 226262 47336
rect 225706 46780 225942 47016
rect 226026 46780 226262 47016
rect 225706 11100 225942 11336
rect 226026 11100 226262 11336
rect 225706 10780 225942 11016
rect 226026 10780 226262 11016
rect 225706 -7300 225942 -7064
rect 226026 -7300 226262 -7064
rect 225706 -7620 225942 -7384
rect 226026 -7620 226262 -7384
rect 253026 704604 253262 704840
rect 253346 704604 253582 704840
rect 253026 704284 253262 704520
rect 253346 704284 253582 704520
rect 253026 686420 253262 686656
rect 253346 686420 253582 686656
rect 253026 686100 253262 686336
rect 253346 686100 253582 686336
rect 253026 650420 253262 650656
rect 253346 650420 253582 650656
rect 253026 650100 253262 650336
rect 253346 650100 253582 650336
rect 253026 614420 253262 614656
rect 253346 614420 253582 614656
rect 253026 614100 253262 614336
rect 253346 614100 253582 614336
rect 253026 578420 253262 578656
rect 253346 578420 253582 578656
rect 253026 578100 253262 578336
rect 253346 578100 253582 578336
rect 253026 542420 253262 542656
rect 253346 542420 253582 542656
rect 253026 542100 253262 542336
rect 253346 542100 253582 542336
rect 253026 506420 253262 506656
rect 253346 506420 253582 506656
rect 253026 506100 253262 506336
rect 253346 506100 253582 506336
rect 253026 470420 253262 470656
rect 253346 470420 253582 470656
rect 253026 470100 253262 470336
rect 253346 470100 253582 470336
rect 253026 434420 253262 434656
rect 253346 434420 253582 434656
rect 253026 434100 253262 434336
rect 253346 434100 253582 434336
rect 253026 398420 253262 398656
rect 253346 398420 253582 398656
rect 253026 398100 253262 398336
rect 253346 398100 253582 398336
rect 253026 362420 253262 362656
rect 253346 362420 253582 362656
rect 253026 362100 253262 362336
rect 253346 362100 253582 362336
rect 253026 326420 253262 326656
rect 253346 326420 253582 326656
rect 253026 326100 253262 326336
rect 253346 326100 253582 326336
rect 253026 290420 253262 290656
rect 253346 290420 253582 290656
rect 253026 290100 253262 290336
rect 253346 290100 253582 290336
rect 253026 254420 253262 254656
rect 253346 254420 253582 254656
rect 253026 254100 253262 254336
rect 253346 254100 253582 254336
rect 253026 218420 253262 218656
rect 253346 218420 253582 218656
rect 253026 218100 253262 218336
rect 253346 218100 253582 218336
rect 253026 182420 253262 182656
rect 253346 182420 253582 182656
rect 253026 182100 253262 182336
rect 253346 182100 253582 182336
rect 253026 146420 253262 146656
rect 253346 146420 253582 146656
rect 253026 146100 253262 146336
rect 253346 146100 253582 146336
rect 253026 110420 253262 110656
rect 253346 110420 253582 110656
rect 253026 110100 253262 110336
rect 253346 110100 253582 110336
rect 253026 74420 253262 74656
rect 253346 74420 253582 74656
rect 253026 74100 253262 74336
rect 253346 74100 253582 74336
rect 253026 38420 253262 38656
rect 253346 38420 253582 38656
rect 253026 38100 253262 38336
rect 253346 38100 253582 38336
rect 253026 2420 253262 2656
rect 253346 2420 253582 2656
rect 253026 2100 253262 2336
rect 253346 2100 253582 2336
rect 253026 -580 253262 -344
rect 253346 -580 253582 -344
rect 253026 -900 253262 -664
rect 253346 -900 253582 -664
rect 254266 705564 254502 705800
rect 254586 705564 254822 705800
rect 254266 705244 254502 705480
rect 254586 705244 254822 705480
rect 254266 687660 254502 687896
rect 254586 687660 254822 687896
rect 254266 687340 254502 687576
rect 254586 687340 254822 687576
rect 254266 651660 254502 651896
rect 254586 651660 254822 651896
rect 254266 651340 254502 651576
rect 254586 651340 254822 651576
rect 254266 615660 254502 615896
rect 254586 615660 254822 615896
rect 254266 615340 254502 615576
rect 254586 615340 254822 615576
rect 254266 579660 254502 579896
rect 254586 579660 254822 579896
rect 254266 579340 254502 579576
rect 254586 579340 254822 579576
rect 254266 543660 254502 543896
rect 254586 543660 254822 543896
rect 254266 543340 254502 543576
rect 254586 543340 254822 543576
rect 254266 507660 254502 507896
rect 254586 507660 254822 507896
rect 254266 507340 254502 507576
rect 254586 507340 254822 507576
rect 254266 471660 254502 471896
rect 254586 471660 254822 471896
rect 254266 471340 254502 471576
rect 254586 471340 254822 471576
rect 254266 435660 254502 435896
rect 254586 435660 254822 435896
rect 254266 435340 254502 435576
rect 254586 435340 254822 435576
rect 254266 399660 254502 399896
rect 254586 399660 254822 399896
rect 254266 399340 254502 399576
rect 254586 399340 254822 399576
rect 254266 363660 254502 363896
rect 254586 363660 254822 363896
rect 254266 363340 254502 363576
rect 254586 363340 254822 363576
rect 254266 327660 254502 327896
rect 254586 327660 254822 327896
rect 254266 327340 254502 327576
rect 254586 327340 254822 327576
rect 254266 291660 254502 291896
rect 254586 291660 254822 291896
rect 254266 291340 254502 291576
rect 254586 291340 254822 291576
rect 254266 255660 254502 255896
rect 254586 255660 254822 255896
rect 254266 255340 254502 255576
rect 254586 255340 254822 255576
rect 254266 219660 254502 219896
rect 254586 219660 254822 219896
rect 254266 219340 254502 219576
rect 254586 219340 254822 219576
rect 254266 183660 254502 183896
rect 254586 183660 254822 183896
rect 254266 183340 254502 183576
rect 254586 183340 254822 183576
rect 254266 147660 254502 147896
rect 254586 147660 254822 147896
rect 254266 147340 254502 147576
rect 254586 147340 254822 147576
rect 254266 111660 254502 111896
rect 254586 111660 254822 111896
rect 254266 111340 254502 111576
rect 254586 111340 254822 111576
rect 254266 75660 254502 75896
rect 254586 75660 254822 75896
rect 254266 75340 254502 75576
rect 254586 75340 254822 75576
rect 254266 39660 254502 39896
rect 254586 39660 254822 39896
rect 254266 39340 254502 39576
rect 254586 39340 254822 39576
rect 254266 3660 254502 3896
rect 254586 3660 254822 3896
rect 254266 3340 254502 3576
rect 254586 3340 254822 3576
rect 254266 -1540 254502 -1304
rect 254586 -1540 254822 -1304
rect 254266 -1860 254502 -1624
rect 254586 -1860 254822 -1624
rect 255506 706524 255742 706760
rect 255826 706524 256062 706760
rect 255506 706204 255742 706440
rect 255826 706204 256062 706440
rect 255506 688900 255742 689136
rect 255826 688900 256062 689136
rect 255506 688580 255742 688816
rect 255826 688580 256062 688816
rect 255506 652900 255742 653136
rect 255826 652900 256062 653136
rect 255506 652580 255742 652816
rect 255826 652580 256062 652816
rect 255506 616900 255742 617136
rect 255826 616900 256062 617136
rect 255506 616580 255742 616816
rect 255826 616580 256062 616816
rect 255506 580900 255742 581136
rect 255826 580900 256062 581136
rect 255506 580580 255742 580816
rect 255826 580580 256062 580816
rect 255506 544900 255742 545136
rect 255826 544900 256062 545136
rect 255506 544580 255742 544816
rect 255826 544580 256062 544816
rect 255506 508900 255742 509136
rect 255826 508900 256062 509136
rect 255506 508580 255742 508816
rect 255826 508580 256062 508816
rect 255506 472900 255742 473136
rect 255826 472900 256062 473136
rect 255506 472580 255742 472816
rect 255826 472580 256062 472816
rect 255506 436900 255742 437136
rect 255826 436900 256062 437136
rect 255506 436580 255742 436816
rect 255826 436580 256062 436816
rect 255506 400900 255742 401136
rect 255826 400900 256062 401136
rect 255506 400580 255742 400816
rect 255826 400580 256062 400816
rect 255506 364900 255742 365136
rect 255826 364900 256062 365136
rect 255506 364580 255742 364816
rect 255826 364580 256062 364816
rect 255506 328900 255742 329136
rect 255826 328900 256062 329136
rect 255506 328580 255742 328816
rect 255826 328580 256062 328816
rect 255506 292900 255742 293136
rect 255826 292900 256062 293136
rect 255506 292580 255742 292816
rect 255826 292580 256062 292816
rect 255506 256900 255742 257136
rect 255826 256900 256062 257136
rect 255506 256580 255742 256816
rect 255826 256580 256062 256816
rect 255506 220900 255742 221136
rect 255826 220900 256062 221136
rect 255506 220580 255742 220816
rect 255826 220580 256062 220816
rect 255506 184900 255742 185136
rect 255826 184900 256062 185136
rect 255506 184580 255742 184816
rect 255826 184580 256062 184816
rect 255506 148900 255742 149136
rect 255826 148900 256062 149136
rect 255506 148580 255742 148816
rect 255826 148580 256062 148816
rect 255506 112900 255742 113136
rect 255826 112900 256062 113136
rect 255506 112580 255742 112816
rect 255826 112580 256062 112816
rect 255506 76900 255742 77136
rect 255826 76900 256062 77136
rect 255506 76580 255742 76816
rect 255826 76580 256062 76816
rect 255506 40900 255742 41136
rect 255826 40900 256062 41136
rect 255506 40580 255742 40816
rect 255826 40580 256062 40816
rect 255506 4900 255742 5136
rect 255826 4900 256062 5136
rect 255506 4580 255742 4816
rect 255826 4580 256062 4816
rect 255506 -2500 255742 -2264
rect 255826 -2500 256062 -2264
rect 255506 -2820 255742 -2584
rect 255826 -2820 256062 -2584
rect 256746 707484 256982 707720
rect 257066 707484 257302 707720
rect 256746 707164 256982 707400
rect 257066 707164 257302 707400
rect 256746 690140 256982 690376
rect 257066 690140 257302 690376
rect 256746 689820 256982 690056
rect 257066 689820 257302 690056
rect 256746 654140 256982 654376
rect 257066 654140 257302 654376
rect 256746 653820 256982 654056
rect 257066 653820 257302 654056
rect 256746 618140 256982 618376
rect 257066 618140 257302 618376
rect 256746 617820 256982 618056
rect 257066 617820 257302 618056
rect 256746 582140 256982 582376
rect 257066 582140 257302 582376
rect 256746 581820 256982 582056
rect 257066 581820 257302 582056
rect 256746 546140 256982 546376
rect 257066 546140 257302 546376
rect 256746 545820 256982 546056
rect 257066 545820 257302 546056
rect 256746 510140 256982 510376
rect 257066 510140 257302 510376
rect 256746 509820 256982 510056
rect 257066 509820 257302 510056
rect 256746 474140 256982 474376
rect 257066 474140 257302 474376
rect 256746 473820 256982 474056
rect 257066 473820 257302 474056
rect 256746 438140 256982 438376
rect 257066 438140 257302 438376
rect 256746 437820 256982 438056
rect 257066 437820 257302 438056
rect 256746 402140 256982 402376
rect 257066 402140 257302 402376
rect 256746 401820 256982 402056
rect 257066 401820 257302 402056
rect 256746 366140 256982 366376
rect 257066 366140 257302 366376
rect 256746 365820 256982 366056
rect 257066 365820 257302 366056
rect 256746 330140 256982 330376
rect 257066 330140 257302 330376
rect 256746 329820 256982 330056
rect 257066 329820 257302 330056
rect 256746 294140 256982 294376
rect 257066 294140 257302 294376
rect 256746 293820 256982 294056
rect 257066 293820 257302 294056
rect 256746 258140 256982 258376
rect 257066 258140 257302 258376
rect 256746 257820 256982 258056
rect 257066 257820 257302 258056
rect 256746 222140 256982 222376
rect 257066 222140 257302 222376
rect 256746 221820 256982 222056
rect 257066 221820 257302 222056
rect 256746 186140 256982 186376
rect 257066 186140 257302 186376
rect 256746 185820 256982 186056
rect 257066 185820 257302 186056
rect 256746 150140 256982 150376
rect 257066 150140 257302 150376
rect 256746 149820 256982 150056
rect 257066 149820 257302 150056
rect 256746 114140 256982 114376
rect 257066 114140 257302 114376
rect 256746 113820 256982 114056
rect 257066 113820 257302 114056
rect 256746 78140 256982 78376
rect 257066 78140 257302 78376
rect 256746 77820 256982 78056
rect 257066 77820 257302 78056
rect 256746 42140 256982 42376
rect 257066 42140 257302 42376
rect 256746 41820 256982 42056
rect 257066 41820 257302 42056
rect 256746 6140 256982 6376
rect 257066 6140 257302 6376
rect 256746 5820 256982 6056
rect 257066 5820 257302 6056
rect 256746 -3460 256982 -3224
rect 257066 -3460 257302 -3224
rect 256746 -3780 256982 -3544
rect 257066 -3780 257302 -3544
rect 257986 708444 258222 708680
rect 258306 708444 258542 708680
rect 257986 708124 258222 708360
rect 258306 708124 258542 708360
rect 257986 691380 258222 691616
rect 258306 691380 258542 691616
rect 257986 691060 258222 691296
rect 258306 691060 258542 691296
rect 257986 655380 258222 655616
rect 258306 655380 258542 655616
rect 257986 655060 258222 655296
rect 258306 655060 258542 655296
rect 257986 619380 258222 619616
rect 258306 619380 258542 619616
rect 257986 619060 258222 619296
rect 258306 619060 258542 619296
rect 257986 583380 258222 583616
rect 258306 583380 258542 583616
rect 257986 583060 258222 583296
rect 258306 583060 258542 583296
rect 257986 547380 258222 547616
rect 258306 547380 258542 547616
rect 257986 547060 258222 547296
rect 258306 547060 258542 547296
rect 257986 511380 258222 511616
rect 258306 511380 258542 511616
rect 257986 511060 258222 511296
rect 258306 511060 258542 511296
rect 257986 475380 258222 475616
rect 258306 475380 258542 475616
rect 257986 475060 258222 475296
rect 258306 475060 258542 475296
rect 257986 439380 258222 439616
rect 258306 439380 258542 439616
rect 257986 439060 258222 439296
rect 258306 439060 258542 439296
rect 257986 403380 258222 403616
rect 258306 403380 258542 403616
rect 257986 403060 258222 403296
rect 258306 403060 258542 403296
rect 257986 367380 258222 367616
rect 258306 367380 258542 367616
rect 257986 367060 258222 367296
rect 258306 367060 258542 367296
rect 257986 331380 258222 331616
rect 258306 331380 258542 331616
rect 257986 331060 258222 331296
rect 258306 331060 258542 331296
rect 257986 295380 258222 295616
rect 258306 295380 258542 295616
rect 257986 295060 258222 295296
rect 258306 295060 258542 295296
rect 257986 259380 258222 259616
rect 258306 259380 258542 259616
rect 257986 259060 258222 259296
rect 258306 259060 258542 259296
rect 257986 223380 258222 223616
rect 258306 223380 258542 223616
rect 257986 223060 258222 223296
rect 258306 223060 258542 223296
rect 257986 187380 258222 187616
rect 258306 187380 258542 187616
rect 257986 187060 258222 187296
rect 258306 187060 258542 187296
rect 257986 151380 258222 151616
rect 258306 151380 258542 151616
rect 257986 151060 258222 151296
rect 258306 151060 258542 151296
rect 257986 115380 258222 115616
rect 258306 115380 258542 115616
rect 257986 115060 258222 115296
rect 258306 115060 258542 115296
rect 257986 79380 258222 79616
rect 258306 79380 258542 79616
rect 257986 79060 258222 79296
rect 258306 79060 258542 79296
rect 257986 43380 258222 43616
rect 258306 43380 258542 43616
rect 257986 43060 258222 43296
rect 258306 43060 258542 43296
rect 257986 7380 258222 7616
rect 258306 7380 258542 7616
rect 257986 7060 258222 7296
rect 258306 7060 258542 7296
rect 257986 -4420 258222 -4184
rect 258306 -4420 258542 -4184
rect 257986 -4740 258222 -4504
rect 258306 -4740 258542 -4504
rect 259226 709404 259462 709640
rect 259546 709404 259782 709640
rect 259226 709084 259462 709320
rect 259546 709084 259782 709320
rect 259226 692620 259462 692856
rect 259546 692620 259782 692856
rect 259226 692300 259462 692536
rect 259546 692300 259782 692536
rect 259226 656620 259462 656856
rect 259546 656620 259782 656856
rect 259226 656300 259462 656536
rect 259546 656300 259782 656536
rect 259226 620620 259462 620856
rect 259546 620620 259782 620856
rect 259226 620300 259462 620536
rect 259546 620300 259782 620536
rect 259226 584620 259462 584856
rect 259546 584620 259782 584856
rect 259226 584300 259462 584536
rect 259546 584300 259782 584536
rect 259226 548620 259462 548856
rect 259546 548620 259782 548856
rect 259226 548300 259462 548536
rect 259546 548300 259782 548536
rect 259226 512620 259462 512856
rect 259546 512620 259782 512856
rect 259226 512300 259462 512536
rect 259546 512300 259782 512536
rect 259226 476620 259462 476856
rect 259546 476620 259782 476856
rect 259226 476300 259462 476536
rect 259546 476300 259782 476536
rect 259226 440620 259462 440856
rect 259546 440620 259782 440856
rect 259226 440300 259462 440536
rect 259546 440300 259782 440536
rect 259226 404620 259462 404856
rect 259546 404620 259782 404856
rect 259226 404300 259462 404536
rect 259546 404300 259782 404536
rect 259226 368620 259462 368856
rect 259546 368620 259782 368856
rect 259226 368300 259462 368536
rect 259546 368300 259782 368536
rect 259226 332620 259462 332856
rect 259546 332620 259782 332856
rect 259226 332300 259462 332536
rect 259546 332300 259782 332536
rect 259226 296620 259462 296856
rect 259546 296620 259782 296856
rect 259226 296300 259462 296536
rect 259546 296300 259782 296536
rect 259226 260620 259462 260856
rect 259546 260620 259782 260856
rect 259226 260300 259462 260536
rect 259546 260300 259782 260536
rect 259226 224620 259462 224856
rect 259546 224620 259782 224856
rect 259226 224300 259462 224536
rect 259546 224300 259782 224536
rect 259226 188620 259462 188856
rect 259546 188620 259782 188856
rect 259226 188300 259462 188536
rect 259546 188300 259782 188536
rect 259226 152620 259462 152856
rect 259546 152620 259782 152856
rect 259226 152300 259462 152536
rect 259546 152300 259782 152536
rect 259226 116620 259462 116856
rect 259546 116620 259782 116856
rect 259226 116300 259462 116536
rect 259546 116300 259782 116536
rect 259226 80620 259462 80856
rect 259546 80620 259782 80856
rect 259226 80300 259462 80536
rect 259546 80300 259782 80536
rect 259226 44620 259462 44856
rect 259546 44620 259782 44856
rect 259226 44300 259462 44536
rect 259546 44300 259782 44536
rect 259226 8620 259462 8856
rect 259546 8620 259782 8856
rect 259226 8300 259462 8536
rect 259546 8300 259782 8536
rect 259226 -5380 259462 -5144
rect 259546 -5380 259782 -5144
rect 259226 -5700 259462 -5464
rect 259546 -5700 259782 -5464
rect 260466 710364 260702 710600
rect 260786 710364 261022 710600
rect 260466 710044 260702 710280
rect 260786 710044 261022 710280
rect 260466 693860 260702 694096
rect 260786 693860 261022 694096
rect 260466 693540 260702 693776
rect 260786 693540 261022 693776
rect 260466 657860 260702 658096
rect 260786 657860 261022 658096
rect 260466 657540 260702 657776
rect 260786 657540 261022 657776
rect 260466 621860 260702 622096
rect 260786 621860 261022 622096
rect 260466 621540 260702 621776
rect 260786 621540 261022 621776
rect 260466 585860 260702 586096
rect 260786 585860 261022 586096
rect 260466 585540 260702 585776
rect 260786 585540 261022 585776
rect 260466 549860 260702 550096
rect 260786 549860 261022 550096
rect 260466 549540 260702 549776
rect 260786 549540 261022 549776
rect 260466 513860 260702 514096
rect 260786 513860 261022 514096
rect 260466 513540 260702 513776
rect 260786 513540 261022 513776
rect 260466 477860 260702 478096
rect 260786 477860 261022 478096
rect 260466 477540 260702 477776
rect 260786 477540 261022 477776
rect 260466 441860 260702 442096
rect 260786 441860 261022 442096
rect 260466 441540 260702 441776
rect 260786 441540 261022 441776
rect 260466 405860 260702 406096
rect 260786 405860 261022 406096
rect 260466 405540 260702 405776
rect 260786 405540 261022 405776
rect 260466 369860 260702 370096
rect 260786 369860 261022 370096
rect 260466 369540 260702 369776
rect 260786 369540 261022 369776
rect 260466 333860 260702 334096
rect 260786 333860 261022 334096
rect 260466 333540 260702 333776
rect 260786 333540 261022 333776
rect 260466 297860 260702 298096
rect 260786 297860 261022 298096
rect 260466 297540 260702 297776
rect 260786 297540 261022 297776
rect 260466 261860 260702 262096
rect 260786 261860 261022 262096
rect 260466 261540 260702 261776
rect 260786 261540 261022 261776
rect 260466 225860 260702 226096
rect 260786 225860 261022 226096
rect 260466 225540 260702 225776
rect 260786 225540 261022 225776
rect 260466 189860 260702 190096
rect 260786 189860 261022 190096
rect 260466 189540 260702 189776
rect 260786 189540 261022 189776
rect 260466 153860 260702 154096
rect 260786 153860 261022 154096
rect 260466 153540 260702 153776
rect 260786 153540 261022 153776
rect 260466 117860 260702 118096
rect 260786 117860 261022 118096
rect 260466 117540 260702 117776
rect 260786 117540 261022 117776
rect 260466 81860 260702 82096
rect 260786 81860 261022 82096
rect 260466 81540 260702 81776
rect 260786 81540 261022 81776
rect 260466 45860 260702 46096
rect 260786 45860 261022 46096
rect 260466 45540 260702 45776
rect 260786 45540 261022 45776
rect 260466 9860 260702 10096
rect 260786 9860 261022 10096
rect 260466 9540 260702 9776
rect 260786 9540 261022 9776
rect 260466 -6340 260702 -6104
rect 260786 -6340 261022 -6104
rect 260466 -6660 260702 -6424
rect 260786 -6660 261022 -6424
rect 261706 711324 261942 711560
rect 262026 711324 262262 711560
rect 261706 711004 261942 711240
rect 262026 711004 262262 711240
rect 261706 695100 261942 695336
rect 262026 695100 262262 695336
rect 261706 694780 261942 695016
rect 262026 694780 262262 695016
rect 261706 659100 261942 659336
rect 262026 659100 262262 659336
rect 261706 658780 261942 659016
rect 262026 658780 262262 659016
rect 261706 623100 261942 623336
rect 262026 623100 262262 623336
rect 261706 622780 261942 623016
rect 262026 622780 262262 623016
rect 261706 587100 261942 587336
rect 262026 587100 262262 587336
rect 261706 586780 261942 587016
rect 262026 586780 262262 587016
rect 261706 551100 261942 551336
rect 262026 551100 262262 551336
rect 261706 550780 261942 551016
rect 262026 550780 262262 551016
rect 261706 515100 261942 515336
rect 262026 515100 262262 515336
rect 261706 514780 261942 515016
rect 262026 514780 262262 515016
rect 261706 479100 261942 479336
rect 262026 479100 262262 479336
rect 261706 478780 261942 479016
rect 262026 478780 262262 479016
rect 261706 443100 261942 443336
rect 262026 443100 262262 443336
rect 261706 442780 261942 443016
rect 262026 442780 262262 443016
rect 261706 407100 261942 407336
rect 262026 407100 262262 407336
rect 261706 406780 261942 407016
rect 262026 406780 262262 407016
rect 261706 371100 261942 371336
rect 262026 371100 262262 371336
rect 261706 370780 261942 371016
rect 262026 370780 262262 371016
rect 261706 335100 261942 335336
rect 262026 335100 262262 335336
rect 261706 334780 261942 335016
rect 262026 334780 262262 335016
rect 261706 299100 261942 299336
rect 262026 299100 262262 299336
rect 261706 298780 261942 299016
rect 262026 298780 262262 299016
rect 261706 263100 261942 263336
rect 262026 263100 262262 263336
rect 261706 262780 261942 263016
rect 262026 262780 262262 263016
rect 261706 227100 261942 227336
rect 262026 227100 262262 227336
rect 261706 226780 261942 227016
rect 262026 226780 262262 227016
rect 261706 191100 261942 191336
rect 262026 191100 262262 191336
rect 261706 190780 261942 191016
rect 262026 190780 262262 191016
rect 261706 155100 261942 155336
rect 262026 155100 262262 155336
rect 261706 154780 261942 155016
rect 262026 154780 262262 155016
rect 261706 119100 261942 119336
rect 262026 119100 262262 119336
rect 261706 118780 261942 119016
rect 262026 118780 262262 119016
rect 261706 83100 261942 83336
rect 262026 83100 262262 83336
rect 261706 82780 261942 83016
rect 262026 82780 262262 83016
rect 261706 47100 261942 47336
rect 262026 47100 262262 47336
rect 261706 46780 261942 47016
rect 262026 46780 262262 47016
rect 261706 11100 261942 11336
rect 262026 11100 262262 11336
rect 261706 10780 261942 11016
rect 262026 10780 262262 11016
rect 261706 -7300 261942 -7064
rect 262026 -7300 262262 -7064
rect 261706 -7620 261942 -7384
rect 262026 -7620 262262 -7384
rect 289026 704604 289262 704840
rect 289346 704604 289582 704840
rect 289026 704284 289262 704520
rect 289346 704284 289582 704520
rect 289026 686420 289262 686656
rect 289346 686420 289582 686656
rect 289026 686100 289262 686336
rect 289346 686100 289582 686336
rect 289026 650420 289262 650656
rect 289346 650420 289582 650656
rect 289026 650100 289262 650336
rect 289346 650100 289582 650336
rect 289026 614420 289262 614656
rect 289346 614420 289582 614656
rect 289026 614100 289262 614336
rect 289346 614100 289582 614336
rect 289026 578420 289262 578656
rect 289346 578420 289582 578656
rect 289026 578100 289262 578336
rect 289346 578100 289582 578336
rect 289026 542420 289262 542656
rect 289346 542420 289582 542656
rect 289026 542100 289262 542336
rect 289346 542100 289582 542336
rect 289026 506420 289262 506656
rect 289346 506420 289582 506656
rect 289026 506100 289262 506336
rect 289346 506100 289582 506336
rect 289026 470420 289262 470656
rect 289346 470420 289582 470656
rect 289026 470100 289262 470336
rect 289346 470100 289582 470336
rect 289026 434420 289262 434656
rect 289346 434420 289582 434656
rect 289026 434100 289262 434336
rect 289346 434100 289582 434336
rect 289026 398420 289262 398656
rect 289346 398420 289582 398656
rect 289026 398100 289262 398336
rect 289346 398100 289582 398336
rect 289026 362420 289262 362656
rect 289346 362420 289582 362656
rect 289026 362100 289262 362336
rect 289346 362100 289582 362336
rect 289026 326420 289262 326656
rect 289346 326420 289582 326656
rect 289026 326100 289262 326336
rect 289346 326100 289582 326336
rect 289026 290420 289262 290656
rect 289346 290420 289582 290656
rect 289026 290100 289262 290336
rect 289346 290100 289582 290336
rect 289026 254420 289262 254656
rect 289346 254420 289582 254656
rect 289026 254100 289262 254336
rect 289346 254100 289582 254336
rect 289026 218420 289262 218656
rect 289346 218420 289582 218656
rect 289026 218100 289262 218336
rect 289346 218100 289582 218336
rect 289026 182420 289262 182656
rect 289346 182420 289582 182656
rect 289026 182100 289262 182336
rect 289346 182100 289582 182336
rect 289026 146420 289262 146656
rect 289346 146420 289582 146656
rect 289026 146100 289262 146336
rect 289346 146100 289582 146336
rect 289026 110420 289262 110656
rect 289346 110420 289582 110656
rect 289026 110100 289262 110336
rect 289346 110100 289582 110336
rect 289026 74420 289262 74656
rect 289346 74420 289582 74656
rect 289026 74100 289262 74336
rect 289346 74100 289582 74336
rect 289026 38420 289262 38656
rect 289346 38420 289582 38656
rect 289026 38100 289262 38336
rect 289346 38100 289582 38336
rect 289026 2420 289262 2656
rect 289346 2420 289582 2656
rect 289026 2100 289262 2336
rect 289346 2100 289582 2336
rect 289026 -580 289262 -344
rect 289346 -580 289582 -344
rect 289026 -900 289262 -664
rect 289346 -900 289582 -664
rect 290266 705564 290502 705800
rect 290586 705564 290822 705800
rect 290266 705244 290502 705480
rect 290586 705244 290822 705480
rect 290266 687660 290502 687896
rect 290586 687660 290822 687896
rect 290266 687340 290502 687576
rect 290586 687340 290822 687576
rect 290266 651660 290502 651896
rect 290586 651660 290822 651896
rect 290266 651340 290502 651576
rect 290586 651340 290822 651576
rect 290266 615660 290502 615896
rect 290586 615660 290822 615896
rect 290266 615340 290502 615576
rect 290586 615340 290822 615576
rect 290266 579660 290502 579896
rect 290586 579660 290822 579896
rect 290266 579340 290502 579576
rect 290586 579340 290822 579576
rect 290266 543660 290502 543896
rect 290586 543660 290822 543896
rect 290266 543340 290502 543576
rect 290586 543340 290822 543576
rect 290266 507660 290502 507896
rect 290586 507660 290822 507896
rect 290266 507340 290502 507576
rect 290586 507340 290822 507576
rect 290266 471660 290502 471896
rect 290586 471660 290822 471896
rect 290266 471340 290502 471576
rect 290586 471340 290822 471576
rect 290266 435660 290502 435896
rect 290586 435660 290822 435896
rect 290266 435340 290502 435576
rect 290586 435340 290822 435576
rect 290266 399660 290502 399896
rect 290586 399660 290822 399896
rect 290266 399340 290502 399576
rect 290586 399340 290822 399576
rect 290266 363660 290502 363896
rect 290586 363660 290822 363896
rect 290266 363340 290502 363576
rect 290586 363340 290822 363576
rect 290266 327660 290502 327896
rect 290586 327660 290822 327896
rect 290266 327340 290502 327576
rect 290586 327340 290822 327576
rect 290266 291660 290502 291896
rect 290586 291660 290822 291896
rect 290266 291340 290502 291576
rect 290586 291340 290822 291576
rect 290266 255660 290502 255896
rect 290586 255660 290822 255896
rect 290266 255340 290502 255576
rect 290586 255340 290822 255576
rect 290266 219660 290502 219896
rect 290586 219660 290822 219896
rect 290266 219340 290502 219576
rect 290586 219340 290822 219576
rect 290266 183660 290502 183896
rect 290586 183660 290822 183896
rect 290266 183340 290502 183576
rect 290586 183340 290822 183576
rect 290266 147660 290502 147896
rect 290586 147660 290822 147896
rect 290266 147340 290502 147576
rect 290586 147340 290822 147576
rect 290266 111660 290502 111896
rect 290586 111660 290822 111896
rect 290266 111340 290502 111576
rect 290586 111340 290822 111576
rect 290266 75660 290502 75896
rect 290586 75660 290822 75896
rect 290266 75340 290502 75576
rect 290586 75340 290822 75576
rect 290266 39660 290502 39896
rect 290586 39660 290822 39896
rect 290266 39340 290502 39576
rect 290586 39340 290822 39576
rect 290266 3660 290502 3896
rect 290586 3660 290822 3896
rect 290266 3340 290502 3576
rect 290586 3340 290822 3576
rect 290266 -1540 290502 -1304
rect 290586 -1540 290822 -1304
rect 290266 -1860 290502 -1624
rect 290586 -1860 290822 -1624
rect 291506 706524 291742 706760
rect 291826 706524 292062 706760
rect 291506 706204 291742 706440
rect 291826 706204 292062 706440
rect 291506 688900 291742 689136
rect 291826 688900 292062 689136
rect 291506 688580 291742 688816
rect 291826 688580 292062 688816
rect 291506 652900 291742 653136
rect 291826 652900 292062 653136
rect 291506 652580 291742 652816
rect 291826 652580 292062 652816
rect 291506 616900 291742 617136
rect 291826 616900 292062 617136
rect 291506 616580 291742 616816
rect 291826 616580 292062 616816
rect 291506 580900 291742 581136
rect 291826 580900 292062 581136
rect 291506 580580 291742 580816
rect 291826 580580 292062 580816
rect 291506 544900 291742 545136
rect 291826 544900 292062 545136
rect 291506 544580 291742 544816
rect 291826 544580 292062 544816
rect 291506 508900 291742 509136
rect 291826 508900 292062 509136
rect 291506 508580 291742 508816
rect 291826 508580 292062 508816
rect 291506 472900 291742 473136
rect 291826 472900 292062 473136
rect 291506 472580 291742 472816
rect 291826 472580 292062 472816
rect 291506 436900 291742 437136
rect 291826 436900 292062 437136
rect 291506 436580 291742 436816
rect 291826 436580 292062 436816
rect 291506 400900 291742 401136
rect 291826 400900 292062 401136
rect 291506 400580 291742 400816
rect 291826 400580 292062 400816
rect 291506 364900 291742 365136
rect 291826 364900 292062 365136
rect 291506 364580 291742 364816
rect 291826 364580 292062 364816
rect 291506 328900 291742 329136
rect 291826 328900 292062 329136
rect 291506 328580 291742 328816
rect 291826 328580 292062 328816
rect 291506 292900 291742 293136
rect 291826 292900 292062 293136
rect 291506 292580 291742 292816
rect 291826 292580 292062 292816
rect 291506 256900 291742 257136
rect 291826 256900 292062 257136
rect 291506 256580 291742 256816
rect 291826 256580 292062 256816
rect 291506 220900 291742 221136
rect 291826 220900 292062 221136
rect 291506 220580 291742 220816
rect 291826 220580 292062 220816
rect 291506 184900 291742 185136
rect 291826 184900 292062 185136
rect 291506 184580 291742 184816
rect 291826 184580 292062 184816
rect 291506 148900 291742 149136
rect 291826 148900 292062 149136
rect 291506 148580 291742 148816
rect 291826 148580 292062 148816
rect 291506 112900 291742 113136
rect 291826 112900 292062 113136
rect 291506 112580 291742 112816
rect 291826 112580 292062 112816
rect 291506 76900 291742 77136
rect 291826 76900 292062 77136
rect 291506 76580 291742 76816
rect 291826 76580 292062 76816
rect 291506 40900 291742 41136
rect 291826 40900 292062 41136
rect 291506 40580 291742 40816
rect 291826 40580 292062 40816
rect 291506 4900 291742 5136
rect 291826 4900 292062 5136
rect 291506 4580 291742 4816
rect 291826 4580 292062 4816
rect 291506 -2500 291742 -2264
rect 291826 -2500 292062 -2264
rect 291506 -2820 291742 -2584
rect 291826 -2820 292062 -2584
rect 292746 707484 292982 707720
rect 293066 707484 293302 707720
rect 292746 707164 292982 707400
rect 293066 707164 293302 707400
rect 292746 690140 292982 690376
rect 293066 690140 293302 690376
rect 292746 689820 292982 690056
rect 293066 689820 293302 690056
rect 292746 654140 292982 654376
rect 293066 654140 293302 654376
rect 292746 653820 292982 654056
rect 293066 653820 293302 654056
rect 292746 618140 292982 618376
rect 293066 618140 293302 618376
rect 292746 617820 292982 618056
rect 293066 617820 293302 618056
rect 292746 582140 292982 582376
rect 293066 582140 293302 582376
rect 292746 581820 292982 582056
rect 293066 581820 293302 582056
rect 292746 546140 292982 546376
rect 293066 546140 293302 546376
rect 292746 545820 292982 546056
rect 293066 545820 293302 546056
rect 292746 510140 292982 510376
rect 293066 510140 293302 510376
rect 292746 509820 292982 510056
rect 293066 509820 293302 510056
rect 292746 474140 292982 474376
rect 293066 474140 293302 474376
rect 292746 473820 292982 474056
rect 293066 473820 293302 474056
rect 292746 438140 292982 438376
rect 293066 438140 293302 438376
rect 292746 437820 292982 438056
rect 293066 437820 293302 438056
rect 292746 402140 292982 402376
rect 293066 402140 293302 402376
rect 292746 401820 292982 402056
rect 293066 401820 293302 402056
rect 292746 366140 292982 366376
rect 293066 366140 293302 366376
rect 292746 365820 292982 366056
rect 293066 365820 293302 366056
rect 292746 330140 292982 330376
rect 293066 330140 293302 330376
rect 292746 329820 292982 330056
rect 293066 329820 293302 330056
rect 292746 294140 292982 294376
rect 293066 294140 293302 294376
rect 292746 293820 292982 294056
rect 293066 293820 293302 294056
rect 292746 258140 292982 258376
rect 293066 258140 293302 258376
rect 292746 257820 292982 258056
rect 293066 257820 293302 258056
rect 292746 222140 292982 222376
rect 293066 222140 293302 222376
rect 292746 221820 292982 222056
rect 293066 221820 293302 222056
rect 292746 186140 292982 186376
rect 293066 186140 293302 186376
rect 292746 185820 292982 186056
rect 293066 185820 293302 186056
rect 292746 150140 292982 150376
rect 293066 150140 293302 150376
rect 292746 149820 292982 150056
rect 293066 149820 293302 150056
rect 292746 114140 292982 114376
rect 293066 114140 293302 114376
rect 292746 113820 292982 114056
rect 293066 113820 293302 114056
rect 292746 78140 292982 78376
rect 293066 78140 293302 78376
rect 292746 77820 292982 78056
rect 293066 77820 293302 78056
rect 292746 42140 292982 42376
rect 293066 42140 293302 42376
rect 292746 41820 292982 42056
rect 293066 41820 293302 42056
rect 292746 6140 292982 6376
rect 293066 6140 293302 6376
rect 292746 5820 292982 6056
rect 293066 5820 293302 6056
rect 292746 -3460 292982 -3224
rect 293066 -3460 293302 -3224
rect 292746 -3780 292982 -3544
rect 293066 -3780 293302 -3544
rect 293986 708444 294222 708680
rect 294306 708444 294542 708680
rect 293986 708124 294222 708360
rect 294306 708124 294542 708360
rect 293986 691380 294222 691616
rect 294306 691380 294542 691616
rect 293986 691060 294222 691296
rect 294306 691060 294542 691296
rect 293986 655380 294222 655616
rect 294306 655380 294542 655616
rect 293986 655060 294222 655296
rect 294306 655060 294542 655296
rect 293986 619380 294222 619616
rect 294306 619380 294542 619616
rect 293986 619060 294222 619296
rect 294306 619060 294542 619296
rect 293986 583380 294222 583616
rect 294306 583380 294542 583616
rect 293986 583060 294222 583296
rect 294306 583060 294542 583296
rect 293986 547380 294222 547616
rect 294306 547380 294542 547616
rect 293986 547060 294222 547296
rect 294306 547060 294542 547296
rect 293986 511380 294222 511616
rect 294306 511380 294542 511616
rect 293986 511060 294222 511296
rect 294306 511060 294542 511296
rect 293986 475380 294222 475616
rect 294306 475380 294542 475616
rect 293986 475060 294222 475296
rect 294306 475060 294542 475296
rect 293986 439380 294222 439616
rect 294306 439380 294542 439616
rect 293986 439060 294222 439296
rect 294306 439060 294542 439296
rect 293986 403380 294222 403616
rect 294306 403380 294542 403616
rect 293986 403060 294222 403296
rect 294306 403060 294542 403296
rect 293986 367380 294222 367616
rect 294306 367380 294542 367616
rect 293986 367060 294222 367296
rect 294306 367060 294542 367296
rect 293986 331380 294222 331616
rect 294306 331380 294542 331616
rect 293986 331060 294222 331296
rect 294306 331060 294542 331296
rect 293986 295380 294222 295616
rect 294306 295380 294542 295616
rect 293986 295060 294222 295296
rect 294306 295060 294542 295296
rect 293986 259380 294222 259616
rect 294306 259380 294542 259616
rect 293986 259060 294222 259296
rect 294306 259060 294542 259296
rect 293986 223380 294222 223616
rect 294306 223380 294542 223616
rect 293986 223060 294222 223296
rect 294306 223060 294542 223296
rect 293986 187380 294222 187616
rect 294306 187380 294542 187616
rect 293986 187060 294222 187296
rect 294306 187060 294542 187296
rect 293986 151380 294222 151616
rect 294306 151380 294542 151616
rect 293986 151060 294222 151296
rect 294306 151060 294542 151296
rect 293986 115380 294222 115616
rect 294306 115380 294542 115616
rect 293986 115060 294222 115296
rect 294306 115060 294542 115296
rect 293986 79380 294222 79616
rect 294306 79380 294542 79616
rect 293986 79060 294222 79296
rect 294306 79060 294542 79296
rect 293986 43380 294222 43616
rect 294306 43380 294542 43616
rect 293986 43060 294222 43296
rect 294306 43060 294542 43296
rect 293986 7380 294222 7616
rect 294306 7380 294542 7616
rect 293986 7060 294222 7296
rect 294306 7060 294542 7296
rect 293986 -4420 294222 -4184
rect 294306 -4420 294542 -4184
rect 293986 -4740 294222 -4504
rect 294306 -4740 294542 -4504
rect 295226 709404 295462 709640
rect 295546 709404 295782 709640
rect 295226 709084 295462 709320
rect 295546 709084 295782 709320
rect 295226 692620 295462 692856
rect 295546 692620 295782 692856
rect 295226 692300 295462 692536
rect 295546 692300 295782 692536
rect 295226 656620 295462 656856
rect 295546 656620 295782 656856
rect 295226 656300 295462 656536
rect 295546 656300 295782 656536
rect 295226 620620 295462 620856
rect 295546 620620 295782 620856
rect 295226 620300 295462 620536
rect 295546 620300 295782 620536
rect 295226 584620 295462 584856
rect 295546 584620 295782 584856
rect 295226 584300 295462 584536
rect 295546 584300 295782 584536
rect 295226 548620 295462 548856
rect 295546 548620 295782 548856
rect 295226 548300 295462 548536
rect 295546 548300 295782 548536
rect 295226 512620 295462 512856
rect 295546 512620 295782 512856
rect 295226 512300 295462 512536
rect 295546 512300 295782 512536
rect 295226 476620 295462 476856
rect 295546 476620 295782 476856
rect 295226 476300 295462 476536
rect 295546 476300 295782 476536
rect 295226 440620 295462 440856
rect 295546 440620 295782 440856
rect 295226 440300 295462 440536
rect 295546 440300 295782 440536
rect 295226 404620 295462 404856
rect 295546 404620 295782 404856
rect 295226 404300 295462 404536
rect 295546 404300 295782 404536
rect 295226 368620 295462 368856
rect 295546 368620 295782 368856
rect 295226 368300 295462 368536
rect 295546 368300 295782 368536
rect 295226 332620 295462 332856
rect 295546 332620 295782 332856
rect 295226 332300 295462 332536
rect 295546 332300 295782 332536
rect 295226 296620 295462 296856
rect 295546 296620 295782 296856
rect 295226 296300 295462 296536
rect 295546 296300 295782 296536
rect 295226 260620 295462 260856
rect 295546 260620 295782 260856
rect 295226 260300 295462 260536
rect 295546 260300 295782 260536
rect 295226 224620 295462 224856
rect 295546 224620 295782 224856
rect 295226 224300 295462 224536
rect 295546 224300 295782 224536
rect 295226 188620 295462 188856
rect 295546 188620 295782 188856
rect 295226 188300 295462 188536
rect 295546 188300 295782 188536
rect 295226 152620 295462 152856
rect 295546 152620 295782 152856
rect 295226 152300 295462 152536
rect 295546 152300 295782 152536
rect 295226 116620 295462 116856
rect 295546 116620 295782 116856
rect 295226 116300 295462 116536
rect 295546 116300 295782 116536
rect 295226 80620 295462 80856
rect 295546 80620 295782 80856
rect 295226 80300 295462 80536
rect 295546 80300 295782 80536
rect 295226 44620 295462 44856
rect 295546 44620 295782 44856
rect 295226 44300 295462 44536
rect 295546 44300 295782 44536
rect 295226 8620 295462 8856
rect 295546 8620 295782 8856
rect 295226 8300 295462 8536
rect 295546 8300 295782 8536
rect 295226 -5380 295462 -5144
rect 295546 -5380 295782 -5144
rect 295226 -5700 295462 -5464
rect 295546 -5700 295782 -5464
rect 296466 710364 296702 710600
rect 296786 710364 297022 710600
rect 296466 710044 296702 710280
rect 296786 710044 297022 710280
rect 296466 693860 296702 694096
rect 296786 693860 297022 694096
rect 296466 693540 296702 693776
rect 296786 693540 297022 693776
rect 296466 657860 296702 658096
rect 296786 657860 297022 658096
rect 296466 657540 296702 657776
rect 296786 657540 297022 657776
rect 296466 621860 296702 622096
rect 296786 621860 297022 622096
rect 296466 621540 296702 621776
rect 296786 621540 297022 621776
rect 296466 585860 296702 586096
rect 296786 585860 297022 586096
rect 296466 585540 296702 585776
rect 296786 585540 297022 585776
rect 296466 549860 296702 550096
rect 296786 549860 297022 550096
rect 296466 549540 296702 549776
rect 296786 549540 297022 549776
rect 296466 513860 296702 514096
rect 296786 513860 297022 514096
rect 296466 513540 296702 513776
rect 296786 513540 297022 513776
rect 296466 477860 296702 478096
rect 296786 477860 297022 478096
rect 296466 477540 296702 477776
rect 296786 477540 297022 477776
rect 296466 441860 296702 442096
rect 296786 441860 297022 442096
rect 296466 441540 296702 441776
rect 296786 441540 297022 441776
rect 296466 405860 296702 406096
rect 296786 405860 297022 406096
rect 296466 405540 296702 405776
rect 296786 405540 297022 405776
rect 296466 369860 296702 370096
rect 296786 369860 297022 370096
rect 296466 369540 296702 369776
rect 296786 369540 297022 369776
rect 296466 333860 296702 334096
rect 296786 333860 297022 334096
rect 296466 333540 296702 333776
rect 296786 333540 297022 333776
rect 296466 297860 296702 298096
rect 296786 297860 297022 298096
rect 296466 297540 296702 297776
rect 296786 297540 297022 297776
rect 296466 261860 296702 262096
rect 296786 261860 297022 262096
rect 296466 261540 296702 261776
rect 296786 261540 297022 261776
rect 296466 225860 296702 226096
rect 296786 225860 297022 226096
rect 296466 225540 296702 225776
rect 296786 225540 297022 225776
rect 296466 189860 296702 190096
rect 296786 189860 297022 190096
rect 296466 189540 296702 189776
rect 296786 189540 297022 189776
rect 296466 153860 296702 154096
rect 296786 153860 297022 154096
rect 296466 153540 296702 153776
rect 296786 153540 297022 153776
rect 296466 117860 296702 118096
rect 296786 117860 297022 118096
rect 296466 117540 296702 117776
rect 296786 117540 297022 117776
rect 296466 81860 296702 82096
rect 296786 81860 297022 82096
rect 296466 81540 296702 81776
rect 296786 81540 297022 81776
rect 296466 45860 296702 46096
rect 296786 45860 297022 46096
rect 296466 45540 296702 45776
rect 296786 45540 297022 45776
rect 296466 9860 296702 10096
rect 296786 9860 297022 10096
rect 296466 9540 296702 9776
rect 296786 9540 297022 9776
rect 296466 -6340 296702 -6104
rect 296786 -6340 297022 -6104
rect 296466 -6660 296702 -6424
rect 296786 -6660 297022 -6424
rect 297706 711324 297942 711560
rect 298026 711324 298262 711560
rect 297706 711004 297942 711240
rect 298026 711004 298262 711240
rect 297706 695100 297942 695336
rect 298026 695100 298262 695336
rect 297706 694780 297942 695016
rect 298026 694780 298262 695016
rect 297706 659100 297942 659336
rect 298026 659100 298262 659336
rect 297706 658780 297942 659016
rect 298026 658780 298262 659016
rect 297706 623100 297942 623336
rect 298026 623100 298262 623336
rect 297706 622780 297942 623016
rect 298026 622780 298262 623016
rect 297706 587100 297942 587336
rect 298026 587100 298262 587336
rect 297706 586780 297942 587016
rect 298026 586780 298262 587016
rect 297706 551100 297942 551336
rect 298026 551100 298262 551336
rect 297706 550780 297942 551016
rect 298026 550780 298262 551016
rect 297706 515100 297942 515336
rect 298026 515100 298262 515336
rect 297706 514780 297942 515016
rect 298026 514780 298262 515016
rect 297706 479100 297942 479336
rect 298026 479100 298262 479336
rect 297706 478780 297942 479016
rect 298026 478780 298262 479016
rect 297706 443100 297942 443336
rect 298026 443100 298262 443336
rect 297706 442780 297942 443016
rect 298026 442780 298262 443016
rect 297706 407100 297942 407336
rect 298026 407100 298262 407336
rect 297706 406780 297942 407016
rect 298026 406780 298262 407016
rect 297706 371100 297942 371336
rect 298026 371100 298262 371336
rect 297706 370780 297942 371016
rect 298026 370780 298262 371016
rect 297706 335100 297942 335336
rect 298026 335100 298262 335336
rect 297706 334780 297942 335016
rect 298026 334780 298262 335016
rect 297706 299100 297942 299336
rect 298026 299100 298262 299336
rect 297706 298780 297942 299016
rect 298026 298780 298262 299016
rect 297706 263100 297942 263336
rect 298026 263100 298262 263336
rect 297706 262780 297942 263016
rect 298026 262780 298262 263016
rect 297706 227100 297942 227336
rect 298026 227100 298262 227336
rect 297706 226780 297942 227016
rect 298026 226780 298262 227016
rect 297706 191100 297942 191336
rect 298026 191100 298262 191336
rect 297706 190780 297942 191016
rect 298026 190780 298262 191016
rect 297706 155100 297942 155336
rect 298026 155100 298262 155336
rect 297706 154780 297942 155016
rect 298026 154780 298262 155016
rect 297706 119100 297942 119336
rect 298026 119100 298262 119336
rect 297706 118780 297942 119016
rect 298026 118780 298262 119016
rect 297706 83100 297942 83336
rect 298026 83100 298262 83336
rect 297706 82780 297942 83016
rect 298026 82780 298262 83016
rect 297706 47100 297942 47336
rect 298026 47100 298262 47336
rect 297706 46780 297942 47016
rect 298026 46780 298262 47016
rect 297706 11100 297942 11336
rect 298026 11100 298262 11336
rect 297706 10780 297942 11016
rect 298026 10780 298262 11016
rect 297706 -7300 297942 -7064
rect 298026 -7300 298262 -7064
rect 297706 -7620 297942 -7384
rect 298026 -7620 298262 -7384
rect 325026 704604 325262 704840
rect 325346 704604 325582 704840
rect 325026 704284 325262 704520
rect 325346 704284 325582 704520
rect 325026 686420 325262 686656
rect 325346 686420 325582 686656
rect 325026 686100 325262 686336
rect 325346 686100 325582 686336
rect 325026 650420 325262 650656
rect 325346 650420 325582 650656
rect 325026 650100 325262 650336
rect 325346 650100 325582 650336
rect 325026 614420 325262 614656
rect 325346 614420 325582 614656
rect 325026 614100 325262 614336
rect 325346 614100 325582 614336
rect 325026 578420 325262 578656
rect 325346 578420 325582 578656
rect 325026 578100 325262 578336
rect 325346 578100 325582 578336
rect 325026 542420 325262 542656
rect 325346 542420 325582 542656
rect 325026 542100 325262 542336
rect 325346 542100 325582 542336
rect 325026 506420 325262 506656
rect 325346 506420 325582 506656
rect 325026 506100 325262 506336
rect 325346 506100 325582 506336
rect 325026 470420 325262 470656
rect 325346 470420 325582 470656
rect 325026 470100 325262 470336
rect 325346 470100 325582 470336
rect 325026 434420 325262 434656
rect 325346 434420 325582 434656
rect 325026 434100 325262 434336
rect 325346 434100 325582 434336
rect 325026 398420 325262 398656
rect 325346 398420 325582 398656
rect 325026 398100 325262 398336
rect 325346 398100 325582 398336
rect 325026 362420 325262 362656
rect 325346 362420 325582 362656
rect 325026 362100 325262 362336
rect 325346 362100 325582 362336
rect 325026 326420 325262 326656
rect 325346 326420 325582 326656
rect 325026 326100 325262 326336
rect 325346 326100 325582 326336
rect 325026 290420 325262 290656
rect 325346 290420 325582 290656
rect 325026 290100 325262 290336
rect 325346 290100 325582 290336
rect 325026 254420 325262 254656
rect 325346 254420 325582 254656
rect 325026 254100 325262 254336
rect 325346 254100 325582 254336
rect 325026 218420 325262 218656
rect 325346 218420 325582 218656
rect 325026 218100 325262 218336
rect 325346 218100 325582 218336
rect 325026 182420 325262 182656
rect 325346 182420 325582 182656
rect 325026 182100 325262 182336
rect 325346 182100 325582 182336
rect 325026 146420 325262 146656
rect 325346 146420 325582 146656
rect 325026 146100 325262 146336
rect 325346 146100 325582 146336
rect 325026 110420 325262 110656
rect 325346 110420 325582 110656
rect 325026 110100 325262 110336
rect 325346 110100 325582 110336
rect 325026 74420 325262 74656
rect 325346 74420 325582 74656
rect 325026 74100 325262 74336
rect 325346 74100 325582 74336
rect 325026 38420 325262 38656
rect 325346 38420 325582 38656
rect 325026 38100 325262 38336
rect 325346 38100 325582 38336
rect 325026 2420 325262 2656
rect 325346 2420 325582 2656
rect 325026 2100 325262 2336
rect 325346 2100 325582 2336
rect 325026 -580 325262 -344
rect 325346 -580 325582 -344
rect 325026 -900 325262 -664
rect 325346 -900 325582 -664
rect 326266 705564 326502 705800
rect 326586 705564 326822 705800
rect 326266 705244 326502 705480
rect 326586 705244 326822 705480
rect 326266 687660 326502 687896
rect 326586 687660 326822 687896
rect 326266 687340 326502 687576
rect 326586 687340 326822 687576
rect 326266 651660 326502 651896
rect 326586 651660 326822 651896
rect 326266 651340 326502 651576
rect 326586 651340 326822 651576
rect 326266 615660 326502 615896
rect 326586 615660 326822 615896
rect 326266 615340 326502 615576
rect 326586 615340 326822 615576
rect 326266 579660 326502 579896
rect 326586 579660 326822 579896
rect 326266 579340 326502 579576
rect 326586 579340 326822 579576
rect 326266 543660 326502 543896
rect 326586 543660 326822 543896
rect 326266 543340 326502 543576
rect 326586 543340 326822 543576
rect 326266 507660 326502 507896
rect 326586 507660 326822 507896
rect 326266 507340 326502 507576
rect 326586 507340 326822 507576
rect 326266 471660 326502 471896
rect 326586 471660 326822 471896
rect 326266 471340 326502 471576
rect 326586 471340 326822 471576
rect 326266 435660 326502 435896
rect 326586 435660 326822 435896
rect 326266 435340 326502 435576
rect 326586 435340 326822 435576
rect 326266 399660 326502 399896
rect 326586 399660 326822 399896
rect 326266 399340 326502 399576
rect 326586 399340 326822 399576
rect 326266 363660 326502 363896
rect 326586 363660 326822 363896
rect 326266 363340 326502 363576
rect 326586 363340 326822 363576
rect 326266 327660 326502 327896
rect 326586 327660 326822 327896
rect 326266 327340 326502 327576
rect 326586 327340 326822 327576
rect 326266 291660 326502 291896
rect 326586 291660 326822 291896
rect 326266 291340 326502 291576
rect 326586 291340 326822 291576
rect 326266 255660 326502 255896
rect 326586 255660 326822 255896
rect 326266 255340 326502 255576
rect 326586 255340 326822 255576
rect 326266 219660 326502 219896
rect 326586 219660 326822 219896
rect 326266 219340 326502 219576
rect 326586 219340 326822 219576
rect 326266 183660 326502 183896
rect 326586 183660 326822 183896
rect 326266 183340 326502 183576
rect 326586 183340 326822 183576
rect 326266 147660 326502 147896
rect 326586 147660 326822 147896
rect 326266 147340 326502 147576
rect 326586 147340 326822 147576
rect 326266 111660 326502 111896
rect 326586 111660 326822 111896
rect 326266 111340 326502 111576
rect 326586 111340 326822 111576
rect 326266 75660 326502 75896
rect 326586 75660 326822 75896
rect 326266 75340 326502 75576
rect 326586 75340 326822 75576
rect 326266 39660 326502 39896
rect 326586 39660 326822 39896
rect 326266 39340 326502 39576
rect 326586 39340 326822 39576
rect 326266 3660 326502 3896
rect 326586 3660 326822 3896
rect 326266 3340 326502 3576
rect 326586 3340 326822 3576
rect 326266 -1540 326502 -1304
rect 326586 -1540 326822 -1304
rect 326266 -1860 326502 -1624
rect 326586 -1860 326822 -1624
rect 327506 706524 327742 706760
rect 327826 706524 328062 706760
rect 327506 706204 327742 706440
rect 327826 706204 328062 706440
rect 327506 688900 327742 689136
rect 327826 688900 328062 689136
rect 327506 688580 327742 688816
rect 327826 688580 328062 688816
rect 327506 652900 327742 653136
rect 327826 652900 328062 653136
rect 327506 652580 327742 652816
rect 327826 652580 328062 652816
rect 327506 616900 327742 617136
rect 327826 616900 328062 617136
rect 327506 616580 327742 616816
rect 327826 616580 328062 616816
rect 327506 580900 327742 581136
rect 327826 580900 328062 581136
rect 327506 580580 327742 580816
rect 327826 580580 328062 580816
rect 327506 544900 327742 545136
rect 327826 544900 328062 545136
rect 327506 544580 327742 544816
rect 327826 544580 328062 544816
rect 327506 508900 327742 509136
rect 327826 508900 328062 509136
rect 327506 508580 327742 508816
rect 327826 508580 328062 508816
rect 327506 472900 327742 473136
rect 327826 472900 328062 473136
rect 327506 472580 327742 472816
rect 327826 472580 328062 472816
rect 327506 436900 327742 437136
rect 327826 436900 328062 437136
rect 327506 436580 327742 436816
rect 327826 436580 328062 436816
rect 327506 400900 327742 401136
rect 327826 400900 328062 401136
rect 327506 400580 327742 400816
rect 327826 400580 328062 400816
rect 327506 364900 327742 365136
rect 327826 364900 328062 365136
rect 327506 364580 327742 364816
rect 327826 364580 328062 364816
rect 327506 328900 327742 329136
rect 327826 328900 328062 329136
rect 327506 328580 327742 328816
rect 327826 328580 328062 328816
rect 327506 292900 327742 293136
rect 327826 292900 328062 293136
rect 327506 292580 327742 292816
rect 327826 292580 328062 292816
rect 327506 256900 327742 257136
rect 327826 256900 328062 257136
rect 327506 256580 327742 256816
rect 327826 256580 328062 256816
rect 327506 220900 327742 221136
rect 327826 220900 328062 221136
rect 327506 220580 327742 220816
rect 327826 220580 328062 220816
rect 327506 184900 327742 185136
rect 327826 184900 328062 185136
rect 327506 184580 327742 184816
rect 327826 184580 328062 184816
rect 327506 148900 327742 149136
rect 327826 148900 328062 149136
rect 327506 148580 327742 148816
rect 327826 148580 328062 148816
rect 327506 112900 327742 113136
rect 327826 112900 328062 113136
rect 327506 112580 327742 112816
rect 327826 112580 328062 112816
rect 327506 76900 327742 77136
rect 327826 76900 328062 77136
rect 327506 76580 327742 76816
rect 327826 76580 328062 76816
rect 327506 40900 327742 41136
rect 327826 40900 328062 41136
rect 327506 40580 327742 40816
rect 327826 40580 328062 40816
rect 327506 4900 327742 5136
rect 327826 4900 328062 5136
rect 327506 4580 327742 4816
rect 327826 4580 328062 4816
rect 327506 -2500 327742 -2264
rect 327826 -2500 328062 -2264
rect 327506 -2820 327742 -2584
rect 327826 -2820 328062 -2584
rect 328746 707484 328982 707720
rect 329066 707484 329302 707720
rect 328746 707164 328982 707400
rect 329066 707164 329302 707400
rect 328746 690140 328982 690376
rect 329066 690140 329302 690376
rect 328746 689820 328982 690056
rect 329066 689820 329302 690056
rect 328746 654140 328982 654376
rect 329066 654140 329302 654376
rect 328746 653820 328982 654056
rect 329066 653820 329302 654056
rect 328746 618140 328982 618376
rect 329066 618140 329302 618376
rect 328746 617820 328982 618056
rect 329066 617820 329302 618056
rect 328746 582140 328982 582376
rect 329066 582140 329302 582376
rect 328746 581820 328982 582056
rect 329066 581820 329302 582056
rect 328746 546140 328982 546376
rect 329066 546140 329302 546376
rect 328746 545820 328982 546056
rect 329066 545820 329302 546056
rect 328746 510140 328982 510376
rect 329066 510140 329302 510376
rect 328746 509820 328982 510056
rect 329066 509820 329302 510056
rect 328746 474140 328982 474376
rect 329066 474140 329302 474376
rect 328746 473820 328982 474056
rect 329066 473820 329302 474056
rect 328746 438140 328982 438376
rect 329066 438140 329302 438376
rect 328746 437820 328982 438056
rect 329066 437820 329302 438056
rect 328746 402140 328982 402376
rect 329066 402140 329302 402376
rect 328746 401820 328982 402056
rect 329066 401820 329302 402056
rect 328746 366140 328982 366376
rect 329066 366140 329302 366376
rect 328746 365820 328982 366056
rect 329066 365820 329302 366056
rect 328746 330140 328982 330376
rect 329066 330140 329302 330376
rect 328746 329820 328982 330056
rect 329066 329820 329302 330056
rect 328746 294140 328982 294376
rect 329066 294140 329302 294376
rect 328746 293820 328982 294056
rect 329066 293820 329302 294056
rect 328746 258140 328982 258376
rect 329066 258140 329302 258376
rect 328746 257820 328982 258056
rect 329066 257820 329302 258056
rect 328746 222140 328982 222376
rect 329066 222140 329302 222376
rect 328746 221820 328982 222056
rect 329066 221820 329302 222056
rect 328746 186140 328982 186376
rect 329066 186140 329302 186376
rect 328746 185820 328982 186056
rect 329066 185820 329302 186056
rect 328746 150140 328982 150376
rect 329066 150140 329302 150376
rect 328746 149820 328982 150056
rect 329066 149820 329302 150056
rect 328746 114140 328982 114376
rect 329066 114140 329302 114376
rect 328746 113820 328982 114056
rect 329066 113820 329302 114056
rect 328746 78140 328982 78376
rect 329066 78140 329302 78376
rect 328746 77820 328982 78056
rect 329066 77820 329302 78056
rect 328746 42140 328982 42376
rect 329066 42140 329302 42376
rect 328746 41820 328982 42056
rect 329066 41820 329302 42056
rect 328746 6140 328982 6376
rect 329066 6140 329302 6376
rect 328746 5820 328982 6056
rect 329066 5820 329302 6056
rect 328746 -3460 328982 -3224
rect 329066 -3460 329302 -3224
rect 328746 -3780 328982 -3544
rect 329066 -3780 329302 -3544
rect 329986 708444 330222 708680
rect 330306 708444 330542 708680
rect 329986 708124 330222 708360
rect 330306 708124 330542 708360
rect 329986 691380 330222 691616
rect 330306 691380 330542 691616
rect 329986 691060 330222 691296
rect 330306 691060 330542 691296
rect 329986 655380 330222 655616
rect 330306 655380 330542 655616
rect 329986 655060 330222 655296
rect 330306 655060 330542 655296
rect 329986 619380 330222 619616
rect 330306 619380 330542 619616
rect 329986 619060 330222 619296
rect 330306 619060 330542 619296
rect 329986 583380 330222 583616
rect 330306 583380 330542 583616
rect 329986 583060 330222 583296
rect 330306 583060 330542 583296
rect 329986 547380 330222 547616
rect 330306 547380 330542 547616
rect 329986 547060 330222 547296
rect 330306 547060 330542 547296
rect 329986 511380 330222 511616
rect 330306 511380 330542 511616
rect 329986 511060 330222 511296
rect 330306 511060 330542 511296
rect 329986 475380 330222 475616
rect 330306 475380 330542 475616
rect 329986 475060 330222 475296
rect 330306 475060 330542 475296
rect 329986 439380 330222 439616
rect 330306 439380 330542 439616
rect 329986 439060 330222 439296
rect 330306 439060 330542 439296
rect 329986 403380 330222 403616
rect 330306 403380 330542 403616
rect 329986 403060 330222 403296
rect 330306 403060 330542 403296
rect 329986 367380 330222 367616
rect 330306 367380 330542 367616
rect 329986 367060 330222 367296
rect 330306 367060 330542 367296
rect 329986 331380 330222 331616
rect 330306 331380 330542 331616
rect 329986 331060 330222 331296
rect 330306 331060 330542 331296
rect 329986 295380 330222 295616
rect 330306 295380 330542 295616
rect 329986 295060 330222 295296
rect 330306 295060 330542 295296
rect 329986 259380 330222 259616
rect 330306 259380 330542 259616
rect 329986 259060 330222 259296
rect 330306 259060 330542 259296
rect 329986 223380 330222 223616
rect 330306 223380 330542 223616
rect 329986 223060 330222 223296
rect 330306 223060 330542 223296
rect 329986 187380 330222 187616
rect 330306 187380 330542 187616
rect 329986 187060 330222 187296
rect 330306 187060 330542 187296
rect 329986 151380 330222 151616
rect 330306 151380 330542 151616
rect 329986 151060 330222 151296
rect 330306 151060 330542 151296
rect 329986 115380 330222 115616
rect 330306 115380 330542 115616
rect 329986 115060 330222 115296
rect 330306 115060 330542 115296
rect 329986 79380 330222 79616
rect 330306 79380 330542 79616
rect 329986 79060 330222 79296
rect 330306 79060 330542 79296
rect 329986 43380 330222 43616
rect 330306 43380 330542 43616
rect 329986 43060 330222 43296
rect 330306 43060 330542 43296
rect 329986 7380 330222 7616
rect 330306 7380 330542 7616
rect 329986 7060 330222 7296
rect 330306 7060 330542 7296
rect 329986 -4420 330222 -4184
rect 330306 -4420 330542 -4184
rect 329986 -4740 330222 -4504
rect 330306 -4740 330542 -4504
rect 331226 709404 331462 709640
rect 331546 709404 331782 709640
rect 331226 709084 331462 709320
rect 331546 709084 331782 709320
rect 331226 692620 331462 692856
rect 331546 692620 331782 692856
rect 331226 692300 331462 692536
rect 331546 692300 331782 692536
rect 331226 656620 331462 656856
rect 331546 656620 331782 656856
rect 331226 656300 331462 656536
rect 331546 656300 331782 656536
rect 331226 620620 331462 620856
rect 331546 620620 331782 620856
rect 331226 620300 331462 620536
rect 331546 620300 331782 620536
rect 331226 584620 331462 584856
rect 331546 584620 331782 584856
rect 331226 584300 331462 584536
rect 331546 584300 331782 584536
rect 331226 548620 331462 548856
rect 331546 548620 331782 548856
rect 331226 548300 331462 548536
rect 331546 548300 331782 548536
rect 331226 512620 331462 512856
rect 331546 512620 331782 512856
rect 331226 512300 331462 512536
rect 331546 512300 331782 512536
rect 331226 476620 331462 476856
rect 331546 476620 331782 476856
rect 331226 476300 331462 476536
rect 331546 476300 331782 476536
rect 331226 440620 331462 440856
rect 331546 440620 331782 440856
rect 331226 440300 331462 440536
rect 331546 440300 331782 440536
rect 331226 404620 331462 404856
rect 331546 404620 331782 404856
rect 331226 404300 331462 404536
rect 331546 404300 331782 404536
rect 331226 368620 331462 368856
rect 331546 368620 331782 368856
rect 331226 368300 331462 368536
rect 331546 368300 331782 368536
rect 331226 332620 331462 332856
rect 331546 332620 331782 332856
rect 331226 332300 331462 332536
rect 331546 332300 331782 332536
rect 331226 296620 331462 296856
rect 331546 296620 331782 296856
rect 331226 296300 331462 296536
rect 331546 296300 331782 296536
rect 331226 260620 331462 260856
rect 331546 260620 331782 260856
rect 331226 260300 331462 260536
rect 331546 260300 331782 260536
rect 331226 224620 331462 224856
rect 331546 224620 331782 224856
rect 331226 224300 331462 224536
rect 331546 224300 331782 224536
rect 331226 188620 331462 188856
rect 331546 188620 331782 188856
rect 331226 188300 331462 188536
rect 331546 188300 331782 188536
rect 331226 152620 331462 152856
rect 331546 152620 331782 152856
rect 331226 152300 331462 152536
rect 331546 152300 331782 152536
rect 331226 116620 331462 116856
rect 331546 116620 331782 116856
rect 331226 116300 331462 116536
rect 331546 116300 331782 116536
rect 331226 80620 331462 80856
rect 331546 80620 331782 80856
rect 331226 80300 331462 80536
rect 331546 80300 331782 80536
rect 331226 44620 331462 44856
rect 331546 44620 331782 44856
rect 331226 44300 331462 44536
rect 331546 44300 331782 44536
rect 331226 8620 331462 8856
rect 331546 8620 331782 8856
rect 331226 8300 331462 8536
rect 331546 8300 331782 8536
rect 331226 -5380 331462 -5144
rect 331546 -5380 331782 -5144
rect 331226 -5700 331462 -5464
rect 331546 -5700 331782 -5464
rect 332466 710364 332702 710600
rect 332786 710364 333022 710600
rect 332466 710044 332702 710280
rect 332786 710044 333022 710280
rect 332466 693860 332702 694096
rect 332786 693860 333022 694096
rect 332466 693540 332702 693776
rect 332786 693540 333022 693776
rect 332466 657860 332702 658096
rect 332786 657860 333022 658096
rect 332466 657540 332702 657776
rect 332786 657540 333022 657776
rect 332466 621860 332702 622096
rect 332786 621860 333022 622096
rect 332466 621540 332702 621776
rect 332786 621540 333022 621776
rect 332466 585860 332702 586096
rect 332786 585860 333022 586096
rect 332466 585540 332702 585776
rect 332786 585540 333022 585776
rect 332466 549860 332702 550096
rect 332786 549860 333022 550096
rect 332466 549540 332702 549776
rect 332786 549540 333022 549776
rect 332466 513860 332702 514096
rect 332786 513860 333022 514096
rect 332466 513540 332702 513776
rect 332786 513540 333022 513776
rect 332466 477860 332702 478096
rect 332786 477860 333022 478096
rect 332466 477540 332702 477776
rect 332786 477540 333022 477776
rect 332466 441860 332702 442096
rect 332786 441860 333022 442096
rect 332466 441540 332702 441776
rect 332786 441540 333022 441776
rect 332466 405860 332702 406096
rect 332786 405860 333022 406096
rect 332466 405540 332702 405776
rect 332786 405540 333022 405776
rect 332466 369860 332702 370096
rect 332786 369860 333022 370096
rect 332466 369540 332702 369776
rect 332786 369540 333022 369776
rect 332466 333860 332702 334096
rect 332786 333860 333022 334096
rect 332466 333540 332702 333776
rect 332786 333540 333022 333776
rect 332466 297860 332702 298096
rect 332786 297860 333022 298096
rect 332466 297540 332702 297776
rect 332786 297540 333022 297776
rect 332466 261860 332702 262096
rect 332786 261860 333022 262096
rect 332466 261540 332702 261776
rect 332786 261540 333022 261776
rect 332466 225860 332702 226096
rect 332786 225860 333022 226096
rect 332466 225540 332702 225776
rect 332786 225540 333022 225776
rect 332466 189860 332702 190096
rect 332786 189860 333022 190096
rect 332466 189540 332702 189776
rect 332786 189540 333022 189776
rect 332466 153860 332702 154096
rect 332786 153860 333022 154096
rect 332466 153540 332702 153776
rect 332786 153540 333022 153776
rect 332466 117860 332702 118096
rect 332786 117860 333022 118096
rect 332466 117540 332702 117776
rect 332786 117540 333022 117776
rect 332466 81860 332702 82096
rect 332786 81860 333022 82096
rect 332466 81540 332702 81776
rect 332786 81540 333022 81776
rect 332466 45860 332702 46096
rect 332786 45860 333022 46096
rect 332466 45540 332702 45776
rect 332786 45540 333022 45776
rect 332466 9860 332702 10096
rect 332786 9860 333022 10096
rect 332466 9540 332702 9776
rect 332786 9540 333022 9776
rect 332466 -6340 332702 -6104
rect 332786 -6340 333022 -6104
rect 332466 -6660 332702 -6424
rect 332786 -6660 333022 -6424
rect 333706 711324 333942 711560
rect 334026 711324 334262 711560
rect 333706 711004 333942 711240
rect 334026 711004 334262 711240
rect 333706 695100 333942 695336
rect 334026 695100 334262 695336
rect 333706 694780 333942 695016
rect 334026 694780 334262 695016
rect 333706 659100 333942 659336
rect 334026 659100 334262 659336
rect 333706 658780 333942 659016
rect 334026 658780 334262 659016
rect 333706 623100 333942 623336
rect 334026 623100 334262 623336
rect 333706 622780 333942 623016
rect 334026 622780 334262 623016
rect 333706 587100 333942 587336
rect 334026 587100 334262 587336
rect 333706 586780 333942 587016
rect 334026 586780 334262 587016
rect 333706 551100 333942 551336
rect 334026 551100 334262 551336
rect 333706 550780 333942 551016
rect 334026 550780 334262 551016
rect 333706 515100 333942 515336
rect 334026 515100 334262 515336
rect 333706 514780 333942 515016
rect 334026 514780 334262 515016
rect 333706 479100 333942 479336
rect 334026 479100 334262 479336
rect 333706 478780 333942 479016
rect 334026 478780 334262 479016
rect 333706 443100 333942 443336
rect 334026 443100 334262 443336
rect 333706 442780 333942 443016
rect 334026 442780 334262 443016
rect 333706 407100 333942 407336
rect 334026 407100 334262 407336
rect 333706 406780 333942 407016
rect 334026 406780 334262 407016
rect 333706 371100 333942 371336
rect 334026 371100 334262 371336
rect 333706 370780 333942 371016
rect 334026 370780 334262 371016
rect 333706 335100 333942 335336
rect 334026 335100 334262 335336
rect 333706 334780 333942 335016
rect 334026 334780 334262 335016
rect 333706 299100 333942 299336
rect 334026 299100 334262 299336
rect 333706 298780 333942 299016
rect 334026 298780 334262 299016
rect 333706 263100 333942 263336
rect 334026 263100 334262 263336
rect 333706 262780 333942 263016
rect 334026 262780 334262 263016
rect 333706 227100 333942 227336
rect 334026 227100 334262 227336
rect 333706 226780 333942 227016
rect 334026 226780 334262 227016
rect 333706 191100 333942 191336
rect 334026 191100 334262 191336
rect 333706 190780 333942 191016
rect 334026 190780 334262 191016
rect 333706 155100 333942 155336
rect 334026 155100 334262 155336
rect 333706 154780 333942 155016
rect 334026 154780 334262 155016
rect 333706 119100 333942 119336
rect 334026 119100 334262 119336
rect 333706 118780 333942 119016
rect 334026 118780 334262 119016
rect 333706 83100 333942 83336
rect 334026 83100 334262 83336
rect 333706 82780 333942 83016
rect 334026 82780 334262 83016
rect 333706 47100 333942 47336
rect 334026 47100 334262 47336
rect 333706 46780 333942 47016
rect 334026 46780 334262 47016
rect 333706 11100 333942 11336
rect 334026 11100 334262 11336
rect 333706 10780 333942 11016
rect 334026 10780 334262 11016
rect 333706 -7300 333942 -7064
rect 334026 -7300 334262 -7064
rect 333706 -7620 333942 -7384
rect 334026 -7620 334262 -7384
rect 361026 704604 361262 704840
rect 361346 704604 361582 704840
rect 361026 704284 361262 704520
rect 361346 704284 361582 704520
rect 361026 686420 361262 686656
rect 361346 686420 361582 686656
rect 361026 686100 361262 686336
rect 361346 686100 361582 686336
rect 361026 650420 361262 650656
rect 361346 650420 361582 650656
rect 361026 650100 361262 650336
rect 361346 650100 361582 650336
rect 361026 614420 361262 614656
rect 361346 614420 361582 614656
rect 361026 614100 361262 614336
rect 361346 614100 361582 614336
rect 361026 578420 361262 578656
rect 361346 578420 361582 578656
rect 361026 578100 361262 578336
rect 361346 578100 361582 578336
rect 361026 542420 361262 542656
rect 361346 542420 361582 542656
rect 361026 542100 361262 542336
rect 361346 542100 361582 542336
rect 361026 506420 361262 506656
rect 361346 506420 361582 506656
rect 361026 506100 361262 506336
rect 361346 506100 361582 506336
rect 361026 470420 361262 470656
rect 361346 470420 361582 470656
rect 361026 470100 361262 470336
rect 361346 470100 361582 470336
rect 361026 434420 361262 434656
rect 361346 434420 361582 434656
rect 361026 434100 361262 434336
rect 361346 434100 361582 434336
rect 361026 398420 361262 398656
rect 361346 398420 361582 398656
rect 361026 398100 361262 398336
rect 361346 398100 361582 398336
rect 361026 362420 361262 362656
rect 361346 362420 361582 362656
rect 361026 362100 361262 362336
rect 361346 362100 361582 362336
rect 361026 326420 361262 326656
rect 361346 326420 361582 326656
rect 361026 326100 361262 326336
rect 361346 326100 361582 326336
rect 361026 290420 361262 290656
rect 361346 290420 361582 290656
rect 361026 290100 361262 290336
rect 361346 290100 361582 290336
rect 361026 254420 361262 254656
rect 361346 254420 361582 254656
rect 361026 254100 361262 254336
rect 361346 254100 361582 254336
rect 361026 218420 361262 218656
rect 361346 218420 361582 218656
rect 361026 218100 361262 218336
rect 361346 218100 361582 218336
rect 361026 182420 361262 182656
rect 361346 182420 361582 182656
rect 361026 182100 361262 182336
rect 361346 182100 361582 182336
rect 361026 146420 361262 146656
rect 361346 146420 361582 146656
rect 361026 146100 361262 146336
rect 361346 146100 361582 146336
rect 361026 110420 361262 110656
rect 361346 110420 361582 110656
rect 361026 110100 361262 110336
rect 361346 110100 361582 110336
rect 361026 74420 361262 74656
rect 361346 74420 361582 74656
rect 361026 74100 361262 74336
rect 361346 74100 361582 74336
rect 361026 38420 361262 38656
rect 361346 38420 361582 38656
rect 361026 38100 361262 38336
rect 361346 38100 361582 38336
rect 361026 2420 361262 2656
rect 361346 2420 361582 2656
rect 361026 2100 361262 2336
rect 361346 2100 361582 2336
rect 361026 -580 361262 -344
rect 361346 -580 361582 -344
rect 361026 -900 361262 -664
rect 361346 -900 361582 -664
rect 362266 705564 362502 705800
rect 362586 705564 362822 705800
rect 362266 705244 362502 705480
rect 362586 705244 362822 705480
rect 362266 687660 362502 687896
rect 362586 687660 362822 687896
rect 362266 687340 362502 687576
rect 362586 687340 362822 687576
rect 362266 651660 362502 651896
rect 362586 651660 362822 651896
rect 362266 651340 362502 651576
rect 362586 651340 362822 651576
rect 362266 615660 362502 615896
rect 362586 615660 362822 615896
rect 362266 615340 362502 615576
rect 362586 615340 362822 615576
rect 362266 579660 362502 579896
rect 362586 579660 362822 579896
rect 362266 579340 362502 579576
rect 362586 579340 362822 579576
rect 362266 543660 362502 543896
rect 362586 543660 362822 543896
rect 362266 543340 362502 543576
rect 362586 543340 362822 543576
rect 362266 507660 362502 507896
rect 362586 507660 362822 507896
rect 362266 507340 362502 507576
rect 362586 507340 362822 507576
rect 362266 471660 362502 471896
rect 362586 471660 362822 471896
rect 362266 471340 362502 471576
rect 362586 471340 362822 471576
rect 362266 435660 362502 435896
rect 362586 435660 362822 435896
rect 362266 435340 362502 435576
rect 362586 435340 362822 435576
rect 362266 399660 362502 399896
rect 362586 399660 362822 399896
rect 362266 399340 362502 399576
rect 362586 399340 362822 399576
rect 362266 363660 362502 363896
rect 362586 363660 362822 363896
rect 362266 363340 362502 363576
rect 362586 363340 362822 363576
rect 362266 327660 362502 327896
rect 362586 327660 362822 327896
rect 362266 327340 362502 327576
rect 362586 327340 362822 327576
rect 362266 291660 362502 291896
rect 362586 291660 362822 291896
rect 362266 291340 362502 291576
rect 362586 291340 362822 291576
rect 362266 255660 362502 255896
rect 362586 255660 362822 255896
rect 362266 255340 362502 255576
rect 362586 255340 362822 255576
rect 362266 219660 362502 219896
rect 362586 219660 362822 219896
rect 362266 219340 362502 219576
rect 362586 219340 362822 219576
rect 362266 183660 362502 183896
rect 362586 183660 362822 183896
rect 362266 183340 362502 183576
rect 362586 183340 362822 183576
rect 362266 147660 362502 147896
rect 362586 147660 362822 147896
rect 362266 147340 362502 147576
rect 362586 147340 362822 147576
rect 362266 111660 362502 111896
rect 362586 111660 362822 111896
rect 362266 111340 362502 111576
rect 362586 111340 362822 111576
rect 362266 75660 362502 75896
rect 362586 75660 362822 75896
rect 362266 75340 362502 75576
rect 362586 75340 362822 75576
rect 362266 39660 362502 39896
rect 362586 39660 362822 39896
rect 362266 39340 362502 39576
rect 362586 39340 362822 39576
rect 362266 3660 362502 3896
rect 362586 3660 362822 3896
rect 362266 3340 362502 3576
rect 362586 3340 362822 3576
rect 362266 -1540 362502 -1304
rect 362586 -1540 362822 -1304
rect 362266 -1860 362502 -1624
rect 362586 -1860 362822 -1624
rect 363506 706524 363742 706760
rect 363826 706524 364062 706760
rect 363506 706204 363742 706440
rect 363826 706204 364062 706440
rect 363506 688900 363742 689136
rect 363826 688900 364062 689136
rect 363506 688580 363742 688816
rect 363826 688580 364062 688816
rect 363506 652900 363742 653136
rect 363826 652900 364062 653136
rect 363506 652580 363742 652816
rect 363826 652580 364062 652816
rect 363506 616900 363742 617136
rect 363826 616900 364062 617136
rect 363506 616580 363742 616816
rect 363826 616580 364062 616816
rect 363506 580900 363742 581136
rect 363826 580900 364062 581136
rect 363506 580580 363742 580816
rect 363826 580580 364062 580816
rect 363506 544900 363742 545136
rect 363826 544900 364062 545136
rect 363506 544580 363742 544816
rect 363826 544580 364062 544816
rect 363506 508900 363742 509136
rect 363826 508900 364062 509136
rect 363506 508580 363742 508816
rect 363826 508580 364062 508816
rect 363506 472900 363742 473136
rect 363826 472900 364062 473136
rect 363506 472580 363742 472816
rect 363826 472580 364062 472816
rect 363506 436900 363742 437136
rect 363826 436900 364062 437136
rect 363506 436580 363742 436816
rect 363826 436580 364062 436816
rect 363506 400900 363742 401136
rect 363826 400900 364062 401136
rect 363506 400580 363742 400816
rect 363826 400580 364062 400816
rect 363506 364900 363742 365136
rect 363826 364900 364062 365136
rect 363506 364580 363742 364816
rect 363826 364580 364062 364816
rect 363506 328900 363742 329136
rect 363826 328900 364062 329136
rect 363506 328580 363742 328816
rect 363826 328580 364062 328816
rect 363506 292900 363742 293136
rect 363826 292900 364062 293136
rect 363506 292580 363742 292816
rect 363826 292580 364062 292816
rect 363506 256900 363742 257136
rect 363826 256900 364062 257136
rect 363506 256580 363742 256816
rect 363826 256580 364062 256816
rect 363506 220900 363742 221136
rect 363826 220900 364062 221136
rect 363506 220580 363742 220816
rect 363826 220580 364062 220816
rect 363506 184900 363742 185136
rect 363826 184900 364062 185136
rect 363506 184580 363742 184816
rect 363826 184580 364062 184816
rect 363506 148900 363742 149136
rect 363826 148900 364062 149136
rect 363506 148580 363742 148816
rect 363826 148580 364062 148816
rect 363506 112900 363742 113136
rect 363826 112900 364062 113136
rect 363506 112580 363742 112816
rect 363826 112580 364062 112816
rect 363506 76900 363742 77136
rect 363826 76900 364062 77136
rect 363506 76580 363742 76816
rect 363826 76580 364062 76816
rect 363506 40900 363742 41136
rect 363826 40900 364062 41136
rect 363506 40580 363742 40816
rect 363826 40580 364062 40816
rect 363506 4900 363742 5136
rect 363826 4900 364062 5136
rect 363506 4580 363742 4816
rect 363826 4580 364062 4816
rect 363506 -2500 363742 -2264
rect 363826 -2500 364062 -2264
rect 363506 -2820 363742 -2584
rect 363826 -2820 364062 -2584
rect 364746 707484 364982 707720
rect 365066 707484 365302 707720
rect 364746 707164 364982 707400
rect 365066 707164 365302 707400
rect 364746 690140 364982 690376
rect 365066 690140 365302 690376
rect 364746 689820 364982 690056
rect 365066 689820 365302 690056
rect 364746 654140 364982 654376
rect 365066 654140 365302 654376
rect 364746 653820 364982 654056
rect 365066 653820 365302 654056
rect 364746 618140 364982 618376
rect 365066 618140 365302 618376
rect 364746 617820 364982 618056
rect 365066 617820 365302 618056
rect 364746 582140 364982 582376
rect 365066 582140 365302 582376
rect 364746 581820 364982 582056
rect 365066 581820 365302 582056
rect 364746 546140 364982 546376
rect 365066 546140 365302 546376
rect 364746 545820 364982 546056
rect 365066 545820 365302 546056
rect 364746 510140 364982 510376
rect 365066 510140 365302 510376
rect 364746 509820 364982 510056
rect 365066 509820 365302 510056
rect 364746 474140 364982 474376
rect 365066 474140 365302 474376
rect 364746 473820 364982 474056
rect 365066 473820 365302 474056
rect 364746 438140 364982 438376
rect 365066 438140 365302 438376
rect 364746 437820 364982 438056
rect 365066 437820 365302 438056
rect 364746 402140 364982 402376
rect 365066 402140 365302 402376
rect 364746 401820 364982 402056
rect 365066 401820 365302 402056
rect 364746 366140 364982 366376
rect 365066 366140 365302 366376
rect 364746 365820 364982 366056
rect 365066 365820 365302 366056
rect 364746 330140 364982 330376
rect 365066 330140 365302 330376
rect 364746 329820 364982 330056
rect 365066 329820 365302 330056
rect 364746 294140 364982 294376
rect 365066 294140 365302 294376
rect 364746 293820 364982 294056
rect 365066 293820 365302 294056
rect 364746 258140 364982 258376
rect 365066 258140 365302 258376
rect 364746 257820 364982 258056
rect 365066 257820 365302 258056
rect 364746 222140 364982 222376
rect 365066 222140 365302 222376
rect 364746 221820 364982 222056
rect 365066 221820 365302 222056
rect 364746 186140 364982 186376
rect 365066 186140 365302 186376
rect 364746 185820 364982 186056
rect 365066 185820 365302 186056
rect 364746 150140 364982 150376
rect 365066 150140 365302 150376
rect 364746 149820 364982 150056
rect 365066 149820 365302 150056
rect 364746 114140 364982 114376
rect 365066 114140 365302 114376
rect 364746 113820 364982 114056
rect 365066 113820 365302 114056
rect 364746 78140 364982 78376
rect 365066 78140 365302 78376
rect 364746 77820 364982 78056
rect 365066 77820 365302 78056
rect 364746 42140 364982 42376
rect 365066 42140 365302 42376
rect 364746 41820 364982 42056
rect 365066 41820 365302 42056
rect 364746 6140 364982 6376
rect 365066 6140 365302 6376
rect 364746 5820 364982 6056
rect 365066 5820 365302 6056
rect 364746 -3460 364982 -3224
rect 365066 -3460 365302 -3224
rect 364746 -3780 364982 -3544
rect 365066 -3780 365302 -3544
rect 365986 708444 366222 708680
rect 366306 708444 366542 708680
rect 365986 708124 366222 708360
rect 366306 708124 366542 708360
rect 365986 691380 366222 691616
rect 366306 691380 366542 691616
rect 365986 691060 366222 691296
rect 366306 691060 366542 691296
rect 365986 655380 366222 655616
rect 366306 655380 366542 655616
rect 365986 655060 366222 655296
rect 366306 655060 366542 655296
rect 365986 619380 366222 619616
rect 366306 619380 366542 619616
rect 365986 619060 366222 619296
rect 366306 619060 366542 619296
rect 365986 583380 366222 583616
rect 366306 583380 366542 583616
rect 365986 583060 366222 583296
rect 366306 583060 366542 583296
rect 365986 547380 366222 547616
rect 366306 547380 366542 547616
rect 365986 547060 366222 547296
rect 366306 547060 366542 547296
rect 365986 511380 366222 511616
rect 366306 511380 366542 511616
rect 365986 511060 366222 511296
rect 366306 511060 366542 511296
rect 365986 475380 366222 475616
rect 366306 475380 366542 475616
rect 365986 475060 366222 475296
rect 366306 475060 366542 475296
rect 365986 439380 366222 439616
rect 366306 439380 366542 439616
rect 365986 439060 366222 439296
rect 366306 439060 366542 439296
rect 365986 403380 366222 403616
rect 366306 403380 366542 403616
rect 365986 403060 366222 403296
rect 366306 403060 366542 403296
rect 365986 367380 366222 367616
rect 366306 367380 366542 367616
rect 365986 367060 366222 367296
rect 366306 367060 366542 367296
rect 365986 331380 366222 331616
rect 366306 331380 366542 331616
rect 365986 331060 366222 331296
rect 366306 331060 366542 331296
rect 365986 295380 366222 295616
rect 366306 295380 366542 295616
rect 365986 295060 366222 295296
rect 366306 295060 366542 295296
rect 365986 259380 366222 259616
rect 366306 259380 366542 259616
rect 365986 259060 366222 259296
rect 366306 259060 366542 259296
rect 365986 223380 366222 223616
rect 366306 223380 366542 223616
rect 365986 223060 366222 223296
rect 366306 223060 366542 223296
rect 365986 187380 366222 187616
rect 366306 187380 366542 187616
rect 365986 187060 366222 187296
rect 366306 187060 366542 187296
rect 365986 151380 366222 151616
rect 366306 151380 366542 151616
rect 365986 151060 366222 151296
rect 366306 151060 366542 151296
rect 365986 115380 366222 115616
rect 366306 115380 366542 115616
rect 365986 115060 366222 115296
rect 366306 115060 366542 115296
rect 365986 79380 366222 79616
rect 366306 79380 366542 79616
rect 365986 79060 366222 79296
rect 366306 79060 366542 79296
rect 365986 43380 366222 43616
rect 366306 43380 366542 43616
rect 365986 43060 366222 43296
rect 366306 43060 366542 43296
rect 365986 7380 366222 7616
rect 366306 7380 366542 7616
rect 365986 7060 366222 7296
rect 366306 7060 366542 7296
rect 365986 -4420 366222 -4184
rect 366306 -4420 366542 -4184
rect 365986 -4740 366222 -4504
rect 366306 -4740 366542 -4504
rect 367226 709404 367462 709640
rect 367546 709404 367782 709640
rect 367226 709084 367462 709320
rect 367546 709084 367782 709320
rect 367226 692620 367462 692856
rect 367546 692620 367782 692856
rect 367226 692300 367462 692536
rect 367546 692300 367782 692536
rect 367226 656620 367462 656856
rect 367546 656620 367782 656856
rect 367226 656300 367462 656536
rect 367546 656300 367782 656536
rect 367226 620620 367462 620856
rect 367546 620620 367782 620856
rect 367226 620300 367462 620536
rect 367546 620300 367782 620536
rect 367226 584620 367462 584856
rect 367546 584620 367782 584856
rect 367226 584300 367462 584536
rect 367546 584300 367782 584536
rect 367226 548620 367462 548856
rect 367546 548620 367782 548856
rect 367226 548300 367462 548536
rect 367546 548300 367782 548536
rect 367226 512620 367462 512856
rect 367546 512620 367782 512856
rect 367226 512300 367462 512536
rect 367546 512300 367782 512536
rect 367226 476620 367462 476856
rect 367546 476620 367782 476856
rect 367226 476300 367462 476536
rect 367546 476300 367782 476536
rect 367226 440620 367462 440856
rect 367546 440620 367782 440856
rect 367226 440300 367462 440536
rect 367546 440300 367782 440536
rect 367226 404620 367462 404856
rect 367546 404620 367782 404856
rect 367226 404300 367462 404536
rect 367546 404300 367782 404536
rect 367226 368620 367462 368856
rect 367546 368620 367782 368856
rect 367226 368300 367462 368536
rect 367546 368300 367782 368536
rect 367226 332620 367462 332856
rect 367546 332620 367782 332856
rect 367226 332300 367462 332536
rect 367546 332300 367782 332536
rect 367226 296620 367462 296856
rect 367546 296620 367782 296856
rect 367226 296300 367462 296536
rect 367546 296300 367782 296536
rect 367226 260620 367462 260856
rect 367546 260620 367782 260856
rect 367226 260300 367462 260536
rect 367546 260300 367782 260536
rect 367226 224620 367462 224856
rect 367546 224620 367782 224856
rect 367226 224300 367462 224536
rect 367546 224300 367782 224536
rect 367226 188620 367462 188856
rect 367546 188620 367782 188856
rect 367226 188300 367462 188536
rect 367546 188300 367782 188536
rect 367226 152620 367462 152856
rect 367546 152620 367782 152856
rect 367226 152300 367462 152536
rect 367546 152300 367782 152536
rect 367226 116620 367462 116856
rect 367546 116620 367782 116856
rect 367226 116300 367462 116536
rect 367546 116300 367782 116536
rect 367226 80620 367462 80856
rect 367546 80620 367782 80856
rect 367226 80300 367462 80536
rect 367546 80300 367782 80536
rect 367226 44620 367462 44856
rect 367546 44620 367782 44856
rect 367226 44300 367462 44536
rect 367546 44300 367782 44536
rect 367226 8620 367462 8856
rect 367546 8620 367782 8856
rect 367226 8300 367462 8536
rect 367546 8300 367782 8536
rect 367226 -5380 367462 -5144
rect 367546 -5380 367782 -5144
rect 367226 -5700 367462 -5464
rect 367546 -5700 367782 -5464
rect 368466 710364 368702 710600
rect 368786 710364 369022 710600
rect 368466 710044 368702 710280
rect 368786 710044 369022 710280
rect 368466 693860 368702 694096
rect 368786 693860 369022 694096
rect 368466 693540 368702 693776
rect 368786 693540 369022 693776
rect 368466 657860 368702 658096
rect 368786 657860 369022 658096
rect 368466 657540 368702 657776
rect 368786 657540 369022 657776
rect 368466 621860 368702 622096
rect 368786 621860 369022 622096
rect 368466 621540 368702 621776
rect 368786 621540 369022 621776
rect 368466 585860 368702 586096
rect 368786 585860 369022 586096
rect 368466 585540 368702 585776
rect 368786 585540 369022 585776
rect 368466 549860 368702 550096
rect 368786 549860 369022 550096
rect 368466 549540 368702 549776
rect 368786 549540 369022 549776
rect 368466 513860 368702 514096
rect 368786 513860 369022 514096
rect 368466 513540 368702 513776
rect 368786 513540 369022 513776
rect 368466 477860 368702 478096
rect 368786 477860 369022 478096
rect 368466 477540 368702 477776
rect 368786 477540 369022 477776
rect 368466 441860 368702 442096
rect 368786 441860 369022 442096
rect 368466 441540 368702 441776
rect 368786 441540 369022 441776
rect 368466 405860 368702 406096
rect 368786 405860 369022 406096
rect 368466 405540 368702 405776
rect 368786 405540 369022 405776
rect 368466 369860 368702 370096
rect 368786 369860 369022 370096
rect 368466 369540 368702 369776
rect 368786 369540 369022 369776
rect 368466 333860 368702 334096
rect 368786 333860 369022 334096
rect 368466 333540 368702 333776
rect 368786 333540 369022 333776
rect 368466 297860 368702 298096
rect 368786 297860 369022 298096
rect 368466 297540 368702 297776
rect 368786 297540 369022 297776
rect 368466 261860 368702 262096
rect 368786 261860 369022 262096
rect 368466 261540 368702 261776
rect 368786 261540 369022 261776
rect 368466 225860 368702 226096
rect 368786 225860 369022 226096
rect 368466 225540 368702 225776
rect 368786 225540 369022 225776
rect 368466 189860 368702 190096
rect 368786 189860 369022 190096
rect 368466 189540 368702 189776
rect 368786 189540 369022 189776
rect 368466 153860 368702 154096
rect 368786 153860 369022 154096
rect 368466 153540 368702 153776
rect 368786 153540 369022 153776
rect 368466 117860 368702 118096
rect 368786 117860 369022 118096
rect 368466 117540 368702 117776
rect 368786 117540 369022 117776
rect 368466 81860 368702 82096
rect 368786 81860 369022 82096
rect 368466 81540 368702 81776
rect 368786 81540 369022 81776
rect 368466 45860 368702 46096
rect 368786 45860 369022 46096
rect 368466 45540 368702 45776
rect 368786 45540 369022 45776
rect 368466 9860 368702 10096
rect 368786 9860 369022 10096
rect 368466 9540 368702 9776
rect 368786 9540 369022 9776
rect 368466 -6340 368702 -6104
rect 368786 -6340 369022 -6104
rect 368466 -6660 368702 -6424
rect 368786 -6660 369022 -6424
rect 369706 711324 369942 711560
rect 370026 711324 370262 711560
rect 369706 711004 369942 711240
rect 370026 711004 370262 711240
rect 369706 695100 369942 695336
rect 370026 695100 370262 695336
rect 369706 694780 369942 695016
rect 370026 694780 370262 695016
rect 369706 659100 369942 659336
rect 370026 659100 370262 659336
rect 369706 658780 369942 659016
rect 370026 658780 370262 659016
rect 369706 623100 369942 623336
rect 370026 623100 370262 623336
rect 369706 622780 369942 623016
rect 370026 622780 370262 623016
rect 369706 587100 369942 587336
rect 370026 587100 370262 587336
rect 369706 586780 369942 587016
rect 370026 586780 370262 587016
rect 369706 551100 369942 551336
rect 370026 551100 370262 551336
rect 369706 550780 369942 551016
rect 370026 550780 370262 551016
rect 369706 515100 369942 515336
rect 370026 515100 370262 515336
rect 369706 514780 369942 515016
rect 370026 514780 370262 515016
rect 369706 479100 369942 479336
rect 370026 479100 370262 479336
rect 369706 478780 369942 479016
rect 370026 478780 370262 479016
rect 369706 443100 369942 443336
rect 370026 443100 370262 443336
rect 369706 442780 369942 443016
rect 370026 442780 370262 443016
rect 369706 407100 369942 407336
rect 370026 407100 370262 407336
rect 369706 406780 369942 407016
rect 370026 406780 370262 407016
rect 369706 371100 369942 371336
rect 370026 371100 370262 371336
rect 369706 370780 369942 371016
rect 370026 370780 370262 371016
rect 369706 335100 369942 335336
rect 370026 335100 370262 335336
rect 369706 334780 369942 335016
rect 370026 334780 370262 335016
rect 369706 299100 369942 299336
rect 370026 299100 370262 299336
rect 369706 298780 369942 299016
rect 370026 298780 370262 299016
rect 369706 263100 369942 263336
rect 370026 263100 370262 263336
rect 369706 262780 369942 263016
rect 370026 262780 370262 263016
rect 369706 227100 369942 227336
rect 370026 227100 370262 227336
rect 369706 226780 369942 227016
rect 370026 226780 370262 227016
rect 369706 191100 369942 191336
rect 370026 191100 370262 191336
rect 369706 190780 369942 191016
rect 370026 190780 370262 191016
rect 369706 155100 369942 155336
rect 370026 155100 370262 155336
rect 369706 154780 369942 155016
rect 370026 154780 370262 155016
rect 369706 119100 369942 119336
rect 370026 119100 370262 119336
rect 369706 118780 369942 119016
rect 370026 118780 370262 119016
rect 369706 83100 369942 83336
rect 370026 83100 370262 83336
rect 369706 82780 369942 83016
rect 370026 82780 370262 83016
rect 369706 47100 369942 47336
rect 370026 47100 370262 47336
rect 369706 46780 369942 47016
rect 370026 46780 370262 47016
rect 369706 11100 369942 11336
rect 370026 11100 370262 11336
rect 369706 10780 369942 11016
rect 370026 10780 370262 11016
rect 369706 -7300 369942 -7064
rect 370026 -7300 370262 -7064
rect 369706 -7620 369942 -7384
rect 370026 -7620 370262 -7384
rect 397026 704604 397262 704840
rect 397346 704604 397582 704840
rect 397026 704284 397262 704520
rect 397346 704284 397582 704520
rect 397026 686420 397262 686656
rect 397346 686420 397582 686656
rect 397026 686100 397262 686336
rect 397346 686100 397582 686336
rect 397026 650420 397262 650656
rect 397346 650420 397582 650656
rect 397026 650100 397262 650336
rect 397346 650100 397582 650336
rect 397026 614420 397262 614656
rect 397346 614420 397582 614656
rect 397026 614100 397262 614336
rect 397346 614100 397582 614336
rect 397026 578420 397262 578656
rect 397346 578420 397582 578656
rect 397026 578100 397262 578336
rect 397346 578100 397582 578336
rect 397026 542420 397262 542656
rect 397346 542420 397582 542656
rect 397026 542100 397262 542336
rect 397346 542100 397582 542336
rect 397026 506420 397262 506656
rect 397346 506420 397582 506656
rect 397026 506100 397262 506336
rect 397346 506100 397582 506336
rect 397026 470420 397262 470656
rect 397346 470420 397582 470656
rect 397026 470100 397262 470336
rect 397346 470100 397582 470336
rect 397026 434420 397262 434656
rect 397346 434420 397582 434656
rect 397026 434100 397262 434336
rect 397346 434100 397582 434336
rect 397026 398420 397262 398656
rect 397346 398420 397582 398656
rect 397026 398100 397262 398336
rect 397346 398100 397582 398336
rect 397026 362420 397262 362656
rect 397346 362420 397582 362656
rect 397026 362100 397262 362336
rect 397346 362100 397582 362336
rect 397026 326420 397262 326656
rect 397346 326420 397582 326656
rect 397026 326100 397262 326336
rect 397346 326100 397582 326336
rect 397026 290420 397262 290656
rect 397346 290420 397582 290656
rect 397026 290100 397262 290336
rect 397346 290100 397582 290336
rect 397026 254420 397262 254656
rect 397346 254420 397582 254656
rect 397026 254100 397262 254336
rect 397346 254100 397582 254336
rect 397026 218420 397262 218656
rect 397346 218420 397582 218656
rect 397026 218100 397262 218336
rect 397346 218100 397582 218336
rect 397026 182420 397262 182656
rect 397346 182420 397582 182656
rect 397026 182100 397262 182336
rect 397346 182100 397582 182336
rect 397026 146420 397262 146656
rect 397346 146420 397582 146656
rect 397026 146100 397262 146336
rect 397346 146100 397582 146336
rect 397026 110420 397262 110656
rect 397346 110420 397582 110656
rect 397026 110100 397262 110336
rect 397346 110100 397582 110336
rect 397026 74420 397262 74656
rect 397346 74420 397582 74656
rect 397026 74100 397262 74336
rect 397346 74100 397582 74336
rect 397026 38420 397262 38656
rect 397346 38420 397582 38656
rect 397026 38100 397262 38336
rect 397346 38100 397582 38336
rect 397026 2420 397262 2656
rect 397346 2420 397582 2656
rect 397026 2100 397262 2336
rect 397346 2100 397582 2336
rect 397026 -580 397262 -344
rect 397346 -580 397582 -344
rect 397026 -900 397262 -664
rect 397346 -900 397582 -664
rect 398266 705564 398502 705800
rect 398586 705564 398822 705800
rect 398266 705244 398502 705480
rect 398586 705244 398822 705480
rect 398266 687660 398502 687896
rect 398586 687660 398822 687896
rect 398266 687340 398502 687576
rect 398586 687340 398822 687576
rect 398266 651660 398502 651896
rect 398586 651660 398822 651896
rect 398266 651340 398502 651576
rect 398586 651340 398822 651576
rect 398266 615660 398502 615896
rect 398586 615660 398822 615896
rect 398266 615340 398502 615576
rect 398586 615340 398822 615576
rect 398266 579660 398502 579896
rect 398586 579660 398822 579896
rect 398266 579340 398502 579576
rect 398586 579340 398822 579576
rect 398266 543660 398502 543896
rect 398586 543660 398822 543896
rect 398266 543340 398502 543576
rect 398586 543340 398822 543576
rect 398266 507660 398502 507896
rect 398586 507660 398822 507896
rect 398266 507340 398502 507576
rect 398586 507340 398822 507576
rect 398266 471660 398502 471896
rect 398586 471660 398822 471896
rect 398266 471340 398502 471576
rect 398586 471340 398822 471576
rect 398266 435660 398502 435896
rect 398586 435660 398822 435896
rect 398266 435340 398502 435576
rect 398586 435340 398822 435576
rect 398266 399660 398502 399896
rect 398586 399660 398822 399896
rect 398266 399340 398502 399576
rect 398586 399340 398822 399576
rect 398266 363660 398502 363896
rect 398586 363660 398822 363896
rect 398266 363340 398502 363576
rect 398586 363340 398822 363576
rect 398266 327660 398502 327896
rect 398586 327660 398822 327896
rect 398266 327340 398502 327576
rect 398586 327340 398822 327576
rect 398266 291660 398502 291896
rect 398586 291660 398822 291896
rect 398266 291340 398502 291576
rect 398586 291340 398822 291576
rect 398266 255660 398502 255896
rect 398586 255660 398822 255896
rect 398266 255340 398502 255576
rect 398586 255340 398822 255576
rect 398266 219660 398502 219896
rect 398586 219660 398822 219896
rect 398266 219340 398502 219576
rect 398586 219340 398822 219576
rect 398266 183660 398502 183896
rect 398586 183660 398822 183896
rect 398266 183340 398502 183576
rect 398586 183340 398822 183576
rect 398266 147660 398502 147896
rect 398586 147660 398822 147896
rect 398266 147340 398502 147576
rect 398586 147340 398822 147576
rect 398266 111660 398502 111896
rect 398586 111660 398822 111896
rect 398266 111340 398502 111576
rect 398586 111340 398822 111576
rect 398266 75660 398502 75896
rect 398586 75660 398822 75896
rect 398266 75340 398502 75576
rect 398586 75340 398822 75576
rect 398266 39660 398502 39896
rect 398586 39660 398822 39896
rect 398266 39340 398502 39576
rect 398586 39340 398822 39576
rect 398266 3660 398502 3896
rect 398586 3660 398822 3896
rect 398266 3340 398502 3576
rect 398586 3340 398822 3576
rect 398266 -1540 398502 -1304
rect 398586 -1540 398822 -1304
rect 398266 -1860 398502 -1624
rect 398586 -1860 398822 -1624
rect 399506 706524 399742 706760
rect 399826 706524 400062 706760
rect 399506 706204 399742 706440
rect 399826 706204 400062 706440
rect 399506 688900 399742 689136
rect 399826 688900 400062 689136
rect 399506 688580 399742 688816
rect 399826 688580 400062 688816
rect 399506 652900 399742 653136
rect 399826 652900 400062 653136
rect 399506 652580 399742 652816
rect 399826 652580 400062 652816
rect 399506 616900 399742 617136
rect 399826 616900 400062 617136
rect 399506 616580 399742 616816
rect 399826 616580 400062 616816
rect 399506 580900 399742 581136
rect 399826 580900 400062 581136
rect 399506 580580 399742 580816
rect 399826 580580 400062 580816
rect 399506 544900 399742 545136
rect 399826 544900 400062 545136
rect 399506 544580 399742 544816
rect 399826 544580 400062 544816
rect 399506 508900 399742 509136
rect 399826 508900 400062 509136
rect 399506 508580 399742 508816
rect 399826 508580 400062 508816
rect 399506 472900 399742 473136
rect 399826 472900 400062 473136
rect 399506 472580 399742 472816
rect 399826 472580 400062 472816
rect 399506 436900 399742 437136
rect 399826 436900 400062 437136
rect 399506 436580 399742 436816
rect 399826 436580 400062 436816
rect 399506 400900 399742 401136
rect 399826 400900 400062 401136
rect 399506 400580 399742 400816
rect 399826 400580 400062 400816
rect 399506 364900 399742 365136
rect 399826 364900 400062 365136
rect 399506 364580 399742 364816
rect 399826 364580 400062 364816
rect 399506 328900 399742 329136
rect 399826 328900 400062 329136
rect 399506 328580 399742 328816
rect 399826 328580 400062 328816
rect 399506 292900 399742 293136
rect 399826 292900 400062 293136
rect 399506 292580 399742 292816
rect 399826 292580 400062 292816
rect 399506 256900 399742 257136
rect 399826 256900 400062 257136
rect 399506 256580 399742 256816
rect 399826 256580 400062 256816
rect 399506 220900 399742 221136
rect 399826 220900 400062 221136
rect 399506 220580 399742 220816
rect 399826 220580 400062 220816
rect 399506 184900 399742 185136
rect 399826 184900 400062 185136
rect 399506 184580 399742 184816
rect 399826 184580 400062 184816
rect 399506 148900 399742 149136
rect 399826 148900 400062 149136
rect 399506 148580 399742 148816
rect 399826 148580 400062 148816
rect 399506 112900 399742 113136
rect 399826 112900 400062 113136
rect 399506 112580 399742 112816
rect 399826 112580 400062 112816
rect 399506 76900 399742 77136
rect 399826 76900 400062 77136
rect 399506 76580 399742 76816
rect 399826 76580 400062 76816
rect 399506 40900 399742 41136
rect 399826 40900 400062 41136
rect 399506 40580 399742 40816
rect 399826 40580 400062 40816
rect 399506 4900 399742 5136
rect 399826 4900 400062 5136
rect 399506 4580 399742 4816
rect 399826 4580 400062 4816
rect 399506 -2500 399742 -2264
rect 399826 -2500 400062 -2264
rect 399506 -2820 399742 -2584
rect 399826 -2820 400062 -2584
rect 400746 707484 400982 707720
rect 401066 707484 401302 707720
rect 400746 707164 400982 707400
rect 401066 707164 401302 707400
rect 400746 690140 400982 690376
rect 401066 690140 401302 690376
rect 400746 689820 400982 690056
rect 401066 689820 401302 690056
rect 400746 654140 400982 654376
rect 401066 654140 401302 654376
rect 400746 653820 400982 654056
rect 401066 653820 401302 654056
rect 400746 618140 400982 618376
rect 401066 618140 401302 618376
rect 400746 617820 400982 618056
rect 401066 617820 401302 618056
rect 400746 582140 400982 582376
rect 401066 582140 401302 582376
rect 400746 581820 400982 582056
rect 401066 581820 401302 582056
rect 400746 546140 400982 546376
rect 401066 546140 401302 546376
rect 400746 545820 400982 546056
rect 401066 545820 401302 546056
rect 400746 510140 400982 510376
rect 401066 510140 401302 510376
rect 400746 509820 400982 510056
rect 401066 509820 401302 510056
rect 400746 474140 400982 474376
rect 401066 474140 401302 474376
rect 400746 473820 400982 474056
rect 401066 473820 401302 474056
rect 400746 438140 400982 438376
rect 401066 438140 401302 438376
rect 400746 437820 400982 438056
rect 401066 437820 401302 438056
rect 400746 402140 400982 402376
rect 401066 402140 401302 402376
rect 400746 401820 400982 402056
rect 401066 401820 401302 402056
rect 400746 366140 400982 366376
rect 401066 366140 401302 366376
rect 400746 365820 400982 366056
rect 401066 365820 401302 366056
rect 400746 330140 400982 330376
rect 401066 330140 401302 330376
rect 400746 329820 400982 330056
rect 401066 329820 401302 330056
rect 400746 294140 400982 294376
rect 401066 294140 401302 294376
rect 400746 293820 400982 294056
rect 401066 293820 401302 294056
rect 400746 258140 400982 258376
rect 401066 258140 401302 258376
rect 400746 257820 400982 258056
rect 401066 257820 401302 258056
rect 400746 222140 400982 222376
rect 401066 222140 401302 222376
rect 400746 221820 400982 222056
rect 401066 221820 401302 222056
rect 400746 186140 400982 186376
rect 401066 186140 401302 186376
rect 400746 185820 400982 186056
rect 401066 185820 401302 186056
rect 400746 150140 400982 150376
rect 401066 150140 401302 150376
rect 400746 149820 400982 150056
rect 401066 149820 401302 150056
rect 400746 114140 400982 114376
rect 401066 114140 401302 114376
rect 400746 113820 400982 114056
rect 401066 113820 401302 114056
rect 400746 78140 400982 78376
rect 401066 78140 401302 78376
rect 400746 77820 400982 78056
rect 401066 77820 401302 78056
rect 400746 42140 400982 42376
rect 401066 42140 401302 42376
rect 400746 41820 400982 42056
rect 401066 41820 401302 42056
rect 400746 6140 400982 6376
rect 401066 6140 401302 6376
rect 400746 5820 400982 6056
rect 401066 5820 401302 6056
rect 400746 -3460 400982 -3224
rect 401066 -3460 401302 -3224
rect 400746 -3780 400982 -3544
rect 401066 -3780 401302 -3544
rect 401986 708444 402222 708680
rect 402306 708444 402542 708680
rect 401986 708124 402222 708360
rect 402306 708124 402542 708360
rect 401986 691380 402222 691616
rect 402306 691380 402542 691616
rect 401986 691060 402222 691296
rect 402306 691060 402542 691296
rect 401986 655380 402222 655616
rect 402306 655380 402542 655616
rect 401986 655060 402222 655296
rect 402306 655060 402542 655296
rect 401986 619380 402222 619616
rect 402306 619380 402542 619616
rect 401986 619060 402222 619296
rect 402306 619060 402542 619296
rect 401986 583380 402222 583616
rect 402306 583380 402542 583616
rect 401986 583060 402222 583296
rect 402306 583060 402542 583296
rect 401986 547380 402222 547616
rect 402306 547380 402542 547616
rect 401986 547060 402222 547296
rect 402306 547060 402542 547296
rect 401986 511380 402222 511616
rect 402306 511380 402542 511616
rect 401986 511060 402222 511296
rect 402306 511060 402542 511296
rect 401986 475380 402222 475616
rect 402306 475380 402542 475616
rect 401986 475060 402222 475296
rect 402306 475060 402542 475296
rect 401986 439380 402222 439616
rect 402306 439380 402542 439616
rect 401986 439060 402222 439296
rect 402306 439060 402542 439296
rect 401986 403380 402222 403616
rect 402306 403380 402542 403616
rect 401986 403060 402222 403296
rect 402306 403060 402542 403296
rect 401986 367380 402222 367616
rect 402306 367380 402542 367616
rect 401986 367060 402222 367296
rect 402306 367060 402542 367296
rect 401986 331380 402222 331616
rect 402306 331380 402542 331616
rect 401986 331060 402222 331296
rect 402306 331060 402542 331296
rect 401986 295380 402222 295616
rect 402306 295380 402542 295616
rect 401986 295060 402222 295296
rect 402306 295060 402542 295296
rect 401986 259380 402222 259616
rect 402306 259380 402542 259616
rect 401986 259060 402222 259296
rect 402306 259060 402542 259296
rect 401986 223380 402222 223616
rect 402306 223380 402542 223616
rect 401986 223060 402222 223296
rect 402306 223060 402542 223296
rect 401986 187380 402222 187616
rect 402306 187380 402542 187616
rect 401986 187060 402222 187296
rect 402306 187060 402542 187296
rect 401986 151380 402222 151616
rect 402306 151380 402542 151616
rect 401986 151060 402222 151296
rect 402306 151060 402542 151296
rect 401986 115380 402222 115616
rect 402306 115380 402542 115616
rect 401986 115060 402222 115296
rect 402306 115060 402542 115296
rect 401986 79380 402222 79616
rect 402306 79380 402542 79616
rect 401986 79060 402222 79296
rect 402306 79060 402542 79296
rect 401986 43380 402222 43616
rect 402306 43380 402542 43616
rect 401986 43060 402222 43296
rect 402306 43060 402542 43296
rect 401986 7380 402222 7616
rect 402306 7380 402542 7616
rect 401986 7060 402222 7296
rect 402306 7060 402542 7296
rect 401986 -4420 402222 -4184
rect 402306 -4420 402542 -4184
rect 401986 -4740 402222 -4504
rect 402306 -4740 402542 -4504
rect 403226 709404 403462 709640
rect 403546 709404 403782 709640
rect 403226 709084 403462 709320
rect 403546 709084 403782 709320
rect 403226 692620 403462 692856
rect 403546 692620 403782 692856
rect 403226 692300 403462 692536
rect 403546 692300 403782 692536
rect 403226 656620 403462 656856
rect 403546 656620 403782 656856
rect 403226 656300 403462 656536
rect 403546 656300 403782 656536
rect 403226 620620 403462 620856
rect 403546 620620 403782 620856
rect 403226 620300 403462 620536
rect 403546 620300 403782 620536
rect 403226 584620 403462 584856
rect 403546 584620 403782 584856
rect 403226 584300 403462 584536
rect 403546 584300 403782 584536
rect 403226 548620 403462 548856
rect 403546 548620 403782 548856
rect 403226 548300 403462 548536
rect 403546 548300 403782 548536
rect 403226 512620 403462 512856
rect 403546 512620 403782 512856
rect 403226 512300 403462 512536
rect 403546 512300 403782 512536
rect 403226 476620 403462 476856
rect 403546 476620 403782 476856
rect 403226 476300 403462 476536
rect 403546 476300 403782 476536
rect 403226 440620 403462 440856
rect 403546 440620 403782 440856
rect 403226 440300 403462 440536
rect 403546 440300 403782 440536
rect 403226 404620 403462 404856
rect 403546 404620 403782 404856
rect 403226 404300 403462 404536
rect 403546 404300 403782 404536
rect 403226 368620 403462 368856
rect 403546 368620 403782 368856
rect 403226 368300 403462 368536
rect 403546 368300 403782 368536
rect 403226 332620 403462 332856
rect 403546 332620 403782 332856
rect 403226 332300 403462 332536
rect 403546 332300 403782 332536
rect 403226 296620 403462 296856
rect 403546 296620 403782 296856
rect 403226 296300 403462 296536
rect 403546 296300 403782 296536
rect 403226 260620 403462 260856
rect 403546 260620 403782 260856
rect 403226 260300 403462 260536
rect 403546 260300 403782 260536
rect 403226 224620 403462 224856
rect 403546 224620 403782 224856
rect 403226 224300 403462 224536
rect 403546 224300 403782 224536
rect 403226 188620 403462 188856
rect 403546 188620 403782 188856
rect 403226 188300 403462 188536
rect 403546 188300 403782 188536
rect 403226 152620 403462 152856
rect 403546 152620 403782 152856
rect 403226 152300 403462 152536
rect 403546 152300 403782 152536
rect 403226 116620 403462 116856
rect 403546 116620 403782 116856
rect 403226 116300 403462 116536
rect 403546 116300 403782 116536
rect 403226 80620 403462 80856
rect 403546 80620 403782 80856
rect 403226 80300 403462 80536
rect 403546 80300 403782 80536
rect 403226 44620 403462 44856
rect 403546 44620 403782 44856
rect 403226 44300 403462 44536
rect 403546 44300 403782 44536
rect 403226 8620 403462 8856
rect 403546 8620 403782 8856
rect 403226 8300 403462 8536
rect 403546 8300 403782 8536
rect 403226 -5380 403462 -5144
rect 403546 -5380 403782 -5144
rect 403226 -5700 403462 -5464
rect 403546 -5700 403782 -5464
rect 404466 710364 404702 710600
rect 404786 710364 405022 710600
rect 404466 710044 404702 710280
rect 404786 710044 405022 710280
rect 404466 693860 404702 694096
rect 404786 693860 405022 694096
rect 404466 693540 404702 693776
rect 404786 693540 405022 693776
rect 404466 657860 404702 658096
rect 404786 657860 405022 658096
rect 404466 657540 404702 657776
rect 404786 657540 405022 657776
rect 404466 621860 404702 622096
rect 404786 621860 405022 622096
rect 404466 621540 404702 621776
rect 404786 621540 405022 621776
rect 404466 585860 404702 586096
rect 404786 585860 405022 586096
rect 404466 585540 404702 585776
rect 404786 585540 405022 585776
rect 404466 549860 404702 550096
rect 404786 549860 405022 550096
rect 404466 549540 404702 549776
rect 404786 549540 405022 549776
rect 404466 513860 404702 514096
rect 404786 513860 405022 514096
rect 404466 513540 404702 513776
rect 404786 513540 405022 513776
rect 404466 477860 404702 478096
rect 404786 477860 405022 478096
rect 404466 477540 404702 477776
rect 404786 477540 405022 477776
rect 404466 441860 404702 442096
rect 404786 441860 405022 442096
rect 404466 441540 404702 441776
rect 404786 441540 405022 441776
rect 404466 405860 404702 406096
rect 404786 405860 405022 406096
rect 404466 405540 404702 405776
rect 404786 405540 405022 405776
rect 404466 369860 404702 370096
rect 404786 369860 405022 370096
rect 404466 369540 404702 369776
rect 404786 369540 405022 369776
rect 404466 333860 404702 334096
rect 404786 333860 405022 334096
rect 404466 333540 404702 333776
rect 404786 333540 405022 333776
rect 404466 297860 404702 298096
rect 404786 297860 405022 298096
rect 404466 297540 404702 297776
rect 404786 297540 405022 297776
rect 404466 261860 404702 262096
rect 404786 261860 405022 262096
rect 404466 261540 404702 261776
rect 404786 261540 405022 261776
rect 404466 225860 404702 226096
rect 404786 225860 405022 226096
rect 404466 225540 404702 225776
rect 404786 225540 405022 225776
rect 404466 189860 404702 190096
rect 404786 189860 405022 190096
rect 404466 189540 404702 189776
rect 404786 189540 405022 189776
rect 404466 153860 404702 154096
rect 404786 153860 405022 154096
rect 404466 153540 404702 153776
rect 404786 153540 405022 153776
rect 404466 117860 404702 118096
rect 404786 117860 405022 118096
rect 404466 117540 404702 117776
rect 404786 117540 405022 117776
rect 404466 81860 404702 82096
rect 404786 81860 405022 82096
rect 404466 81540 404702 81776
rect 404786 81540 405022 81776
rect 404466 45860 404702 46096
rect 404786 45860 405022 46096
rect 404466 45540 404702 45776
rect 404786 45540 405022 45776
rect 404466 9860 404702 10096
rect 404786 9860 405022 10096
rect 404466 9540 404702 9776
rect 404786 9540 405022 9776
rect 404466 -6340 404702 -6104
rect 404786 -6340 405022 -6104
rect 404466 -6660 404702 -6424
rect 404786 -6660 405022 -6424
rect 405706 711324 405942 711560
rect 406026 711324 406262 711560
rect 405706 711004 405942 711240
rect 406026 711004 406262 711240
rect 405706 695100 405942 695336
rect 406026 695100 406262 695336
rect 405706 694780 405942 695016
rect 406026 694780 406262 695016
rect 405706 659100 405942 659336
rect 406026 659100 406262 659336
rect 405706 658780 405942 659016
rect 406026 658780 406262 659016
rect 405706 623100 405942 623336
rect 406026 623100 406262 623336
rect 405706 622780 405942 623016
rect 406026 622780 406262 623016
rect 405706 587100 405942 587336
rect 406026 587100 406262 587336
rect 405706 586780 405942 587016
rect 406026 586780 406262 587016
rect 405706 551100 405942 551336
rect 406026 551100 406262 551336
rect 405706 550780 405942 551016
rect 406026 550780 406262 551016
rect 405706 515100 405942 515336
rect 406026 515100 406262 515336
rect 405706 514780 405942 515016
rect 406026 514780 406262 515016
rect 405706 479100 405942 479336
rect 406026 479100 406262 479336
rect 405706 478780 405942 479016
rect 406026 478780 406262 479016
rect 405706 443100 405942 443336
rect 406026 443100 406262 443336
rect 405706 442780 405942 443016
rect 406026 442780 406262 443016
rect 405706 407100 405942 407336
rect 406026 407100 406262 407336
rect 405706 406780 405942 407016
rect 406026 406780 406262 407016
rect 405706 371100 405942 371336
rect 406026 371100 406262 371336
rect 405706 370780 405942 371016
rect 406026 370780 406262 371016
rect 405706 335100 405942 335336
rect 406026 335100 406262 335336
rect 405706 334780 405942 335016
rect 406026 334780 406262 335016
rect 405706 299100 405942 299336
rect 406026 299100 406262 299336
rect 405706 298780 405942 299016
rect 406026 298780 406262 299016
rect 405706 263100 405942 263336
rect 406026 263100 406262 263336
rect 405706 262780 405942 263016
rect 406026 262780 406262 263016
rect 405706 227100 405942 227336
rect 406026 227100 406262 227336
rect 405706 226780 405942 227016
rect 406026 226780 406262 227016
rect 405706 191100 405942 191336
rect 406026 191100 406262 191336
rect 405706 190780 405942 191016
rect 406026 190780 406262 191016
rect 405706 155100 405942 155336
rect 406026 155100 406262 155336
rect 405706 154780 405942 155016
rect 406026 154780 406262 155016
rect 405706 119100 405942 119336
rect 406026 119100 406262 119336
rect 405706 118780 405942 119016
rect 406026 118780 406262 119016
rect 405706 83100 405942 83336
rect 406026 83100 406262 83336
rect 405706 82780 405942 83016
rect 406026 82780 406262 83016
rect 405706 47100 405942 47336
rect 406026 47100 406262 47336
rect 405706 46780 405942 47016
rect 406026 46780 406262 47016
rect 405706 11100 405942 11336
rect 406026 11100 406262 11336
rect 405706 10780 405942 11016
rect 406026 10780 406262 11016
rect 405706 -7300 405942 -7064
rect 406026 -7300 406262 -7064
rect 405706 -7620 405942 -7384
rect 406026 -7620 406262 -7384
rect 433026 704604 433262 704840
rect 433346 704604 433582 704840
rect 433026 704284 433262 704520
rect 433346 704284 433582 704520
rect 433026 686420 433262 686656
rect 433346 686420 433582 686656
rect 433026 686100 433262 686336
rect 433346 686100 433582 686336
rect 433026 650420 433262 650656
rect 433346 650420 433582 650656
rect 433026 650100 433262 650336
rect 433346 650100 433582 650336
rect 433026 614420 433262 614656
rect 433346 614420 433582 614656
rect 433026 614100 433262 614336
rect 433346 614100 433582 614336
rect 433026 578420 433262 578656
rect 433346 578420 433582 578656
rect 433026 578100 433262 578336
rect 433346 578100 433582 578336
rect 433026 542420 433262 542656
rect 433346 542420 433582 542656
rect 433026 542100 433262 542336
rect 433346 542100 433582 542336
rect 433026 506420 433262 506656
rect 433346 506420 433582 506656
rect 433026 506100 433262 506336
rect 433346 506100 433582 506336
rect 433026 470420 433262 470656
rect 433346 470420 433582 470656
rect 433026 470100 433262 470336
rect 433346 470100 433582 470336
rect 433026 434420 433262 434656
rect 433346 434420 433582 434656
rect 433026 434100 433262 434336
rect 433346 434100 433582 434336
rect 433026 398420 433262 398656
rect 433346 398420 433582 398656
rect 433026 398100 433262 398336
rect 433346 398100 433582 398336
rect 433026 362420 433262 362656
rect 433346 362420 433582 362656
rect 433026 362100 433262 362336
rect 433346 362100 433582 362336
rect 433026 326420 433262 326656
rect 433346 326420 433582 326656
rect 433026 326100 433262 326336
rect 433346 326100 433582 326336
rect 433026 290420 433262 290656
rect 433346 290420 433582 290656
rect 433026 290100 433262 290336
rect 433346 290100 433582 290336
rect 433026 254420 433262 254656
rect 433346 254420 433582 254656
rect 433026 254100 433262 254336
rect 433346 254100 433582 254336
rect 433026 218420 433262 218656
rect 433346 218420 433582 218656
rect 433026 218100 433262 218336
rect 433346 218100 433582 218336
rect 433026 182420 433262 182656
rect 433346 182420 433582 182656
rect 433026 182100 433262 182336
rect 433346 182100 433582 182336
rect 433026 146420 433262 146656
rect 433346 146420 433582 146656
rect 433026 146100 433262 146336
rect 433346 146100 433582 146336
rect 433026 110420 433262 110656
rect 433346 110420 433582 110656
rect 433026 110100 433262 110336
rect 433346 110100 433582 110336
rect 433026 74420 433262 74656
rect 433346 74420 433582 74656
rect 433026 74100 433262 74336
rect 433346 74100 433582 74336
rect 433026 38420 433262 38656
rect 433346 38420 433582 38656
rect 433026 38100 433262 38336
rect 433346 38100 433582 38336
rect 433026 2420 433262 2656
rect 433346 2420 433582 2656
rect 433026 2100 433262 2336
rect 433346 2100 433582 2336
rect 433026 -580 433262 -344
rect 433346 -580 433582 -344
rect 433026 -900 433262 -664
rect 433346 -900 433582 -664
rect 434266 705564 434502 705800
rect 434586 705564 434822 705800
rect 434266 705244 434502 705480
rect 434586 705244 434822 705480
rect 434266 687660 434502 687896
rect 434586 687660 434822 687896
rect 434266 687340 434502 687576
rect 434586 687340 434822 687576
rect 434266 651660 434502 651896
rect 434586 651660 434822 651896
rect 434266 651340 434502 651576
rect 434586 651340 434822 651576
rect 434266 615660 434502 615896
rect 434586 615660 434822 615896
rect 434266 615340 434502 615576
rect 434586 615340 434822 615576
rect 434266 579660 434502 579896
rect 434586 579660 434822 579896
rect 434266 579340 434502 579576
rect 434586 579340 434822 579576
rect 434266 543660 434502 543896
rect 434586 543660 434822 543896
rect 434266 543340 434502 543576
rect 434586 543340 434822 543576
rect 434266 507660 434502 507896
rect 434586 507660 434822 507896
rect 434266 507340 434502 507576
rect 434586 507340 434822 507576
rect 434266 471660 434502 471896
rect 434586 471660 434822 471896
rect 434266 471340 434502 471576
rect 434586 471340 434822 471576
rect 434266 435660 434502 435896
rect 434586 435660 434822 435896
rect 434266 435340 434502 435576
rect 434586 435340 434822 435576
rect 434266 399660 434502 399896
rect 434586 399660 434822 399896
rect 434266 399340 434502 399576
rect 434586 399340 434822 399576
rect 434266 363660 434502 363896
rect 434586 363660 434822 363896
rect 434266 363340 434502 363576
rect 434586 363340 434822 363576
rect 434266 327660 434502 327896
rect 434586 327660 434822 327896
rect 434266 327340 434502 327576
rect 434586 327340 434822 327576
rect 434266 291660 434502 291896
rect 434586 291660 434822 291896
rect 434266 291340 434502 291576
rect 434586 291340 434822 291576
rect 434266 255660 434502 255896
rect 434586 255660 434822 255896
rect 434266 255340 434502 255576
rect 434586 255340 434822 255576
rect 434266 219660 434502 219896
rect 434586 219660 434822 219896
rect 434266 219340 434502 219576
rect 434586 219340 434822 219576
rect 434266 183660 434502 183896
rect 434586 183660 434822 183896
rect 434266 183340 434502 183576
rect 434586 183340 434822 183576
rect 434266 147660 434502 147896
rect 434586 147660 434822 147896
rect 434266 147340 434502 147576
rect 434586 147340 434822 147576
rect 434266 111660 434502 111896
rect 434586 111660 434822 111896
rect 434266 111340 434502 111576
rect 434586 111340 434822 111576
rect 434266 75660 434502 75896
rect 434586 75660 434822 75896
rect 434266 75340 434502 75576
rect 434586 75340 434822 75576
rect 434266 39660 434502 39896
rect 434586 39660 434822 39896
rect 434266 39340 434502 39576
rect 434586 39340 434822 39576
rect 434266 3660 434502 3896
rect 434586 3660 434822 3896
rect 434266 3340 434502 3576
rect 434586 3340 434822 3576
rect 434266 -1540 434502 -1304
rect 434586 -1540 434822 -1304
rect 434266 -1860 434502 -1624
rect 434586 -1860 434822 -1624
rect 435506 706524 435742 706760
rect 435826 706524 436062 706760
rect 435506 706204 435742 706440
rect 435826 706204 436062 706440
rect 435506 688900 435742 689136
rect 435826 688900 436062 689136
rect 435506 688580 435742 688816
rect 435826 688580 436062 688816
rect 435506 652900 435742 653136
rect 435826 652900 436062 653136
rect 435506 652580 435742 652816
rect 435826 652580 436062 652816
rect 435506 616900 435742 617136
rect 435826 616900 436062 617136
rect 435506 616580 435742 616816
rect 435826 616580 436062 616816
rect 435506 580900 435742 581136
rect 435826 580900 436062 581136
rect 435506 580580 435742 580816
rect 435826 580580 436062 580816
rect 435506 544900 435742 545136
rect 435826 544900 436062 545136
rect 435506 544580 435742 544816
rect 435826 544580 436062 544816
rect 435506 508900 435742 509136
rect 435826 508900 436062 509136
rect 435506 508580 435742 508816
rect 435826 508580 436062 508816
rect 435506 472900 435742 473136
rect 435826 472900 436062 473136
rect 435506 472580 435742 472816
rect 435826 472580 436062 472816
rect 435506 436900 435742 437136
rect 435826 436900 436062 437136
rect 435506 436580 435742 436816
rect 435826 436580 436062 436816
rect 435506 400900 435742 401136
rect 435826 400900 436062 401136
rect 435506 400580 435742 400816
rect 435826 400580 436062 400816
rect 435506 364900 435742 365136
rect 435826 364900 436062 365136
rect 435506 364580 435742 364816
rect 435826 364580 436062 364816
rect 435506 328900 435742 329136
rect 435826 328900 436062 329136
rect 435506 328580 435742 328816
rect 435826 328580 436062 328816
rect 435506 292900 435742 293136
rect 435826 292900 436062 293136
rect 435506 292580 435742 292816
rect 435826 292580 436062 292816
rect 435506 256900 435742 257136
rect 435826 256900 436062 257136
rect 435506 256580 435742 256816
rect 435826 256580 436062 256816
rect 435506 220900 435742 221136
rect 435826 220900 436062 221136
rect 435506 220580 435742 220816
rect 435826 220580 436062 220816
rect 435506 184900 435742 185136
rect 435826 184900 436062 185136
rect 435506 184580 435742 184816
rect 435826 184580 436062 184816
rect 435506 148900 435742 149136
rect 435826 148900 436062 149136
rect 435506 148580 435742 148816
rect 435826 148580 436062 148816
rect 435506 112900 435742 113136
rect 435826 112900 436062 113136
rect 435506 112580 435742 112816
rect 435826 112580 436062 112816
rect 435506 76900 435742 77136
rect 435826 76900 436062 77136
rect 435506 76580 435742 76816
rect 435826 76580 436062 76816
rect 435506 40900 435742 41136
rect 435826 40900 436062 41136
rect 435506 40580 435742 40816
rect 435826 40580 436062 40816
rect 435506 4900 435742 5136
rect 435826 4900 436062 5136
rect 435506 4580 435742 4816
rect 435826 4580 436062 4816
rect 435506 -2500 435742 -2264
rect 435826 -2500 436062 -2264
rect 435506 -2820 435742 -2584
rect 435826 -2820 436062 -2584
rect 436746 707484 436982 707720
rect 437066 707484 437302 707720
rect 436746 707164 436982 707400
rect 437066 707164 437302 707400
rect 436746 690140 436982 690376
rect 437066 690140 437302 690376
rect 436746 689820 436982 690056
rect 437066 689820 437302 690056
rect 436746 654140 436982 654376
rect 437066 654140 437302 654376
rect 436746 653820 436982 654056
rect 437066 653820 437302 654056
rect 436746 618140 436982 618376
rect 437066 618140 437302 618376
rect 436746 617820 436982 618056
rect 437066 617820 437302 618056
rect 436746 582140 436982 582376
rect 437066 582140 437302 582376
rect 436746 581820 436982 582056
rect 437066 581820 437302 582056
rect 436746 546140 436982 546376
rect 437066 546140 437302 546376
rect 436746 545820 436982 546056
rect 437066 545820 437302 546056
rect 436746 510140 436982 510376
rect 437066 510140 437302 510376
rect 436746 509820 436982 510056
rect 437066 509820 437302 510056
rect 436746 474140 436982 474376
rect 437066 474140 437302 474376
rect 436746 473820 436982 474056
rect 437066 473820 437302 474056
rect 436746 438140 436982 438376
rect 437066 438140 437302 438376
rect 436746 437820 436982 438056
rect 437066 437820 437302 438056
rect 436746 402140 436982 402376
rect 437066 402140 437302 402376
rect 436746 401820 436982 402056
rect 437066 401820 437302 402056
rect 436746 366140 436982 366376
rect 437066 366140 437302 366376
rect 436746 365820 436982 366056
rect 437066 365820 437302 366056
rect 436746 330140 436982 330376
rect 437066 330140 437302 330376
rect 436746 329820 436982 330056
rect 437066 329820 437302 330056
rect 436746 294140 436982 294376
rect 437066 294140 437302 294376
rect 436746 293820 436982 294056
rect 437066 293820 437302 294056
rect 436746 258140 436982 258376
rect 437066 258140 437302 258376
rect 436746 257820 436982 258056
rect 437066 257820 437302 258056
rect 436746 222140 436982 222376
rect 437066 222140 437302 222376
rect 436746 221820 436982 222056
rect 437066 221820 437302 222056
rect 436746 186140 436982 186376
rect 437066 186140 437302 186376
rect 436746 185820 436982 186056
rect 437066 185820 437302 186056
rect 436746 150140 436982 150376
rect 437066 150140 437302 150376
rect 436746 149820 436982 150056
rect 437066 149820 437302 150056
rect 436746 114140 436982 114376
rect 437066 114140 437302 114376
rect 436746 113820 436982 114056
rect 437066 113820 437302 114056
rect 436746 78140 436982 78376
rect 437066 78140 437302 78376
rect 436746 77820 436982 78056
rect 437066 77820 437302 78056
rect 436746 42140 436982 42376
rect 437066 42140 437302 42376
rect 436746 41820 436982 42056
rect 437066 41820 437302 42056
rect 436746 6140 436982 6376
rect 437066 6140 437302 6376
rect 436746 5820 436982 6056
rect 437066 5820 437302 6056
rect 436746 -3460 436982 -3224
rect 437066 -3460 437302 -3224
rect 436746 -3780 436982 -3544
rect 437066 -3780 437302 -3544
rect 437986 708444 438222 708680
rect 438306 708444 438542 708680
rect 437986 708124 438222 708360
rect 438306 708124 438542 708360
rect 437986 691380 438222 691616
rect 438306 691380 438542 691616
rect 437986 691060 438222 691296
rect 438306 691060 438542 691296
rect 437986 655380 438222 655616
rect 438306 655380 438542 655616
rect 437986 655060 438222 655296
rect 438306 655060 438542 655296
rect 437986 619380 438222 619616
rect 438306 619380 438542 619616
rect 437986 619060 438222 619296
rect 438306 619060 438542 619296
rect 437986 583380 438222 583616
rect 438306 583380 438542 583616
rect 437986 583060 438222 583296
rect 438306 583060 438542 583296
rect 437986 547380 438222 547616
rect 438306 547380 438542 547616
rect 437986 547060 438222 547296
rect 438306 547060 438542 547296
rect 437986 511380 438222 511616
rect 438306 511380 438542 511616
rect 437986 511060 438222 511296
rect 438306 511060 438542 511296
rect 437986 475380 438222 475616
rect 438306 475380 438542 475616
rect 437986 475060 438222 475296
rect 438306 475060 438542 475296
rect 437986 439380 438222 439616
rect 438306 439380 438542 439616
rect 437986 439060 438222 439296
rect 438306 439060 438542 439296
rect 437986 403380 438222 403616
rect 438306 403380 438542 403616
rect 437986 403060 438222 403296
rect 438306 403060 438542 403296
rect 437986 367380 438222 367616
rect 438306 367380 438542 367616
rect 437986 367060 438222 367296
rect 438306 367060 438542 367296
rect 437986 331380 438222 331616
rect 438306 331380 438542 331616
rect 437986 331060 438222 331296
rect 438306 331060 438542 331296
rect 437986 295380 438222 295616
rect 438306 295380 438542 295616
rect 437986 295060 438222 295296
rect 438306 295060 438542 295296
rect 437986 259380 438222 259616
rect 438306 259380 438542 259616
rect 437986 259060 438222 259296
rect 438306 259060 438542 259296
rect 437986 223380 438222 223616
rect 438306 223380 438542 223616
rect 437986 223060 438222 223296
rect 438306 223060 438542 223296
rect 437986 187380 438222 187616
rect 438306 187380 438542 187616
rect 437986 187060 438222 187296
rect 438306 187060 438542 187296
rect 437986 151380 438222 151616
rect 438306 151380 438542 151616
rect 437986 151060 438222 151296
rect 438306 151060 438542 151296
rect 437986 115380 438222 115616
rect 438306 115380 438542 115616
rect 437986 115060 438222 115296
rect 438306 115060 438542 115296
rect 437986 79380 438222 79616
rect 438306 79380 438542 79616
rect 437986 79060 438222 79296
rect 438306 79060 438542 79296
rect 437986 43380 438222 43616
rect 438306 43380 438542 43616
rect 437986 43060 438222 43296
rect 438306 43060 438542 43296
rect 437986 7380 438222 7616
rect 438306 7380 438542 7616
rect 437986 7060 438222 7296
rect 438306 7060 438542 7296
rect 437986 -4420 438222 -4184
rect 438306 -4420 438542 -4184
rect 437986 -4740 438222 -4504
rect 438306 -4740 438542 -4504
rect 439226 709404 439462 709640
rect 439546 709404 439782 709640
rect 439226 709084 439462 709320
rect 439546 709084 439782 709320
rect 439226 692620 439462 692856
rect 439546 692620 439782 692856
rect 439226 692300 439462 692536
rect 439546 692300 439782 692536
rect 439226 656620 439462 656856
rect 439546 656620 439782 656856
rect 439226 656300 439462 656536
rect 439546 656300 439782 656536
rect 439226 620620 439462 620856
rect 439546 620620 439782 620856
rect 439226 620300 439462 620536
rect 439546 620300 439782 620536
rect 439226 584620 439462 584856
rect 439546 584620 439782 584856
rect 439226 584300 439462 584536
rect 439546 584300 439782 584536
rect 439226 548620 439462 548856
rect 439546 548620 439782 548856
rect 439226 548300 439462 548536
rect 439546 548300 439782 548536
rect 439226 512620 439462 512856
rect 439546 512620 439782 512856
rect 439226 512300 439462 512536
rect 439546 512300 439782 512536
rect 439226 476620 439462 476856
rect 439546 476620 439782 476856
rect 439226 476300 439462 476536
rect 439546 476300 439782 476536
rect 439226 440620 439462 440856
rect 439546 440620 439782 440856
rect 439226 440300 439462 440536
rect 439546 440300 439782 440536
rect 439226 404620 439462 404856
rect 439546 404620 439782 404856
rect 439226 404300 439462 404536
rect 439546 404300 439782 404536
rect 439226 368620 439462 368856
rect 439546 368620 439782 368856
rect 439226 368300 439462 368536
rect 439546 368300 439782 368536
rect 439226 332620 439462 332856
rect 439546 332620 439782 332856
rect 439226 332300 439462 332536
rect 439546 332300 439782 332536
rect 439226 296620 439462 296856
rect 439546 296620 439782 296856
rect 439226 296300 439462 296536
rect 439546 296300 439782 296536
rect 439226 260620 439462 260856
rect 439546 260620 439782 260856
rect 439226 260300 439462 260536
rect 439546 260300 439782 260536
rect 439226 224620 439462 224856
rect 439546 224620 439782 224856
rect 439226 224300 439462 224536
rect 439546 224300 439782 224536
rect 439226 188620 439462 188856
rect 439546 188620 439782 188856
rect 439226 188300 439462 188536
rect 439546 188300 439782 188536
rect 439226 152620 439462 152856
rect 439546 152620 439782 152856
rect 439226 152300 439462 152536
rect 439546 152300 439782 152536
rect 439226 116620 439462 116856
rect 439546 116620 439782 116856
rect 439226 116300 439462 116536
rect 439546 116300 439782 116536
rect 439226 80620 439462 80856
rect 439546 80620 439782 80856
rect 439226 80300 439462 80536
rect 439546 80300 439782 80536
rect 439226 44620 439462 44856
rect 439546 44620 439782 44856
rect 439226 44300 439462 44536
rect 439546 44300 439782 44536
rect 439226 8620 439462 8856
rect 439546 8620 439782 8856
rect 439226 8300 439462 8536
rect 439546 8300 439782 8536
rect 439226 -5380 439462 -5144
rect 439546 -5380 439782 -5144
rect 439226 -5700 439462 -5464
rect 439546 -5700 439782 -5464
rect 440466 710364 440702 710600
rect 440786 710364 441022 710600
rect 440466 710044 440702 710280
rect 440786 710044 441022 710280
rect 440466 693860 440702 694096
rect 440786 693860 441022 694096
rect 440466 693540 440702 693776
rect 440786 693540 441022 693776
rect 440466 657860 440702 658096
rect 440786 657860 441022 658096
rect 440466 657540 440702 657776
rect 440786 657540 441022 657776
rect 440466 621860 440702 622096
rect 440786 621860 441022 622096
rect 440466 621540 440702 621776
rect 440786 621540 441022 621776
rect 440466 585860 440702 586096
rect 440786 585860 441022 586096
rect 440466 585540 440702 585776
rect 440786 585540 441022 585776
rect 440466 549860 440702 550096
rect 440786 549860 441022 550096
rect 440466 549540 440702 549776
rect 440786 549540 441022 549776
rect 440466 513860 440702 514096
rect 440786 513860 441022 514096
rect 440466 513540 440702 513776
rect 440786 513540 441022 513776
rect 440466 477860 440702 478096
rect 440786 477860 441022 478096
rect 440466 477540 440702 477776
rect 440786 477540 441022 477776
rect 440466 441860 440702 442096
rect 440786 441860 441022 442096
rect 440466 441540 440702 441776
rect 440786 441540 441022 441776
rect 440466 405860 440702 406096
rect 440786 405860 441022 406096
rect 440466 405540 440702 405776
rect 440786 405540 441022 405776
rect 440466 369860 440702 370096
rect 440786 369860 441022 370096
rect 440466 369540 440702 369776
rect 440786 369540 441022 369776
rect 440466 333860 440702 334096
rect 440786 333860 441022 334096
rect 440466 333540 440702 333776
rect 440786 333540 441022 333776
rect 440466 297860 440702 298096
rect 440786 297860 441022 298096
rect 440466 297540 440702 297776
rect 440786 297540 441022 297776
rect 440466 261860 440702 262096
rect 440786 261860 441022 262096
rect 440466 261540 440702 261776
rect 440786 261540 441022 261776
rect 440466 225860 440702 226096
rect 440786 225860 441022 226096
rect 440466 225540 440702 225776
rect 440786 225540 441022 225776
rect 440466 189860 440702 190096
rect 440786 189860 441022 190096
rect 440466 189540 440702 189776
rect 440786 189540 441022 189776
rect 440466 153860 440702 154096
rect 440786 153860 441022 154096
rect 440466 153540 440702 153776
rect 440786 153540 441022 153776
rect 440466 117860 440702 118096
rect 440786 117860 441022 118096
rect 440466 117540 440702 117776
rect 440786 117540 441022 117776
rect 440466 81860 440702 82096
rect 440786 81860 441022 82096
rect 440466 81540 440702 81776
rect 440786 81540 441022 81776
rect 440466 45860 440702 46096
rect 440786 45860 441022 46096
rect 440466 45540 440702 45776
rect 440786 45540 441022 45776
rect 440466 9860 440702 10096
rect 440786 9860 441022 10096
rect 440466 9540 440702 9776
rect 440786 9540 441022 9776
rect 440466 -6340 440702 -6104
rect 440786 -6340 441022 -6104
rect 440466 -6660 440702 -6424
rect 440786 -6660 441022 -6424
rect 441706 711324 441942 711560
rect 442026 711324 442262 711560
rect 441706 711004 441942 711240
rect 442026 711004 442262 711240
rect 441706 695100 441942 695336
rect 442026 695100 442262 695336
rect 441706 694780 441942 695016
rect 442026 694780 442262 695016
rect 441706 659100 441942 659336
rect 442026 659100 442262 659336
rect 441706 658780 441942 659016
rect 442026 658780 442262 659016
rect 441706 623100 441942 623336
rect 442026 623100 442262 623336
rect 441706 622780 441942 623016
rect 442026 622780 442262 623016
rect 441706 587100 441942 587336
rect 442026 587100 442262 587336
rect 441706 586780 441942 587016
rect 442026 586780 442262 587016
rect 441706 551100 441942 551336
rect 442026 551100 442262 551336
rect 441706 550780 441942 551016
rect 442026 550780 442262 551016
rect 441706 515100 441942 515336
rect 442026 515100 442262 515336
rect 441706 514780 441942 515016
rect 442026 514780 442262 515016
rect 441706 479100 441942 479336
rect 442026 479100 442262 479336
rect 441706 478780 441942 479016
rect 442026 478780 442262 479016
rect 441706 443100 441942 443336
rect 442026 443100 442262 443336
rect 441706 442780 441942 443016
rect 442026 442780 442262 443016
rect 441706 407100 441942 407336
rect 442026 407100 442262 407336
rect 441706 406780 441942 407016
rect 442026 406780 442262 407016
rect 441706 371100 441942 371336
rect 442026 371100 442262 371336
rect 441706 370780 441942 371016
rect 442026 370780 442262 371016
rect 441706 335100 441942 335336
rect 442026 335100 442262 335336
rect 441706 334780 441942 335016
rect 442026 334780 442262 335016
rect 441706 299100 441942 299336
rect 442026 299100 442262 299336
rect 441706 298780 441942 299016
rect 442026 298780 442262 299016
rect 441706 263100 441942 263336
rect 442026 263100 442262 263336
rect 441706 262780 441942 263016
rect 442026 262780 442262 263016
rect 441706 227100 441942 227336
rect 442026 227100 442262 227336
rect 441706 226780 441942 227016
rect 442026 226780 442262 227016
rect 441706 191100 441942 191336
rect 442026 191100 442262 191336
rect 441706 190780 441942 191016
rect 442026 190780 442262 191016
rect 441706 155100 441942 155336
rect 442026 155100 442262 155336
rect 441706 154780 441942 155016
rect 442026 154780 442262 155016
rect 441706 119100 441942 119336
rect 442026 119100 442262 119336
rect 441706 118780 441942 119016
rect 442026 118780 442262 119016
rect 441706 83100 441942 83336
rect 442026 83100 442262 83336
rect 441706 82780 441942 83016
rect 442026 82780 442262 83016
rect 441706 47100 441942 47336
rect 442026 47100 442262 47336
rect 441706 46780 441942 47016
rect 442026 46780 442262 47016
rect 441706 11100 441942 11336
rect 442026 11100 442262 11336
rect 441706 10780 441942 11016
rect 442026 10780 442262 11016
rect 441706 -7300 441942 -7064
rect 442026 -7300 442262 -7064
rect 441706 -7620 441942 -7384
rect 442026 -7620 442262 -7384
rect 469026 704604 469262 704840
rect 469346 704604 469582 704840
rect 469026 704284 469262 704520
rect 469346 704284 469582 704520
rect 469026 686420 469262 686656
rect 469346 686420 469582 686656
rect 469026 686100 469262 686336
rect 469346 686100 469582 686336
rect 469026 650420 469262 650656
rect 469346 650420 469582 650656
rect 469026 650100 469262 650336
rect 469346 650100 469582 650336
rect 469026 614420 469262 614656
rect 469346 614420 469582 614656
rect 469026 614100 469262 614336
rect 469346 614100 469582 614336
rect 469026 578420 469262 578656
rect 469346 578420 469582 578656
rect 469026 578100 469262 578336
rect 469346 578100 469582 578336
rect 469026 542420 469262 542656
rect 469346 542420 469582 542656
rect 469026 542100 469262 542336
rect 469346 542100 469582 542336
rect 469026 506420 469262 506656
rect 469346 506420 469582 506656
rect 469026 506100 469262 506336
rect 469346 506100 469582 506336
rect 469026 470420 469262 470656
rect 469346 470420 469582 470656
rect 469026 470100 469262 470336
rect 469346 470100 469582 470336
rect 469026 434420 469262 434656
rect 469346 434420 469582 434656
rect 469026 434100 469262 434336
rect 469346 434100 469582 434336
rect 469026 398420 469262 398656
rect 469346 398420 469582 398656
rect 469026 398100 469262 398336
rect 469346 398100 469582 398336
rect 469026 362420 469262 362656
rect 469346 362420 469582 362656
rect 469026 362100 469262 362336
rect 469346 362100 469582 362336
rect 469026 326420 469262 326656
rect 469346 326420 469582 326656
rect 469026 326100 469262 326336
rect 469346 326100 469582 326336
rect 469026 290420 469262 290656
rect 469346 290420 469582 290656
rect 469026 290100 469262 290336
rect 469346 290100 469582 290336
rect 469026 254420 469262 254656
rect 469346 254420 469582 254656
rect 469026 254100 469262 254336
rect 469346 254100 469582 254336
rect 469026 218420 469262 218656
rect 469346 218420 469582 218656
rect 469026 218100 469262 218336
rect 469346 218100 469582 218336
rect 469026 182420 469262 182656
rect 469346 182420 469582 182656
rect 469026 182100 469262 182336
rect 469346 182100 469582 182336
rect 469026 146420 469262 146656
rect 469346 146420 469582 146656
rect 469026 146100 469262 146336
rect 469346 146100 469582 146336
rect 469026 110420 469262 110656
rect 469346 110420 469582 110656
rect 469026 110100 469262 110336
rect 469346 110100 469582 110336
rect 469026 74420 469262 74656
rect 469346 74420 469582 74656
rect 469026 74100 469262 74336
rect 469346 74100 469582 74336
rect 469026 38420 469262 38656
rect 469346 38420 469582 38656
rect 469026 38100 469262 38336
rect 469346 38100 469582 38336
rect 469026 2420 469262 2656
rect 469346 2420 469582 2656
rect 469026 2100 469262 2336
rect 469346 2100 469582 2336
rect 469026 -580 469262 -344
rect 469346 -580 469582 -344
rect 469026 -900 469262 -664
rect 469346 -900 469582 -664
rect 470266 705564 470502 705800
rect 470586 705564 470822 705800
rect 470266 705244 470502 705480
rect 470586 705244 470822 705480
rect 470266 687660 470502 687896
rect 470586 687660 470822 687896
rect 470266 687340 470502 687576
rect 470586 687340 470822 687576
rect 470266 651660 470502 651896
rect 470586 651660 470822 651896
rect 470266 651340 470502 651576
rect 470586 651340 470822 651576
rect 470266 615660 470502 615896
rect 470586 615660 470822 615896
rect 470266 615340 470502 615576
rect 470586 615340 470822 615576
rect 470266 579660 470502 579896
rect 470586 579660 470822 579896
rect 470266 579340 470502 579576
rect 470586 579340 470822 579576
rect 470266 543660 470502 543896
rect 470586 543660 470822 543896
rect 470266 543340 470502 543576
rect 470586 543340 470822 543576
rect 470266 507660 470502 507896
rect 470586 507660 470822 507896
rect 470266 507340 470502 507576
rect 470586 507340 470822 507576
rect 470266 471660 470502 471896
rect 470586 471660 470822 471896
rect 470266 471340 470502 471576
rect 470586 471340 470822 471576
rect 470266 435660 470502 435896
rect 470586 435660 470822 435896
rect 470266 435340 470502 435576
rect 470586 435340 470822 435576
rect 470266 399660 470502 399896
rect 470586 399660 470822 399896
rect 470266 399340 470502 399576
rect 470586 399340 470822 399576
rect 470266 363660 470502 363896
rect 470586 363660 470822 363896
rect 470266 363340 470502 363576
rect 470586 363340 470822 363576
rect 470266 327660 470502 327896
rect 470586 327660 470822 327896
rect 470266 327340 470502 327576
rect 470586 327340 470822 327576
rect 470266 291660 470502 291896
rect 470586 291660 470822 291896
rect 470266 291340 470502 291576
rect 470586 291340 470822 291576
rect 470266 255660 470502 255896
rect 470586 255660 470822 255896
rect 470266 255340 470502 255576
rect 470586 255340 470822 255576
rect 470266 219660 470502 219896
rect 470586 219660 470822 219896
rect 470266 219340 470502 219576
rect 470586 219340 470822 219576
rect 470266 183660 470502 183896
rect 470586 183660 470822 183896
rect 470266 183340 470502 183576
rect 470586 183340 470822 183576
rect 470266 147660 470502 147896
rect 470586 147660 470822 147896
rect 470266 147340 470502 147576
rect 470586 147340 470822 147576
rect 470266 111660 470502 111896
rect 470586 111660 470822 111896
rect 470266 111340 470502 111576
rect 470586 111340 470822 111576
rect 470266 75660 470502 75896
rect 470586 75660 470822 75896
rect 470266 75340 470502 75576
rect 470586 75340 470822 75576
rect 470266 39660 470502 39896
rect 470586 39660 470822 39896
rect 470266 39340 470502 39576
rect 470586 39340 470822 39576
rect 470266 3660 470502 3896
rect 470586 3660 470822 3896
rect 470266 3340 470502 3576
rect 470586 3340 470822 3576
rect 470266 -1540 470502 -1304
rect 470586 -1540 470822 -1304
rect 470266 -1860 470502 -1624
rect 470586 -1860 470822 -1624
rect 471506 706524 471742 706760
rect 471826 706524 472062 706760
rect 471506 706204 471742 706440
rect 471826 706204 472062 706440
rect 471506 688900 471742 689136
rect 471826 688900 472062 689136
rect 471506 688580 471742 688816
rect 471826 688580 472062 688816
rect 471506 652900 471742 653136
rect 471826 652900 472062 653136
rect 471506 652580 471742 652816
rect 471826 652580 472062 652816
rect 471506 616900 471742 617136
rect 471826 616900 472062 617136
rect 471506 616580 471742 616816
rect 471826 616580 472062 616816
rect 471506 580900 471742 581136
rect 471826 580900 472062 581136
rect 471506 580580 471742 580816
rect 471826 580580 472062 580816
rect 471506 544900 471742 545136
rect 471826 544900 472062 545136
rect 471506 544580 471742 544816
rect 471826 544580 472062 544816
rect 471506 508900 471742 509136
rect 471826 508900 472062 509136
rect 471506 508580 471742 508816
rect 471826 508580 472062 508816
rect 471506 472900 471742 473136
rect 471826 472900 472062 473136
rect 471506 472580 471742 472816
rect 471826 472580 472062 472816
rect 471506 436900 471742 437136
rect 471826 436900 472062 437136
rect 471506 436580 471742 436816
rect 471826 436580 472062 436816
rect 471506 400900 471742 401136
rect 471826 400900 472062 401136
rect 471506 400580 471742 400816
rect 471826 400580 472062 400816
rect 471506 364900 471742 365136
rect 471826 364900 472062 365136
rect 471506 364580 471742 364816
rect 471826 364580 472062 364816
rect 472746 707484 472982 707720
rect 473066 707484 473302 707720
rect 472746 707164 472982 707400
rect 473066 707164 473302 707400
rect 472746 690140 472982 690376
rect 473066 690140 473302 690376
rect 472746 689820 472982 690056
rect 473066 689820 473302 690056
rect 472746 654140 472982 654376
rect 473066 654140 473302 654376
rect 472746 653820 472982 654056
rect 473066 653820 473302 654056
rect 472746 618140 472982 618376
rect 473066 618140 473302 618376
rect 472746 617820 472982 618056
rect 473066 617820 473302 618056
rect 472746 582140 472982 582376
rect 473066 582140 473302 582376
rect 472746 581820 472982 582056
rect 473066 581820 473302 582056
rect 472746 546140 472982 546376
rect 473066 546140 473302 546376
rect 472746 545820 472982 546056
rect 473066 545820 473302 546056
rect 472746 510140 472982 510376
rect 473066 510140 473302 510376
rect 472746 509820 472982 510056
rect 473066 509820 473302 510056
rect 472746 474140 472982 474376
rect 473066 474140 473302 474376
rect 472746 473820 472982 474056
rect 473066 473820 473302 474056
rect 473986 708444 474222 708680
rect 474306 708444 474542 708680
rect 473986 708124 474222 708360
rect 474306 708124 474542 708360
rect 473986 691380 474222 691616
rect 474306 691380 474542 691616
rect 473986 691060 474222 691296
rect 474306 691060 474542 691296
rect 473986 655380 474222 655616
rect 474306 655380 474542 655616
rect 473986 655060 474222 655296
rect 474306 655060 474542 655296
rect 473986 619380 474222 619616
rect 474306 619380 474542 619616
rect 473986 619060 474222 619296
rect 474306 619060 474542 619296
rect 473986 583380 474222 583616
rect 474306 583380 474542 583616
rect 473986 583060 474222 583296
rect 474306 583060 474542 583296
rect 473986 547380 474222 547616
rect 474306 547380 474542 547616
rect 473986 547060 474222 547296
rect 474306 547060 474542 547296
rect 473986 511380 474222 511616
rect 474306 511380 474542 511616
rect 473986 511060 474222 511296
rect 474306 511060 474542 511296
rect 473986 475380 474222 475616
rect 474306 475380 474542 475616
rect 473986 475060 474222 475296
rect 474306 475060 474542 475296
rect 472746 438140 472982 438376
rect 473066 438140 473302 438376
rect 472746 437820 472982 438056
rect 473066 437820 473302 438056
rect 473986 439380 474222 439616
rect 474306 439380 474542 439616
rect 473986 439060 474222 439296
rect 474306 439060 474542 439296
rect 472746 402140 472982 402376
rect 473066 402140 473302 402376
rect 472746 401820 472982 402056
rect 473066 401820 473302 402056
rect 473986 403380 474222 403616
rect 474306 403380 474542 403616
rect 473986 403060 474222 403296
rect 474306 403060 474542 403296
rect 472746 366140 472982 366376
rect 473066 366140 473302 366376
rect 472746 365820 472982 366056
rect 473066 365820 473302 366056
rect 475226 709404 475462 709640
rect 475546 709404 475782 709640
rect 475226 709084 475462 709320
rect 475546 709084 475782 709320
rect 475226 692620 475462 692856
rect 475546 692620 475782 692856
rect 475226 692300 475462 692536
rect 475546 692300 475782 692536
rect 475226 656620 475462 656856
rect 475546 656620 475782 656856
rect 475226 656300 475462 656536
rect 475546 656300 475782 656536
rect 475226 620620 475462 620856
rect 475546 620620 475782 620856
rect 475226 620300 475462 620536
rect 475546 620300 475782 620536
rect 475226 584620 475462 584856
rect 475546 584620 475782 584856
rect 475226 584300 475462 584536
rect 475546 584300 475782 584536
rect 475226 548620 475462 548856
rect 475546 548620 475782 548856
rect 475226 548300 475462 548536
rect 475546 548300 475782 548536
rect 475226 512620 475462 512856
rect 475546 512620 475782 512856
rect 475226 512300 475462 512536
rect 475546 512300 475782 512536
rect 475226 476620 475462 476856
rect 475546 476620 475782 476856
rect 475226 476300 475462 476536
rect 475546 476300 475782 476536
rect 475226 440620 475462 440856
rect 475546 440620 475782 440856
rect 475226 440300 475462 440536
rect 475546 440300 475782 440536
rect 475226 404620 475462 404856
rect 475546 404620 475782 404856
rect 475226 404300 475462 404536
rect 475546 404300 475782 404536
rect 473986 367380 474222 367616
rect 474306 367380 474542 367616
rect 473986 367060 474222 367296
rect 474306 367060 474542 367296
rect 475226 368620 475462 368856
rect 475546 368620 475782 368856
rect 475226 368300 475462 368536
rect 475546 368300 475782 368536
rect 476466 710364 476702 710600
rect 476786 710364 477022 710600
rect 476466 710044 476702 710280
rect 476786 710044 477022 710280
rect 476466 693860 476702 694096
rect 476786 693860 477022 694096
rect 476466 693540 476702 693776
rect 476786 693540 477022 693776
rect 476466 657860 476702 658096
rect 476786 657860 477022 658096
rect 476466 657540 476702 657776
rect 476786 657540 477022 657776
rect 476466 621860 476702 622096
rect 476786 621860 477022 622096
rect 476466 621540 476702 621776
rect 476786 621540 477022 621776
rect 476466 585860 476702 586096
rect 476786 585860 477022 586096
rect 476466 585540 476702 585776
rect 476786 585540 477022 585776
rect 476466 549860 476702 550096
rect 476786 549860 477022 550096
rect 476466 549540 476702 549776
rect 476786 549540 477022 549776
rect 476466 513860 476702 514096
rect 476786 513860 477022 514096
rect 476466 513540 476702 513776
rect 476786 513540 477022 513776
rect 476466 477860 476702 478096
rect 476786 477860 477022 478096
rect 476466 477540 476702 477776
rect 476786 477540 477022 477776
rect 476466 441860 476702 442096
rect 476786 441860 477022 442096
rect 476466 441540 476702 441776
rect 476786 441540 477022 441776
rect 476466 405860 476702 406096
rect 476786 405860 477022 406096
rect 476466 405540 476702 405776
rect 476786 405540 477022 405776
rect 476466 369860 476702 370096
rect 476786 369860 477022 370096
rect 476466 369540 476702 369776
rect 476786 369540 477022 369776
rect 477706 711324 477942 711560
rect 478026 711324 478262 711560
rect 477706 711004 477942 711240
rect 478026 711004 478262 711240
rect 477706 695100 477942 695336
rect 478026 695100 478262 695336
rect 477706 694780 477942 695016
rect 478026 694780 478262 695016
rect 477706 659100 477942 659336
rect 478026 659100 478262 659336
rect 477706 658780 477942 659016
rect 478026 658780 478262 659016
rect 477706 623100 477942 623336
rect 478026 623100 478262 623336
rect 477706 622780 477942 623016
rect 478026 622780 478262 623016
rect 477706 587100 477942 587336
rect 478026 587100 478262 587336
rect 477706 586780 477942 587016
rect 478026 586780 478262 587016
rect 477706 551100 477942 551336
rect 478026 551100 478262 551336
rect 477706 550780 477942 551016
rect 478026 550780 478262 551016
rect 477706 515100 477942 515336
rect 478026 515100 478262 515336
rect 477706 514780 477942 515016
rect 478026 514780 478262 515016
rect 477706 479100 477942 479336
rect 478026 479100 478262 479336
rect 477706 478780 477942 479016
rect 478026 478780 478262 479016
rect 505026 704604 505262 704840
rect 505346 704604 505582 704840
rect 505026 704284 505262 704520
rect 505346 704284 505582 704520
rect 505026 686420 505262 686656
rect 505346 686420 505582 686656
rect 505026 686100 505262 686336
rect 505346 686100 505582 686336
rect 505026 650420 505262 650656
rect 505346 650420 505582 650656
rect 505026 650100 505262 650336
rect 505346 650100 505582 650336
rect 505026 614420 505262 614656
rect 505346 614420 505582 614656
rect 505026 614100 505262 614336
rect 505346 614100 505582 614336
rect 505026 578420 505262 578656
rect 505346 578420 505582 578656
rect 505026 578100 505262 578336
rect 505346 578100 505582 578336
rect 505026 542420 505262 542656
rect 505346 542420 505582 542656
rect 505026 542100 505262 542336
rect 505346 542100 505582 542336
rect 505026 506420 505262 506656
rect 505346 506420 505582 506656
rect 505026 506100 505262 506336
rect 505346 506100 505582 506336
rect 505026 470420 505262 470656
rect 505346 470420 505582 470656
rect 505026 470100 505262 470336
rect 505346 470100 505582 470336
rect 477706 443100 477942 443336
rect 478026 443100 478262 443336
rect 477706 442780 477942 443016
rect 478026 442780 478262 443016
rect 477706 407100 477942 407336
rect 478026 407100 478262 407336
rect 477706 406780 477942 407016
rect 478026 406780 478262 407016
rect 505026 434420 505262 434656
rect 505346 434420 505582 434656
rect 505026 434100 505262 434336
rect 505346 434100 505582 434336
rect 477706 371100 477942 371336
rect 478026 371100 478262 371336
rect 477706 370780 477942 371016
rect 478026 370780 478262 371016
rect 471506 328900 471742 329136
rect 471826 328900 472062 329136
rect 471506 328580 471742 328816
rect 471826 328580 472062 328816
rect 471506 292900 471742 293136
rect 471826 292900 472062 293136
rect 471506 292580 471742 292816
rect 471826 292580 472062 292816
rect 472746 330140 472982 330376
rect 473066 330140 473302 330376
rect 472746 329820 472982 330056
rect 473066 329820 473302 330056
rect 473986 331380 474222 331616
rect 474306 331380 474542 331616
rect 473986 331060 474222 331296
rect 474306 331060 474542 331296
rect 472746 294140 472982 294376
rect 473066 294140 473302 294376
rect 472746 293820 472982 294056
rect 473066 293820 473302 294056
rect 473986 295380 474222 295616
rect 474306 295380 474542 295616
rect 473986 295060 474222 295296
rect 474306 295060 474542 295296
rect 475226 332620 475462 332856
rect 475546 332620 475782 332856
rect 475226 332300 475462 332536
rect 475546 332300 475782 332536
rect 475226 296620 475462 296856
rect 475546 296620 475782 296856
rect 475226 296300 475462 296536
rect 475546 296300 475782 296536
rect 476466 333860 476702 334096
rect 476786 333860 477022 334096
rect 476466 333540 476702 333776
rect 476786 333540 477022 333776
rect 476466 297860 476702 298096
rect 476786 297860 477022 298096
rect 476466 297540 476702 297776
rect 476786 297540 477022 297776
rect 477706 335100 477942 335336
rect 478026 335100 478262 335336
rect 477706 334780 477942 335016
rect 478026 334780 478262 335016
rect 505026 398420 505262 398656
rect 505346 398420 505582 398656
rect 505026 398100 505262 398336
rect 505346 398100 505582 398336
rect 505026 362420 505262 362656
rect 505346 362420 505582 362656
rect 505026 362100 505262 362336
rect 505346 362100 505582 362336
rect 505026 326420 505262 326656
rect 505346 326420 505582 326656
rect 505026 326100 505262 326336
rect 505346 326100 505582 326336
rect 477706 299100 477942 299336
rect 478026 299100 478262 299336
rect 477706 298780 477942 299016
rect 478026 298780 478262 299016
rect 505026 290420 505262 290656
rect 505346 290420 505582 290656
rect 505026 290100 505262 290336
rect 505346 290100 505582 290336
rect 471506 256900 471742 257136
rect 471826 256900 472062 257136
rect 471506 256580 471742 256816
rect 471826 256580 472062 256816
rect 471506 220900 471742 221136
rect 471826 220900 472062 221136
rect 471506 220580 471742 220816
rect 471826 220580 472062 220816
rect 471506 184900 471742 185136
rect 471826 184900 472062 185136
rect 471506 184580 471742 184816
rect 471826 184580 472062 184816
rect 471506 148900 471742 149136
rect 471826 148900 472062 149136
rect 471506 148580 471742 148816
rect 471826 148580 472062 148816
rect 471506 112900 471742 113136
rect 471826 112900 472062 113136
rect 471506 112580 471742 112816
rect 471826 112580 472062 112816
rect 471506 76900 471742 77136
rect 471826 76900 472062 77136
rect 471506 76580 471742 76816
rect 471826 76580 472062 76816
rect 471506 40900 471742 41136
rect 471826 40900 472062 41136
rect 471506 40580 471742 40816
rect 471826 40580 472062 40816
rect 471506 4900 471742 5136
rect 471826 4900 472062 5136
rect 471506 4580 471742 4816
rect 471826 4580 472062 4816
rect 471506 -2500 471742 -2264
rect 471826 -2500 472062 -2264
rect 471506 -2820 471742 -2584
rect 471826 -2820 472062 -2584
rect 472746 258140 472982 258376
rect 473066 258140 473302 258376
rect 472746 257820 472982 258056
rect 473066 257820 473302 258056
rect 472746 222140 472982 222376
rect 473066 222140 473302 222376
rect 472746 221820 472982 222056
rect 473066 221820 473302 222056
rect 472746 186140 472982 186376
rect 473066 186140 473302 186376
rect 472746 185820 472982 186056
rect 473066 185820 473302 186056
rect 472746 150140 472982 150376
rect 473066 150140 473302 150376
rect 472746 149820 472982 150056
rect 473066 149820 473302 150056
rect 472746 114140 472982 114376
rect 473066 114140 473302 114376
rect 472746 113820 472982 114056
rect 473066 113820 473302 114056
rect 472746 78140 472982 78376
rect 473066 78140 473302 78376
rect 472746 77820 472982 78056
rect 473066 77820 473302 78056
rect 472746 42140 472982 42376
rect 473066 42140 473302 42376
rect 472746 41820 472982 42056
rect 473066 41820 473302 42056
rect 472746 6140 472982 6376
rect 473066 6140 473302 6376
rect 472746 5820 472982 6056
rect 473066 5820 473302 6056
rect 472746 -3460 472982 -3224
rect 473066 -3460 473302 -3224
rect 472746 -3780 472982 -3544
rect 473066 -3780 473302 -3544
rect 473986 259380 474222 259616
rect 474306 259380 474542 259616
rect 473986 259060 474222 259296
rect 474306 259060 474542 259296
rect 473986 223380 474222 223616
rect 474306 223380 474542 223616
rect 473986 223060 474222 223296
rect 474306 223060 474542 223296
rect 473986 187380 474222 187616
rect 474306 187380 474542 187616
rect 473986 187060 474222 187296
rect 474306 187060 474542 187296
rect 473986 151380 474222 151616
rect 474306 151380 474542 151616
rect 473986 151060 474222 151296
rect 474306 151060 474542 151296
rect 473986 115380 474222 115616
rect 474306 115380 474542 115616
rect 473986 115060 474222 115296
rect 474306 115060 474542 115296
rect 473986 79380 474222 79616
rect 474306 79380 474542 79616
rect 473986 79060 474222 79296
rect 474306 79060 474542 79296
rect 473986 43380 474222 43616
rect 474306 43380 474542 43616
rect 473986 43060 474222 43296
rect 474306 43060 474542 43296
rect 473986 7380 474222 7616
rect 474306 7380 474542 7616
rect 473986 7060 474222 7296
rect 474306 7060 474542 7296
rect 473986 -4420 474222 -4184
rect 474306 -4420 474542 -4184
rect 473986 -4740 474222 -4504
rect 474306 -4740 474542 -4504
rect 475226 260620 475462 260856
rect 475546 260620 475782 260856
rect 475226 260300 475462 260536
rect 475546 260300 475782 260536
rect 475226 224620 475462 224856
rect 475546 224620 475782 224856
rect 475226 224300 475462 224536
rect 475546 224300 475782 224536
rect 475226 188620 475462 188856
rect 475546 188620 475782 188856
rect 475226 188300 475462 188536
rect 475546 188300 475782 188536
rect 475226 152620 475462 152856
rect 475546 152620 475782 152856
rect 475226 152300 475462 152536
rect 475546 152300 475782 152536
rect 475226 116620 475462 116856
rect 475546 116620 475782 116856
rect 475226 116300 475462 116536
rect 475546 116300 475782 116536
rect 475226 80620 475462 80856
rect 475546 80620 475782 80856
rect 475226 80300 475462 80536
rect 475546 80300 475782 80536
rect 475226 44620 475462 44856
rect 475546 44620 475782 44856
rect 475226 44300 475462 44536
rect 475546 44300 475782 44536
rect 475226 8620 475462 8856
rect 475546 8620 475782 8856
rect 475226 8300 475462 8536
rect 475546 8300 475782 8536
rect 475226 -5380 475462 -5144
rect 475546 -5380 475782 -5144
rect 475226 -5700 475462 -5464
rect 475546 -5700 475782 -5464
rect 476466 261860 476702 262096
rect 476786 261860 477022 262096
rect 476466 261540 476702 261776
rect 476786 261540 477022 261776
rect 476466 225860 476702 226096
rect 476786 225860 477022 226096
rect 476466 225540 476702 225776
rect 476786 225540 477022 225776
rect 477706 263100 477942 263336
rect 478026 263100 478262 263336
rect 477706 262780 477942 263016
rect 478026 262780 478262 263016
rect 505026 254420 505262 254656
rect 505346 254420 505582 254656
rect 505026 254100 505262 254336
rect 505346 254100 505582 254336
rect 477706 227100 477942 227336
rect 478026 227100 478262 227336
rect 477706 226780 477942 227016
rect 478026 226780 478262 227016
rect 476466 189860 476702 190096
rect 476786 189860 477022 190096
rect 476466 189540 476702 189776
rect 476786 189540 477022 189776
rect 476466 153860 476702 154096
rect 476786 153860 477022 154096
rect 476466 153540 476702 153776
rect 476786 153540 477022 153776
rect 476466 117860 476702 118096
rect 476786 117860 477022 118096
rect 476466 117540 476702 117776
rect 476786 117540 477022 117776
rect 476466 81860 476702 82096
rect 476786 81860 477022 82096
rect 476466 81540 476702 81776
rect 476786 81540 477022 81776
rect 476466 45860 476702 46096
rect 476786 45860 477022 46096
rect 476466 45540 476702 45776
rect 476786 45540 477022 45776
rect 476466 9860 476702 10096
rect 476786 9860 477022 10096
rect 476466 9540 476702 9776
rect 476786 9540 477022 9776
rect 476466 -6340 476702 -6104
rect 476786 -6340 477022 -6104
rect 476466 -6660 476702 -6424
rect 476786 -6660 477022 -6424
rect 477706 191100 477942 191336
rect 478026 191100 478262 191336
rect 477706 190780 477942 191016
rect 478026 190780 478262 191016
rect 477706 155100 477942 155336
rect 478026 155100 478262 155336
rect 477706 154780 477942 155016
rect 478026 154780 478262 155016
rect 477706 119100 477942 119336
rect 478026 119100 478262 119336
rect 477706 118780 477942 119016
rect 478026 118780 478262 119016
rect 477706 83100 477942 83336
rect 478026 83100 478262 83336
rect 477706 82780 477942 83016
rect 478026 82780 478262 83016
rect 477706 47100 477942 47336
rect 478026 47100 478262 47336
rect 477706 46780 477942 47016
rect 478026 46780 478262 47016
rect 477706 11100 477942 11336
rect 478026 11100 478262 11336
rect 477706 10780 477942 11016
rect 478026 10780 478262 11016
rect 477706 -7300 477942 -7064
rect 478026 -7300 478262 -7064
rect 477706 -7620 477942 -7384
rect 478026 -7620 478262 -7384
rect 505026 218420 505262 218656
rect 505346 218420 505582 218656
rect 505026 218100 505262 218336
rect 505346 218100 505582 218336
rect 505026 182420 505262 182656
rect 505346 182420 505582 182656
rect 505026 182100 505262 182336
rect 505346 182100 505582 182336
rect 505026 146420 505262 146656
rect 505346 146420 505582 146656
rect 505026 146100 505262 146336
rect 505346 146100 505582 146336
rect 505026 110420 505262 110656
rect 505346 110420 505582 110656
rect 505026 110100 505262 110336
rect 505346 110100 505582 110336
rect 505026 74420 505262 74656
rect 505346 74420 505582 74656
rect 505026 74100 505262 74336
rect 505346 74100 505582 74336
rect 505026 38420 505262 38656
rect 505346 38420 505582 38656
rect 505026 38100 505262 38336
rect 505346 38100 505582 38336
rect 505026 2420 505262 2656
rect 505346 2420 505582 2656
rect 505026 2100 505262 2336
rect 505346 2100 505582 2336
rect 505026 -580 505262 -344
rect 505346 -580 505582 -344
rect 505026 -900 505262 -664
rect 505346 -900 505582 -664
rect 506266 705564 506502 705800
rect 506586 705564 506822 705800
rect 506266 705244 506502 705480
rect 506586 705244 506822 705480
rect 506266 687660 506502 687896
rect 506586 687660 506822 687896
rect 506266 687340 506502 687576
rect 506586 687340 506822 687576
rect 506266 651660 506502 651896
rect 506586 651660 506822 651896
rect 506266 651340 506502 651576
rect 506586 651340 506822 651576
rect 506266 615660 506502 615896
rect 506586 615660 506822 615896
rect 506266 615340 506502 615576
rect 506586 615340 506822 615576
rect 506266 579660 506502 579896
rect 506586 579660 506822 579896
rect 506266 579340 506502 579576
rect 506586 579340 506822 579576
rect 506266 543660 506502 543896
rect 506586 543660 506822 543896
rect 506266 543340 506502 543576
rect 506586 543340 506822 543576
rect 506266 507660 506502 507896
rect 506586 507660 506822 507896
rect 506266 507340 506502 507576
rect 506586 507340 506822 507576
rect 506266 471660 506502 471896
rect 506586 471660 506822 471896
rect 506266 471340 506502 471576
rect 506586 471340 506822 471576
rect 506266 435660 506502 435896
rect 506586 435660 506822 435896
rect 506266 435340 506502 435576
rect 506586 435340 506822 435576
rect 506266 399660 506502 399896
rect 506586 399660 506822 399896
rect 506266 399340 506502 399576
rect 506586 399340 506822 399576
rect 506266 363660 506502 363896
rect 506586 363660 506822 363896
rect 506266 363340 506502 363576
rect 506586 363340 506822 363576
rect 506266 327660 506502 327896
rect 506586 327660 506822 327896
rect 506266 327340 506502 327576
rect 506586 327340 506822 327576
rect 506266 291660 506502 291896
rect 506586 291660 506822 291896
rect 506266 291340 506502 291576
rect 506586 291340 506822 291576
rect 506266 255660 506502 255896
rect 506586 255660 506822 255896
rect 506266 255340 506502 255576
rect 506586 255340 506822 255576
rect 506266 219660 506502 219896
rect 506586 219660 506822 219896
rect 506266 219340 506502 219576
rect 506586 219340 506822 219576
rect 506266 183660 506502 183896
rect 506586 183660 506822 183896
rect 506266 183340 506502 183576
rect 506586 183340 506822 183576
rect 506266 147660 506502 147896
rect 506586 147660 506822 147896
rect 506266 147340 506502 147576
rect 506586 147340 506822 147576
rect 506266 111660 506502 111896
rect 506586 111660 506822 111896
rect 506266 111340 506502 111576
rect 506586 111340 506822 111576
rect 506266 75660 506502 75896
rect 506586 75660 506822 75896
rect 506266 75340 506502 75576
rect 506586 75340 506822 75576
rect 506266 39660 506502 39896
rect 506586 39660 506822 39896
rect 506266 39340 506502 39576
rect 506586 39340 506822 39576
rect 506266 3660 506502 3896
rect 506586 3660 506822 3896
rect 506266 3340 506502 3576
rect 506586 3340 506822 3576
rect 506266 -1540 506502 -1304
rect 506586 -1540 506822 -1304
rect 506266 -1860 506502 -1624
rect 506586 -1860 506822 -1624
rect 507506 706524 507742 706760
rect 507826 706524 508062 706760
rect 507506 706204 507742 706440
rect 507826 706204 508062 706440
rect 507506 688900 507742 689136
rect 507826 688900 508062 689136
rect 507506 688580 507742 688816
rect 507826 688580 508062 688816
rect 507506 652900 507742 653136
rect 507826 652900 508062 653136
rect 507506 652580 507742 652816
rect 507826 652580 508062 652816
rect 507506 616900 507742 617136
rect 507826 616900 508062 617136
rect 507506 616580 507742 616816
rect 507826 616580 508062 616816
rect 507506 580900 507742 581136
rect 507826 580900 508062 581136
rect 507506 580580 507742 580816
rect 507826 580580 508062 580816
rect 507506 544900 507742 545136
rect 507826 544900 508062 545136
rect 507506 544580 507742 544816
rect 507826 544580 508062 544816
rect 507506 508900 507742 509136
rect 507826 508900 508062 509136
rect 507506 508580 507742 508816
rect 507826 508580 508062 508816
rect 507506 472900 507742 473136
rect 507826 472900 508062 473136
rect 507506 472580 507742 472816
rect 507826 472580 508062 472816
rect 507506 436900 507742 437136
rect 507826 436900 508062 437136
rect 507506 436580 507742 436816
rect 507826 436580 508062 436816
rect 507506 400900 507742 401136
rect 507826 400900 508062 401136
rect 507506 400580 507742 400816
rect 507826 400580 508062 400816
rect 507506 364900 507742 365136
rect 507826 364900 508062 365136
rect 507506 364580 507742 364816
rect 507826 364580 508062 364816
rect 507506 328900 507742 329136
rect 507826 328900 508062 329136
rect 507506 328580 507742 328816
rect 507826 328580 508062 328816
rect 507506 292900 507742 293136
rect 507826 292900 508062 293136
rect 507506 292580 507742 292816
rect 507826 292580 508062 292816
rect 507506 256900 507742 257136
rect 507826 256900 508062 257136
rect 507506 256580 507742 256816
rect 507826 256580 508062 256816
rect 507506 220900 507742 221136
rect 507826 220900 508062 221136
rect 507506 220580 507742 220816
rect 507826 220580 508062 220816
rect 507506 184900 507742 185136
rect 507826 184900 508062 185136
rect 507506 184580 507742 184816
rect 507826 184580 508062 184816
rect 507506 148900 507742 149136
rect 507826 148900 508062 149136
rect 507506 148580 507742 148816
rect 507826 148580 508062 148816
rect 507506 112900 507742 113136
rect 507826 112900 508062 113136
rect 507506 112580 507742 112816
rect 507826 112580 508062 112816
rect 507506 76900 507742 77136
rect 507826 76900 508062 77136
rect 507506 76580 507742 76816
rect 507826 76580 508062 76816
rect 507506 40900 507742 41136
rect 507826 40900 508062 41136
rect 507506 40580 507742 40816
rect 507826 40580 508062 40816
rect 507506 4900 507742 5136
rect 507826 4900 508062 5136
rect 507506 4580 507742 4816
rect 507826 4580 508062 4816
rect 507506 -2500 507742 -2264
rect 507826 -2500 508062 -2264
rect 507506 -2820 507742 -2584
rect 507826 -2820 508062 -2584
rect 508746 707484 508982 707720
rect 509066 707484 509302 707720
rect 508746 707164 508982 707400
rect 509066 707164 509302 707400
rect 508746 690140 508982 690376
rect 509066 690140 509302 690376
rect 508746 689820 508982 690056
rect 509066 689820 509302 690056
rect 508746 654140 508982 654376
rect 509066 654140 509302 654376
rect 508746 653820 508982 654056
rect 509066 653820 509302 654056
rect 508746 618140 508982 618376
rect 509066 618140 509302 618376
rect 508746 617820 508982 618056
rect 509066 617820 509302 618056
rect 508746 582140 508982 582376
rect 509066 582140 509302 582376
rect 508746 581820 508982 582056
rect 509066 581820 509302 582056
rect 508746 546140 508982 546376
rect 509066 546140 509302 546376
rect 508746 545820 508982 546056
rect 509066 545820 509302 546056
rect 508746 510140 508982 510376
rect 509066 510140 509302 510376
rect 508746 509820 508982 510056
rect 509066 509820 509302 510056
rect 508746 474140 508982 474376
rect 509066 474140 509302 474376
rect 508746 473820 508982 474056
rect 509066 473820 509302 474056
rect 508746 438140 508982 438376
rect 509066 438140 509302 438376
rect 508746 437820 508982 438056
rect 509066 437820 509302 438056
rect 508746 402140 508982 402376
rect 509066 402140 509302 402376
rect 508746 401820 508982 402056
rect 509066 401820 509302 402056
rect 508746 366140 508982 366376
rect 509066 366140 509302 366376
rect 508746 365820 508982 366056
rect 509066 365820 509302 366056
rect 508746 330140 508982 330376
rect 509066 330140 509302 330376
rect 508746 329820 508982 330056
rect 509066 329820 509302 330056
rect 508746 294140 508982 294376
rect 509066 294140 509302 294376
rect 508746 293820 508982 294056
rect 509066 293820 509302 294056
rect 508746 258140 508982 258376
rect 509066 258140 509302 258376
rect 508746 257820 508982 258056
rect 509066 257820 509302 258056
rect 508746 222140 508982 222376
rect 509066 222140 509302 222376
rect 508746 221820 508982 222056
rect 509066 221820 509302 222056
rect 508746 186140 508982 186376
rect 509066 186140 509302 186376
rect 508746 185820 508982 186056
rect 509066 185820 509302 186056
rect 508746 150140 508982 150376
rect 509066 150140 509302 150376
rect 508746 149820 508982 150056
rect 509066 149820 509302 150056
rect 508746 114140 508982 114376
rect 509066 114140 509302 114376
rect 508746 113820 508982 114056
rect 509066 113820 509302 114056
rect 508746 78140 508982 78376
rect 509066 78140 509302 78376
rect 508746 77820 508982 78056
rect 509066 77820 509302 78056
rect 508746 42140 508982 42376
rect 509066 42140 509302 42376
rect 508746 41820 508982 42056
rect 509066 41820 509302 42056
rect 508746 6140 508982 6376
rect 509066 6140 509302 6376
rect 508746 5820 508982 6056
rect 509066 5820 509302 6056
rect 508746 -3460 508982 -3224
rect 509066 -3460 509302 -3224
rect 508746 -3780 508982 -3544
rect 509066 -3780 509302 -3544
rect 509986 708444 510222 708680
rect 510306 708444 510542 708680
rect 509986 708124 510222 708360
rect 510306 708124 510542 708360
rect 509986 691380 510222 691616
rect 510306 691380 510542 691616
rect 509986 691060 510222 691296
rect 510306 691060 510542 691296
rect 509986 655380 510222 655616
rect 510306 655380 510542 655616
rect 509986 655060 510222 655296
rect 510306 655060 510542 655296
rect 509986 619380 510222 619616
rect 510306 619380 510542 619616
rect 509986 619060 510222 619296
rect 510306 619060 510542 619296
rect 509986 583380 510222 583616
rect 510306 583380 510542 583616
rect 509986 583060 510222 583296
rect 510306 583060 510542 583296
rect 509986 547380 510222 547616
rect 510306 547380 510542 547616
rect 509986 547060 510222 547296
rect 510306 547060 510542 547296
rect 509986 511380 510222 511616
rect 510306 511380 510542 511616
rect 509986 511060 510222 511296
rect 510306 511060 510542 511296
rect 509986 475380 510222 475616
rect 510306 475380 510542 475616
rect 509986 475060 510222 475296
rect 510306 475060 510542 475296
rect 509986 439380 510222 439616
rect 510306 439380 510542 439616
rect 509986 439060 510222 439296
rect 510306 439060 510542 439296
rect 509986 403380 510222 403616
rect 510306 403380 510542 403616
rect 509986 403060 510222 403296
rect 510306 403060 510542 403296
rect 509986 367380 510222 367616
rect 510306 367380 510542 367616
rect 509986 367060 510222 367296
rect 510306 367060 510542 367296
rect 509986 331380 510222 331616
rect 510306 331380 510542 331616
rect 509986 331060 510222 331296
rect 510306 331060 510542 331296
rect 509986 295380 510222 295616
rect 510306 295380 510542 295616
rect 509986 295060 510222 295296
rect 510306 295060 510542 295296
rect 509986 259380 510222 259616
rect 510306 259380 510542 259616
rect 509986 259060 510222 259296
rect 510306 259060 510542 259296
rect 509986 223380 510222 223616
rect 510306 223380 510542 223616
rect 509986 223060 510222 223296
rect 510306 223060 510542 223296
rect 509986 187380 510222 187616
rect 510306 187380 510542 187616
rect 509986 187060 510222 187296
rect 510306 187060 510542 187296
rect 509986 151380 510222 151616
rect 510306 151380 510542 151616
rect 509986 151060 510222 151296
rect 510306 151060 510542 151296
rect 509986 115380 510222 115616
rect 510306 115380 510542 115616
rect 509986 115060 510222 115296
rect 510306 115060 510542 115296
rect 509986 79380 510222 79616
rect 510306 79380 510542 79616
rect 509986 79060 510222 79296
rect 510306 79060 510542 79296
rect 509986 43380 510222 43616
rect 510306 43380 510542 43616
rect 509986 43060 510222 43296
rect 510306 43060 510542 43296
rect 509986 7380 510222 7616
rect 510306 7380 510542 7616
rect 509986 7060 510222 7296
rect 510306 7060 510542 7296
rect 509986 -4420 510222 -4184
rect 510306 -4420 510542 -4184
rect 509986 -4740 510222 -4504
rect 510306 -4740 510542 -4504
rect 511226 709404 511462 709640
rect 511546 709404 511782 709640
rect 511226 709084 511462 709320
rect 511546 709084 511782 709320
rect 511226 692620 511462 692856
rect 511546 692620 511782 692856
rect 511226 692300 511462 692536
rect 511546 692300 511782 692536
rect 511226 656620 511462 656856
rect 511546 656620 511782 656856
rect 511226 656300 511462 656536
rect 511546 656300 511782 656536
rect 511226 620620 511462 620856
rect 511546 620620 511782 620856
rect 511226 620300 511462 620536
rect 511546 620300 511782 620536
rect 511226 584620 511462 584856
rect 511546 584620 511782 584856
rect 511226 584300 511462 584536
rect 511546 584300 511782 584536
rect 511226 548620 511462 548856
rect 511546 548620 511782 548856
rect 511226 548300 511462 548536
rect 511546 548300 511782 548536
rect 511226 512620 511462 512856
rect 511546 512620 511782 512856
rect 511226 512300 511462 512536
rect 511546 512300 511782 512536
rect 511226 476620 511462 476856
rect 511546 476620 511782 476856
rect 511226 476300 511462 476536
rect 511546 476300 511782 476536
rect 511226 440620 511462 440856
rect 511546 440620 511782 440856
rect 511226 440300 511462 440536
rect 511546 440300 511782 440536
rect 511226 404620 511462 404856
rect 511546 404620 511782 404856
rect 511226 404300 511462 404536
rect 511546 404300 511782 404536
rect 511226 368620 511462 368856
rect 511546 368620 511782 368856
rect 511226 368300 511462 368536
rect 511546 368300 511782 368536
rect 511226 332620 511462 332856
rect 511546 332620 511782 332856
rect 511226 332300 511462 332536
rect 511546 332300 511782 332536
rect 511226 296620 511462 296856
rect 511546 296620 511782 296856
rect 511226 296300 511462 296536
rect 511546 296300 511782 296536
rect 511226 260620 511462 260856
rect 511546 260620 511782 260856
rect 511226 260300 511462 260536
rect 511546 260300 511782 260536
rect 511226 224620 511462 224856
rect 511546 224620 511782 224856
rect 511226 224300 511462 224536
rect 511546 224300 511782 224536
rect 511226 188620 511462 188856
rect 511546 188620 511782 188856
rect 511226 188300 511462 188536
rect 511546 188300 511782 188536
rect 511226 152620 511462 152856
rect 511546 152620 511782 152856
rect 511226 152300 511462 152536
rect 511546 152300 511782 152536
rect 511226 116620 511462 116856
rect 511546 116620 511782 116856
rect 511226 116300 511462 116536
rect 511546 116300 511782 116536
rect 511226 80620 511462 80856
rect 511546 80620 511782 80856
rect 511226 80300 511462 80536
rect 511546 80300 511782 80536
rect 511226 44620 511462 44856
rect 511546 44620 511782 44856
rect 511226 44300 511462 44536
rect 511546 44300 511782 44536
rect 511226 8620 511462 8856
rect 511546 8620 511782 8856
rect 511226 8300 511462 8536
rect 511546 8300 511782 8536
rect 511226 -5380 511462 -5144
rect 511546 -5380 511782 -5144
rect 511226 -5700 511462 -5464
rect 511546 -5700 511782 -5464
rect 512466 710364 512702 710600
rect 512786 710364 513022 710600
rect 512466 710044 512702 710280
rect 512786 710044 513022 710280
rect 512466 693860 512702 694096
rect 512786 693860 513022 694096
rect 512466 693540 512702 693776
rect 512786 693540 513022 693776
rect 512466 657860 512702 658096
rect 512786 657860 513022 658096
rect 512466 657540 512702 657776
rect 512786 657540 513022 657776
rect 512466 621860 512702 622096
rect 512786 621860 513022 622096
rect 512466 621540 512702 621776
rect 512786 621540 513022 621776
rect 512466 585860 512702 586096
rect 512786 585860 513022 586096
rect 512466 585540 512702 585776
rect 512786 585540 513022 585776
rect 512466 549860 512702 550096
rect 512786 549860 513022 550096
rect 512466 549540 512702 549776
rect 512786 549540 513022 549776
rect 512466 513860 512702 514096
rect 512786 513860 513022 514096
rect 512466 513540 512702 513776
rect 512786 513540 513022 513776
rect 512466 477860 512702 478096
rect 512786 477860 513022 478096
rect 512466 477540 512702 477776
rect 512786 477540 513022 477776
rect 512466 441860 512702 442096
rect 512786 441860 513022 442096
rect 512466 441540 512702 441776
rect 512786 441540 513022 441776
rect 512466 405860 512702 406096
rect 512786 405860 513022 406096
rect 512466 405540 512702 405776
rect 512786 405540 513022 405776
rect 512466 369860 512702 370096
rect 512786 369860 513022 370096
rect 512466 369540 512702 369776
rect 512786 369540 513022 369776
rect 512466 333860 512702 334096
rect 512786 333860 513022 334096
rect 512466 333540 512702 333776
rect 512786 333540 513022 333776
rect 512466 297860 512702 298096
rect 512786 297860 513022 298096
rect 512466 297540 512702 297776
rect 512786 297540 513022 297776
rect 512466 261860 512702 262096
rect 512786 261860 513022 262096
rect 512466 261540 512702 261776
rect 512786 261540 513022 261776
rect 512466 225860 512702 226096
rect 512786 225860 513022 226096
rect 512466 225540 512702 225776
rect 512786 225540 513022 225776
rect 512466 189860 512702 190096
rect 512786 189860 513022 190096
rect 512466 189540 512702 189776
rect 512786 189540 513022 189776
rect 512466 153860 512702 154096
rect 512786 153860 513022 154096
rect 512466 153540 512702 153776
rect 512786 153540 513022 153776
rect 512466 117860 512702 118096
rect 512786 117860 513022 118096
rect 512466 117540 512702 117776
rect 512786 117540 513022 117776
rect 512466 81860 512702 82096
rect 512786 81860 513022 82096
rect 512466 81540 512702 81776
rect 512786 81540 513022 81776
rect 512466 45860 512702 46096
rect 512786 45860 513022 46096
rect 512466 45540 512702 45776
rect 512786 45540 513022 45776
rect 512466 9860 512702 10096
rect 512786 9860 513022 10096
rect 512466 9540 512702 9776
rect 512786 9540 513022 9776
rect 512466 -6340 512702 -6104
rect 512786 -6340 513022 -6104
rect 512466 -6660 512702 -6424
rect 512786 -6660 513022 -6424
rect 513706 711324 513942 711560
rect 514026 711324 514262 711560
rect 513706 711004 513942 711240
rect 514026 711004 514262 711240
rect 513706 695100 513942 695336
rect 514026 695100 514262 695336
rect 513706 694780 513942 695016
rect 514026 694780 514262 695016
rect 513706 659100 513942 659336
rect 514026 659100 514262 659336
rect 513706 658780 513942 659016
rect 514026 658780 514262 659016
rect 513706 623100 513942 623336
rect 514026 623100 514262 623336
rect 513706 622780 513942 623016
rect 514026 622780 514262 623016
rect 513706 587100 513942 587336
rect 514026 587100 514262 587336
rect 513706 586780 513942 587016
rect 514026 586780 514262 587016
rect 513706 551100 513942 551336
rect 514026 551100 514262 551336
rect 513706 550780 513942 551016
rect 514026 550780 514262 551016
rect 513706 515100 513942 515336
rect 514026 515100 514262 515336
rect 513706 514780 513942 515016
rect 514026 514780 514262 515016
rect 513706 479100 513942 479336
rect 514026 479100 514262 479336
rect 513706 478780 513942 479016
rect 514026 478780 514262 479016
rect 541026 704604 541262 704840
rect 541346 704604 541582 704840
rect 541026 704284 541262 704520
rect 541346 704284 541582 704520
rect 541026 686420 541262 686656
rect 541346 686420 541582 686656
rect 541026 686100 541262 686336
rect 541346 686100 541582 686336
rect 541026 650420 541262 650656
rect 541346 650420 541582 650656
rect 541026 650100 541262 650336
rect 541346 650100 541582 650336
rect 541026 614420 541262 614656
rect 541346 614420 541582 614656
rect 541026 614100 541262 614336
rect 541346 614100 541582 614336
rect 541026 578420 541262 578656
rect 541346 578420 541582 578656
rect 541026 578100 541262 578336
rect 541346 578100 541582 578336
rect 541026 542420 541262 542656
rect 541346 542420 541582 542656
rect 541026 542100 541262 542336
rect 541346 542100 541582 542336
rect 541026 506420 541262 506656
rect 541346 506420 541582 506656
rect 541026 506100 541262 506336
rect 541346 506100 541582 506336
rect 541026 470420 541262 470656
rect 541346 470420 541582 470656
rect 541026 470100 541262 470336
rect 541346 470100 541582 470336
rect 542266 705564 542502 705800
rect 542586 705564 542822 705800
rect 542266 705244 542502 705480
rect 542586 705244 542822 705480
rect 542266 687660 542502 687896
rect 542586 687660 542822 687896
rect 542266 687340 542502 687576
rect 542586 687340 542822 687576
rect 542266 651660 542502 651896
rect 542586 651660 542822 651896
rect 542266 651340 542502 651576
rect 542586 651340 542822 651576
rect 542266 615660 542502 615896
rect 542586 615660 542822 615896
rect 542266 615340 542502 615576
rect 542586 615340 542822 615576
rect 542266 579660 542502 579896
rect 542586 579660 542822 579896
rect 542266 579340 542502 579576
rect 542586 579340 542822 579576
rect 542266 543660 542502 543896
rect 542586 543660 542822 543896
rect 542266 543340 542502 543576
rect 542586 543340 542822 543576
rect 542266 507660 542502 507896
rect 542586 507660 542822 507896
rect 542266 507340 542502 507576
rect 542586 507340 542822 507576
rect 542266 471660 542502 471896
rect 542586 471660 542822 471896
rect 542266 471340 542502 471576
rect 542586 471340 542822 471576
rect 543506 706524 543742 706760
rect 543826 706524 544062 706760
rect 543506 706204 543742 706440
rect 543826 706204 544062 706440
rect 543506 688900 543742 689136
rect 543826 688900 544062 689136
rect 543506 688580 543742 688816
rect 543826 688580 544062 688816
rect 543506 652900 543742 653136
rect 543826 652900 544062 653136
rect 543506 652580 543742 652816
rect 543826 652580 544062 652816
rect 543506 616900 543742 617136
rect 543826 616900 544062 617136
rect 543506 616580 543742 616816
rect 543826 616580 544062 616816
rect 543506 580900 543742 581136
rect 543826 580900 544062 581136
rect 543506 580580 543742 580816
rect 543826 580580 544062 580816
rect 543506 544900 543742 545136
rect 543826 544900 544062 545136
rect 543506 544580 543742 544816
rect 543826 544580 544062 544816
rect 543506 508900 543742 509136
rect 543826 508900 544062 509136
rect 543506 508580 543742 508816
rect 543826 508580 544062 508816
rect 543506 472900 543742 473136
rect 543826 472900 544062 473136
rect 543506 472580 543742 472816
rect 543826 472580 544062 472816
rect 544746 707484 544982 707720
rect 545066 707484 545302 707720
rect 544746 707164 544982 707400
rect 545066 707164 545302 707400
rect 544746 690140 544982 690376
rect 545066 690140 545302 690376
rect 544746 689820 544982 690056
rect 545066 689820 545302 690056
rect 544746 654140 544982 654376
rect 545066 654140 545302 654376
rect 544746 653820 544982 654056
rect 545066 653820 545302 654056
rect 544746 618140 544982 618376
rect 545066 618140 545302 618376
rect 544746 617820 544982 618056
rect 545066 617820 545302 618056
rect 544746 582140 544982 582376
rect 545066 582140 545302 582376
rect 544746 581820 544982 582056
rect 545066 581820 545302 582056
rect 544746 546140 544982 546376
rect 545066 546140 545302 546376
rect 544746 545820 544982 546056
rect 545066 545820 545302 546056
rect 544746 510140 544982 510376
rect 545066 510140 545302 510376
rect 544746 509820 544982 510056
rect 545066 509820 545302 510056
rect 544746 474140 544982 474376
rect 545066 474140 545302 474376
rect 544746 473820 544982 474056
rect 545066 473820 545302 474056
rect 513706 443100 513942 443336
rect 514026 443100 514262 443336
rect 513706 442780 513942 443016
rect 514026 442780 514262 443016
rect 540918 435660 541154 435896
rect 540918 435340 541154 435576
rect 539952 434420 540188 434656
rect 539952 434100 540188 434336
rect 542850 435660 543086 435896
rect 542850 435340 543086 435576
rect 541884 434420 542120 434656
rect 541884 434100 542120 434336
rect 543816 434420 544052 434656
rect 543816 434100 544052 434336
rect 545986 708444 546222 708680
rect 546306 708444 546542 708680
rect 545986 708124 546222 708360
rect 546306 708124 546542 708360
rect 545986 691380 546222 691616
rect 546306 691380 546542 691616
rect 545986 691060 546222 691296
rect 546306 691060 546542 691296
rect 545986 655380 546222 655616
rect 546306 655380 546542 655616
rect 545986 655060 546222 655296
rect 546306 655060 546542 655296
rect 545986 619380 546222 619616
rect 546306 619380 546542 619616
rect 545986 619060 546222 619296
rect 546306 619060 546542 619296
rect 545986 583380 546222 583616
rect 546306 583380 546542 583616
rect 545986 583060 546222 583296
rect 546306 583060 546542 583296
rect 545986 547380 546222 547616
rect 546306 547380 546542 547616
rect 545986 547060 546222 547296
rect 546306 547060 546542 547296
rect 545986 511380 546222 511616
rect 546306 511380 546542 511616
rect 545986 511060 546222 511296
rect 546306 511060 546542 511296
rect 545986 475380 546222 475616
rect 546306 475380 546542 475616
rect 545986 475060 546222 475296
rect 546306 475060 546542 475296
rect 547226 709404 547462 709640
rect 547546 709404 547782 709640
rect 547226 709084 547462 709320
rect 547546 709084 547782 709320
rect 547226 692620 547462 692856
rect 547546 692620 547782 692856
rect 547226 692300 547462 692536
rect 547546 692300 547782 692536
rect 547226 656620 547462 656856
rect 547546 656620 547782 656856
rect 547226 656300 547462 656536
rect 547546 656300 547782 656536
rect 547226 620620 547462 620856
rect 547546 620620 547782 620856
rect 547226 620300 547462 620536
rect 547546 620300 547782 620536
rect 547226 584620 547462 584856
rect 547546 584620 547782 584856
rect 547226 584300 547462 584536
rect 547546 584300 547782 584536
rect 547226 548620 547462 548856
rect 547546 548620 547782 548856
rect 547226 548300 547462 548536
rect 547546 548300 547782 548536
rect 547226 512620 547462 512856
rect 547546 512620 547782 512856
rect 547226 512300 547462 512536
rect 547546 512300 547782 512536
rect 547226 476620 547462 476856
rect 547546 476620 547782 476856
rect 547226 476300 547462 476536
rect 547546 476300 547782 476536
rect 547226 440620 547462 440856
rect 547546 440620 547782 440856
rect 547226 440300 547462 440536
rect 547546 440300 547782 440536
rect 544782 435660 545018 435896
rect 544782 435340 545018 435576
rect 546714 435660 546950 435896
rect 546714 435340 546950 435576
rect 545748 434420 545984 434656
rect 545748 434100 545984 434336
rect 513706 407100 513942 407336
rect 514026 407100 514262 407336
rect 513706 406780 513942 407016
rect 514026 406780 514262 407016
rect 540918 399660 541154 399896
rect 540918 399340 541154 399576
rect 539952 398420 540188 398656
rect 539952 398100 540188 398336
rect 542850 399660 543086 399896
rect 542850 399340 543086 399576
rect 541884 398420 542120 398656
rect 541884 398100 542120 398336
rect 543816 398420 544052 398656
rect 543816 398100 544052 398336
rect 547226 404620 547462 404856
rect 547546 404620 547782 404856
rect 547226 404300 547462 404536
rect 547546 404300 547782 404536
rect 544782 399660 545018 399896
rect 544782 399340 545018 399576
rect 546714 399660 546950 399896
rect 546714 399340 546950 399576
rect 545748 398420 545984 398656
rect 545748 398100 545984 398336
rect 513706 371100 513942 371336
rect 514026 371100 514262 371336
rect 513706 370780 513942 371016
rect 514026 370780 514262 371016
rect 540918 363660 541154 363896
rect 540918 363340 541154 363576
rect 539952 362420 540188 362656
rect 539952 362100 540188 362336
rect 542850 363660 543086 363896
rect 542850 363340 543086 363576
rect 541884 362420 542120 362656
rect 541884 362100 542120 362336
rect 543816 362420 544052 362656
rect 543816 362100 544052 362336
rect 547226 368620 547462 368856
rect 547546 368620 547782 368856
rect 547226 368300 547462 368536
rect 547546 368300 547782 368536
rect 544782 363660 545018 363896
rect 544782 363340 545018 363576
rect 546714 363660 546950 363896
rect 546714 363340 546950 363576
rect 545748 362420 545984 362656
rect 545748 362100 545984 362336
rect 513706 335100 513942 335336
rect 514026 335100 514262 335336
rect 513706 334780 513942 335016
rect 514026 334780 514262 335016
rect 540918 327660 541154 327896
rect 540918 327340 541154 327576
rect 539952 326420 540188 326656
rect 539952 326100 540188 326336
rect 542850 327660 543086 327896
rect 542850 327340 543086 327576
rect 541884 326420 542120 326656
rect 541884 326100 542120 326336
rect 543816 326420 544052 326656
rect 543816 326100 544052 326336
rect 547226 332620 547462 332856
rect 547546 332620 547782 332856
rect 547226 332300 547462 332536
rect 547546 332300 547782 332536
rect 544782 327660 545018 327896
rect 544782 327340 545018 327576
rect 546714 327660 546950 327896
rect 546714 327340 546950 327576
rect 545748 326420 545984 326656
rect 545748 326100 545984 326336
rect 513706 299100 513942 299336
rect 514026 299100 514262 299336
rect 513706 298780 513942 299016
rect 514026 298780 514262 299016
rect 547226 296620 547462 296856
rect 547546 296620 547782 296856
rect 547226 296300 547462 296536
rect 547546 296300 547782 296536
rect 540918 291660 541154 291896
rect 540918 291340 541154 291576
rect 542850 291660 543086 291896
rect 542850 291340 543086 291576
rect 544782 291660 545018 291896
rect 544782 291340 545018 291576
rect 546714 291660 546950 291896
rect 546714 291340 546950 291576
rect 539952 290420 540188 290656
rect 539952 290100 540188 290336
rect 541884 290420 542120 290656
rect 541884 290100 542120 290336
rect 543816 290420 544052 290656
rect 543816 290100 544052 290336
rect 545748 290420 545984 290656
rect 545748 290100 545984 290336
rect 513706 263100 513942 263336
rect 514026 263100 514262 263336
rect 513706 262780 513942 263016
rect 514026 262780 514262 263016
rect 513706 227100 513942 227336
rect 514026 227100 514262 227336
rect 513706 226780 513942 227016
rect 514026 226780 514262 227016
rect 513706 191100 513942 191336
rect 514026 191100 514262 191336
rect 513706 190780 513942 191016
rect 514026 190780 514262 191016
rect 513706 155100 513942 155336
rect 514026 155100 514262 155336
rect 513706 154780 513942 155016
rect 514026 154780 514262 155016
rect 513706 119100 513942 119336
rect 514026 119100 514262 119336
rect 513706 118780 513942 119016
rect 514026 118780 514262 119016
rect 513706 83100 513942 83336
rect 514026 83100 514262 83336
rect 513706 82780 513942 83016
rect 514026 82780 514262 83016
rect 513706 47100 513942 47336
rect 514026 47100 514262 47336
rect 513706 46780 513942 47016
rect 514026 46780 514262 47016
rect 513706 11100 513942 11336
rect 514026 11100 514262 11336
rect 513706 10780 513942 11016
rect 514026 10780 514262 11016
rect 513706 -7300 513942 -7064
rect 514026 -7300 514262 -7064
rect 513706 -7620 513942 -7384
rect 514026 -7620 514262 -7384
rect 541026 254420 541262 254656
rect 541346 254420 541582 254656
rect 541026 254100 541262 254336
rect 541346 254100 541582 254336
rect 541026 218420 541262 218656
rect 541346 218420 541582 218656
rect 541026 218100 541262 218336
rect 541346 218100 541582 218336
rect 541026 182420 541262 182656
rect 541346 182420 541582 182656
rect 541026 182100 541262 182336
rect 541346 182100 541582 182336
rect 541026 146420 541262 146656
rect 541346 146420 541582 146656
rect 541026 146100 541262 146336
rect 541346 146100 541582 146336
rect 541026 110420 541262 110656
rect 541346 110420 541582 110656
rect 541026 110100 541262 110336
rect 541346 110100 541582 110336
rect 541026 74420 541262 74656
rect 541346 74420 541582 74656
rect 541026 74100 541262 74336
rect 541346 74100 541582 74336
rect 541026 38420 541262 38656
rect 541346 38420 541582 38656
rect 541026 38100 541262 38336
rect 541346 38100 541582 38336
rect 541026 2420 541262 2656
rect 541346 2420 541582 2656
rect 541026 2100 541262 2336
rect 541346 2100 541582 2336
rect 541026 -580 541262 -344
rect 541346 -580 541582 -344
rect 541026 -900 541262 -664
rect 541346 -900 541582 -664
rect 542266 255660 542502 255896
rect 542586 255660 542822 255896
rect 542266 255340 542502 255576
rect 542586 255340 542822 255576
rect 542266 219660 542502 219896
rect 542586 219660 542822 219896
rect 542266 219340 542502 219576
rect 542586 219340 542822 219576
rect 542266 183660 542502 183896
rect 542586 183660 542822 183896
rect 542266 183340 542502 183576
rect 542586 183340 542822 183576
rect 542266 147660 542502 147896
rect 542586 147660 542822 147896
rect 542266 147340 542502 147576
rect 542586 147340 542822 147576
rect 542266 111660 542502 111896
rect 542586 111660 542822 111896
rect 542266 111340 542502 111576
rect 542586 111340 542822 111576
rect 542266 75660 542502 75896
rect 542586 75660 542822 75896
rect 542266 75340 542502 75576
rect 542586 75340 542822 75576
rect 542266 39660 542502 39896
rect 542586 39660 542822 39896
rect 542266 39340 542502 39576
rect 542586 39340 542822 39576
rect 542266 3660 542502 3896
rect 542586 3660 542822 3896
rect 542266 3340 542502 3576
rect 542586 3340 542822 3576
rect 542266 -1540 542502 -1304
rect 542586 -1540 542822 -1304
rect 542266 -1860 542502 -1624
rect 542586 -1860 542822 -1624
rect 543506 256900 543742 257136
rect 543826 256900 544062 257136
rect 543506 256580 543742 256816
rect 543826 256580 544062 256816
rect 543506 220900 543742 221136
rect 543826 220900 544062 221136
rect 543506 220580 543742 220816
rect 543826 220580 544062 220816
rect 543506 184900 543742 185136
rect 543826 184900 544062 185136
rect 543506 184580 543742 184816
rect 543826 184580 544062 184816
rect 543506 148900 543742 149136
rect 543826 148900 544062 149136
rect 543506 148580 543742 148816
rect 543826 148580 544062 148816
rect 543506 112900 543742 113136
rect 543826 112900 544062 113136
rect 543506 112580 543742 112816
rect 543826 112580 544062 112816
rect 543506 76900 543742 77136
rect 543826 76900 544062 77136
rect 543506 76580 543742 76816
rect 543826 76580 544062 76816
rect 543506 40900 543742 41136
rect 543826 40900 544062 41136
rect 543506 40580 543742 40816
rect 543826 40580 544062 40816
rect 543506 4900 543742 5136
rect 543826 4900 544062 5136
rect 543506 4580 543742 4816
rect 543826 4580 544062 4816
rect 543506 -2500 543742 -2264
rect 543826 -2500 544062 -2264
rect 543506 -2820 543742 -2584
rect 543826 -2820 544062 -2584
rect 544746 258140 544982 258376
rect 545066 258140 545302 258376
rect 544746 257820 544982 258056
rect 545066 257820 545302 258056
rect 544746 222140 544982 222376
rect 545066 222140 545302 222376
rect 544746 221820 544982 222056
rect 545066 221820 545302 222056
rect 544746 186140 544982 186376
rect 545066 186140 545302 186376
rect 544746 185820 544982 186056
rect 545066 185820 545302 186056
rect 544746 150140 544982 150376
rect 545066 150140 545302 150376
rect 544746 149820 544982 150056
rect 545066 149820 545302 150056
rect 544746 114140 544982 114376
rect 545066 114140 545302 114376
rect 544746 113820 544982 114056
rect 545066 113820 545302 114056
rect 544746 78140 544982 78376
rect 545066 78140 545302 78376
rect 544746 77820 544982 78056
rect 545066 77820 545302 78056
rect 544746 42140 544982 42376
rect 545066 42140 545302 42376
rect 544746 41820 544982 42056
rect 545066 41820 545302 42056
rect 544746 6140 544982 6376
rect 545066 6140 545302 6376
rect 544746 5820 544982 6056
rect 545066 5820 545302 6056
rect 544746 -3460 544982 -3224
rect 545066 -3460 545302 -3224
rect 544746 -3780 544982 -3544
rect 545066 -3780 545302 -3544
rect 545986 259380 546222 259616
rect 546306 259380 546542 259616
rect 545986 259060 546222 259296
rect 546306 259060 546542 259296
rect 545986 223380 546222 223616
rect 546306 223380 546542 223616
rect 545986 223060 546222 223296
rect 546306 223060 546542 223296
rect 545986 187380 546222 187616
rect 546306 187380 546542 187616
rect 545986 187060 546222 187296
rect 546306 187060 546542 187296
rect 545986 151380 546222 151616
rect 546306 151380 546542 151616
rect 545986 151060 546222 151296
rect 546306 151060 546542 151296
rect 545986 115380 546222 115616
rect 546306 115380 546542 115616
rect 545986 115060 546222 115296
rect 546306 115060 546542 115296
rect 545986 79380 546222 79616
rect 546306 79380 546542 79616
rect 545986 79060 546222 79296
rect 546306 79060 546542 79296
rect 545986 43380 546222 43616
rect 546306 43380 546542 43616
rect 545986 43060 546222 43296
rect 546306 43060 546542 43296
rect 545986 7380 546222 7616
rect 546306 7380 546542 7616
rect 545986 7060 546222 7296
rect 546306 7060 546542 7296
rect 545986 -4420 546222 -4184
rect 546306 -4420 546542 -4184
rect 545986 -4740 546222 -4504
rect 546306 -4740 546542 -4504
rect 547226 260620 547462 260856
rect 547546 260620 547782 260856
rect 547226 260300 547462 260536
rect 547546 260300 547782 260536
rect 547226 224620 547462 224856
rect 547546 224620 547782 224856
rect 547226 224300 547462 224536
rect 547546 224300 547782 224536
rect 547226 188620 547462 188856
rect 547546 188620 547782 188856
rect 547226 188300 547462 188536
rect 547546 188300 547782 188536
rect 547226 152620 547462 152856
rect 547546 152620 547782 152856
rect 547226 152300 547462 152536
rect 547546 152300 547782 152536
rect 547226 116620 547462 116856
rect 547546 116620 547782 116856
rect 547226 116300 547462 116536
rect 547546 116300 547782 116536
rect 547226 80620 547462 80856
rect 547546 80620 547782 80856
rect 547226 80300 547462 80536
rect 547546 80300 547782 80536
rect 547226 44620 547462 44856
rect 547546 44620 547782 44856
rect 547226 44300 547462 44536
rect 547546 44300 547782 44536
rect 547226 8620 547462 8856
rect 547546 8620 547782 8856
rect 547226 8300 547462 8536
rect 547546 8300 547782 8536
rect 547226 -5380 547462 -5144
rect 547546 -5380 547782 -5144
rect 547226 -5700 547462 -5464
rect 547546 -5700 547782 -5464
rect 548466 710364 548702 710600
rect 548786 710364 549022 710600
rect 548466 710044 548702 710280
rect 548786 710044 549022 710280
rect 548466 693860 548702 694096
rect 548786 693860 549022 694096
rect 548466 693540 548702 693776
rect 548786 693540 549022 693776
rect 548466 657860 548702 658096
rect 548786 657860 549022 658096
rect 548466 657540 548702 657776
rect 548786 657540 549022 657776
rect 548466 621860 548702 622096
rect 548786 621860 549022 622096
rect 548466 621540 548702 621776
rect 548786 621540 549022 621776
rect 548466 585860 548702 586096
rect 548786 585860 549022 586096
rect 548466 585540 548702 585776
rect 548786 585540 549022 585776
rect 548466 549860 548702 550096
rect 548786 549860 549022 550096
rect 548466 549540 548702 549776
rect 548786 549540 549022 549776
rect 548466 513860 548702 514096
rect 548786 513860 549022 514096
rect 548466 513540 548702 513776
rect 548786 513540 549022 513776
rect 548466 477860 548702 478096
rect 548786 477860 549022 478096
rect 548466 477540 548702 477776
rect 548786 477540 549022 477776
rect 548466 441860 548702 442096
rect 548786 441860 549022 442096
rect 548466 441540 548702 441776
rect 548786 441540 549022 441776
rect 548466 405860 548702 406096
rect 548786 405860 549022 406096
rect 548466 405540 548702 405776
rect 548786 405540 549022 405776
rect 548466 369860 548702 370096
rect 548786 369860 549022 370096
rect 548466 369540 548702 369776
rect 548786 369540 549022 369776
rect 548466 333860 548702 334096
rect 548786 333860 549022 334096
rect 548466 333540 548702 333776
rect 548786 333540 549022 333776
rect 548466 297860 548702 298096
rect 548786 297860 549022 298096
rect 548466 297540 548702 297776
rect 548786 297540 549022 297776
rect 548466 261860 548702 262096
rect 548786 261860 549022 262096
rect 548466 261540 548702 261776
rect 548786 261540 549022 261776
rect 548466 225860 548702 226096
rect 548786 225860 549022 226096
rect 548466 225540 548702 225776
rect 548786 225540 549022 225776
rect 548466 189860 548702 190096
rect 548786 189860 549022 190096
rect 548466 189540 548702 189776
rect 548786 189540 549022 189776
rect 548466 153860 548702 154096
rect 548786 153860 549022 154096
rect 548466 153540 548702 153776
rect 548786 153540 549022 153776
rect 548466 117860 548702 118096
rect 548786 117860 549022 118096
rect 548466 117540 548702 117776
rect 548786 117540 549022 117776
rect 548466 81860 548702 82096
rect 548786 81860 549022 82096
rect 548466 81540 548702 81776
rect 548786 81540 549022 81776
rect 548466 45860 548702 46096
rect 548786 45860 549022 46096
rect 548466 45540 548702 45776
rect 548786 45540 549022 45776
rect 548466 9860 548702 10096
rect 548786 9860 549022 10096
rect 548466 9540 548702 9776
rect 548786 9540 549022 9776
rect 548466 -6340 548702 -6104
rect 548786 -6340 549022 -6104
rect 548466 -6660 548702 -6424
rect 548786 -6660 549022 -6424
rect 549706 711324 549942 711560
rect 550026 711324 550262 711560
rect 549706 711004 549942 711240
rect 550026 711004 550262 711240
rect 549706 695100 549942 695336
rect 550026 695100 550262 695336
rect 549706 694780 549942 695016
rect 550026 694780 550262 695016
rect 549706 659100 549942 659336
rect 550026 659100 550262 659336
rect 549706 658780 549942 659016
rect 550026 658780 550262 659016
rect 549706 623100 549942 623336
rect 550026 623100 550262 623336
rect 549706 622780 549942 623016
rect 550026 622780 550262 623016
rect 549706 587100 549942 587336
rect 550026 587100 550262 587336
rect 549706 586780 549942 587016
rect 550026 586780 550262 587016
rect 549706 551100 549942 551336
rect 550026 551100 550262 551336
rect 549706 550780 549942 551016
rect 550026 550780 550262 551016
rect 549706 515100 549942 515336
rect 550026 515100 550262 515336
rect 549706 514780 549942 515016
rect 550026 514780 550262 515016
rect 549706 479100 549942 479336
rect 550026 479100 550262 479336
rect 549706 478780 549942 479016
rect 550026 478780 550262 479016
rect 549706 443100 549942 443336
rect 550026 443100 550262 443336
rect 549706 442780 549942 443016
rect 550026 442780 550262 443016
rect 549706 407100 549942 407336
rect 550026 407100 550262 407336
rect 549706 406780 549942 407016
rect 550026 406780 550262 407016
rect 549706 371100 549942 371336
rect 550026 371100 550262 371336
rect 549706 370780 549942 371016
rect 550026 370780 550262 371016
rect 549706 335100 549942 335336
rect 550026 335100 550262 335336
rect 549706 334780 549942 335016
rect 550026 334780 550262 335016
rect 549706 299100 549942 299336
rect 550026 299100 550262 299336
rect 549706 298780 549942 299016
rect 550026 298780 550262 299016
rect 549706 263100 549942 263336
rect 550026 263100 550262 263336
rect 549706 262780 549942 263016
rect 550026 262780 550262 263016
rect 549706 227100 549942 227336
rect 550026 227100 550262 227336
rect 549706 226780 549942 227016
rect 550026 226780 550262 227016
rect 549706 191100 549942 191336
rect 550026 191100 550262 191336
rect 549706 190780 549942 191016
rect 550026 190780 550262 191016
rect 549706 155100 549942 155336
rect 550026 155100 550262 155336
rect 549706 154780 549942 155016
rect 550026 154780 550262 155016
rect 549706 119100 549942 119336
rect 550026 119100 550262 119336
rect 549706 118780 549942 119016
rect 550026 118780 550262 119016
rect 549706 83100 549942 83336
rect 550026 83100 550262 83336
rect 549706 82780 549942 83016
rect 550026 82780 550262 83016
rect 549706 47100 549942 47336
rect 550026 47100 550262 47336
rect 549706 46780 549942 47016
rect 550026 46780 550262 47016
rect 549706 11100 549942 11336
rect 550026 11100 550262 11336
rect 549706 10780 549942 11016
rect 550026 10780 550262 11016
rect 549706 -7300 549942 -7064
rect 550026 -7300 550262 -7064
rect 549706 -7620 549942 -7384
rect 550026 -7620 550262 -7384
rect 577026 704604 577262 704840
rect 577346 704604 577582 704840
rect 577026 704284 577262 704520
rect 577346 704284 577582 704520
rect 577026 686420 577262 686656
rect 577346 686420 577582 686656
rect 577026 686100 577262 686336
rect 577346 686100 577582 686336
rect 577026 650420 577262 650656
rect 577346 650420 577582 650656
rect 577026 650100 577262 650336
rect 577346 650100 577582 650336
rect 577026 614420 577262 614656
rect 577346 614420 577582 614656
rect 577026 614100 577262 614336
rect 577346 614100 577582 614336
rect 577026 578420 577262 578656
rect 577346 578420 577582 578656
rect 577026 578100 577262 578336
rect 577346 578100 577582 578336
rect 577026 542420 577262 542656
rect 577346 542420 577582 542656
rect 577026 542100 577262 542336
rect 577346 542100 577582 542336
rect 577026 506420 577262 506656
rect 577346 506420 577582 506656
rect 577026 506100 577262 506336
rect 577346 506100 577582 506336
rect 577026 470420 577262 470656
rect 577346 470420 577582 470656
rect 577026 470100 577262 470336
rect 577346 470100 577582 470336
rect 577026 434420 577262 434656
rect 577346 434420 577582 434656
rect 577026 434100 577262 434336
rect 577346 434100 577582 434336
rect 577026 398420 577262 398656
rect 577346 398420 577582 398656
rect 577026 398100 577262 398336
rect 577346 398100 577582 398336
rect 577026 362420 577262 362656
rect 577346 362420 577582 362656
rect 577026 362100 577262 362336
rect 577346 362100 577582 362336
rect 577026 326420 577262 326656
rect 577346 326420 577582 326656
rect 577026 326100 577262 326336
rect 577346 326100 577582 326336
rect 577026 290420 577262 290656
rect 577346 290420 577582 290656
rect 577026 290100 577262 290336
rect 577346 290100 577582 290336
rect 577026 254420 577262 254656
rect 577346 254420 577582 254656
rect 577026 254100 577262 254336
rect 577346 254100 577582 254336
rect 577026 218420 577262 218656
rect 577346 218420 577582 218656
rect 577026 218100 577262 218336
rect 577346 218100 577582 218336
rect 577026 182420 577262 182656
rect 577346 182420 577582 182656
rect 577026 182100 577262 182336
rect 577346 182100 577582 182336
rect 577026 146420 577262 146656
rect 577346 146420 577582 146656
rect 577026 146100 577262 146336
rect 577346 146100 577582 146336
rect 577026 110420 577262 110656
rect 577346 110420 577582 110656
rect 577026 110100 577262 110336
rect 577346 110100 577582 110336
rect 577026 74420 577262 74656
rect 577346 74420 577582 74656
rect 577026 74100 577262 74336
rect 577346 74100 577582 74336
rect 577026 38420 577262 38656
rect 577346 38420 577582 38656
rect 577026 38100 577262 38336
rect 577346 38100 577582 38336
rect 577026 2420 577262 2656
rect 577346 2420 577582 2656
rect 577026 2100 577262 2336
rect 577346 2100 577582 2336
rect 577026 -580 577262 -344
rect 577346 -580 577582 -344
rect 577026 -900 577262 -664
rect 577346 -900 577582 -664
rect 578266 705564 578502 705800
rect 578586 705564 578822 705800
rect 578266 705244 578502 705480
rect 578586 705244 578822 705480
rect 578266 687660 578502 687896
rect 578586 687660 578822 687896
rect 578266 687340 578502 687576
rect 578586 687340 578822 687576
rect 578266 651660 578502 651896
rect 578586 651660 578822 651896
rect 578266 651340 578502 651576
rect 578586 651340 578822 651576
rect 578266 615660 578502 615896
rect 578586 615660 578822 615896
rect 578266 615340 578502 615576
rect 578586 615340 578822 615576
rect 578266 579660 578502 579896
rect 578586 579660 578822 579896
rect 578266 579340 578502 579576
rect 578586 579340 578822 579576
rect 578266 543660 578502 543896
rect 578586 543660 578822 543896
rect 578266 543340 578502 543576
rect 578586 543340 578822 543576
rect 578266 507660 578502 507896
rect 578586 507660 578822 507896
rect 578266 507340 578502 507576
rect 578586 507340 578822 507576
rect 578266 471660 578502 471896
rect 578586 471660 578822 471896
rect 578266 471340 578502 471576
rect 578586 471340 578822 471576
rect 578266 435660 578502 435896
rect 578586 435660 578822 435896
rect 578266 435340 578502 435576
rect 578586 435340 578822 435576
rect 578266 399660 578502 399896
rect 578586 399660 578822 399896
rect 578266 399340 578502 399576
rect 578586 399340 578822 399576
rect 578266 363660 578502 363896
rect 578586 363660 578822 363896
rect 578266 363340 578502 363576
rect 578586 363340 578822 363576
rect 578266 327660 578502 327896
rect 578586 327660 578822 327896
rect 578266 327340 578502 327576
rect 578586 327340 578822 327576
rect 578266 291660 578502 291896
rect 578586 291660 578822 291896
rect 578266 291340 578502 291576
rect 578586 291340 578822 291576
rect 578266 255660 578502 255896
rect 578586 255660 578822 255896
rect 578266 255340 578502 255576
rect 578586 255340 578822 255576
rect 578266 219660 578502 219896
rect 578586 219660 578822 219896
rect 578266 219340 578502 219576
rect 578586 219340 578822 219576
rect 578266 183660 578502 183896
rect 578586 183660 578822 183896
rect 578266 183340 578502 183576
rect 578586 183340 578822 183576
rect 578266 147660 578502 147896
rect 578586 147660 578822 147896
rect 578266 147340 578502 147576
rect 578586 147340 578822 147576
rect 578266 111660 578502 111896
rect 578586 111660 578822 111896
rect 578266 111340 578502 111576
rect 578586 111340 578822 111576
rect 578266 75660 578502 75896
rect 578586 75660 578822 75896
rect 578266 75340 578502 75576
rect 578586 75340 578822 75576
rect 578266 39660 578502 39896
rect 578586 39660 578822 39896
rect 578266 39340 578502 39576
rect 578586 39340 578822 39576
rect 578266 3660 578502 3896
rect 578586 3660 578822 3896
rect 578266 3340 578502 3576
rect 578586 3340 578822 3576
rect 578266 -1540 578502 -1304
rect 578586 -1540 578822 -1304
rect 578266 -1860 578502 -1624
rect 578586 -1860 578822 -1624
rect 579506 706524 579742 706760
rect 579826 706524 580062 706760
rect 579506 706204 579742 706440
rect 579826 706204 580062 706440
rect 579506 688900 579742 689136
rect 579826 688900 580062 689136
rect 579506 688580 579742 688816
rect 579826 688580 580062 688816
rect 579506 652900 579742 653136
rect 579826 652900 580062 653136
rect 579506 652580 579742 652816
rect 579826 652580 580062 652816
rect 579506 616900 579742 617136
rect 579826 616900 580062 617136
rect 579506 616580 579742 616816
rect 579826 616580 580062 616816
rect 579506 580900 579742 581136
rect 579826 580900 580062 581136
rect 579506 580580 579742 580816
rect 579826 580580 580062 580816
rect 579506 544900 579742 545136
rect 579826 544900 580062 545136
rect 579506 544580 579742 544816
rect 579826 544580 580062 544816
rect 579506 508900 579742 509136
rect 579826 508900 580062 509136
rect 579506 508580 579742 508816
rect 579826 508580 580062 508816
rect 579506 472900 579742 473136
rect 579826 472900 580062 473136
rect 579506 472580 579742 472816
rect 579826 472580 580062 472816
rect 579506 436900 579742 437136
rect 579826 436900 580062 437136
rect 579506 436580 579742 436816
rect 579826 436580 580062 436816
rect 579506 400900 579742 401136
rect 579826 400900 580062 401136
rect 579506 400580 579742 400816
rect 579826 400580 580062 400816
rect 579506 364900 579742 365136
rect 579826 364900 580062 365136
rect 579506 364580 579742 364816
rect 579826 364580 580062 364816
rect 579506 328900 579742 329136
rect 579826 328900 580062 329136
rect 579506 328580 579742 328816
rect 579826 328580 580062 328816
rect 579506 292900 579742 293136
rect 579826 292900 580062 293136
rect 579506 292580 579742 292816
rect 579826 292580 580062 292816
rect 579506 256900 579742 257136
rect 579826 256900 580062 257136
rect 579506 256580 579742 256816
rect 579826 256580 580062 256816
rect 579506 220900 579742 221136
rect 579826 220900 580062 221136
rect 579506 220580 579742 220816
rect 579826 220580 580062 220816
rect 579506 184900 579742 185136
rect 579826 184900 580062 185136
rect 579506 184580 579742 184816
rect 579826 184580 580062 184816
rect 579506 148900 579742 149136
rect 579826 148900 580062 149136
rect 579506 148580 579742 148816
rect 579826 148580 580062 148816
rect 579506 112900 579742 113136
rect 579826 112900 580062 113136
rect 579506 112580 579742 112816
rect 579826 112580 580062 112816
rect 579506 76900 579742 77136
rect 579826 76900 580062 77136
rect 579506 76580 579742 76816
rect 579826 76580 580062 76816
rect 579506 40900 579742 41136
rect 579826 40900 580062 41136
rect 579506 40580 579742 40816
rect 579826 40580 580062 40816
rect 579506 4900 579742 5136
rect 579826 4900 580062 5136
rect 579506 4580 579742 4816
rect 579826 4580 580062 4816
rect 579506 -2500 579742 -2264
rect 579826 -2500 580062 -2264
rect 579506 -2820 579742 -2584
rect 579826 -2820 580062 -2584
rect 580746 707484 580982 707720
rect 581066 707484 581302 707720
rect 580746 707164 580982 707400
rect 581066 707164 581302 707400
rect 580746 690140 580982 690376
rect 581066 690140 581302 690376
rect 580746 689820 580982 690056
rect 581066 689820 581302 690056
rect 580746 654140 580982 654376
rect 581066 654140 581302 654376
rect 580746 653820 580982 654056
rect 581066 653820 581302 654056
rect 580746 618140 580982 618376
rect 581066 618140 581302 618376
rect 580746 617820 580982 618056
rect 581066 617820 581302 618056
rect 580746 582140 580982 582376
rect 581066 582140 581302 582376
rect 580746 581820 580982 582056
rect 581066 581820 581302 582056
rect 580746 546140 580982 546376
rect 581066 546140 581302 546376
rect 580746 545820 580982 546056
rect 581066 545820 581302 546056
rect 580746 510140 580982 510376
rect 581066 510140 581302 510376
rect 580746 509820 580982 510056
rect 581066 509820 581302 510056
rect 580746 474140 580982 474376
rect 581066 474140 581302 474376
rect 580746 473820 580982 474056
rect 581066 473820 581302 474056
rect 580746 438140 580982 438376
rect 581066 438140 581302 438376
rect 580746 437820 580982 438056
rect 581066 437820 581302 438056
rect 580746 402140 580982 402376
rect 581066 402140 581302 402376
rect 580746 401820 580982 402056
rect 581066 401820 581302 402056
rect 580746 366140 580982 366376
rect 581066 366140 581302 366376
rect 580746 365820 580982 366056
rect 581066 365820 581302 366056
rect 580746 330140 580982 330376
rect 581066 330140 581302 330376
rect 580746 329820 580982 330056
rect 581066 329820 581302 330056
rect 580746 294140 580982 294376
rect 581066 294140 581302 294376
rect 580746 293820 580982 294056
rect 581066 293820 581302 294056
rect 580746 258140 580982 258376
rect 581066 258140 581302 258376
rect 580746 257820 580982 258056
rect 581066 257820 581302 258056
rect 580746 222140 580982 222376
rect 581066 222140 581302 222376
rect 580746 221820 580982 222056
rect 581066 221820 581302 222056
rect 580746 186140 580982 186376
rect 581066 186140 581302 186376
rect 580746 185820 580982 186056
rect 581066 185820 581302 186056
rect 580746 150140 580982 150376
rect 581066 150140 581302 150376
rect 580746 149820 580982 150056
rect 581066 149820 581302 150056
rect 580746 114140 580982 114376
rect 581066 114140 581302 114376
rect 580746 113820 580982 114056
rect 581066 113820 581302 114056
rect 580746 78140 580982 78376
rect 581066 78140 581302 78376
rect 580746 77820 580982 78056
rect 581066 77820 581302 78056
rect 580746 42140 580982 42376
rect 581066 42140 581302 42376
rect 580746 41820 580982 42056
rect 581066 41820 581302 42056
rect 580746 6140 580982 6376
rect 581066 6140 581302 6376
rect 580746 5820 580982 6056
rect 581066 5820 581302 6056
rect 580746 -3460 580982 -3224
rect 581066 -3460 581302 -3224
rect 580746 -3780 580982 -3544
rect 581066 -3780 581302 -3544
rect 592062 711324 592298 711560
rect 592382 711324 592618 711560
rect 592062 711004 592298 711240
rect 592382 711004 592618 711240
rect 591102 710364 591338 710600
rect 591422 710364 591658 710600
rect 591102 710044 591338 710280
rect 591422 710044 591658 710280
rect 590142 709404 590378 709640
rect 590462 709404 590698 709640
rect 590142 709084 590378 709320
rect 590462 709084 590698 709320
rect 581986 708444 582222 708680
rect 582306 708444 582542 708680
rect 581986 708124 582222 708360
rect 582306 708124 582542 708360
rect 589182 708444 589418 708680
rect 589502 708444 589738 708680
rect 589182 708124 589418 708360
rect 589502 708124 589738 708360
rect 588222 707484 588458 707720
rect 588542 707484 588778 707720
rect 588222 707164 588458 707400
rect 588542 707164 588778 707400
rect 587262 706524 587498 706760
rect 587582 706524 587818 706760
rect 587262 706204 587498 706440
rect 587582 706204 587818 706440
rect 586302 705564 586538 705800
rect 586622 705564 586858 705800
rect 586302 705244 586538 705480
rect 586622 705244 586858 705480
rect 581986 691380 582222 691616
rect 582306 691380 582542 691616
rect 581986 691060 582222 691296
rect 582306 691060 582542 691296
rect 581986 655380 582222 655616
rect 582306 655380 582542 655616
rect 581986 655060 582222 655296
rect 582306 655060 582542 655296
rect 581986 619380 582222 619616
rect 582306 619380 582542 619616
rect 581986 619060 582222 619296
rect 582306 619060 582542 619296
rect 581986 583380 582222 583616
rect 582306 583380 582542 583616
rect 581986 583060 582222 583296
rect 582306 583060 582542 583296
rect 581986 547380 582222 547616
rect 582306 547380 582542 547616
rect 581986 547060 582222 547296
rect 582306 547060 582542 547296
rect 581986 511380 582222 511616
rect 582306 511380 582542 511616
rect 581986 511060 582222 511296
rect 582306 511060 582542 511296
rect 581986 475380 582222 475616
rect 582306 475380 582542 475616
rect 581986 475060 582222 475296
rect 582306 475060 582542 475296
rect 581986 439380 582222 439616
rect 582306 439380 582542 439616
rect 581986 439060 582222 439296
rect 582306 439060 582542 439296
rect 581986 403380 582222 403616
rect 582306 403380 582542 403616
rect 581986 403060 582222 403296
rect 582306 403060 582542 403296
rect 581986 367380 582222 367616
rect 582306 367380 582542 367616
rect 581986 367060 582222 367296
rect 582306 367060 582542 367296
rect 581986 331380 582222 331616
rect 582306 331380 582542 331616
rect 581986 331060 582222 331296
rect 582306 331060 582542 331296
rect 581986 295380 582222 295616
rect 582306 295380 582542 295616
rect 581986 295060 582222 295296
rect 582306 295060 582542 295296
rect 581986 259380 582222 259616
rect 582306 259380 582542 259616
rect 581986 259060 582222 259296
rect 582306 259060 582542 259296
rect 581986 223380 582222 223616
rect 582306 223380 582542 223616
rect 581986 223060 582222 223296
rect 582306 223060 582542 223296
rect 581986 187380 582222 187616
rect 582306 187380 582542 187616
rect 581986 187060 582222 187296
rect 582306 187060 582542 187296
rect 581986 151380 582222 151616
rect 582306 151380 582542 151616
rect 581986 151060 582222 151296
rect 582306 151060 582542 151296
rect 581986 115380 582222 115616
rect 582306 115380 582542 115616
rect 581986 115060 582222 115296
rect 582306 115060 582542 115296
rect 581986 79380 582222 79616
rect 582306 79380 582542 79616
rect 581986 79060 582222 79296
rect 582306 79060 582542 79296
rect 581986 43380 582222 43616
rect 582306 43380 582542 43616
rect 581986 43060 582222 43296
rect 582306 43060 582542 43296
rect 581986 7380 582222 7616
rect 582306 7380 582542 7616
rect 581986 7060 582222 7296
rect 582306 7060 582542 7296
rect 585342 704604 585578 704840
rect 585662 704604 585898 704840
rect 585342 704284 585578 704520
rect 585662 704284 585898 704520
rect 585342 686420 585578 686656
rect 585662 686420 585898 686656
rect 585342 686100 585578 686336
rect 585662 686100 585898 686336
rect 585342 650420 585578 650656
rect 585662 650420 585898 650656
rect 585342 650100 585578 650336
rect 585662 650100 585898 650336
rect 585342 614420 585578 614656
rect 585662 614420 585898 614656
rect 585342 614100 585578 614336
rect 585662 614100 585898 614336
rect 585342 578420 585578 578656
rect 585662 578420 585898 578656
rect 585342 578100 585578 578336
rect 585662 578100 585898 578336
rect 585342 542420 585578 542656
rect 585662 542420 585898 542656
rect 585342 542100 585578 542336
rect 585662 542100 585898 542336
rect 585342 506420 585578 506656
rect 585662 506420 585898 506656
rect 585342 506100 585578 506336
rect 585662 506100 585898 506336
rect 585342 470420 585578 470656
rect 585662 470420 585898 470656
rect 585342 470100 585578 470336
rect 585662 470100 585898 470336
rect 585342 434420 585578 434656
rect 585662 434420 585898 434656
rect 585342 434100 585578 434336
rect 585662 434100 585898 434336
rect 585342 398420 585578 398656
rect 585662 398420 585898 398656
rect 585342 398100 585578 398336
rect 585662 398100 585898 398336
rect 585342 362420 585578 362656
rect 585662 362420 585898 362656
rect 585342 362100 585578 362336
rect 585662 362100 585898 362336
rect 585342 326420 585578 326656
rect 585662 326420 585898 326656
rect 585342 326100 585578 326336
rect 585662 326100 585898 326336
rect 585342 290420 585578 290656
rect 585662 290420 585898 290656
rect 585342 290100 585578 290336
rect 585662 290100 585898 290336
rect 585342 254420 585578 254656
rect 585662 254420 585898 254656
rect 585342 254100 585578 254336
rect 585662 254100 585898 254336
rect 585342 218420 585578 218656
rect 585662 218420 585898 218656
rect 585342 218100 585578 218336
rect 585662 218100 585898 218336
rect 585342 182420 585578 182656
rect 585662 182420 585898 182656
rect 585342 182100 585578 182336
rect 585662 182100 585898 182336
rect 585342 146420 585578 146656
rect 585662 146420 585898 146656
rect 585342 146100 585578 146336
rect 585662 146100 585898 146336
rect 585342 110420 585578 110656
rect 585662 110420 585898 110656
rect 585342 110100 585578 110336
rect 585662 110100 585898 110336
rect 585342 74420 585578 74656
rect 585662 74420 585898 74656
rect 585342 74100 585578 74336
rect 585662 74100 585898 74336
rect 585342 38420 585578 38656
rect 585662 38420 585898 38656
rect 585342 38100 585578 38336
rect 585662 38100 585898 38336
rect 585342 2420 585578 2656
rect 585662 2420 585898 2656
rect 585342 2100 585578 2336
rect 585662 2100 585898 2336
rect 585342 -580 585578 -344
rect 585662 -580 585898 -344
rect 585342 -900 585578 -664
rect 585662 -900 585898 -664
rect 586302 687660 586538 687896
rect 586622 687660 586858 687896
rect 586302 687340 586538 687576
rect 586622 687340 586858 687576
rect 586302 651660 586538 651896
rect 586622 651660 586858 651896
rect 586302 651340 586538 651576
rect 586622 651340 586858 651576
rect 586302 615660 586538 615896
rect 586622 615660 586858 615896
rect 586302 615340 586538 615576
rect 586622 615340 586858 615576
rect 586302 579660 586538 579896
rect 586622 579660 586858 579896
rect 586302 579340 586538 579576
rect 586622 579340 586858 579576
rect 586302 543660 586538 543896
rect 586622 543660 586858 543896
rect 586302 543340 586538 543576
rect 586622 543340 586858 543576
rect 586302 507660 586538 507896
rect 586622 507660 586858 507896
rect 586302 507340 586538 507576
rect 586622 507340 586858 507576
rect 586302 471660 586538 471896
rect 586622 471660 586858 471896
rect 586302 471340 586538 471576
rect 586622 471340 586858 471576
rect 586302 435660 586538 435896
rect 586622 435660 586858 435896
rect 586302 435340 586538 435576
rect 586622 435340 586858 435576
rect 586302 399660 586538 399896
rect 586622 399660 586858 399896
rect 586302 399340 586538 399576
rect 586622 399340 586858 399576
rect 586302 363660 586538 363896
rect 586622 363660 586858 363896
rect 586302 363340 586538 363576
rect 586622 363340 586858 363576
rect 586302 327660 586538 327896
rect 586622 327660 586858 327896
rect 586302 327340 586538 327576
rect 586622 327340 586858 327576
rect 586302 291660 586538 291896
rect 586622 291660 586858 291896
rect 586302 291340 586538 291576
rect 586622 291340 586858 291576
rect 586302 255660 586538 255896
rect 586622 255660 586858 255896
rect 586302 255340 586538 255576
rect 586622 255340 586858 255576
rect 586302 219660 586538 219896
rect 586622 219660 586858 219896
rect 586302 219340 586538 219576
rect 586622 219340 586858 219576
rect 586302 183660 586538 183896
rect 586622 183660 586858 183896
rect 586302 183340 586538 183576
rect 586622 183340 586858 183576
rect 586302 147660 586538 147896
rect 586622 147660 586858 147896
rect 586302 147340 586538 147576
rect 586622 147340 586858 147576
rect 586302 111660 586538 111896
rect 586622 111660 586858 111896
rect 586302 111340 586538 111576
rect 586622 111340 586858 111576
rect 586302 75660 586538 75896
rect 586622 75660 586858 75896
rect 586302 75340 586538 75576
rect 586622 75340 586858 75576
rect 586302 39660 586538 39896
rect 586622 39660 586858 39896
rect 586302 39340 586538 39576
rect 586622 39340 586858 39576
rect 586302 3660 586538 3896
rect 586622 3660 586858 3896
rect 586302 3340 586538 3576
rect 586622 3340 586858 3576
rect 586302 -1540 586538 -1304
rect 586622 -1540 586858 -1304
rect 586302 -1860 586538 -1624
rect 586622 -1860 586858 -1624
rect 587262 688900 587498 689136
rect 587582 688900 587818 689136
rect 587262 688580 587498 688816
rect 587582 688580 587818 688816
rect 587262 652900 587498 653136
rect 587582 652900 587818 653136
rect 587262 652580 587498 652816
rect 587582 652580 587818 652816
rect 587262 616900 587498 617136
rect 587582 616900 587818 617136
rect 587262 616580 587498 616816
rect 587582 616580 587818 616816
rect 587262 580900 587498 581136
rect 587582 580900 587818 581136
rect 587262 580580 587498 580816
rect 587582 580580 587818 580816
rect 587262 544900 587498 545136
rect 587582 544900 587818 545136
rect 587262 544580 587498 544816
rect 587582 544580 587818 544816
rect 587262 508900 587498 509136
rect 587582 508900 587818 509136
rect 587262 508580 587498 508816
rect 587582 508580 587818 508816
rect 587262 472900 587498 473136
rect 587582 472900 587818 473136
rect 587262 472580 587498 472816
rect 587582 472580 587818 472816
rect 587262 436900 587498 437136
rect 587582 436900 587818 437136
rect 587262 436580 587498 436816
rect 587582 436580 587818 436816
rect 587262 400900 587498 401136
rect 587582 400900 587818 401136
rect 587262 400580 587498 400816
rect 587582 400580 587818 400816
rect 587262 364900 587498 365136
rect 587582 364900 587818 365136
rect 587262 364580 587498 364816
rect 587582 364580 587818 364816
rect 587262 328900 587498 329136
rect 587582 328900 587818 329136
rect 587262 328580 587498 328816
rect 587582 328580 587818 328816
rect 587262 292900 587498 293136
rect 587582 292900 587818 293136
rect 587262 292580 587498 292816
rect 587582 292580 587818 292816
rect 587262 256900 587498 257136
rect 587582 256900 587818 257136
rect 587262 256580 587498 256816
rect 587582 256580 587818 256816
rect 587262 220900 587498 221136
rect 587582 220900 587818 221136
rect 587262 220580 587498 220816
rect 587582 220580 587818 220816
rect 587262 184900 587498 185136
rect 587582 184900 587818 185136
rect 587262 184580 587498 184816
rect 587582 184580 587818 184816
rect 587262 148900 587498 149136
rect 587582 148900 587818 149136
rect 587262 148580 587498 148816
rect 587582 148580 587818 148816
rect 587262 112900 587498 113136
rect 587582 112900 587818 113136
rect 587262 112580 587498 112816
rect 587582 112580 587818 112816
rect 587262 76900 587498 77136
rect 587582 76900 587818 77136
rect 587262 76580 587498 76816
rect 587582 76580 587818 76816
rect 587262 40900 587498 41136
rect 587582 40900 587818 41136
rect 587262 40580 587498 40816
rect 587582 40580 587818 40816
rect 587262 4900 587498 5136
rect 587582 4900 587818 5136
rect 587262 4580 587498 4816
rect 587582 4580 587818 4816
rect 587262 -2500 587498 -2264
rect 587582 -2500 587818 -2264
rect 587262 -2820 587498 -2584
rect 587582 -2820 587818 -2584
rect 588222 690140 588458 690376
rect 588542 690140 588778 690376
rect 588222 689820 588458 690056
rect 588542 689820 588778 690056
rect 588222 654140 588458 654376
rect 588542 654140 588778 654376
rect 588222 653820 588458 654056
rect 588542 653820 588778 654056
rect 588222 618140 588458 618376
rect 588542 618140 588778 618376
rect 588222 617820 588458 618056
rect 588542 617820 588778 618056
rect 588222 582140 588458 582376
rect 588542 582140 588778 582376
rect 588222 581820 588458 582056
rect 588542 581820 588778 582056
rect 588222 546140 588458 546376
rect 588542 546140 588778 546376
rect 588222 545820 588458 546056
rect 588542 545820 588778 546056
rect 588222 510140 588458 510376
rect 588542 510140 588778 510376
rect 588222 509820 588458 510056
rect 588542 509820 588778 510056
rect 588222 474140 588458 474376
rect 588542 474140 588778 474376
rect 588222 473820 588458 474056
rect 588542 473820 588778 474056
rect 588222 438140 588458 438376
rect 588542 438140 588778 438376
rect 588222 437820 588458 438056
rect 588542 437820 588778 438056
rect 588222 402140 588458 402376
rect 588542 402140 588778 402376
rect 588222 401820 588458 402056
rect 588542 401820 588778 402056
rect 588222 366140 588458 366376
rect 588542 366140 588778 366376
rect 588222 365820 588458 366056
rect 588542 365820 588778 366056
rect 588222 330140 588458 330376
rect 588542 330140 588778 330376
rect 588222 329820 588458 330056
rect 588542 329820 588778 330056
rect 588222 294140 588458 294376
rect 588542 294140 588778 294376
rect 588222 293820 588458 294056
rect 588542 293820 588778 294056
rect 588222 258140 588458 258376
rect 588542 258140 588778 258376
rect 588222 257820 588458 258056
rect 588542 257820 588778 258056
rect 588222 222140 588458 222376
rect 588542 222140 588778 222376
rect 588222 221820 588458 222056
rect 588542 221820 588778 222056
rect 588222 186140 588458 186376
rect 588542 186140 588778 186376
rect 588222 185820 588458 186056
rect 588542 185820 588778 186056
rect 588222 150140 588458 150376
rect 588542 150140 588778 150376
rect 588222 149820 588458 150056
rect 588542 149820 588778 150056
rect 588222 114140 588458 114376
rect 588542 114140 588778 114376
rect 588222 113820 588458 114056
rect 588542 113820 588778 114056
rect 588222 78140 588458 78376
rect 588542 78140 588778 78376
rect 588222 77820 588458 78056
rect 588542 77820 588778 78056
rect 588222 42140 588458 42376
rect 588542 42140 588778 42376
rect 588222 41820 588458 42056
rect 588542 41820 588778 42056
rect 588222 6140 588458 6376
rect 588542 6140 588778 6376
rect 588222 5820 588458 6056
rect 588542 5820 588778 6056
rect 588222 -3460 588458 -3224
rect 588542 -3460 588778 -3224
rect 588222 -3780 588458 -3544
rect 588542 -3780 588778 -3544
rect 589182 691380 589418 691616
rect 589502 691380 589738 691616
rect 589182 691060 589418 691296
rect 589502 691060 589738 691296
rect 589182 655380 589418 655616
rect 589502 655380 589738 655616
rect 589182 655060 589418 655296
rect 589502 655060 589738 655296
rect 589182 619380 589418 619616
rect 589502 619380 589738 619616
rect 589182 619060 589418 619296
rect 589502 619060 589738 619296
rect 589182 583380 589418 583616
rect 589502 583380 589738 583616
rect 589182 583060 589418 583296
rect 589502 583060 589738 583296
rect 589182 547380 589418 547616
rect 589502 547380 589738 547616
rect 589182 547060 589418 547296
rect 589502 547060 589738 547296
rect 589182 511380 589418 511616
rect 589502 511380 589738 511616
rect 589182 511060 589418 511296
rect 589502 511060 589738 511296
rect 589182 475380 589418 475616
rect 589502 475380 589738 475616
rect 589182 475060 589418 475296
rect 589502 475060 589738 475296
rect 589182 439380 589418 439616
rect 589502 439380 589738 439616
rect 589182 439060 589418 439296
rect 589502 439060 589738 439296
rect 589182 403380 589418 403616
rect 589502 403380 589738 403616
rect 589182 403060 589418 403296
rect 589502 403060 589738 403296
rect 589182 367380 589418 367616
rect 589502 367380 589738 367616
rect 589182 367060 589418 367296
rect 589502 367060 589738 367296
rect 589182 331380 589418 331616
rect 589502 331380 589738 331616
rect 589182 331060 589418 331296
rect 589502 331060 589738 331296
rect 589182 295380 589418 295616
rect 589502 295380 589738 295616
rect 589182 295060 589418 295296
rect 589502 295060 589738 295296
rect 589182 259380 589418 259616
rect 589502 259380 589738 259616
rect 589182 259060 589418 259296
rect 589502 259060 589738 259296
rect 589182 223380 589418 223616
rect 589502 223380 589738 223616
rect 589182 223060 589418 223296
rect 589502 223060 589738 223296
rect 589182 187380 589418 187616
rect 589502 187380 589738 187616
rect 589182 187060 589418 187296
rect 589502 187060 589738 187296
rect 589182 151380 589418 151616
rect 589502 151380 589738 151616
rect 589182 151060 589418 151296
rect 589502 151060 589738 151296
rect 589182 115380 589418 115616
rect 589502 115380 589738 115616
rect 589182 115060 589418 115296
rect 589502 115060 589738 115296
rect 589182 79380 589418 79616
rect 589502 79380 589738 79616
rect 589182 79060 589418 79296
rect 589502 79060 589738 79296
rect 589182 43380 589418 43616
rect 589502 43380 589738 43616
rect 589182 43060 589418 43296
rect 589502 43060 589738 43296
rect 589182 7380 589418 7616
rect 589502 7380 589738 7616
rect 589182 7060 589418 7296
rect 589502 7060 589738 7296
rect 581986 -4420 582222 -4184
rect 582306 -4420 582542 -4184
rect 581986 -4740 582222 -4504
rect 582306 -4740 582542 -4504
rect 589182 -4420 589418 -4184
rect 589502 -4420 589738 -4184
rect 589182 -4740 589418 -4504
rect 589502 -4740 589738 -4504
rect 590142 692620 590378 692856
rect 590462 692620 590698 692856
rect 590142 692300 590378 692536
rect 590462 692300 590698 692536
rect 590142 656620 590378 656856
rect 590462 656620 590698 656856
rect 590142 656300 590378 656536
rect 590462 656300 590698 656536
rect 590142 620620 590378 620856
rect 590462 620620 590698 620856
rect 590142 620300 590378 620536
rect 590462 620300 590698 620536
rect 590142 584620 590378 584856
rect 590462 584620 590698 584856
rect 590142 584300 590378 584536
rect 590462 584300 590698 584536
rect 590142 548620 590378 548856
rect 590462 548620 590698 548856
rect 590142 548300 590378 548536
rect 590462 548300 590698 548536
rect 590142 512620 590378 512856
rect 590462 512620 590698 512856
rect 590142 512300 590378 512536
rect 590462 512300 590698 512536
rect 590142 476620 590378 476856
rect 590462 476620 590698 476856
rect 590142 476300 590378 476536
rect 590462 476300 590698 476536
rect 590142 440620 590378 440856
rect 590462 440620 590698 440856
rect 590142 440300 590378 440536
rect 590462 440300 590698 440536
rect 590142 404620 590378 404856
rect 590462 404620 590698 404856
rect 590142 404300 590378 404536
rect 590462 404300 590698 404536
rect 590142 368620 590378 368856
rect 590462 368620 590698 368856
rect 590142 368300 590378 368536
rect 590462 368300 590698 368536
rect 590142 332620 590378 332856
rect 590462 332620 590698 332856
rect 590142 332300 590378 332536
rect 590462 332300 590698 332536
rect 590142 296620 590378 296856
rect 590462 296620 590698 296856
rect 590142 296300 590378 296536
rect 590462 296300 590698 296536
rect 590142 260620 590378 260856
rect 590462 260620 590698 260856
rect 590142 260300 590378 260536
rect 590462 260300 590698 260536
rect 590142 224620 590378 224856
rect 590462 224620 590698 224856
rect 590142 224300 590378 224536
rect 590462 224300 590698 224536
rect 590142 188620 590378 188856
rect 590462 188620 590698 188856
rect 590142 188300 590378 188536
rect 590462 188300 590698 188536
rect 590142 152620 590378 152856
rect 590462 152620 590698 152856
rect 590142 152300 590378 152536
rect 590462 152300 590698 152536
rect 590142 116620 590378 116856
rect 590462 116620 590698 116856
rect 590142 116300 590378 116536
rect 590462 116300 590698 116536
rect 590142 80620 590378 80856
rect 590462 80620 590698 80856
rect 590142 80300 590378 80536
rect 590462 80300 590698 80536
rect 590142 44620 590378 44856
rect 590462 44620 590698 44856
rect 590142 44300 590378 44536
rect 590462 44300 590698 44536
rect 590142 8620 590378 8856
rect 590462 8620 590698 8856
rect 590142 8300 590378 8536
rect 590462 8300 590698 8536
rect 590142 -5380 590378 -5144
rect 590462 -5380 590698 -5144
rect 590142 -5700 590378 -5464
rect 590462 -5700 590698 -5464
rect 591102 693860 591338 694096
rect 591422 693860 591658 694096
rect 591102 693540 591338 693776
rect 591422 693540 591658 693776
rect 591102 657860 591338 658096
rect 591422 657860 591658 658096
rect 591102 657540 591338 657776
rect 591422 657540 591658 657776
rect 591102 621860 591338 622096
rect 591422 621860 591658 622096
rect 591102 621540 591338 621776
rect 591422 621540 591658 621776
rect 591102 585860 591338 586096
rect 591422 585860 591658 586096
rect 591102 585540 591338 585776
rect 591422 585540 591658 585776
rect 591102 549860 591338 550096
rect 591422 549860 591658 550096
rect 591102 549540 591338 549776
rect 591422 549540 591658 549776
rect 591102 513860 591338 514096
rect 591422 513860 591658 514096
rect 591102 513540 591338 513776
rect 591422 513540 591658 513776
rect 591102 477860 591338 478096
rect 591422 477860 591658 478096
rect 591102 477540 591338 477776
rect 591422 477540 591658 477776
rect 591102 441860 591338 442096
rect 591422 441860 591658 442096
rect 591102 441540 591338 441776
rect 591422 441540 591658 441776
rect 591102 405860 591338 406096
rect 591422 405860 591658 406096
rect 591102 405540 591338 405776
rect 591422 405540 591658 405776
rect 591102 369860 591338 370096
rect 591422 369860 591658 370096
rect 591102 369540 591338 369776
rect 591422 369540 591658 369776
rect 591102 333860 591338 334096
rect 591422 333860 591658 334096
rect 591102 333540 591338 333776
rect 591422 333540 591658 333776
rect 591102 297860 591338 298096
rect 591422 297860 591658 298096
rect 591102 297540 591338 297776
rect 591422 297540 591658 297776
rect 591102 261860 591338 262096
rect 591422 261860 591658 262096
rect 591102 261540 591338 261776
rect 591422 261540 591658 261776
rect 591102 225860 591338 226096
rect 591422 225860 591658 226096
rect 591102 225540 591338 225776
rect 591422 225540 591658 225776
rect 591102 189860 591338 190096
rect 591422 189860 591658 190096
rect 591102 189540 591338 189776
rect 591422 189540 591658 189776
rect 591102 153860 591338 154096
rect 591422 153860 591658 154096
rect 591102 153540 591338 153776
rect 591422 153540 591658 153776
rect 591102 117860 591338 118096
rect 591422 117860 591658 118096
rect 591102 117540 591338 117776
rect 591422 117540 591658 117776
rect 591102 81860 591338 82096
rect 591422 81860 591658 82096
rect 591102 81540 591338 81776
rect 591422 81540 591658 81776
rect 591102 45860 591338 46096
rect 591422 45860 591658 46096
rect 591102 45540 591338 45776
rect 591422 45540 591658 45776
rect 591102 9860 591338 10096
rect 591422 9860 591658 10096
rect 591102 9540 591338 9776
rect 591422 9540 591658 9776
rect 591102 -6340 591338 -6104
rect 591422 -6340 591658 -6104
rect 591102 -6660 591338 -6424
rect 591422 -6660 591658 -6424
rect 592062 695100 592298 695336
rect 592382 695100 592618 695336
rect 592062 694780 592298 695016
rect 592382 694780 592618 695016
rect 592062 659100 592298 659336
rect 592382 659100 592618 659336
rect 592062 658780 592298 659016
rect 592382 658780 592618 659016
rect 592062 623100 592298 623336
rect 592382 623100 592618 623336
rect 592062 622780 592298 623016
rect 592382 622780 592618 623016
rect 592062 587100 592298 587336
rect 592382 587100 592618 587336
rect 592062 586780 592298 587016
rect 592382 586780 592618 587016
rect 592062 551100 592298 551336
rect 592382 551100 592618 551336
rect 592062 550780 592298 551016
rect 592382 550780 592618 551016
rect 592062 515100 592298 515336
rect 592382 515100 592618 515336
rect 592062 514780 592298 515016
rect 592382 514780 592618 515016
rect 592062 479100 592298 479336
rect 592382 479100 592618 479336
rect 592062 478780 592298 479016
rect 592382 478780 592618 479016
rect 592062 443100 592298 443336
rect 592382 443100 592618 443336
rect 592062 442780 592298 443016
rect 592382 442780 592618 443016
rect 592062 407100 592298 407336
rect 592382 407100 592618 407336
rect 592062 406780 592298 407016
rect 592382 406780 592618 407016
rect 592062 371100 592298 371336
rect 592382 371100 592618 371336
rect 592062 370780 592298 371016
rect 592382 370780 592618 371016
rect 592062 335100 592298 335336
rect 592382 335100 592618 335336
rect 592062 334780 592298 335016
rect 592382 334780 592618 335016
rect 592062 299100 592298 299336
rect 592382 299100 592618 299336
rect 592062 298780 592298 299016
rect 592382 298780 592618 299016
rect 592062 263100 592298 263336
rect 592382 263100 592618 263336
rect 592062 262780 592298 263016
rect 592382 262780 592618 263016
rect 592062 227100 592298 227336
rect 592382 227100 592618 227336
rect 592062 226780 592298 227016
rect 592382 226780 592618 227016
rect 592062 191100 592298 191336
rect 592382 191100 592618 191336
rect 592062 190780 592298 191016
rect 592382 190780 592618 191016
rect 592062 155100 592298 155336
rect 592382 155100 592618 155336
rect 592062 154780 592298 155016
rect 592382 154780 592618 155016
rect 592062 119100 592298 119336
rect 592382 119100 592618 119336
rect 592062 118780 592298 119016
rect 592382 118780 592618 119016
rect 592062 83100 592298 83336
rect 592382 83100 592618 83336
rect 592062 82780 592298 83016
rect 592382 82780 592618 83016
rect 592062 47100 592298 47336
rect 592382 47100 592618 47336
rect 592062 46780 592298 47016
rect 592382 46780 592618 47016
rect 592062 11100 592298 11336
rect 592382 11100 592618 11336
rect 592062 10780 592298 11016
rect 592382 10780 592618 11016
rect 592062 -7300 592298 -7064
rect 592382 -7300 592618 -7064
rect 592062 -7620 592298 -7384
rect 592382 -7620 592618 -7384
<< metal5 >>
rect -8726 711560 592650 711592
rect -8726 711324 -8694 711560
rect -8458 711324 -8374 711560
rect -8138 711324 9706 711560
rect 9942 711324 10026 711560
rect 10262 711324 45706 711560
rect 45942 711324 46026 711560
rect 46262 711324 81706 711560
rect 81942 711324 82026 711560
rect 82262 711324 117706 711560
rect 117942 711324 118026 711560
rect 118262 711324 153706 711560
rect 153942 711324 154026 711560
rect 154262 711324 189706 711560
rect 189942 711324 190026 711560
rect 190262 711324 225706 711560
rect 225942 711324 226026 711560
rect 226262 711324 261706 711560
rect 261942 711324 262026 711560
rect 262262 711324 297706 711560
rect 297942 711324 298026 711560
rect 298262 711324 333706 711560
rect 333942 711324 334026 711560
rect 334262 711324 369706 711560
rect 369942 711324 370026 711560
rect 370262 711324 405706 711560
rect 405942 711324 406026 711560
rect 406262 711324 441706 711560
rect 441942 711324 442026 711560
rect 442262 711324 477706 711560
rect 477942 711324 478026 711560
rect 478262 711324 513706 711560
rect 513942 711324 514026 711560
rect 514262 711324 549706 711560
rect 549942 711324 550026 711560
rect 550262 711324 592062 711560
rect 592298 711324 592382 711560
rect 592618 711324 592650 711560
rect -8726 711240 592650 711324
rect -8726 711004 -8694 711240
rect -8458 711004 -8374 711240
rect -8138 711004 9706 711240
rect 9942 711004 10026 711240
rect 10262 711004 45706 711240
rect 45942 711004 46026 711240
rect 46262 711004 81706 711240
rect 81942 711004 82026 711240
rect 82262 711004 117706 711240
rect 117942 711004 118026 711240
rect 118262 711004 153706 711240
rect 153942 711004 154026 711240
rect 154262 711004 189706 711240
rect 189942 711004 190026 711240
rect 190262 711004 225706 711240
rect 225942 711004 226026 711240
rect 226262 711004 261706 711240
rect 261942 711004 262026 711240
rect 262262 711004 297706 711240
rect 297942 711004 298026 711240
rect 298262 711004 333706 711240
rect 333942 711004 334026 711240
rect 334262 711004 369706 711240
rect 369942 711004 370026 711240
rect 370262 711004 405706 711240
rect 405942 711004 406026 711240
rect 406262 711004 441706 711240
rect 441942 711004 442026 711240
rect 442262 711004 477706 711240
rect 477942 711004 478026 711240
rect 478262 711004 513706 711240
rect 513942 711004 514026 711240
rect 514262 711004 549706 711240
rect 549942 711004 550026 711240
rect 550262 711004 592062 711240
rect 592298 711004 592382 711240
rect 592618 711004 592650 711240
rect -8726 710972 592650 711004
rect -7766 710600 591690 710632
rect -7766 710364 -7734 710600
rect -7498 710364 -7414 710600
rect -7178 710364 8466 710600
rect 8702 710364 8786 710600
rect 9022 710364 44466 710600
rect 44702 710364 44786 710600
rect 45022 710364 80466 710600
rect 80702 710364 80786 710600
rect 81022 710364 116466 710600
rect 116702 710364 116786 710600
rect 117022 710364 152466 710600
rect 152702 710364 152786 710600
rect 153022 710364 188466 710600
rect 188702 710364 188786 710600
rect 189022 710364 224466 710600
rect 224702 710364 224786 710600
rect 225022 710364 260466 710600
rect 260702 710364 260786 710600
rect 261022 710364 296466 710600
rect 296702 710364 296786 710600
rect 297022 710364 332466 710600
rect 332702 710364 332786 710600
rect 333022 710364 368466 710600
rect 368702 710364 368786 710600
rect 369022 710364 404466 710600
rect 404702 710364 404786 710600
rect 405022 710364 440466 710600
rect 440702 710364 440786 710600
rect 441022 710364 476466 710600
rect 476702 710364 476786 710600
rect 477022 710364 512466 710600
rect 512702 710364 512786 710600
rect 513022 710364 548466 710600
rect 548702 710364 548786 710600
rect 549022 710364 591102 710600
rect 591338 710364 591422 710600
rect 591658 710364 591690 710600
rect -7766 710280 591690 710364
rect -7766 710044 -7734 710280
rect -7498 710044 -7414 710280
rect -7178 710044 8466 710280
rect 8702 710044 8786 710280
rect 9022 710044 44466 710280
rect 44702 710044 44786 710280
rect 45022 710044 80466 710280
rect 80702 710044 80786 710280
rect 81022 710044 116466 710280
rect 116702 710044 116786 710280
rect 117022 710044 152466 710280
rect 152702 710044 152786 710280
rect 153022 710044 188466 710280
rect 188702 710044 188786 710280
rect 189022 710044 224466 710280
rect 224702 710044 224786 710280
rect 225022 710044 260466 710280
rect 260702 710044 260786 710280
rect 261022 710044 296466 710280
rect 296702 710044 296786 710280
rect 297022 710044 332466 710280
rect 332702 710044 332786 710280
rect 333022 710044 368466 710280
rect 368702 710044 368786 710280
rect 369022 710044 404466 710280
rect 404702 710044 404786 710280
rect 405022 710044 440466 710280
rect 440702 710044 440786 710280
rect 441022 710044 476466 710280
rect 476702 710044 476786 710280
rect 477022 710044 512466 710280
rect 512702 710044 512786 710280
rect 513022 710044 548466 710280
rect 548702 710044 548786 710280
rect 549022 710044 591102 710280
rect 591338 710044 591422 710280
rect 591658 710044 591690 710280
rect -7766 710012 591690 710044
rect -6806 709640 590730 709672
rect -6806 709404 -6774 709640
rect -6538 709404 -6454 709640
rect -6218 709404 7226 709640
rect 7462 709404 7546 709640
rect 7782 709404 43226 709640
rect 43462 709404 43546 709640
rect 43782 709404 79226 709640
rect 79462 709404 79546 709640
rect 79782 709404 115226 709640
rect 115462 709404 115546 709640
rect 115782 709404 151226 709640
rect 151462 709404 151546 709640
rect 151782 709404 187226 709640
rect 187462 709404 187546 709640
rect 187782 709404 223226 709640
rect 223462 709404 223546 709640
rect 223782 709404 259226 709640
rect 259462 709404 259546 709640
rect 259782 709404 295226 709640
rect 295462 709404 295546 709640
rect 295782 709404 331226 709640
rect 331462 709404 331546 709640
rect 331782 709404 367226 709640
rect 367462 709404 367546 709640
rect 367782 709404 403226 709640
rect 403462 709404 403546 709640
rect 403782 709404 439226 709640
rect 439462 709404 439546 709640
rect 439782 709404 475226 709640
rect 475462 709404 475546 709640
rect 475782 709404 511226 709640
rect 511462 709404 511546 709640
rect 511782 709404 547226 709640
rect 547462 709404 547546 709640
rect 547782 709404 590142 709640
rect 590378 709404 590462 709640
rect 590698 709404 590730 709640
rect -6806 709320 590730 709404
rect -6806 709084 -6774 709320
rect -6538 709084 -6454 709320
rect -6218 709084 7226 709320
rect 7462 709084 7546 709320
rect 7782 709084 43226 709320
rect 43462 709084 43546 709320
rect 43782 709084 79226 709320
rect 79462 709084 79546 709320
rect 79782 709084 115226 709320
rect 115462 709084 115546 709320
rect 115782 709084 151226 709320
rect 151462 709084 151546 709320
rect 151782 709084 187226 709320
rect 187462 709084 187546 709320
rect 187782 709084 223226 709320
rect 223462 709084 223546 709320
rect 223782 709084 259226 709320
rect 259462 709084 259546 709320
rect 259782 709084 295226 709320
rect 295462 709084 295546 709320
rect 295782 709084 331226 709320
rect 331462 709084 331546 709320
rect 331782 709084 367226 709320
rect 367462 709084 367546 709320
rect 367782 709084 403226 709320
rect 403462 709084 403546 709320
rect 403782 709084 439226 709320
rect 439462 709084 439546 709320
rect 439782 709084 475226 709320
rect 475462 709084 475546 709320
rect 475782 709084 511226 709320
rect 511462 709084 511546 709320
rect 511782 709084 547226 709320
rect 547462 709084 547546 709320
rect 547782 709084 590142 709320
rect 590378 709084 590462 709320
rect 590698 709084 590730 709320
rect -6806 709052 590730 709084
rect -5846 708680 589770 708712
rect -5846 708444 -5814 708680
rect -5578 708444 -5494 708680
rect -5258 708444 5986 708680
rect 6222 708444 6306 708680
rect 6542 708444 41986 708680
rect 42222 708444 42306 708680
rect 42542 708444 77986 708680
rect 78222 708444 78306 708680
rect 78542 708444 113986 708680
rect 114222 708444 114306 708680
rect 114542 708444 149986 708680
rect 150222 708444 150306 708680
rect 150542 708444 185986 708680
rect 186222 708444 186306 708680
rect 186542 708444 221986 708680
rect 222222 708444 222306 708680
rect 222542 708444 257986 708680
rect 258222 708444 258306 708680
rect 258542 708444 293986 708680
rect 294222 708444 294306 708680
rect 294542 708444 329986 708680
rect 330222 708444 330306 708680
rect 330542 708444 365986 708680
rect 366222 708444 366306 708680
rect 366542 708444 401986 708680
rect 402222 708444 402306 708680
rect 402542 708444 437986 708680
rect 438222 708444 438306 708680
rect 438542 708444 473986 708680
rect 474222 708444 474306 708680
rect 474542 708444 509986 708680
rect 510222 708444 510306 708680
rect 510542 708444 545986 708680
rect 546222 708444 546306 708680
rect 546542 708444 581986 708680
rect 582222 708444 582306 708680
rect 582542 708444 589182 708680
rect 589418 708444 589502 708680
rect 589738 708444 589770 708680
rect -5846 708360 589770 708444
rect -5846 708124 -5814 708360
rect -5578 708124 -5494 708360
rect -5258 708124 5986 708360
rect 6222 708124 6306 708360
rect 6542 708124 41986 708360
rect 42222 708124 42306 708360
rect 42542 708124 77986 708360
rect 78222 708124 78306 708360
rect 78542 708124 113986 708360
rect 114222 708124 114306 708360
rect 114542 708124 149986 708360
rect 150222 708124 150306 708360
rect 150542 708124 185986 708360
rect 186222 708124 186306 708360
rect 186542 708124 221986 708360
rect 222222 708124 222306 708360
rect 222542 708124 257986 708360
rect 258222 708124 258306 708360
rect 258542 708124 293986 708360
rect 294222 708124 294306 708360
rect 294542 708124 329986 708360
rect 330222 708124 330306 708360
rect 330542 708124 365986 708360
rect 366222 708124 366306 708360
rect 366542 708124 401986 708360
rect 402222 708124 402306 708360
rect 402542 708124 437986 708360
rect 438222 708124 438306 708360
rect 438542 708124 473986 708360
rect 474222 708124 474306 708360
rect 474542 708124 509986 708360
rect 510222 708124 510306 708360
rect 510542 708124 545986 708360
rect 546222 708124 546306 708360
rect 546542 708124 581986 708360
rect 582222 708124 582306 708360
rect 582542 708124 589182 708360
rect 589418 708124 589502 708360
rect 589738 708124 589770 708360
rect -5846 708092 589770 708124
rect -4886 707720 588810 707752
rect -4886 707484 -4854 707720
rect -4618 707484 -4534 707720
rect -4298 707484 4746 707720
rect 4982 707484 5066 707720
rect 5302 707484 40746 707720
rect 40982 707484 41066 707720
rect 41302 707484 76746 707720
rect 76982 707484 77066 707720
rect 77302 707484 112746 707720
rect 112982 707484 113066 707720
rect 113302 707484 148746 707720
rect 148982 707484 149066 707720
rect 149302 707484 184746 707720
rect 184982 707484 185066 707720
rect 185302 707484 220746 707720
rect 220982 707484 221066 707720
rect 221302 707484 256746 707720
rect 256982 707484 257066 707720
rect 257302 707484 292746 707720
rect 292982 707484 293066 707720
rect 293302 707484 328746 707720
rect 328982 707484 329066 707720
rect 329302 707484 364746 707720
rect 364982 707484 365066 707720
rect 365302 707484 400746 707720
rect 400982 707484 401066 707720
rect 401302 707484 436746 707720
rect 436982 707484 437066 707720
rect 437302 707484 472746 707720
rect 472982 707484 473066 707720
rect 473302 707484 508746 707720
rect 508982 707484 509066 707720
rect 509302 707484 544746 707720
rect 544982 707484 545066 707720
rect 545302 707484 580746 707720
rect 580982 707484 581066 707720
rect 581302 707484 588222 707720
rect 588458 707484 588542 707720
rect 588778 707484 588810 707720
rect -4886 707400 588810 707484
rect -4886 707164 -4854 707400
rect -4618 707164 -4534 707400
rect -4298 707164 4746 707400
rect 4982 707164 5066 707400
rect 5302 707164 40746 707400
rect 40982 707164 41066 707400
rect 41302 707164 76746 707400
rect 76982 707164 77066 707400
rect 77302 707164 112746 707400
rect 112982 707164 113066 707400
rect 113302 707164 148746 707400
rect 148982 707164 149066 707400
rect 149302 707164 184746 707400
rect 184982 707164 185066 707400
rect 185302 707164 220746 707400
rect 220982 707164 221066 707400
rect 221302 707164 256746 707400
rect 256982 707164 257066 707400
rect 257302 707164 292746 707400
rect 292982 707164 293066 707400
rect 293302 707164 328746 707400
rect 328982 707164 329066 707400
rect 329302 707164 364746 707400
rect 364982 707164 365066 707400
rect 365302 707164 400746 707400
rect 400982 707164 401066 707400
rect 401302 707164 436746 707400
rect 436982 707164 437066 707400
rect 437302 707164 472746 707400
rect 472982 707164 473066 707400
rect 473302 707164 508746 707400
rect 508982 707164 509066 707400
rect 509302 707164 544746 707400
rect 544982 707164 545066 707400
rect 545302 707164 580746 707400
rect 580982 707164 581066 707400
rect 581302 707164 588222 707400
rect 588458 707164 588542 707400
rect 588778 707164 588810 707400
rect -4886 707132 588810 707164
rect -3926 706760 587850 706792
rect -3926 706524 -3894 706760
rect -3658 706524 -3574 706760
rect -3338 706524 3506 706760
rect 3742 706524 3826 706760
rect 4062 706524 39506 706760
rect 39742 706524 39826 706760
rect 40062 706524 75506 706760
rect 75742 706524 75826 706760
rect 76062 706524 111506 706760
rect 111742 706524 111826 706760
rect 112062 706524 147506 706760
rect 147742 706524 147826 706760
rect 148062 706524 183506 706760
rect 183742 706524 183826 706760
rect 184062 706524 219506 706760
rect 219742 706524 219826 706760
rect 220062 706524 255506 706760
rect 255742 706524 255826 706760
rect 256062 706524 291506 706760
rect 291742 706524 291826 706760
rect 292062 706524 327506 706760
rect 327742 706524 327826 706760
rect 328062 706524 363506 706760
rect 363742 706524 363826 706760
rect 364062 706524 399506 706760
rect 399742 706524 399826 706760
rect 400062 706524 435506 706760
rect 435742 706524 435826 706760
rect 436062 706524 471506 706760
rect 471742 706524 471826 706760
rect 472062 706524 507506 706760
rect 507742 706524 507826 706760
rect 508062 706524 543506 706760
rect 543742 706524 543826 706760
rect 544062 706524 579506 706760
rect 579742 706524 579826 706760
rect 580062 706524 587262 706760
rect 587498 706524 587582 706760
rect 587818 706524 587850 706760
rect -3926 706440 587850 706524
rect -3926 706204 -3894 706440
rect -3658 706204 -3574 706440
rect -3338 706204 3506 706440
rect 3742 706204 3826 706440
rect 4062 706204 39506 706440
rect 39742 706204 39826 706440
rect 40062 706204 75506 706440
rect 75742 706204 75826 706440
rect 76062 706204 111506 706440
rect 111742 706204 111826 706440
rect 112062 706204 147506 706440
rect 147742 706204 147826 706440
rect 148062 706204 183506 706440
rect 183742 706204 183826 706440
rect 184062 706204 219506 706440
rect 219742 706204 219826 706440
rect 220062 706204 255506 706440
rect 255742 706204 255826 706440
rect 256062 706204 291506 706440
rect 291742 706204 291826 706440
rect 292062 706204 327506 706440
rect 327742 706204 327826 706440
rect 328062 706204 363506 706440
rect 363742 706204 363826 706440
rect 364062 706204 399506 706440
rect 399742 706204 399826 706440
rect 400062 706204 435506 706440
rect 435742 706204 435826 706440
rect 436062 706204 471506 706440
rect 471742 706204 471826 706440
rect 472062 706204 507506 706440
rect 507742 706204 507826 706440
rect 508062 706204 543506 706440
rect 543742 706204 543826 706440
rect 544062 706204 579506 706440
rect 579742 706204 579826 706440
rect 580062 706204 587262 706440
rect 587498 706204 587582 706440
rect 587818 706204 587850 706440
rect -3926 706172 587850 706204
rect -2966 705800 586890 705832
rect -2966 705564 -2934 705800
rect -2698 705564 -2614 705800
rect -2378 705564 2266 705800
rect 2502 705564 2586 705800
rect 2822 705564 38266 705800
rect 38502 705564 38586 705800
rect 38822 705564 74266 705800
rect 74502 705564 74586 705800
rect 74822 705564 110266 705800
rect 110502 705564 110586 705800
rect 110822 705564 146266 705800
rect 146502 705564 146586 705800
rect 146822 705564 182266 705800
rect 182502 705564 182586 705800
rect 182822 705564 218266 705800
rect 218502 705564 218586 705800
rect 218822 705564 254266 705800
rect 254502 705564 254586 705800
rect 254822 705564 290266 705800
rect 290502 705564 290586 705800
rect 290822 705564 326266 705800
rect 326502 705564 326586 705800
rect 326822 705564 362266 705800
rect 362502 705564 362586 705800
rect 362822 705564 398266 705800
rect 398502 705564 398586 705800
rect 398822 705564 434266 705800
rect 434502 705564 434586 705800
rect 434822 705564 470266 705800
rect 470502 705564 470586 705800
rect 470822 705564 506266 705800
rect 506502 705564 506586 705800
rect 506822 705564 542266 705800
rect 542502 705564 542586 705800
rect 542822 705564 578266 705800
rect 578502 705564 578586 705800
rect 578822 705564 586302 705800
rect 586538 705564 586622 705800
rect 586858 705564 586890 705800
rect -2966 705480 586890 705564
rect -2966 705244 -2934 705480
rect -2698 705244 -2614 705480
rect -2378 705244 2266 705480
rect 2502 705244 2586 705480
rect 2822 705244 38266 705480
rect 38502 705244 38586 705480
rect 38822 705244 74266 705480
rect 74502 705244 74586 705480
rect 74822 705244 110266 705480
rect 110502 705244 110586 705480
rect 110822 705244 146266 705480
rect 146502 705244 146586 705480
rect 146822 705244 182266 705480
rect 182502 705244 182586 705480
rect 182822 705244 218266 705480
rect 218502 705244 218586 705480
rect 218822 705244 254266 705480
rect 254502 705244 254586 705480
rect 254822 705244 290266 705480
rect 290502 705244 290586 705480
rect 290822 705244 326266 705480
rect 326502 705244 326586 705480
rect 326822 705244 362266 705480
rect 362502 705244 362586 705480
rect 362822 705244 398266 705480
rect 398502 705244 398586 705480
rect 398822 705244 434266 705480
rect 434502 705244 434586 705480
rect 434822 705244 470266 705480
rect 470502 705244 470586 705480
rect 470822 705244 506266 705480
rect 506502 705244 506586 705480
rect 506822 705244 542266 705480
rect 542502 705244 542586 705480
rect 542822 705244 578266 705480
rect 578502 705244 578586 705480
rect 578822 705244 586302 705480
rect 586538 705244 586622 705480
rect 586858 705244 586890 705480
rect -2966 705212 586890 705244
rect -2006 704840 585930 704872
rect -2006 704604 -1974 704840
rect -1738 704604 -1654 704840
rect -1418 704604 1026 704840
rect 1262 704604 1346 704840
rect 1582 704604 37026 704840
rect 37262 704604 37346 704840
rect 37582 704604 73026 704840
rect 73262 704604 73346 704840
rect 73582 704604 109026 704840
rect 109262 704604 109346 704840
rect 109582 704604 145026 704840
rect 145262 704604 145346 704840
rect 145582 704604 181026 704840
rect 181262 704604 181346 704840
rect 181582 704604 217026 704840
rect 217262 704604 217346 704840
rect 217582 704604 253026 704840
rect 253262 704604 253346 704840
rect 253582 704604 289026 704840
rect 289262 704604 289346 704840
rect 289582 704604 325026 704840
rect 325262 704604 325346 704840
rect 325582 704604 361026 704840
rect 361262 704604 361346 704840
rect 361582 704604 397026 704840
rect 397262 704604 397346 704840
rect 397582 704604 433026 704840
rect 433262 704604 433346 704840
rect 433582 704604 469026 704840
rect 469262 704604 469346 704840
rect 469582 704604 505026 704840
rect 505262 704604 505346 704840
rect 505582 704604 541026 704840
rect 541262 704604 541346 704840
rect 541582 704604 577026 704840
rect 577262 704604 577346 704840
rect 577582 704604 585342 704840
rect 585578 704604 585662 704840
rect 585898 704604 585930 704840
rect -2006 704520 585930 704604
rect -2006 704284 -1974 704520
rect -1738 704284 -1654 704520
rect -1418 704284 1026 704520
rect 1262 704284 1346 704520
rect 1582 704284 37026 704520
rect 37262 704284 37346 704520
rect 37582 704284 73026 704520
rect 73262 704284 73346 704520
rect 73582 704284 109026 704520
rect 109262 704284 109346 704520
rect 109582 704284 145026 704520
rect 145262 704284 145346 704520
rect 145582 704284 181026 704520
rect 181262 704284 181346 704520
rect 181582 704284 217026 704520
rect 217262 704284 217346 704520
rect 217582 704284 253026 704520
rect 253262 704284 253346 704520
rect 253582 704284 289026 704520
rect 289262 704284 289346 704520
rect 289582 704284 325026 704520
rect 325262 704284 325346 704520
rect 325582 704284 361026 704520
rect 361262 704284 361346 704520
rect 361582 704284 397026 704520
rect 397262 704284 397346 704520
rect 397582 704284 433026 704520
rect 433262 704284 433346 704520
rect 433582 704284 469026 704520
rect 469262 704284 469346 704520
rect 469582 704284 505026 704520
rect 505262 704284 505346 704520
rect 505582 704284 541026 704520
rect 541262 704284 541346 704520
rect 541582 704284 577026 704520
rect 577262 704284 577346 704520
rect 577582 704284 585342 704520
rect 585578 704284 585662 704520
rect 585898 704284 585930 704520
rect -2006 704252 585930 704284
rect -8726 695336 592650 695368
rect -8726 695100 -8694 695336
rect -8458 695100 -8374 695336
rect -8138 695100 9706 695336
rect 9942 695100 10026 695336
rect 10262 695100 45706 695336
rect 45942 695100 46026 695336
rect 46262 695100 81706 695336
rect 81942 695100 82026 695336
rect 82262 695100 117706 695336
rect 117942 695100 118026 695336
rect 118262 695100 153706 695336
rect 153942 695100 154026 695336
rect 154262 695100 189706 695336
rect 189942 695100 190026 695336
rect 190262 695100 225706 695336
rect 225942 695100 226026 695336
rect 226262 695100 261706 695336
rect 261942 695100 262026 695336
rect 262262 695100 297706 695336
rect 297942 695100 298026 695336
rect 298262 695100 333706 695336
rect 333942 695100 334026 695336
rect 334262 695100 369706 695336
rect 369942 695100 370026 695336
rect 370262 695100 405706 695336
rect 405942 695100 406026 695336
rect 406262 695100 441706 695336
rect 441942 695100 442026 695336
rect 442262 695100 477706 695336
rect 477942 695100 478026 695336
rect 478262 695100 513706 695336
rect 513942 695100 514026 695336
rect 514262 695100 549706 695336
rect 549942 695100 550026 695336
rect 550262 695100 592062 695336
rect 592298 695100 592382 695336
rect 592618 695100 592650 695336
rect -8726 695016 592650 695100
rect -8726 694780 -8694 695016
rect -8458 694780 -8374 695016
rect -8138 694780 9706 695016
rect 9942 694780 10026 695016
rect 10262 694780 45706 695016
rect 45942 694780 46026 695016
rect 46262 694780 81706 695016
rect 81942 694780 82026 695016
rect 82262 694780 117706 695016
rect 117942 694780 118026 695016
rect 118262 694780 153706 695016
rect 153942 694780 154026 695016
rect 154262 694780 189706 695016
rect 189942 694780 190026 695016
rect 190262 694780 225706 695016
rect 225942 694780 226026 695016
rect 226262 694780 261706 695016
rect 261942 694780 262026 695016
rect 262262 694780 297706 695016
rect 297942 694780 298026 695016
rect 298262 694780 333706 695016
rect 333942 694780 334026 695016
rect 334262 694780 369706 695016
rect 369942 694780 370026 695016
rect 370262 694780 405706 695016
rect 405942 694780 406026 695016
rect 406262 694780 441706 695016
rect 441942 694780 442026 695016
rect 442262 694780 477706 695016
rect 477942 694780 478026 695016
rect 478262 694780 513706 695016
rect 513942 694780 514026 695016
rect 514262 694780 549706 695016
rect 549942 694780 550026 695016
rect 550262 694780 592062 695016
rect 592298 694780 592382 695016
rect 592618 694780 592650 695016
rect -8726 694748 592650 694780
rect -8726 694096 592650 694128
rect -8726 693860 -7734 694096
rect -7498 693860 -7414 694096
rect -7178 693860 8466 694096
rect 8702 693860 8786 694096
rect 9022 693860 44466 694096
rect 44702 693860 44786 694096
rect 45022 693860 80466 694096
rect 80702 693860 80786 694096
rect 81022 693860 116466 694096
rect 116702 693860 116786 694096
rect 117022 693860 152466 694096
rect 152702 693860 152786 694096
rect 153022 693860 188466 694096
rect 188702 693860 188786 694096
rect 189022 693860 224466 694096
rect 224702 693860 224786 694096
rect 225022 693860 260466 694096
rect 260702 693860 260786 694096
rect 261022 693860 296466 694096
rect 296702 693860 296786 694096
rect 297022 693860 332466 694096
rect 332702 693860 332786 694096
rect 333022 693860 368466 694096
rect 368702 693860 368786 694096
rect 369022 693860 404466 694096
rect 404702 693860 404786 694096
rect 405022 693860 440466 694096
rect 440702 693860 440786 694096
rect 441022 693860 476466 694096
rect 476702 693860 476786 694096
rect 477022 693860 512466 694096
rect 512702 693860 512786 694096
rect 513022 693860 548466 694096
rect 548702 693860 548786 694096
rect 549022 693860 591102 694096
rect 591338 693860 591422 694096
rect 591658 693860 592650 694096
rect -8726 693776 592650 693860
rect -8726 693540 -7734 693776
rect -7498 693540 -7414 693776
rect -7178 693540 8466 693776
rect 8702 693540 8786 693776
rect 9022 693540 44466 693776
rect 44702 693540 44786 693776
rect 45022 693540 80466 693776
rect 80702 693540 80786 693776
rect 81022 693540 116466 693776
rect 116702 693540 116786 693776
rect 117022 693540 152466 693776
rect 152702 693540 152786 693776
rect 153022 693540 188466 693776
rect 188702 693540 188786 693776
rect 189022 693540 224466 693776
rect 224702 693540 224786 693776
rect 225022 693540 260466 693776
rect 260702 693540 260786 693776
rect 261022 693540 296466 693776
rect 296702 693540 296786 693776
rect 297022 693540 332466 693776
rect 332702 693540 332786 693776
rect 333022 693540 368466 693776
rect 368702 693540 368786 693776
rect 369022 693540 404466 693776
rect 404702 693540 404786 693776
rect 405022 693540 440466 693776
rect 440702 693540 440786 693776
rect 441022 693540 476466 693776
rect 476702 693540 476786 693776
rect 477022 693540 512466 693776
rect 512702 693540 512786 693776
rect 513022 693540 548466 693776
rect 548702 693540 548786 693776
rect 549022 693540 591102 693776
rect 591338 693540 591422 693776
rect 591658 693540 592650 693776
rect -8726 693508 592650 693540
rect -8726 692856 592650 692888
rect -8726 692620 -6774 692856
rect -6538 692620 -6454 692856
rect -6218 692620 7226 692856
rect 7462 692620 7546 692856
rect 7782 692620 43226 692856
rect 43462 692620 43546 692856
rect 43782 692620 79226 692856
rect 79462 692620 79546 692856
rect 79782 692620 115226 692856
rect 115462 692620 115546 692856
rect 115782 692620 151226 692856
rect 151462 692620 151546 692856
rect 151782 692620 187226 692856
rect 187462 692620 187546 692856
rect 187782 692620 223226 692856
rect 223462 692620 223546 692856
rect 223782 692620 259226 692856
rect 259462 692620 259546 692856
rect 259782 692620 295226 692856
rect 295462 692620 295546 692856
rect 295782 692620 331226 692856
rect 331462 692620 331546 692856
rect 331782 692620 367226 692856
rect 367462 692620 367546 692856
rect 367782 692620 403226 692856
rect 403462 692620 403546 692856
rect 403782 692620 439226 692856
rect 439462 692620 439546 692856
rect 439782 692620 475226 692856
rect 475462 692620 475546 692856
rect 475782 692620 511226 692856
rect 511462 692620 511546 692856
rect 511782 692620 547226 692856
rect 547462 692620 547546 692856
rect 547782 692620 590142 692856
rect 590378 692620 590462 692856
rect 590698 692620 592650 692856
rect -8726 692536 592650 692620
rect -8726 692300 -6774 692536
rect -6538 692300 -6454 692536
rect -6218 692300 7226 692536
rect 7462 692300 7546 692536
rect 7782 692300 43226 692536
rect 43462 692300 43546 692536
rect 43782 692300 79226 692536
rect 79462 692300 79546 692536
rect 79782 692300 115226 692536
rect 115462 692300 115546 692536
rect 115782 692300 151226 692536
rect 151462 692300 151546 692536
rect 151782 692300 187226 692536
rect 187462 692300 187546 692536
rect 187782 692300 223226 692536
rect 223462 692300 223546 692536
rect 223782 692300 259226 692536
rect 259462 692300 259546 692536
rect 259782 692300 295226 692536
rect 295462 692300 295546 692536
rect 295782 692300 331226 692536
rect 331462 692300 331546 692536
rect 331782 692300 367226 692536
rect 367462 692300 367546 692536
rect 367782 692300 403226 692536
rect 403462 692300 403546 692536
rect 403782 692300 439226 692536
rect 439462 692300 439546 692536
rect 439782 692300 475226 692536
rect 475462 692300 475546 692536
rect 475782 692300 511226 692536
rect 511462 692300 511546 692536
rect 511782 692300 547226 692536
rect 547462 692300 547546 692536
rect 547782 692300 590142 692536
rect 590378 692300 590462 692536
rect 590698 692300 592650 692536
rect -8726 692268 592650 692300
rect -8726 691616 592650 691648
rect -8726 691380 -5814 691616
rect -5578 691380 -5494 691616
rect -5258 691380 5986 691616
rect 6222 691380 6306 691616
rect 6542 691380 41986 691616
rect 42222 691380 42306 691616
rect 42542 691380 77986 691616
rect 78222 691380 78306 691616
rect 78542 691380 113986 691616
rect 114222 691380 114306 691616
rect 114542 691380 149986 691616
rect 150222 691380 150306 691616
rect 150542 691380 185986 691616
rect 186222 691380 186306 691616
rect 186542 691380 221986 691616
rect 222222 691380 222306 691616
rect 222542 691380 257986 691616
rect 258222 691380 258306 691616
rect 258542 691380 293986 691616
rect 294222 691380 294306 691616
rect 294542 691380 329986 691616
rect 330222 691380 330306 691616
rect 330542 691380 365986 691616
rect 366222 691380 366306 691616
rect 366542 691380 401986 691616
rect 402222 691380 402306 691616
rect 402542 691380 437986 691616
rect 438222 691380 438306 691616
rect 438542 691380 473986 691616
rect 474222 691380 474306 691616
rect 474542 691380 509986 691616
rect 510222 691380 510306 691616
rect 510542 691380 545986 691616
rect 546222 691380 546306 691616
rect 546542 691380 581986 691616
rect 582222 691380 582306 691616
rect 582542 691380 589182 691616
rect 589418 691380 589502 691616
rect 589738 691380 592650 691616
rect -8726 691296 592650 691380
rect -8726 691060 -5814 691296
rect -5578 691060 -5494 691296
rect -5258 691060 5986 691296
rect 6222 691060 6306 691296
rect 6542 691060 41986 691296
rect 42222 691060 42306 691296
rect 42542 691060 77986 691296
rect 78222 691060 78306 691296
rect 78542 691060 113986 691296
rect 114222 691060 114306 691296
rect 114542 691060 149986 691296
rect 150222 691060 150306 691296
rect 150542 691060 185986 691296
rect 186222 691060 186306 691296
rect 186542 691060 221986 691296
rect 222222 691060 222306 691296
rect 222542 691060 257986 691296
rect 258222 691060 258306 691296
rect 258542 691060 293986 691296
rect 294222 691060 294306 691296
rect 294542 691060 329986 691296
rect 330222 691060 330306 691296
rect 330542 691060 365986 691296
rect 366222 691060 366306 691296
rect 366542 691060 401986 691296
rect 402222 691060 402306 691296
rect 402542 691060 437986 691296
rect 438222 691060 438306 691296
rect 438542 691060 473986 691296
rect 474222 691060 474306 691296
rect 474542 691060 509986 691296
rect 510222 691060 510306 691296
rect 510542 691060 545986 691296
rect 546222 691060 546306 691296
rect 546542 691060 581986 691296
rect 582222 691060 582306 691296
rect 582542 691060 589182 691296
rect 589418 691060 589502 691296
rect 589738 691060 592650 691296
rect -8726 691028 592650 691060
rect -8726 690376 592650 690408
rect -8726 690140 -4854 690376
rect -4618 690140 -4534 690376
rect -4298 690140 4746 690376
rect 4982 690140 5066 690376
rect 5302 690140 40746 690376
rect 40982 690140 41066 690376
rect 41302 690140 76746 690376
rect 76982 690140 77066 690376
rect 77302 690140 112746 690376
rect 112982 690140 113066 690376
rect 113302 690140 148746 690376
rect 148982 690140 149066 690376
rect 149302 690140 184746 690376
rect 184982 690140 185066 690376
rect 185302 690140 220746 690376
rect 220982 690140 221066 690376
rect 221302 690140 256746 690376
rect 256982 690140 257066 690376
rect 257302 690140 292746 690376
rect 292982 690140 293066 690376
rect 293302 690140 328746 690376
rect 328982 690140 329066 690376
rect 329302 690140 364746 690376
rect 364982 690140 365066 690376
rect 365302 690140 400746 690376
rect 400982 690140 401066 690376
rect 401302 690140 436746 690376
rect 436982 690140 437066 690376
rect 437302 690140 472746 690376
rect 472982 690140 473066 690376
rect 473302 690140 508746 690376
rect 508982 690140 509066 690376
rect 509302 690140 544746 690376
rect 544982 690140 545066 690376
rect 545302 690140 580746 690376
rect 580982 690140 581066 690376
rect 581302 690140 588222 690376
rect 588458 690140 588542 690376
rect 588778 690140 592650 690376
rect -8726 690056 592650 690140
rect -8726 689820 -4854 690056
rect -4618 689820 -4534 690056
rect -4298 689820 4746 690056
rect 4982 689820 5066 690056
rect 5302 689820 40746 690056
rect 40982 689820 41066 690056
rect 41302 689820 76746 690056
rect 76982 689820 77066 690056
rect 77302 689820 112746 690056
rect 112982 689820 113066 690056
rect 113302 689820 148746 690056
rect 148982 689820 149066 690056
rect 149302 689820 184746 690056
rect 184982 689820 185066 690056
rect 185302 689820 220746 690056
rect 220982 689820 221066 690056
rect 221302 689820 256746 690056
rect 256982 689820 257066 690056
rect 257302 689820 292746 690056
rect 292982 689820 293066 690056
rect 293302 689820 328746 690056
rect 328982 689820 329066 690056
rect 329302 689820 364746 690056
rect 364982 689820 365066 690056
rect 365302 689820 400746 690056
rect 400982 689820 401066 690056
rect 401302 689820 436746 690056
rect 436982 689820 437066 690056
rect 437302 689820 472746 690056
rect 472982 689820 473066 690056
rect 473302 689820 508746 690056
rect 508982 689820 509066 690056
rect 509302 689820 544746 690056
rect 544982 689820 545066 690056
rect 545302 689820 580746 690056
rect 580982 689820 581066 690056
rect 581302 689820 588222 690056
rect 588458 689820 588542 690056
rect 588778 689820 592650 690056
rect -8726 689788 592650 689820
rect -8726 689136 592650 689168
rect -8726 688900 -3894 689136
rect -3658 688900 -3574 689136
rect -3338 688900 3506 689136
rect 3742 688900 3826 689136
rect 4062 688900 39506 689136
rect 39742 688900 39826 689136
rect 40062 688900 75506 689136
rect 75742 688900 75826 689136
rect 76062 688900 111506 689136
rect 111742 688900 111826 689136
rect 112062 688900 147506 689136
rect 147742 688900 147826 689136
rect 148062 688900 183506 689136
rect 183742 688900 183826 689136
rect 184062 688900 219506 689136
rect 219742 688900 219826 689136
rect 220062 688900 255506 689136
rect 255742 688900 255826 689136
rect 256062 688900 291506 689136
rect 291742 688900 291826 689136
rect 292062 688900 327506 689136
rect 327742 688900 327826 689136
rect 328062 688900 363506 689136
rect 363742 688900 363826 689136
rect 364062 688900 399506 689136
rect 399742 688900 399826 689136
rect 400062 688900 435506 689136
rect 435742 688900 435826 689136
rect 436062 688900 471506 689136
rect 471742 688900 471826 689136
rect 472062 688900 507506 689136
rect 507742 688900 507826 689136
rect 508062 688900 543506 689136
rect 543742 688900 543826 689136
rect 544062 688900 579506 689136
rect 579742 688900 579826 689136
rect 580062 688900 587262 689136
rect 587498 688900 587582 689136
rect 587818 688900 592650 689136
rect -8726 688816 592650 688900
rect -8726 688580 -3894 688816
rect -3658 688580 -3574 688816
rect -3338 688580 3506 688816
rect 3742 688580 3826 688816
rect 4062 688580 39506 688816
rect 39742 688580 39826 688816
rect 40062 688580 75506 688816
rect 75742 688580 75826 688816
rect 76062 688580 111506 688816
rect 111742 688580 111826 688816
rect 112062 688580 147506 688816
rect 147742 688580 147826 688816
rect 148062 688580 183506 688816
rect 183742 688580 183826 688816
rect 184062 688580 219506 688816
rect 219742 688580 219826 688816
rect 220062 688580 255506 688816
rect 255742 688580 255826 688816
rect 256062 688580 291506 688816
rect 291742 688580 291826 688816
rect 292062 688580 327506 688816
rect 327742 688580 327826 688816
rect 328062 688580 363506 688816
rect 363742 688580 363826 688816
rect 364062 688580 399506 688816
rect 399742 688580 399826 688816
rect 400062 688580 435506 688816
rect 435742 688580 435826 688816
rect 436062 688580 471506 688816
rect 471742 688580 471826 688816
rect 472062 688580 507506 688816
rect 507742 688580 507826 688816
rect 508062 688580 543506 688816
rect 543742 688580 543826 688816
rect 544062 688580 579506 688816
rect 579742 688580 579826 688816
rect 580062 688580 587262 688816
rect 587498 688580 587582 688816
rect 587818 688580 592650 688816
rect -8726 688548 592650 688580
rect -8726 687896 592650 687928
rect -8726 687660 -2934 687896
rect -2698 687660 -2614 687896
rect -2378 687660 2266 687896
rect 2502 687660 2586 687896
rect 2822 687660 38266 687896
rect 38502 687660 38586 687896
rect 38822 687660 74266 687896
rect 74502 687660 74586 687896
rect 74822 687660 110266 687896
rect 110502 687660 110586 687896
rect 110822 687660 146266 687896
rect 146502 687660 146586 687896
rect 146822 687660 182266 687896
rect 182502 687660 182586 687896
rect 182822 687660 218266 687896
rect 218502 687660 218586 687896
rect 218822 687660 254266 687896
rect 254502 687660 254586 687896
rect 254822 687660 290266 687896
rect 290502 687660 290586 687896
rect 290822 687660 326266 687896
rect 326502 687660 326586 687896
rect 326822 687660 362266 687896
rect 362502 687660 362586 687896
rect 362822 687660 398266 687896
rect 398502 687660 398586 687896
rect 398822 687660 434266 687896
rect 434502 687660 434586 687896
rect 434822 687660 470266 687896
rect 470502 687660 470586 687896
rect 470822 687660 506266 687896
rect 506502 687660 506586 687896
rect 506822 687660 542266 687896
rect 542502 687660 542586 687896
rect 542822 687660 578266 687896
rect 578502 687660 578586 687896
rect 578822 687660 586302 687896
rect 586538 687660 586622 687896
rect 586858 687660 592650 687896
rect -8726 687576 592650 687660
rect -8726 687340 -2934 687576
rect -2698 687340 -2614 687576
rect -2378 687340 2266 687576
rect 2502 687340 2586 687576
rect 2822 687340 38266 687576
rect 38502 687340 38586 687576
rect 38822 687340 74266 687576
rect 74502 687340 74586 687576
rect 74822 687340 110266 687576
rect 110502 687340 110586 687576
rect 110822 687340 146266 687576
rect 146502 687340 146586 687576
rect 146822 687340 182266 687576
rect 182502 687340 182586 687576
rect 182822 687340 218266 687576
rect 218502 687340 218586 687576
rect 218822 687340 254266 687576
rect 254502 687340 254586 687576
rect 254822 687340 290266 687576
rect 290502 687340 290586 687576
rect 290822 687340 326266 687576
rect 326502 687340 326586 687576
rect 326822 687340 362266 687576
rect 362502 687340 362586 687576
rect 362822 687340 398266 687576
rect 398502 687340 398586 687576
rect 398822 687340 434266 687576
rect 434502 687340 434586 687576
rect 434822 687340 470266 687576
rect 470502 687340 470586 687576
rect 470822 687340 506266 687576
rect 506502 687340 506586 687576
rect 506822 687340 542266 687576
rect 542502 687340 542586 687576
rect 542822 687340 578266 687576
rect 578502 687340 578586 687576
rect 578822 687340 586302 687576
rect 586538 687340 586622 687576
rect 586858 687340 592650 687576
rect -8726 687308 592650 687340
rect -8726 686656 592650 686688
rect -8726 686420 -1974 686656
rect -1738 686420 -1654 686656
rect -1418 686420 1026 686656
rect 1262 686420 1346 686656
rect 1582 686420 37026 686656
rect 37262 686420 37346 686656
rect 37582 686420 73026 686656
rect 73262 686420 73346 686656
rect 73582 686420 109026 686656
rect 109262 686420 109346 686656
rect 109582 686420 145026 686656
rect 145262 686420 145346 686656
rect 145582 686420 181026 686656
rect 181262 686420 181346 686656
rect 181582 686420 217026 686656
rect 217262 686420 217346 686656
rect 217582 686420 253026 686656
rect 253262 686420 253346 686656
rect 253582 686420 289026 686656
rect 289262 686420 289346 686656
rect 289582 686420 325026 686656
rect 325262 686420 325346 686656
rect 325582 686420 361026 686656
rect 361262 686420 361346 686656
rect 361582 686420 397026 686656
rect 397262 686420 397346 686656
rect 397582 686420 433026 686656
rect 433262 686420 433346 686656
rect 433582 686420 469026 686656
rect 469262 686420 469346 686656
rect 469582 686420 505026 686656
rect 505262 686420 505346 686656
rect 505582 686420 541026 686656
rect 541262 686420 541346 686656
rect 541582 686420 577026 686656
rect 577262 686420 577346 686656
rect 577582 686420 585342 686656
rect 585578 686420 585662 686656
rect 585898 686420 592650 686656
rect -8726 686336 592650 686420
rect -8726 686100 -1974 686336
rect -1738 686100 -1654 686336
rect -1418 686100 1026 686336
rect 1262 686100 1346 686336
rect 1582 686100 37026 686336
rect 37262 686100 37346 686336
rect 37582 686100 73026 686336
rect 73262 686100 73346 686336
rect 73582 686100 109026 686336
rect 109262 686100 109346 686336
rect 109582 686100 145026 686336
rect 145262 686100 145346 686336
rect 145582 686100 181026 686336
rect 181262 686100 181346 686336
rect 181582 686100 217026 686336
rect 217262 686100 217346 686336
rect 217582 686100 253026 686336
rect 253262 686100 253346 686336
rect 253582 686100 289026 686336
rect 289262 686100 289346 686336
rect 289582 686100 325026 686336
rect 325262 686100 325346 686336
rect 325582 686100 361026 686336
rect 361262 686100 361346 686336
rect 361582 686100 397026 686336
rect 397262 686100 397346 686336
rect 397582 686100 433026 686336
rect 433262 686100 433346 686336
rect 433582 686100 469026 686336
rect 469262 686100 469346 686336
rect 469582 686100 505026 686336
rect 505262 686100 505346 686336
rect 505582 686100 541026 686336
rect 541262 686100 541346 686336
rect 541582 686100 577026 686336
rect 577262 686100 577346 686336
rect 577582 686100 585342 686336
rect 585578 686100 585662 686336
rect 585898 686100 592650 686336
rect -8726 686068 592650 686100
rect -8726 659336 592650 659368
rect -8726 659100 -8694 659336
rect -8458 659100 -8374 659336
rect -8138 659100 9706 659336
rect 9942 659100 10026 659336
rect 10262 659100 45706 659336
rect 45942 659100 46026 659336
rect 46262 659100 81706 659336
rect 81942 659100 82026 659336
rect 82262 659100 117706 659336
rect 117942 659100 118026 659336
rect 118262 659100 153706 659336
rect 153942 659100 154026 659336
rect 154262 659100 189706 659336
rect 189942 659100 190026 659336
rect 190262 659100 225706 659336
rect 225942 659100 226026 659336
rect 226262 659100 261706 659336
rect 261942 659100 262026 659336
rect 262262 659100 297706 659336
rect 297942 659100 298026 659336
rect 298262 659100 333706 659336
rect 333942 659100 334026 659336
rect 334262 659100 369706 659336
rect 369942 659100 370026 659336
rect 370262 659100 405706 659336
rect 405942 659100 406026 659336
rect 406262 659100 441706 659336
rect 441942 659100 442026 659336
rect 442262 659100 477706 659336
rect 477942 659100 478026 659336
rect 478262 659100 513706 659336
rect 513942 659100 514026 659336
rect 514262 659100 549706 659336
rect 549942 659100 550026 659336
rect 550262 659100 592062 659336
rect 592298 659100 592382 659336
rect 592618 659100 592650 659336
rect -8726 659016 592650 659100
rect -8726 658780 -8694 659016
rect -8458 658780 -8374 659016
rect -8138 658780 9706 659016
rect 9942 658780 10026 659016
rect 10262 658780 45706 659016
rect 45942 658780 46026 659016
rect 46262 658780 81706 659016
rect 81942 658780 82026 659016
rect 82262 658780 117706 659016
rect 117942 658780 118026 659016
rect 118262 658780 153706 659016
rect 153942 658780 154026 659016
rect 154262 658780 189706 659016
rect 189942 658780 190026 659016
rect 190262 658780 225706 659016
rect 225942 658780 226026 659016
rect 226262 658780 261706 659016
rect 261942 658780 262026 659016
rect 262262 658780 297706 659016
rect 297942 658780 298026 659016
rect 298262 658780 333706 659016
rect 333942 658780 334026 659016
rect 334262 658780 369706 659016
rect 369942 658780 370026 659016
rect 370262 658780 405706 659016
rect 405942 658780 406026 659016
rect 406262 658780 441706 659016
rect 441942 658780 442026 659016
rect 442262 658780 477706 659016
rect 477942 658780 478026 659016
rect 478262 658780 513706 659016
rect 513942 658780 514026 659016
rect 514262 658780 549706 659016
rect 549942 658780 550026 659016
rect 550262 658780 592062 659016
rect 592298 658780 592382 659016
rect 592618 658780 592650 659016
rect -8726 658748 592650 658780
rect -8726 658096 592650 658128
rect -8726 657860 -7734 658096
rect -7498 657860 -7414 658096
rect -7178 657860 8466 658096
rect 8702 657860 8786 658096
rect 9022 657860 44466 658096
rect 44702 657860 44786 658096
rect 45022 657860 80466 658096
rect 80702 657860 80786 658096
rect 81022 657860 116466 658096
rect 116702 657860 116786 658096
rect 117022 657860 152466 658096
rect 152702 657860 152786 658096
rect 153022 657860 188466 658096
rect 188702 657860 188786 658096
rect 189022 657860 224466 658096
rect 224702 657860 224786 658096
rect 225022 657860 260466 658096
rect 260702 657860 260786 658096
rect 261022 657860 296466 658096
rect 296702 657860 296786 658096
rect 297022 657860 332466 658096
rect 332702 657860 332786 658096
rect 333022 657860 368466 658096
rect 368702 657860 368786 658096
rect 369022 657860 404466 658096
rect 404702 657860 404786 658096
rect 405022 657860 440466 658096
rect 440702 657860 440786 658096
rect 441022 657860 476466 658096
rect 476702 657860 476786 658096
rect 477022 657860 512466 658096
rect 512702 657860 512786 658096
rect 513022 657860 548466 658096
rect 548702 657860 548786 658096
rect 549022 657860 591102 658096
rect 591338 657860 591422 658096
rect 591658 657860 592650 658096
rect -8726 657776 592650 657860
rect -8726 657540 -7734 657776
rect -7498 657540 -7414 657776
rect -7178 657540 8466 657776
rect 8702 657540 8786 657776
rect 9022 657540 44466 657776
rect 44702 657540 44786 657776
rect 45022 657540 80466 657776
rect 80702 657540 80786 657776
rect 81022 657540 116466 657776
rect 116702 657540 116786 657776
rect 117022 657540 152466 657776
rect 152702 657540 152786 657776
rect 153022 657540 188466 657776
rect 188702 657540 188786 657776
rect 189022 657540 224466 657776
rect 224702 657540 224786 657776
rect 225022 657540 260466 657776
rect 260702 657540 260786 657776
rect 261022 657540 296466 657776
rect 296702 657540 296786 657776
rect 297022 657540 332466 657776
rect 332702 657540 332786 657776
rect 333022 657540 368466 657776
rect 368702 657540 368786 657776
rect 369022 657540 404466 657776
rect 404702 657540 404786 657776
rect 405022 657540 440466 657776
rect 440702 657540 440786 657776
rect 441022 657540 476466 657776
rect 476702 657540 476786 657776
rect 477022 657540 512466 657776
rect 512702 657540 512786 657776
rect 513022 657540 548466 657776
rect 548702 657540 548786 657776
rect 549022 657540 591102 657776
rect 591338 657540 591422 657776
rect 591658 657540 592650 657776
rect -8726 657508 592650 657540
rect -8726 656856 592650 656888
rect -8726 656620 -6774 656856
rect -6538 656620 -6454 656856
rect -6218 656620 7226 656856
rect 7462 656620 7546 656856
rect 7782 656620 43226 656856
rect 43462 656620 43546 656856
rect 43782 656620 79226 656856
rect 79462 656620 79546 656856
rect 79782 656620 115226 656856
rect 115462 656620 115546 656856
rect 115782 656620 151226 656856
rect 151462 656620 151546 656856
rect 151782 656620 187226 656856
rect 187462 656620 187546 656856
rect 187782 656620 223226 656856
rect 223462 656620 223546 656856
rect 223782 656620 259226 656856
rect 259462 656620 259546 656856
rect 259782 656620 295226 656856
rect 295462 656620 295546 656856
rect 295782 656620 331226 656856
rect 331462 656620 331546 656856
rect 331782 656620 367226 656856
rect 367462 656620 367546 656856
rect 367782 656620 403226 656856
rect 403462 656620 403546 656856
rect 403782 656620 439226 656856
rect 439462 656620 439546 656856
rect 439782 656620 475226 656856
rect 475462 656620 475546 656856
rect 475782 656620 511226 656856
rect 511462 656620 511546 656856
rect 511782 656620 547226 656856
rect 547462 656620 547546 656856
rect 547782 656620 590142 656856
rect 590378 656620 590462 656856
rect 590698 656620 592650 656856
rect -8726 656536 592650 656620
rect -8726 656300 -6774 656536
rect -6538 656300 -6454 656536
rect -6218 656300 7226 656536
rect 7462 656300 7546 656536
rect 7782 656300 43226 656536
rect 43462 656300 43546 656536
rect 43782 656300 79226 656536
rect 79462 656300 79546 656536
rect 79782 656300 115226 656536
rect 115462 656300 115546 656536
rect 115782 656300 151226 656536
rect 151462 656300 151546 656536
rect 151782 656300 187226 656536
rect 187462 656300 187546 656536
rect 187782 656300 223226 656536
rect 223462 656300 223546 656536
rect 223782 656300 259226 656536
rect 259462 656300 259546 656536
rect 259782 656300 295226 656536
rect 295462 656300 295546 656536
rect 295782 656300 331226 656536
rect 331462 656300 331546 656536
rect 331782 656300 367226 656536
rect 367462 656300 367546 656536
rect 367782 656300 403226 656536
rect 403462 656300 403546 656536
rect 403782 656300 439226 656536
rect 439462 656300 439546 656536
rect 439782 656300 475226 656536
rect 475462 656300 475546 656536
rect 475782 656300 511226 656536
rect 511462 656300 511546 656536
rect 511782 656300 547226 656536
rect 547462 656300 547546 656536
rect 547782 656300 590142 656536
rect 590378 656300 590462 656536
rect 590698 656300 592650 656536
rect -8726 656268 592650 656300
rect -8726 655616 592650 655648
rect -8726 655380 -5814 655616
rect -5578 655380 -5494 655616
rect -5258 655380 5986 655616
rect 6222 655380 6306 655616
rect 6542 655380 41986 655616
rect 42222 655380 42306 655616
rect 42542 655380 77986 655616
rect 78222 655380 78306 655616
rect 78542 655380 113986 655616
rect 114222 655380 114306 655616
rect 114542 655380 149986 655616
rect 150222 655380 150306 655616
rect 150542 655380 185986 655616
rect 186222 655380 186306 655616
rect 186542 655380 221986 655616
rect 222222 655380 222306 655616
rect 222542 655380 257986 655616
rect 258222 655380 258306 655616
rect 258542 655380 293986 655616
rect 294222 655380 294306 655616
rect 294542 655380 329986 655616
rect 330222 655380 330306 655616
rect 330542 655380 365986 655616
rect 366222 655380 366306 655616
rect 366542 655380 401986 655616
rect 402222 655380 402306 655616
rect 402542 655380 437986 655616
rect 438222 655380 438306 655616
rect 438542 655380 473986 655616
rect 474222 655380 474306 655616
rect 474542 655380 509986 655616
rect 510222 655380 510306 655616
rect 510542 655380 545986 655616
rect 546222 655380 546306 655616
rect 546542 655380 581986 655616
rect 582222 655380 582306 655616
rect 582542 655380 589182 655616
rect 589418 655380 589502 655616
rect 589738 655380 592650 655616
rect -8726 655296 592650 655380
rect -8726 655060 -5814 655296
rect -5578 655060 -5494 655296
rect -5258 655060 5986 655296
rect 6222 655060 6306 655296
rect 6542 655060 41986 655296
rect 42222 655060 42306 655296
rect 42542 655060 77986 655296
rect 78222 655060 78306 655296
rect 78542 655060 113986 655296
rect 114222 655060 114306 655296
rect 114542 655060 149986 655296
rect 150222 655060 150306 655296
rect 150542 655060 185986 655296
rect 186222 655060 186306 655296
rect 186542 655060 221986 655296
rect 222222 655060 222306 655296
rect 222542 655060 257986 655296
rect 258222 655060 258306 655296
rect 258542 655060 293986 655296
rect 294222 655060 294306 655296
rect 294542 655060 329986 655296
rect 330222 655060 330306 655296
rect 330542 655060 365986 655296
rect 366222 655060 366306 655296
rect 366542 655060 401986 655296
rect 402222 655060 402306 655296
rect 402542 655060 437986 655296
rect 438222 655060 438306 655296
rect 438542 655060 473986 655296
rect 474222 655060 474306 655296
rect 474542 655060 509986 655296
rect 510222 655060 510306 655296
rect 510542 655060 545986 655296
rect 546222 655060 546306 655296
rect 546542 655060 581986 655296
rect 582222 655060 582306 655296
rect 582542 655060 589182 655296
rect 589418 655060 589502 655296
rect 589738 655060 592650 655296
rect -8726 655028 592650 655060
rect -8726 654376 592650 654408
rect -8726 654140 -4854 654376
rect -4618 654140 -4534 654376
rect -4298 654140 4746 654376
rect 4982 654140 5066 654376
rect 5302 654140 40746 654376
rect 40982 654140 41066 654376
rect 41302 654140 76746 654376
rect 76982 654140 77066 654376
rect 77302 654140 112746 654376
rect 112982 654140 113066 654376
rect 113302 654140 148746 654376
rect 148982 654140 149066 654376
rect 149302 654140 184746 654376
rect 184982 654140 185066 654376
rect 185302 654140 220746 654376
rect 220982 654140 221066 654376
rect 221302 654140 256746 654376
rect 256982 654140 257066 654376
rect 257302 654140 292746 654376
rect 292982 654140 293066 654376
rect 293302 654140 328746 654376
rect 328982 654140 329066 654376
rect 329302 654140 364746 654376
rect 364982 654140 365066 654376
rect 365302 654140 400746 654376
rect 400982 654140 401066 654376
rect 401302 654140 436746 654376
rect 436982 654140 437066 654376
rect 437302 654140 472746 654376
rect 472982 654140 473066 654376
rect 473302 654140 508746 654376
rect 508982 654140 509066 654376
rect 509302 654140 544746 654376
rect 544982 654140 545066 654376
rect 545302 654140 580746 654376
rect 580982 654140 581066 654376
rect 581302 654140 588222 654376
rect 588458 654140 588542 654376
rect 588778 654140 592650 654376
rect -8726 654056 592650 654140
rect -8726 653820 -4854 654056
rect -4618 653820 -4534 654056
rect -4298 653820 4746 654056
rect 4982 653820 5066 654056
rect 5302 653820 40746 654056
rect 40982 653820 41066 654056
rect 41302 653820 76746 654056
rect 76982 653820 77066 654056
rect 77302 653820 112746 654056
rect 112982 653820 113066 654056
rect 113302 653820 148746 654056
rect 148982 653820 149066 654056
rect 149302 653820 184746 654056
rect 184982 653820 185066 654056
rect 185302 653820 220746 654056
rect 220982 653820 221066 654056
rect 221302 653820 256746 654056
rect 256982 653820 257066 654056
rect 257302 653820 292746 654056
rect 292982 653820 293066 654056
rect 293302 653820 328746 654056
rect 328982 653820 329066 654056
rect 329302 653820 364746 654056
rect 364982 653820 365066 654056
rect 365302 653820 400746 654056
rect 400982 653820 401066 654056
rect 401302 653820 436746 654056
rect 436982 653820 437066 654056
rect 437302 653820 472746 654056
rect 472982 653820 473066 654056
rect 473302 653820 508746 654056
rect 508982 653820 509066 654056
rect 509302 653820 544746 654056
rect 544982 653820 545066 654056
rect 545302 653820 580746 654056
rect 580982 653820 581066 654056
rect 581302 653820 588222 654056
rect 588458 653820 588542 654056
rect 588778 653820 592650 654056
rect -8726 653788 592650 653820
rect -8726 653136 592650 653168
rect -8726 652900 -3894 653136
rect -3658 652900 -3574 653136
rect -3338 652900 3506 653136
rect 3742 652900 3826 653136
rect 4062 652900 39506 653136
rect 39742 652900 39826 653136
rect 40062 652900 75506 653136
rect 75742 652900 75826 653136
rect 76062 652900 111506 653136
rect 111742 652900 111826 653136
rect 112062 652900 147506 653136
rect 147742 652900 147826 653136
rect 148062 652900 183506 653136
rect 183742 652900 183826 653136
rect 184062 652900 219506 653136
rect 219742 652900 219826 653136
rect 220062 652900 255506 653136
rect 255742 652900 255826 653136
rect 256062 652900 291506 653136
rect 291742 652900 291826 653136
rect 292062 652900 327506 653136
rect 327742 652900 327826 653136
rect 328062 652900 363506 653136
rect 363742 652900 363826 653136
rect 364062 652900 399506 653136
rect 399742 652900 399826 653136
rect 400062 652900 435506 653136
rect 435742 652900 435826 653136
rect 436062 652900 471506 653136
rect 471742 652900 471826 653136
rect 472062 652900 507506 653136
rect 507742 652900 507826 653136
rect 508062 652900 543506 653136
rect 543742 652900 543826 653136
rect 544062 652900 579506 653136
rect 579742 652900 579826 653136
rect 580062 652900 587262 653136
rect 587498 652900 587582 653136
rect 587818 652900 592650 653136
rect -8726 652816 592650 652900
rect -8726 652580 -3894 652816
rect -3658 652580 -3574 652816
rect -3338 652580 3506 652816
rect 3742 652580 3826 652816
rect 4062 652580 39506 652816
rect 39742 652580 39826 652816
rect 40062 652580 75506 652816
rect 75742 652580 75826 652816
rect 76062 652580 111506 652816
rect 111742 652580 111826 652816
rect 112062 652580 147506 652816
rect 147742 652580 147826 652816
rect 148062 652580 183506 652816
rect 183742 652580 183826 652816
rect 184062 652580 219506 652816
rect 219742 652580 219826 652816
rect 220062 652580 255506 652816
rect 255742 652580 255826 652816
rect 256062 652580 291506 652816
rect 291742 652580 291826 652816
rect 292062 652580 327506 652816
rect 327742 652580 327826 652816
rect 328062 652580 363506 652816
rect 363742 652580 363826 652816
rect 364062 652580 399506 652816
rect 399742 652580 399826 652816
rect 400062 652580 435506 652816
rect 435742 652580 435826 652816
rect 436062 652580 471506 652816
rect 471742 652580 471826 652816
rect 472062 652580 507506 652816
rect 507742 652580 507826 652816
rect 508062 652580 543506 652816
rect 543742 652580 543826 652816
rect 544062 652580 579506 652816
rect 579742 652580 579826 652816
rect 580062 652580 587262 652816
rect 587498 652580 587582 652816
rect 587818 652580 592650 652816
rect -8726 652548 592650 652580
rect -8726 651896 592650 651928
rect -8726 651660 -2934 651896
rect -2698 651660 -2614 651896
rect -2378 651660 2266 651896
rect 2502 651660 2586 651896
rect 2822 651660 38266 651896
rect 38502 651660 38586 651896
rect 38822 651660 74266 651896
rect 74502 651660 74586 651896
rect 74822 651660 110266 651896
rect 110502 651660 110586 651896
rect 110822 651660 146266 651896
rect 146502 651660 146586 651896
rect 146822 651660 182266 651896
rect 182502 651660 182586 651896
rect 182822 651660 218266 651896
rect 218502 651660 218586 651896
rect 218822 651660 254266 651896
rect 254502 651660 254586 651896
rect 254822 651660 290266 651896
rect 290502 651660 290586 651896
rect 290822 651660 326266 651896
rect 326502 651660 326586 651896
rect 326822 651660 362266 651896
rect 362502 651660 362586 651896
rect 362822 651660 398266 651896
rect 398502 651660 398586 651896
rect 398822 651660 434266 651896
rect 434502 651660 434586 651896
rect 434822 651660 470266 651896
rect 470502 651660 470586 651896
rect 470822 651660 506266 651896
rect 506502 651660 506586 651896
rect 506822 651660 542266 651896
rect 542502 651660 542586 651896
rect 542822 651660 578266 651896
rect 578502 651660 578586 651896
rect 578822 651660 586302 651896
rect 586538 651660 586622 651896
rect 586858 651660 592650 651896
rect -8726 651576 592650 651660
rect -8726 651340 -2934 651576
rect -2698 651340 -2614 651576
rect -2378 651340 2266 651576
rect 2502 651340 2586 651576
rect 2822 651340 38266 651576
rect 38502 651340 38586 651576
rect 38822 651340 74266 651576
rect 74502 651340 74586 651576
rect 74822 651340 110266 651576
rect 110502 651340 110586 651576
rect 110822 651340 146266 651576
rect 146502 651340 146586 651576
rect 146822 651340 182266 651576
rect 182502 651340 182586 651576
rect 182822 651340 218266 651576
rect 218502 651340 218586 651576
rect 218822 651340 254266 651576
rect 254502 651340 254586 651576
rect 254822 651340 290266 651576
rect 290502 651340 290586 651576
rect 290822 651340 326266 651576
rect 326502 651340 326586 651576
rect 326822 651340 362266 651576
rect 362502 651340 362586 651576
rect 362822 651340 398266 651576
rect 398502 651340 398586 651576
rect 398822 651340 434266 651576
rect 434502 651340 434586 651576
rect 434822 651340 470266 651576
rect 470502 651340 470586 651576
rect 470822 651340 506266 651576
rect 506502 651340 506586 651576
rect 506822 651340 542266 651576
rect 542502 651340 542586 651576
rect 542822 651340 578266 651576
rect 578502 651340 578586 651576
rect 578822 651340 586302 651576
rect 586538 651340 586622 651576
rect 586858 651340 592650 651576
rect -8726 651308 592650 651340
rect -8726 650656 592650 650688
rect -8726 650420 -1974 650656
rect -1738 650420 -1654 650656
rect -1418 650420 1026 650656
rect 1262 650420 1346 650656
rect 1582 650420 37026 650656
rect 37262 650420 37346 650656
rect 37582 650420 73026 650656
rect 73262 650420 73346 650656
rect 73582 650420 109026 650656
rect 109262 650420 109346 650656
rect 109582 650420 145026 650656
rect 145262 650420 145346 650656
rect 145582 650420 181026 650656
rect 181262 650420 181346 650656
rect 181582 650420 217026 650656
rect 217262 650420 217346 650656
rect 217582 650420 253026 650656
rect 253262 650420 253346 650656
rect 253582 650420 289026 650656
rect 289262 650420 289346 650656
rect 289582 650420 325026 650656
rect 325262 650420 325346 650656
rect 325582 650420 361026 650656
rect 361262 650420 361346 650656
rect 361582 650420 397026 650656
rect 397262 650420 397346 650656
rect 397582 650420 433026 650656
rect 433262 650420 433346 650656
rect 433582 650420 469026 650656
rect 469262 650420 469346 650656
rect 469582 650420 505026 650656
rect 505262 650420 505346 650656
rect 505582 650420 541026 650656
rect 541262 650420 541346 650656
rect 541582 650420 577026 650656
rect 577262 650420 577346 650656
rect 577582 650420 585342 650656
rect 585578 650420 585662 650656
rect 585898 650420 592650 650656
rect -8726 650336 592650 650420
rect -8726 650100 -1974 650336
rect -1738 650100 -1654 650336
rect -1418 650100 1026 650336
rect 1262 650100 1346 650336
rect 1582 650100 37026 650336
rect 37262 650100 37346 650336
rect 37582 650100 73026 650336
rect 73262 650100 73346 650336
rect 73582 650100 109026 650336
rect 109262 650100 109346 650336
rect 109582 650100 145026 650336
rect 145262 650100 145346 650336
rect 145582 650100 181026 650336
rect 181262 650100 181346 650336
rect 181582 650100 217026 650336
rect 217262 650100 217346 650336
rect 217582 650100 253026 650336
rect 253262 650100 253346 650336
rect 253582 650100 289026 650336
rect 289262 650100 289346 650336
rect 289582 650100 325026 650336
rect 325262 650100 325346 650336
rect 325582 650100 361026 650336
rect 361262 650100 361346 650336
rect 361582 650100 397026 650336
rect 397262 650100 397346 650336
rect 397582 650100 433026 650336
rect 433262 650100 433346 650336
rect 433582 650100 469026 650336
rect 469262 650100 469346 650336
rect 469582 650100 505026 650336
rect 505262 650100 505346 650336
rect 505582 650100 541026 650336
rect 541262 650100 541346 650336
rect 541582 650100 577026 650336
rect 577262 650100 577346 650336
rect 577582 650100 585342 650336
rect 585578 650100 585662 650336
rect 585898 650100 592650 650336
rect -8726 650068 592650 650100
rect -8726 623336 592650 623368
rect -8726 623100 -8694 623336
rect -8458 623100 -8374 623336
rect -8138 623100 9706 623336
rect 9942 623100 10026 623336
rect 10262 623100 45706 623336
rect 45942 623100 46026 623336
rect 46262 623100 81706 623336
rect 81942 623100 82026 623336
rect 82262 623100 117706 623336
rect 117942 623100 118026 623336
rect 118262 623100 153706 623336
rect 153942 623100 154026 623336
rect 154262 623100 189706 623336
rect 189942 623100 190026 623336
rect 190262 623100 225706 623336
rect 225942 623100 226026 623336
rect 226262 623100 261706 623336
rect 261942 623100 262026 623336
rect 262262 623100 297706 623336
rect 297942 623100 298026 623336
rect 298262 623100 333706 623336
rect 333942 623100 334026 623336
rect 334262 623100 369706 623336
rect 369942 623100 370026 623336
rect 370262 623100 405706 623336
rect 405942 623100 406026 623336
rect 406262 623100 441706 623336
rect 441942 623100 442026 623336
rect 442262 623100 477706 623336
rect 477942 623100 478026 623336
rect 478262 623100 513706 623336
rect 513942 623100 514026 623336
rect 514262 623100 549706 623336
rect 549942 623100 550026 623336
rect 550262 623100 592062 623336
rect 592298 623100 592382 623336
rect 592618 623100 592650 623336
rect -8726 623016 592650 623100
rect -8726 622780 -8694 623016
rect -8458 622780 -8374 623016
rect -8138 622780 9706 623016
rect 9942 622780 10026 623016
rect 10262 622780 45706 623016
rect 45942 622780 46026 623016
rect 46262 622780 81706 623016
rect 81942 622780 82026 623016
rect 82262 622780 117706 623016
rect 117942 622780 118026 623016
rect 118262 622780 153706 623016
rect 153942 622780 154026 623016
rect 154262 622780 189706 623016
rect 189942 622780 190026 623016
rect 190262 622780 225706 623016
rect 225942 622780 226026 623016
rect 226262 622780 261706 623016
rect 261942 622780 262026 623016
rect 262262 622780 297706 623016
rect 297942 622780 298026 623016
rect 298262 622780 333706 623016
rect 333942 622780 334026 623016
rect 334262 622780 369706 623016
rect 369942 622780 370026 623016
rect 370262 622780 405706 623016
rect 405942 622780 406026 623016
rect 406262 622780 441706 623016
rect 441942 622780 442026 623016
rect 442262 622780 477706 623016
rect 477942 622780 478026 623016
rect 478262 622780 513706 623016
rect 513942 622780 514026 623016
rect 514262 622780 549706 623016
rect 549942 622780 550026 623016
rect 550262 622780 592062 623016
rect 592298 622780 592382 623016
rect 592618 622780 592650 623016
rect -8726 622748 592650 622780
rect -8726 622096 592650 622128
rect -8726 621860 -7734 622096
rect -7498 621860 -7414 622096
rect -7178 621860 8466 622096
rect 8702 621860 8786 622096
rect 9022 621860 44466 622096
rect 44702 621860 44786 622096
rect 45022 621860 80466 622096
rect 80702 621860 80786 622096
rect 81022 621860 116466 622096
rect 116702 621860 116786 622096
rect 117022 621860 152466 622096
rect 152702 621860 152786 622096
rect 153022 621860 188466 622096
rect 188702 621860 188786 622096
rect 189022 621860 224466 622096
rect 224702 621860 224786 622096
rect 225022 621860 260466 622096
rect 260702 621860 260786 622096
rect 261022 621860 296466 622096
rect 296702 621860 296786 622096
rect 297022 621860 332466 622096
rect 332702 621860 332786 622096
rect 333022 621860 368466 622096
rect 368702 621860 368786 622096
rect 369022 621860 404466 622096
rect 404702 621860 404786 622096
rect 405022 621860 440466 622096
rect 440702 621860 440786 622096
rect 441022 621860 476466 622096
rect 476702 621860 476786 622096
rect 477022 621860 512466 622096
rect 512702 621860 512786 622096
rect 513022 621860 548466 622096
rect 548702 621860 548786 622096
rect 549022 621860 591102 622096
rect 591338 621860 591422 622096
rect 591658 621860 592650 622096
rect -8726 621776 592650 621860
rect -8726 621540 -7734 621776
rect -7498 621540 -7414 621776
rect -7178 621540 8466 621776
rect 8702 621540 8786 621776
rect 9022 621540 44466 621776
rect 44702 621540 44786 621776
rect 45022 621540 80466 621776
rect 80702 621540 80786 621776
rect 81022 621540 116466 621776
rect 116702 621540 116786 621776
rect 117022 621540 152466 621776
rect 152702 621540 152786 621776
rect 153022 621540 188466 621776
rect 188702 621540 188786 621776
rect 189022 621540 224466 621776
rect 224702 621540 224786 621776
rect 225022 621540 260466 621776
rect 260702 621540 260786 621776
rect 261022 621540 296466 621776
rect 296702 621540 296786 621776
rect 297022 621540 332466 621776
rect 332702 621540 332786 621776
rect 333022 621540 368466 621776
rect 368702 621540 368786 621776
rect 369022 621540 404466 621776
rect 404702 621540 404786 621776
rect 405022 621540 440466 621776
rect 440702 621540 440786 621776
rect 441022 621540 476466 621776
rect 476702 621540 476786 621776
rect 477022 621540 512466 621776
rect 512702 621540 512786 621776
rect 513022 621540 548466 621776
rect 548702 621540 548786 621776
rect 549022 621540 591102 621776
rect 591338 621540 591422 621776
rect 591658 621540 592650 621776
rect -8726 621508 592650 621540
rect -8726 620856 592650 620888
rect -8726 620620 -6774 620856
rect -6538 620620 -6454 620856
rect -6218 620620 7226 620856
rect 7462 620620 7546 620856
rect 7782 620620 43226 620856
rect 43462 620620 43546 620856
rect 43782 620620 79226 620856
rect 79462 620620 79546 620856
rect 79782 620620 115226 620856
rect 115462 620620 115546 620856
rect 115782 620620 151226 620856
rect 151462 620620 151546 620856
rect 151782 620620 187226 620856
rect 187462 620620 187546 620856
rect 187782 620620 223226 620856
rect 223462 620620 223546 620856
rect 223782 620620 259226 620856
rect 259462 620620 259546 620856
rect 259782 620620 295226 620856
rect 295462 620620 295546 620856
rect 295782 620620 331226 620856
rect 331462 620620 331546 620856
rect 331782 620620 367226 620856
rect 367462 620620 367546 620856
rect 367782 620620 403226 620856
rect 403462 620620 403546 620856
rect 403782 620620 439226 620856
rect 439462 620620 439546 620856
rect 439782 620620 475226 620856
rect 475462 620620 475546 620856
rect 475782 620620 511226 620856
rect 511462 620620 511546 620856
rect 511782 620620 547226 620856
rect 547462 620620 547546 620856
rect 547782 620620 590142 620856
rect 590378 620620 590462 620856
rect 590698 620620 592650 620856
rect -8726 620536 592650 620620
rect -8726 620300 -6774 620536
rect -6538 620300 -6454 620536
rect -6218 620300 7226 620536
rect 7462 620300 7546 620536
rect 7782 620300 43226 620536
rect 43462 620300 43546 620536
rect 43782 620300 79226 620536
rect 79462 620300 79546 620536
rect 79782 620300 115226 620536
rect 115462 620300 115546 620536
rect 115782 620300 151226 620536
rect 151462 620300 151546 620536
rect 151782 620300 187226 620536
rect 187462 620300 187546 620536
rect 187782 620300 223226 620536
rect 223462 620300 223546 620536
rect 223782 620300 259226 620536
rect 259462 620300 259546 620536
rect 259782 620300 295226 620536
rect 295462 620300 295546 620536
rect 295782 620300 331226 620536
rect 331462 620300 331546 620536
rect 331782 620300 367226 620536
rect 367462 620300 367546 620536
rect 367782 620300 403226 620536
rect 403462 620300 403546 620536
rect 403782 620300 439226 620536
rect 439462 620300 439546 620536
rect 439782 620300 475226 620536
rect 475462 620300 475546 620536
rect 475782 620300 511226 620536
rect 511462 620300 511546 620536
rect 511782 620300 547226 620536
rect 547462 620300 547546 620536
rect 547782 620300 590142 620536
rect 590378 620300 590462 620536
rect 590698 620300 592650 620536
rect -8726 620268 592650 620300
rect -8726 619616 592650 619648
rect -8726 619380 -5814 619616
rect -5578 619380 -5494 619616
rect -5258 619380 5986 619616
rect 6222 619380 6306 619616
rect 6542 619380 41986 619616
rect 42222 619380 42306 619616
rect 42542 619380 77986 619616
rect 78222 619380 78306 619616
rect 78542 619380 113986 619616
rect 114222 619380 114306 619616
rect 114542 619380 149986 619616
rect 150222 619380 150306 619616
rect 150542 619380 185986 619616
rect 186222 619380 186306 619616
rect 186542 619380 221986 619616
rect 222222 619380 222306 619616
rect 222542 619380 257986 619616
rect 258222 619380 258306 619616
rect 258542 619380 293986 619616
rect 294222 619380 294306 619616
rect 294542 619380 329986 619616
rect 330222 619380 330306 619616
rect 330542 619380 365986 619616
rect 366222 619380 366306 619616
rect 366542 619380 401986 619616
rect 402222 619380 402306 619616
rect 402542 619380 437986 619616
rect 438222 619380 438306 619616
rect 438542 619380 473986 619616
rect 474222 619380 474306 619616
rect 474542 619380 509986 619616
rect 510222 619380 510306 619616
rect 510542 619380 545986 619616
rect 546222 619380 546306 619616
rect 546542 619380 581986 619616
rect 582222 619380 582306 619616
rect 582542 619380 589182 619616
rect 589418 619380 589502 619616
rect 589738 619380 592650 619616
rect -8726 619296 592650 619380
rect -8726 619060 -5814 619296
rect -5578 619060 -5494 619296
rect -5258 619060 5986 619296
rect 6222 619060 6306 619296
rect 6542 619060 41986 619296
rect 42222 619060 42306 619296
rect 42542 619060 77986 619296
rect 78222 619060 78306 619296
rect 78542 619060 113986 619296
rect 114222 619060 114306 619296
rect 114542 619060 149986 619296
rect 150222 619060 150306 619296
rect 150542 619060 185986 619296
rect 186222 619060 186306 619296
rect 186542 619060 221986 619296
rect 222222 619060 222306 619296
rect 222542 619060 257986 619296
rect 258222 619060 258306 619296
rect 258542 619060 293986 619296
rect 294222 619060 294306 619296
rect 294542 619060 329986 619296
rect 330222 619060 330306 619296
rect 330542 619060 365986 619296
rect 366222 619060 366306 619296
rect 366542 619060 401986 619296
rect 402222 619060 402306 619296
rect 402542 619060 437986 619296
rect 438222 619060 438306 619296
rect 438542 619060 473986 619296
rect 474222 619060 474306 619296
rect 474542 619060 509986 619296
rect 510222 619060 510306 619296
rect 510542 619060 545986 619296
rect 546222 619060 546306 619296
rect 546542 619060 581986 619296
rect 582222 619060 582306 619296
rect 582542 619060 589182 619296
rect 589418 619060 589502 619296
rect 589738 619060 592650 619296
rect -8726 619028 592650 619060
rect -8726 618376 592650 618408
rect -8726 618140 -4854 618376
rect -4618 618140 -4534 618376
rect -4298 618140 4746 618376
rect 4982 618140 5066 618376
rect 5302 618140 40746 618376
rect 40982 618140 41066 618376
rect 41302 618140 76746 618376
rect 76982 618140 77066 618376
rect 77302 618140 112746 618376
rect 112982 618140 113066 618376
rect 113302 618140 148746 618376
rect 148982 618140 149066 618376
rect 149302 618140 184746 618376
rect 184982 618140 185066 618376
rect 185302 618140 220746 618376
rect 220982 618140 221066 618376
rect 221302 618140 256746 618376
rect 256982 618140 257066 618376
rect 257302 618140 292746 618376
rect 292982 618140 293066 618376
rect 293302 618140 328746 618376
rect 328982 618140 329066 618376
rect 329302 618140 364746 618376
rect 364982 618140 365066 618376
rect 365302 618140 400746 618376
rect 400982 618140 401066 618376
rect 401302 618140 436746 618376
rect 436982 618140 437066 618376
rect 437302 618140 472746 618376
rect 472982 618140 473066 618376
rect 473302 618140 508746 618376
rect 508982 618140 509066 618376
rect 509302 618140 544746 618376
rect 544982 618140 545066 618376
rect 545302 618140 580746 618376
rect 580982 618140 581066 618376
rect 581302 618140 588222 618376
rect 588458 618140 588542 618376
rect 588778 618140 592650 618376
rect -8726 618056 592650 618140
rect -8726 617820 -4854 618056
rect -4618 617820 -4534 618056
rect -4298 617820 4746 618056
rect 4982 617820 5066 618056
rect 5302 617820 40746 618056
rect 40982 617820 41066 618056
rect 41302 617820 76746 618056
rect 76982 617820 77066 618056
rect 77302 617820 112746 618056
rect 112982 617820 113066 618056
rect 113302 617820 148746 618056
rect 148982 617820 149066 618056
rect 149302 617820 184746 618056
rect 184982 617820 185066 618056
rect 185302 617820 220746 618056
rect 220982 617820 221066 618056
rect 221302 617820 256746 618056
rect 256982 617820 257066 618056
rect 257302 617820 292746 618056
rect 292982 617820 293066 618056
rect 293302 617820 328746 618056
rect 328982 617820 329066 618056
rect 329302 617820 364746 618056
rect 364982 617820 365066 618056
rect 365302 617820 400746 618056
rect 400982 617820 401066 618056
rect 401302 617820 436746 618056
rect 436982 617820 437066 618056
rect 437302 617820 472746 618056
rect 472982 617820 473066 618056
rect 473302 617820 508746 618056
rect 508982 617820 509066 618056
rect 509302 617820 544746 618056
rect 544982 617820 545066 618056
rect 545302 617820 580746 618056
rect 580982 617820 581066 618056
rect 581302 617820 588222 618056
rect 588458 617820 588542 618056
rect 588778 617820 592650 618056
rect -8726 617788 592650 617820
rect -8726 617136 592650 617168
rect -8726 616900 -3894 617136
rect -3658 616900 -3574 617136
rect -3338 616900 3506 617136
rect 3742 616900 3826 617136
rect 4062 616900 39506 617136
rect 39742 616900 39826 617136
rect 40062 616900 75506 617136
rect 75742 616900 75826 617136
rect 76062 616900 111506 617136
rect 111742 616900 111826 617136
rect 112062 616900 147506 617136
rect 147742 616900 147826 617136
rect 148062 616900 183506 617136
rect 183742 616900 183826 617136
rect 184062 616900 219506 617136
rect 219742 616900 219826 617136
rect 220062 616900 255506 617136
rect 255742 616900 255826 617136
rect 256062 616900 291506 617136
rect 291742 616900 291826 617136
rect 292062 616900 327506 617136
rect 327742 616900 327826 617136
rect 328062 616900 363506 617136
rect 363742 616900 363826 617136
rect 364062 616900 399506 617136
rect 399742 616900 399826 617136
rect 400062 616900 435506 617136
rect 435742 616900 435826 617136
rect 436062 616900 471506 617136
rect 471742 616900 471826 617136
rect 472062 616900 507506 617136
rect 507742 616900 507826 617136
rect 508062 616900 543506 617136
rect 543742 616900 543826 617136
rect 544062 616900 579506 617136
rect 579742 616900 579826 617136
rect 580062 616900 587262 617136
rect 587498 616900 587582 617136
rect 587818 616900 592650 617136
rect -8726 616816 592650 616900
rect -8726 616580 -3894 616816
rect -3658 616580 -3574 616816
rect -3338 616580 3506 616816
rect 3742 616580 3826 616816
rect 4062 616580 39506 616816
rect 39742 616580 39826 616816
rect 40062 616580 75506 616816
rect 75742 616580 75826 616816
rect 76062 616580 111506 616816
rect 111742 616580 111826 616816
rect 112062 616580 147506 616816
rect 147742 616580 147826 616816
rect 148062 616580 183506 616816
rect 183742 616580 183826 616816
rect 184062 616580 219506 616816
rect 219742 616580 219826 616816
rect 220062 616580 255506 616816
rect 255742 616580 255826 616816
rect 256062 616580 291506 616816
rect 291742 616580 291826 616816
rect 292062 616580 327506 616816
rect 327742 616580 327826 616816
rect 328062 616580 363506 616816
rect 363742 616580 363826 616816
rect 364062 616580 399506 616816
rect 399742 616580 399826 616816
rect 400062 616580 435506 616816
rect 435742 616580 435826 616816
rect 436062 616580 471506 616816
rect 471742 616580 471826 616816
rect 472062 616580 507506 616816
rect 507742 616580 507826 616816
rect 508062 616580 543506 616816
rect 543742 616580 543826 616816
rect 544062 616580 579506 616816
rect 579742 616580 579826 616816
rect 580062 616580 587262 616816
rect 587498 616580 587582 616816
rect 587818 616580 592650 616816
rect -8726 616548 592650 616580
rect -8726 615896 592650 615928
rect -8726 615660 -2934 615896
rect -2698 615660 -2614 615896
rect -2378 615660 2266 615896
rect 2502 615660 2586 615896
rect 2822 615660 38266 615896
rect 38502 615660 38586 615896
rect 38822 615660 74266 615896
rect 74502 615660 74586 615896
rect 74822 615660 110266 615896
rect 110502 615660 110586 615896
rect 110822 615660 146266 615896
rect 146502 615660 146586 615896
rect 146822 615660 182266 615896
rect 182502 615660 182586 615896
rect 182822 615660 218266 615896
rect 218502 615660 218586 615896
rect 218822 615660 254266 615896
rect 254502 615660 254586 615896
rect 254822 615660 290266 615896
rect 290502 615660 290586 615896
rect 290822 615660 326266 615896
rect 326502 615660 326586 615896
rect 326822 615660 362266 615896
rect 362502 615660 362586 615896
rect 362822 615660 398266 615896
rect 398502 615660 398586 615896
rect 398822 615660 434266 615896
rect 434502 615660 434586 615896
rect 434822 615660 470266 615896
rect 470502 615660 470586 615896
rect 470822 615660 506266 615896
rect 506502 615660 506586 615896
rect 506822 615660 542266 615896
rect 542502 615660 542586 615896
rect 542822 615660 578266 615896
rect 578502 615660 578586 615896
rect 578822 615660 586302 615896
rect 586538 615660 586622 615896
rect 586858 615660 592650 615896
rect -8726 615576 592650 615660
rect -8726 615340 -2934 615576
rect -2698 615340 -2614 615576
rect -2378 615340 2266 615576
rect 2502 615340 2586 615576
rect 2822 615340 38266 615576
rect 38502 615340 38586 615576
rect 38822 615340 74266 615576
rect 74502 615340 74586 615576
rect 74822 615340 110266 615576
rect 110502 615340 110586 615576
rect 110822 615340 146266 615576
rect 146502 615340 146586 615576
rect 146822 615340 182266 615576
rect 182502 615340 182586 615576
rect 182822 615340 218266 615576
rect 218502 615340 218586 615576
rect 218822 615340 254266 615576
rect 254502 615340 254586 615576
rect 254822 615340 290266 615576
rect 290502 615340 290586 615576
rect 290822 615340 326266 615576
rect 326502 615340 326586 615576
rect 326822 615340 362266 615576
rect 362502 615340 362586 615576
rect 362822 615340 398266 615576
rect 398502 615340 398586 615576
rect 398822 615340 434266 615576
rect 434502 615340 434586 615576
rect 434822 615340 470266 615576
rect 470502 615340 470586 615576
rect 470822 615340 506266 615576
rect 506502 615340 506586 615576
rect 506822 615340 542266 615576
rect 542502 615340 542586 615576
rect 542822 615340 578266 615576
rect 578502 615340 578586 615576
rect 578822 615340 586302 615576
rect 586538 615340 586622 615576
rect 586858 615340 592650 615576
rect -8726 615308 592650 615340
rect -8726 614656 592650 614688
rect -8726 614420 -1974 614656
rect -1738 614420 -1654 614656
rect -1418 614420 1026 614656
rect 1262 614420 1346 614656
rect 1582 614420 37026 614656
rect 37262 614420 37346 614656
rect 37582 614420 73026 614656
rect 73262 614420 73346 614656
rect 73582 614420 109026 614656
rect 109262 614420 109346 614656
rect 109582 614420 145026 614656
rect 145262 614420 145346 614656
rect 145582 614420 181026 614656
rect 181262 614420 181346 614656
rect 181582 614420 217026 614656
rect 217262 614420 217346 614656
rect 217582 614420 253026 614656
rect 253262 614420 253346 614656
rect 253582 614420 289026 614656
rect 289262 614420 289346 614656
rect 289582 614420 325026 614656
rect 325262 614420 325346 614656
rect 325582 614420 361026 614656
rect 361262 614420 361346 614656
rect 361582 614420 397026 614656
rect 397262 614420 397346 614656
rect 397582 614420 433026 614656
rect 433262 614420 433346 614656
rect 433582 614420 469026 614656
rect 469262 614420 469346 614656
rect 469582 614420 505026 614656
rect 505262 614420 505346 614656
rect 505582 614420 541026 614656
rect 541262 614420 541346 614656
rect 541582 614420 577026 614656
rect 577262 614420 577346 614656
rect 577582 614420 585342 614656
rect 585578 614420 585662 614656
rect 585898 614420 592650 614656
rect -8726 614336 592650 614420
rect -8726 614100 -1974 614336
rect -1738 614100 -1654 614336
rect -1418 614100 1026 614336
rect 1262 614100 1346 614336
rect 1582 614100 37026 614336
rect 37262 614100 37346 614336
rect 37582 614100 73026 614336
rect 73262 614100 73346 614336
rect 73582 614100 109026 614336
rect 109262 614100 109346 614336
rect 109582 614100 145026 614336
rect 145262 614100 145346 614336
rect 145582 614100 181026 614336
rect 181262 614100 181346 614336
rect 181582 614100 217026 614336
rect 217262 614100 217346 614336
rect 217582 614100 253026 614336
rect 253262 614100 253346 614336
rect 253582 614100 289026 614336
rect 289262 614100 289346 614336
rect 289582 614100 325026 614336
rect 325262 614100 325346 614336
rect 325582 614100 361026 614336
rect 361262 614100 361346 614336
rect 361582 614100 397026 614336
rect 397262 614100 397346 614336
rect 397582 614100 433026 614336
rect 433262 614100 433346 614336
rect 433582 614100 469026 614336
rect 469262 614100 469346 614336
rect 469582 614100 505026 614336
rect 505262 614100 505346 614336
rect 505582 614100 541026 614336
rect 541262 614100 541346 614336
rect 541582 614100 577026 614336
rect 577262 614100 577346 614336
rect 577582 614100 585342 614336
rect 585578 614100 585662 614336
rect 585898 614100 592650 614336
rect -8726 614068 592650 614100
rect -8726 587336 592650 587368
rect -8726 587100 -8694 587336
rect -8458 587100 -8374 587336
rect -8138 587100 9706 587336
rect 9942 587100 10026 587336
rect 10262 587100 45706 587336
rect 45942 587100 46026 587336
rect 46262 587100 81706 587336
rect 81942 587100 82026 587336
rect 82262 587100 117706 587336
rect 117942 587100 118026 587336
rect 118262 587100 153706 587336
rect 153942 587100 154026 587336
rect 154262 587100 189706 587336
rect 189942 587100 190026 587336
rect 190262 587100 225706 587336
rect 225942 587100 226026 587336
rect 226262 587100 261706 587336
rect 261942 587100 262026 587336
rect 262262 587100 297706 587336
rect 297942 587100 298026 587336
rect 298262 587100 333706 587336
rect 333942 587100 334026 587336
rect 334262 587100 369706 587336
rect 369942 587100 370026 587336
rect 370262 587100 405706 587336
rect 405942 587100 406026 587336
rect 406262 587100 441706 587336
rect 441942 587100 442026 587336
rect 442262 587100 477706 587336
rect 477942 587100 478026 587336
rect 478262 587100 513706 587336
rect 513942 587100 514026 587336
rect 514262 587100 549706 587336
rect 549942 587100 550026 587336
rect 550262 587100 592062 587336
rect 592298 587100 592382 587336
rect 592618 587100 592650 587336
rect -8726 587016 592650 587100
rect -8726 586780 -8694 587016
rect -8458 586780 -8374 587016
rect -8138 586780 9706 587016
rect 9942 586780 10026 587016
rect 10262 586780 45706 587016
rect 45942 586780 46026 587016
rect 46262 586780 81706 587016
rect 81942 586780 82026 587016
rect 82262 586780 117706 587016
rect 117942 586780 118026 587016
rect 118262 586780 153706 587016
rect 153942 586780 154026 587016
rect 154262 586780 189706 587016
rect 189942 586780 190026 587016
rect 190262 586780 225706 587016
rect 225942 586780 226026 587016
rect 226262 586780 261706 587016
rect 261942 586780 262026 587016
rect 262262 586780 297706 587016
rect 297942 586780 298026 587016
rect 298262 586780 333706 587016
rect 333942 586780 334026 587016
rect 334262 586780 369706 587016
rect 369942 586780 370026 587016
rect 370262 586780 405706 587016
rect 405942 586780 406026 587016
rect 406262 586780 441706 587016
rect 441942 586780 442026 587016
rect 442262 586780 477706 587016
rect 477942 586780 478026 587016
rect 478262 586780 513706 587016
rect 513942 586780 514026 587016
rect 514262 586780 549706 587016
rect 549942 586780 550026 587016
rect 550262 586780 592062 587016
rect 592298 586780 592382 587016
rect 592618 586780 592650 587016
rect -8726 586748 592650 586780
rect -8726 586096 592650 586128
rect -8726 585860 -7734 586096
rect -7498 585860 -7414 586096
rect -7178 585860 8466 586096
rect 8702 585860 8786 586096
rect 9022 585860 44466 586096
rect 44702 585860 44786 586096
rect 45022 585860 80466 586096
rect 80702 585860 80786 586096
rect 81022 585860 116466 586096
rect 116702 585860 116786 586096
rect 117022 585860 152466 586096
rect 152702 585860 152786 586096
rect 153022 585860 188466 586096
rect 188702 585860 188786 586096
rect 189022 585860 224466 586096
rect 224702 585860 224786 586096
rect 225022 585860 260466 586096
rect 260702 585860 260786 586096
rect 261022 585860 296466 586096
rect 296702 585860 296786 586096
rect 297022 585860 332466 586096
rect 332702 585860 332786 586096
rect 333022 585860 368466 586096
rect 368702 585860 368786 586096
rect 369022 585860 404466 586096
rect 404702 585860 404786 586096
rect 405022 585860 440466 586096
rect 440702 585860 440786 586096
rect 441022 585860 476466 586096
rect 476702 585860 476786 586096
rect 477022 585860 512466 586096
rect 512702 585860 512786 586096
rect 513022 585860 548466 586096
rect 548702 585860 548786 586096
rect 549022 585860 591102 586096
rect 591338 585860 591422 586096
rect 591658 585860 592650 586096
rect -8726 585776 592650 585860
rect -8726 585540 -7734 585776
rect -7498 585540 -7414 585776
rect -7178 585540 8466 585776
rect 8702 585540 8786 585776
rect 9022 585540 44466 585776
rect 44702 585540 44786 585776
rect 45022 585540 80466 585776
rect 80702 585540 80786 585776
rect 81022 585540 116466 585776
rect 116702 585540 116786 585776
rect 117022 585540 152466 585776
rect 152702 585540 152786 585776
rect 153022 585540 188466 585776
rect 188702 585540 188786 585776
rect 189022 585540 224466 585776
rect 224702 585540 224786 585776
rect 225022 585540 260466 585776
rect 260702 585540 260786 585776
rect 261022 585540 296466 585776
rect 296702 585540 296786 585776
rect 297022 585540 332466 585776
rect 332702 585540 332786 585776
rect 333022 585540 368466 585776
rect 368702 585540 368786 585776
rect 369022 585540 404466 585776
rect 404702 585540 404786 585776
rect 405022 585540 440466 585776
rect 440702 585540 440786 585776
rect 441022 585540 476466 585776
rect 476702 585540 476786 585776
rect 477022 585540 512466 585776
rect 512702 585540 512786 585776
rect 513022 585540 548466 585776
rect 548702 585540 548786 585776
rect 549022 585540 591102 585776
rect 591338 585540 591422 585776
rect 591658 585540 592650 585776
rect -8726 585508 592650 585540
rect -8726 584856 592650 584888
rect -8726 584620 -6774 584856
rect -6538 584620 -6454 584856
rect -6218 584620 7226 584856
rect 7462 584620 7546 584856
rect 7782 584620 43226 584856
rect 43462 584620 43546 584856
rect 43782 584620 79226 584856
rect 79462 584620 79546 584856
rect 79782 584620 115226 584856
rect 115462 584620 115546 584856
rect 115782 584620 151226 584856
rect 151462 584620 151546 584856
rect 151782 584620 187226 584856
rect 187462 584620 187546 584856
rect 187782 584620 223226 584856
rect 223462 584620 223546 584856
rect 223782 584620 259226 584856
rect 259462 584620 259546 584856
rect 259782 584620 295226 584856
rect 295462 584620 295546 584856
rect 295782 584620 331226 584856
rect 331462 584620 331546 584856
rect 331782 584620 367226 584856
rect 367462 584620 367546 584856
rect 367782 584620 403226 584856
rect 403462 584620 403546 584856
rect 403782 584620 439226 584856
rect 439462 584620 439546 584856
rect 439782 584620 475226 584856
rect 475462 584620 475546 584856
rect 475782 584620 511226 584856
rect 511462 584620 511546 584856
rect 511782 584620 547226 584856
rect 547462 584620 547546 584856
rect 547782 584620 590142 584856
rect 590378 584620 590462 584856
rect 590698 584620 592650 584856
rect -8726 584536 592650 584620
rect -8726 584300 -6774 584536
rect -6538 584300 -6454 584536
rect -6218 584300 7226 584536
rect 7462 584300 7546 584536
rect 7782 584300 43226 584536
rect 43462 584300 43546 584536
rect 43782 584300 79226 584536
rect 79462 584300 79546 584536
rect 79782 584300 115226 584536
rect 115462 584300 115546 584536
rect 115782 584300 151226 584536
rect 151462 584300 151546 584536
rect 151782 584300 187226 584536
rect 187462 584300 187546 584536
rect 187782 584300 223226 584536
rect 223462 584300 223546 584536
rect 223782 584300 259226 584536
rect 259462 584300 259546 584536
rect 259782 584300 295226 584536
rect 295462 584300 295546 584536
rect 295782 584300 331226 584536
rect 331462 584300 331546 584536
rect 331782 584300 367226 584536
rect 367462 584300 367546 584536
rect 367782 584300 403226 584536
rect 403462 584300 403546 584536
rect 403782 584300 439226 584536
rect 439462 584300 439546 584536
rect 439782 584300 475226 584536
rect 475462 584300 475546 584536
rect 475782 584300 511226 584536
rect 511462 584300 511546 584536
rect 511782 584300 547226 584536
rect 547462 584300 547546 584536
rect 547782 584300 590142 584536
rect 590378 584300 590462 584536
rect 590698 584300 592650 584536
rect -8726 584268 592650 584300
rect -8726 583616 592650 583648
rect -8726 583380 -5814 583616
rect -5578 583380 -5494 583616
rect -5258 583380 5986 583616
rect 6222 583380 6306 583616
rect 6542 583380 41986 583616
rect 42222 583380 42306 583616
rect 42542 583380 77986 583616
rect 78222 583380 78306 583616
rect 78542 583380 113986 583616
rect 114222 583380 114306 583616
rect 114542 583380 149986 583616
rect 150222 583380 150306 583616
rect 150542 583380 185986 583616
rect 186222 583380 186306 583616
rect 186542 583380 221986 583616
rect 222222 583380 222306 583616
rect 222542 583380 257986 583616
rect 258222 583380 258306 583616
rect 258542 583380 293986 583616
rect 294222 583380 294306 583616
rect 294542 583380 329986 583616
rect 330222 583380 330306 583616
rect 330542 583380 365986 583616
rect 366222 583380 366306 583616
rect 366542 583380 401986 583616
rect 402222 583380 402306 583616
rect 402542 583380 437986 583616
rect 438222 583380 438306 583616
rect 438542 583380 473986 583616
rect 474222 583380 474306 583616
rect 474542 583380 509986 583616
rect 510222 583380 510306 583616
rect 510542 583380 545986 583616
rect 546222 583380 546306 583616
rect 546542 583380 581986 583616
rect 582222 583380 582306 583616
rect 582542 583380 589182 583616
rect 589418 583380 589502 583616
rect 589738 583380 592650 583616
rect -8726 583296 592650 583380
rect -8726 583060 -5814 583296
rect -5578 583060 -5494 583296
rect -5258 583060 5986 583296
rect 6222 583060 6306 583296
rect 6542 583060 41986 583296
rect 42222 583060 42306 583296
rect 42542 583060 77986 583296
rect 78222 583060 78306 583296
rect 78542 583060 113986 583296
rect 114222 583060 114306 583296
rect 114542 583060 149986 583296
rect 150222 583060 150306 583296
rect 150542 583060 185986 583296
rect 186222 583060 186306 583296
rect 186542 583060 221986 583296
rect 222222 583060 222306 583296
rect 222542 583060 257986 583296
rect 258222 583060 258306 583296
rect 258542 583060 293986 583296
rect 294222 583060 294306 583296
rect 294542 583060 329986 583296
rect 330222 583060 330306 583296
rect 330542 583060 365986 583296
rect 366222 583060 366306 583296
rect 366542 583060 401986 583296
rect 402222 583060 402306 583296
rect 402542 583060 437986 583296
rect 438222 583060 438306 583296
rect 438542 583060 473986 583296
rect 474222 583060 474306 583296
rect 474542 583060 509986 583296
rect 510222 583060 510306 583296
rect 510542 583060 545986 583296
rect 546222 583060 546306 583296
rect 546542 583060 581986 583296
rect 582222 583060 582306 583296
rect 582542 583060 589182 583296
rect 589418 583060 589502 583296
rect 589738 583060 592650 583296
rect -8726 583028 592650 583060
rect -8726 582376 592650 582408
rect -8726 582140 -4854 582376
rect -4618 582140 -4534 582376
rect -4298 582140 4746 582376
rect 4982 582140 5066 582376
rect 5302 582140 40746 582376
rect 40982 582140 41066 582376
rect 41302 582140 76746 582376
rect 76982 582140 77066 582376
rect 77302 582140 112746 582376
rect 112982 582140 113066 582376
rect 113302 582140 148746 582376
rect 148982 582140 149066 582376
rect 149302 582140 184746 582376
rect 184982 582140 185066 582376
rect 185302 582140 220746 582376
rect 220982 582140 221066 582376
rect 221302 582140 256746 582376
rect 256982 582140 257066 582376
rect 257302 582140 292746 582376
rect 292982 582140 293066 582376
rect 293302 582140 328746 582376
rect 328982 582140 329066 582376
rect 329302 582140 364746 582376
rect 364982 582140 365066 582376
rect 365302 582140 400746 582376
rect 400982 582140 401066 582376
rect 401302 582140 436746 582376
rect 436982 582140 437066 582376
rect 437302 582140 472746 582376
rect 472982 582140 473066 582376
rect 473302 582140 508746 582376
rect 508982 582140 509066 582376
rect 509302 582140 544746 582376
rect 544982 582140 545066 582376
rect 545302 582140 580746 582376
rect 580982 582140 581066 582376
rect 581302 582140 588222 582376
rect 588458 582140 588542 582376
rect 588778 582140 592650 582376
rect -8726 582056 592650 582140
rect -8726 581820 -4854 582056
rect -4618 581820 -4534 582056
rect -4298 581820 4746 582056
rect 4982 581820 5066 582056
rect 5302 581820 40746 582056
rect 40982 581820 41066 582056
rect 41302 581820 76746 582056
rect 76982 581820 77066 582056
rect 77302 581820 112746 582056
rect 112982 581820 113066 582056
rect 113302 581820 148746 582056
rect 148982 581820 149066 582056
rect 149302 581820 184746 582056
rect 184982 581820 185066 582056
rect 185302 581820 220746 582056
rect 220982 581820 221066 582056
rect 221302 581820 256746 582056
rect 256982 581820 257066 582056
rect 257302 581820 292746 582056
rect 292982 581820 293066 582056
rect 293302 581820 328746 582056
rect 328982 581820 329066 582056
rect 329302 581820 364746 582056
rect 364982 581820 365066 582056
rect 365302 581820 400746 582056
rect 400982 581820 401066 582056
rect 401302 581820 436746 582056
rect 436982 581820 437066 582056
rect 437302 581820 472746 582056
rect 472982 581820 473066 582056
rect 473302 581820 508746 582056
rect 508982 581820 509066 582056
rect 509302 581820 544746 582056
rect 544982 581820 545066 582056
rect 545302 581820 580746 582056
rect 580982 581820 581066 582056
rect 581302 581820 588222 582056
rect 588458 581820 588542 582056
rect 588778 581820 592650 582056
rect -8726 581788 592650 581820
rect -8726 581136 592650 581168
rect -8726 580900 -3894 581136
rect -3658 580900 -3574 581136
rect -3338 580900 3506 581136
rect 3742 580900 3826 581136
rect 4062 580900 39506 581136
rect 39742 580900 39826 581136
rect 40062 580900 75506 581136
rect 75742 580900 75826 581136
rect 76062 580900 111506 581136
rect 111742 580900 111826 581136
rect 112062 580900 147506 581136
rect 147742 580900 147826 581136
rect 148062 580900 183506 581136
rect 183742 580900 183826 581136
rect 184062 580900 219506 581136
rect 219742 580900 219826 581136
rect 220062 580900 255506 581136
rect 255742 580900 255826 581136
rect 256062 580900 291506 581136
rect 291742 580900 291826 581136
rect 292062 580900 327506 581136
rect 327742 580900 327826 581136
rect 328062 580900 363506 581136
rect 363742 580900 363826 581136
rect 364062 580900 399506 581136
rect 399742 580900 399826 581136
rect 400062 580900 435506 581136
rect 435742 580900 435826 581136
rect 436062 580900 471506 581136
rect 471742 580900 471826 581136
rect 472062 580900 507506 581136
rect 507742 580900 507826 581136
rect 508062 580900 543506 581136
rect 543742 580900 543826 581136
rect 544062 580900 579506 581136
rect 579742 580900 579826 581136
rect 580062 580900 587262 581136
rect 587498 580900 587582 581136
rect 587818 580900 592650 581136
rect -8726 580816 592650 580900
rect -8726 580580 -3894 580816
rect -3658 580580 -3574 580816
rect -3338 580580 3506 580816
rect 3742 580580 3826 580816
rect 4062 580580 39506 580816
rect 39742 580580 39826 580816
rect 40062 580580 75506 580816
rect 75742 580580 75826 580816
rect 76062 580580 111506 580816
rect 111742 580580 111826 580816
rect 112062 580580 147506 580816
rect 147742 580580 147826 580816
rect 148062 580580 183506 580816
rect 183742 580580 183826 580816
rect 184062 580580 219506 580816
rect 219742 580580 219826 580816
rect 220062 580580 255506 580816
rect 255742 580580 255826 580816
rect 256062 580580 291506 580816
rect 291742 580580 291826 580816
rect 292062 580580 327506 580816
rect 327742 580580 327826 580816
rect 328062 580580 363506 580816
rect 363742 580580 363826 580816
rect 364062 580580 399506 580816
rect 399742 580580 399826 580816
rect 400062 580580 435506 580816
rect 435742 580580 435826 580816
rect 436062 580580 471506 580816
rect 471742 580580 471826 580816
rect 472062 580580 507506 580816
rect 507742 580580 507826 580816
rect 508062 580580 543506 580816
rect 543742 580580 543826 580816
rect 544062 580580 579506 580816
rect 579742 580580 579826 580816
rect 580062 580580 587262 580816
rect 587498 580580 587582 580816
rect 587818 580580 592650 580816
rect -8726 580548 592650 580580
rect -8726 579896 592650 579928
rect -8726 579660 -2934 579896
rect -2698 579660 -2614 579896
rect -2378 579660 2266 579896
rect 2502 579660 2586 579896
rect 2822 579660 38266 579896
rect 38502 579660 38586 579896
rect 38822 579660 74266 579896
rect 74502 579660 74586 579896
rect 74822 579660 110266 579896
rect 110502 579660 110586 579896
rect 110822 579660 146266 579896
rect 146502 579660 146586 579896
rect 146822 579660 182266 579896
rect 182502 579660 182586 579896
rect 182822 579660 218266 579896
rect 218502 579660 218586 579896
rect 218822 579660 254266 579896
rect 254502 579660 254586 579896
rect 254822 579660 290266 579896
rect 290502 579660 290586 579896
rect 290822 579660 326266 579896
rect 326502 579660 326586 579896
rect 326822 579660 362266 579896
rect 362502 579660 362586 579896
rect 362822 579660 398266 579896
rect 398502 579660 398586 579896
rect 398822 579660 434266 579896
rect 434502 579660 434586 579896
rect 434822 579660 470266 579896
rect 470502 579660 470586 579896
rect 470822 579660 506266 579896
rect 506502 579660 506586 579896
rect 506822 579660 542266 579896
rect 542502 579660 542586 579896
rect 542822 579660 578266 579896
rect 578502 579660 578586 579896
rect 578822 579660 586302 579896
rect 586538 579660 586622 579896
rect 586858 579660 592650 579896
rect -8726 579576 592650 579660
rect -8726 579340 -2934 579576
rect -2698 579340 -2614 579576
rect -2378 579340 2266 579576
rect 2502 579340 2586 579576
rect 2822 579340 38266 579576
rect 38502 579340 38586 579576
rect 38822 579340 74266 579576
rect 74502 579340 74586 579576
rect 74822 579340 110266 579576
rect 110502 579340 110586 579576
rect 110822 579340 146266 579576
rect 146502 579340 146586 579576
rect 146822 579340 182266 579576
rect 182502 579340 182586 579576
rect 182822 579340 218266 579576
rect 218502 579340 218586 579576
rect 218822 579340 254266 579576
rect 254502 579340 254586 579576
rect 254822 579340 290266 579576
rect 290502 579340 290586 579576
rect 290822 579340 326266 579576
rect 326502 579340 326586 579576
rect 326822 579340 362266 579576
rect 362502 579340 362586 579576
rect 362822 579340 398266 579576
rect 398502 579340 398586 579576
rect 398822 579340 434266 579576
rect 434502 579340 434586 579576
rect 434822 579340 470266 579576
rect 470502 579340 470586 579576
rect 470822 579340 506266 579576
rect 506502 579340 506586 579576
rect 506822 579340 542266 579576
rect 542502 579340 542586 579576
rect 542822 579340 578266 579576
rect 578502 579340 578586 579576
rect 578822 579340 586302 579576
rect 586538 579340 586622 579576
rect 586858 579340 592650 579576
rect -8726 579308 592650 579340
rect -8726 578656 592650 578688
rect -8726 578420 -1974 578656
rect -1738 578420 -1654 578656
rect -1418 578420 1026 578656
rect 1262 578420 1346 578656
rect 1582 578420 37026 578656
rect 37262 578420 37346 578656
rect 37582 578420 73026 578656
rect 73262 578420 73346 578656
rect 73582 578420 109026 578656
rect 109262 578420 109346 578656
rect 109582 578420 145026 578656
rect 145262 578420 145346 578656
rect 145582 578420 181026 578656
rect 181262 578420 181346 578656
rect 181582 578420 217026 578656
rect 217262 578420 217346 578656
rect 217582 578420 253026 578656
rect 253262 578420 253346 578656
rect 253582 578420 289026 578656
rect 289262 578420 289346 578656
rect 289582 578420 325026 578656
rect 325262 578420 325346 578656
rect 325582 578420 361026 578656
rect 361262 578420 361346 578656
rect 361582 578420 397026 578656
rect 397262 578420 397346 578656
rect 397582 578420 433026 578656
rect 433262 578420 433346 578656
rect 433582 578420 469026 578656
rect 469262 578420 469346 578656
rect 469582 578420 505026 578656
rect 505262 578420 505346 578656
rect 505582 578420 541026 578656
rect 541262 578420 541346 578656
rect 541582 578420 577026 578656
rect 577262 578420 577346 578656
rect 577582 578420 585342 578656
rect 585578 578420 585662 578656
rect 585898 578420 592650 578656
rect -8726 578336 592650 578420
rect -8726 578100 -1974 578336
rect -1738 578100 -1654 578336
rect -1418 578100 1026 578336
rect 1262 578100 1346 578336
rect 1582 578100 37026 578336
rect 37262 578100 37346 578336
rect 37582 578100 73026 578336
rect 73262 578100 73346 578336
rect 73582 578100 109026 578336
rect 109262 578100 109346 578336
rect 109582 578100 145026 578336
rect 145262 578100 145346 578336
rect 145582 578100 181026 578336
rect 181262 578100 181346 578336
rect 181582 578100 217026 578336
rect 217262 578100 217346 578336
rect 217582 578100 253026 578336
rect 253262 578100 253346 578336
rect 253582 578100 289026 578336
rect 289262 578100 289346 578336
rect 289582 578100 325026 578336
rect 325262 578100 325346 578336
rect 325582 578100 361026 578336
rect 361262 578100 361346 578336
rect 361582 578100 397026 578336
rect 397262 578100 397346 578336
rect 397582 578100 433026 578336
rect 433262 578100 433346 578336
rect 433582 578100 469026 578336
rect 469262 578100 469346 578336
rect 469582 578100 505026 578336
rect 505262 578100 505346 578336
rect 505582 578100 541026 578336
rect 541262 578100 541346 578336
rect 541582 578100 577026 578336
rect 577262 578100 577346 578336
rect 577582 578100 585342 578336
rect 585578 578100 585662 578336
rect 585898 578100 592650 578336
rect -8726 578068 592650 578100
rect -8726 551336 592650 551368
rect -8726 551100 -8694 551336
rect -8458 551100 -8374 551336
rect -8138 551100 9706 551336
rect 9942 551100 10026 551336
rect 10262 551100 45706 551336
rect 45942 551100 46026 551336
rect 46262 551100 81706 551336
rect 81942 551100 82026 551336
rect 82262 551100 117706 551336
rect 117942 551100 118026 551336
rect 118262 551100 153706 551336
rect 153942 551100 154026 551336
rect 154262 551100 189706 551336
rect 189942 551100 190026 551336
rect 190262 551100 225706 551336
rect 225942 551100 226026 551336
rect 226262 551100 261706 551336
rect 261942 551100 262026 551336
rect 262262 551100 297706 551336
rect 297942 551100 298026 551336
rect 298262 551100 333706 551336
rect 333942 551100 334026 551336
rect 334262 551100 369706 551336
rect 369942 551100 370026 551336
rect 370262 551100 405706 551336
rect 405942 551100 406026 551336
rect 406262 551100 441706 551336
rect 441942 551100 442026 551336
rect 442262 551100 477706 551336
rect 477942 551100 478026 551336
rect 478262 551100 513706 551336
rect 513942 551100 514026 551336
rect 514262 551100 549706 551336
rect 549942 551100 550026 551336
rect 550262 551100 592062 551336
rect 592298 551100 592382 551336
rect 592618 551100 592650 551336
rect -8726 551016 592650 551100
rect -8726 550780 -8694 551016
rect -8458 550780 -8374 551016
rect -8138 550780 9706 551016
rect 9942 550780 10026 551016
rect 10262 550780 45706 551016
rect 45942 550780 46026 551016
rect 46262 550780 81706 551016
rect 81942 550780 82026 551016
rect 82262 550780 117706 551016
rect 117942 550780 118026 551016
rect 118262 550780 153706 551016
rect 153942 550780 154026 551016
rect 154262 550780 189706 551016
rect 189942 550780 190026 551016
rect 190262 550780 225706 551016
rect 225942 550780 226026 551016
rect 226262 550780 261706 551016
rect 261942 550780 262026 551016
rect 262262 550780 297706 551016
rect 297942 550780 298026 551016
rect 298262 550780 333706 551016
rect 333942 550780 334026 551016
rect 334262 550780 369706 551016
rect 369942 550780 370026 551016
rect 370262 550780 405706 551016
rect 405942 550780 406026 551016
rect 406262 550780 441706 551016
rect 441942 550780 442026 551016
rect 442262 550780 477706 551016
rect 477942 550780 478026 551016
rect 478262 550780 513706 551016
rect 513942 550780 514026 551016
rect 514262 550780 549706 551016
rect 549942 550780 550026 551016
rect 550262 550780 592062 551016
rect 592298 550780 592382 551016
rect 592618 550780 592650 551016
rect -8726 550748 592650 550780
rect -8726 550096 592650 550128
rect -8726 549860 -7734 550096
rect -7498 549860 -7414 550096
rect -7178 549860 8466 550096
rect 8702 549860 8786 550096
rect 9022 549860 44466 550096
rect 44702 549860 44786 550096
rect 45022 549860 80466 550096
rect 80702 549860 80786 550096
rect 81022 549860 116466 550096
rect 116702 549860 116786 550096
rect 117022 549860 152466 550096
rect 152702 549860 152786 550096
rect 153022 549860 188466 550096
rect 188702 549860 188786 550096
rect 189022 549860 224466 550096
rect 224702 549860 224786 550096
rect 225022 549860 260466 550096
rect 260702 549860 260786 550096
rect 261022 549860 296466 550096
rect 296702 549860 296786 550096
rect 297022 549860 332466 550096
rect 332702 549860 332786 550096
rect 333022 549860 368466 550096
rect 368702 549860 368786 550096
rect 369022 549860 404466 550096
rect 404702 549860 404786 550096
rect 405022 549860 440466 550096
rect 440702 549860 440786 550096
rect 441022 549860 476466 550096
rect 476702 549860 476786 550096
rect 477022 549860 512466 550096
rect 512702 549860 512786 550096
rect 513022 549860 548466 550096
rect 548702 549860 548786 550096
rect 549022 549860 591102 550096
rect 591338 549860 591422 550096
rect 591658 549860 592650 550096
rect -8726 549776 592650 549860
rect -8726 549540 -7734 549776
rect -7498 549540 -7414 549776
rect -7178 549540 8466 549776
rect 8702 549540 8786 549776
rect 9022 549540 44466 549776
rect 44702 549540 44786 549776
rect 45022 549540 80466 549776
rect 80702 549540 80786 549776
rect 81022 549540 116466 549776
rect 116702 549540 116786 549776
rect 117022 549540 152466 549776
rect 152702 549540 152786 549776
rect 153022 549540 188466 549776
rect 188702 549540 188786 549776
rect 189022 549540 224466 549776
rect 224702 549540 224786 549776
rect 225022 549540 260466 549776
rect 260702 549540 260786 549776
rect 261022 549540 296466 549776
rect 296702 549540 296786 549776
rect 297022 549540 332466 549776
rect 332702 549540 332786 549776
rect 333022 549540 368466 549776
rect 368702 549540 368786 549776
rect 369022 549540 404466 549776
rect 404702 549540 404786 549776
rect 405022 549540 440466 549776
rect 440702 549540 440786 549776
rect 441022 549540 476466 549776
rect 476702 549540 476786 549776
rect 477022 549540 512466 549776
rect 512702 549540 512786 549776
rect 513022 549540 548466 549776
rect 548702 549540 548786 549776
rect 549022 549540 591102 549776
rect 591338 549540 591422 549776
rect 591658 549540 592650 549776
rect -8726 549508 592650 549540
rect -8726 548856 592650 548888
rect -8726 548620 -6774 548856
rect -6538 548620 -6454 548856
rect -6218 548620 7226 548856
rect 7462 548620 7546 548856
rect 7782 548620 43226 548856
rect 43462 548620 43546 548856
rect 43782 548620 79226 548856
rect 79462 548620 79546 548856
rect 79782 548620 115226 548856
rect 115462 548620 115546 548856
rect 115782 548620 151226 548856
rect 151462 548620 151546 548856
rect 151782 548620 187226 548856
rect 187462 548620 187546 548856
rect 187782 548620 223226 548856
rect 223462 548620 223546 548856
rect 223782 548620 259226 548856
rect 259462 548620 259546 548856
rect 259782 548620 295226 548856
rect 295462 548620 295546 548856
rect 295782 548620 331226 548856
rect 331462 548620 331546 548856
rect 331782 548620 367226 548856
rect 367462 548620 367546 548856
rect 367782 548620 403226 548856
rect 403462 548620 403546 548856
rect 403782 548620 439226 548856
rect 439462 548620 439546 548856
rect 439782 548620 475226 548856
rect 475462 548620 475546 548856
rect 475782 548620 511226 548856
rect 511462 548620 511546 548856
rect 511782 548620 547226 548856
rect 547462 548620 547546 548856
rect 547782 548620 590142 548856
rect 590378 548620 590462 548856
rect 590698 548620 592650 548856
rect -8726 548536 592650 548620
rect -8726 548300 -6774 548536
rect -6538 548300 -6454 548536
rect -6218 548300 7226 548536
rect 7462 548300 7546 548536
rect 7782 548300 43226 548536
rect 43462 548300 43546 548536
rect 43782 548300 79226 548536
rect 79462 548300 79546 548536
rect 79782 548300 115226 548536
rect 115462 548300 115546 548536
rect 115782 548300 151226 548536
rect 151462 548300 151546 548536
rect 151782 548300 187226 548536
rect 187462 548300 187546 548536
rect 187782 548300 223226 548536
rect 223462 548300 223546 548536
rect 223782 548300 259226 548536
rect 259462 548300 259546 548536
rect 259782 548300 295226 548536
rect 295462 548300 295546 548536
rect 295782 548300 331226 548536
rect 331462 548300 331546 548536
rect 331782 548300 367226 548536
rect 367462 548300 367546 548536
rect 367782 548300 403226 548536
rect 403462 548300 403546 548536
rect 403782 548300 439226 548536
rect 439462 548300 439546 548536
rect 439782 548300 475226 548536
rect 475462 548300 475546 548536
rect 475782 548300 511226 548536
rect 511462 548300 511546 548536
rect 511782 548300 547226 548536
rect 547462 548300 547546 548536
rect 547782 548300 590142 548536
rect 590378 548300 590462 548536
rect 590698 548300 592650 548536
rect -8726 548268 592650 548300
rect -8726 547616 592650 547648
rect -8726 547380 -5814 547616
rect -5578 547380 -5494 547616
rect -5258 547380 5986 547616
rect 6222 547380 6306 547616
rect 6542 547380 41986 547616
rect 42222 547380 42306 547616
rect 42542 547380 77986 547616
rect 78222 547380 78306 547616
rect 78542 547380 113986 547616
rect 114222 547380 114306 547616
rect 114542 547380 149986 547616
rect 150222 547380 150306 547616
rect 150542 547380 185986 547616
rect 186222 547380 186306 547616
rect 186542 547380 221986 547616
rect 222222 547380 222306 547616
rect 222542 547380 257986 547616
rect 258222 547380 258306 547616
rect 258542 547380 293986 547616
rect 294222 547380 294306 547616
rect 294542 547380 329986 547616
rect 330222 547380 330306 547616
rect 330542 547380 365986 547616
rect 366222 547380 366306 547616
rect 366542 547380 401986 547616
rect 402222 547380 402306 547616
rect 402542 547380 437986 547616
rect 438222 547380 438306 547616
rect 438542 547380 473986 547616
rect 474222 547380 474306 547616
rect 474542 547380 509986 547616
rect 510222 547380 510306 547616
rect 510542 547380 545986 547616
rect 546222 547380 546306 547616
rect 546542 547380 581986 547616
rect 582222 547380 582306 547616
rect 582542 547380 589182 547616
rect 589418 547380 589502 547616
rect 589738 547380 592650 547616
rect -8726 547296 592650 547380
rect -8726 547060 -5814 547296
rect -5578 547060 -5494 547296
rect -5258 547060 5986 547296
rect 6222 547060 6306 547296
rect 6542 547060 41986 547296
rect 42222 547060 42306 547296
rect 42542 547060 77986 547296
rect 78222 547060 78306 547296
rect 78542 547060 113986 547296
rect 114222 547060 114306 547296
rect 114542 547060 149986 547296
rect 150222 547060 150306 547296
rect 150542 547060 185986 547296
rect 186222 547060 186306 547296
rect 186542 547060 221986 547296
rect 222222 547060 222306 547296
rect 222542 547060 257986 547296
rect 258222 547060 258306 547296
rect 258542 547060 293986 547296
rect 294222 547060 294306 547296
rect 294542 547060 329986 547296
rect 330222 547060 330306 547296
rect 330542 547060 365986 547296
rect 366222 547060 366306 547296
rect 366542 547060 401986 547296
rect 402222 547060 402306 547296
rect 402542 547060 437986 547296
rect 438222 547060 438306 547296
rect 438542 547060 473986 547296
rect 474222 547060 474306 547296
rect 474542 547060 509986 547296
rect 510222 547060 510306 547296
rect 510542 547060 545986 547296
rect 546222 547060 546306 547296
rect 546542 547060 581986 547296
rect 582222 547060 582306 547296
rect 582542 547060 589182 547296
rect 589418 547060 589502 547296
rect 589738 547060 592650 547296
rect -8726 547028 592650 547060
rect -8726 546376 592650 546408
rect -8726 546140 -4854 546376
rect -4618 546140 -4534 546376
rect -4298 546140 4746 546376
rect 4982 546140 5066 546376
rect 5302 546140 40746 546376
rect 40982 546140 41066 546376
rect 41302 546140 76746 546376
rect 76982 546140 77066 546376
rect 77302 546140 112746 546376
rect 112982 546140 113066 546376
rect 113302 546140 148746 546376
rect 148982 546140 149066 546376
rect 149302 546140 184746 546376
rect 184982 546140 185066 546376
rect 185302 546140 220746 546376
rect 220982 546140 221066 546376
rect 221302 546140 256746 546376
rect 256982 546140 257066 546376
rect 257302 546140 292746 546376
rect 292982 546140 293066 546376
rect 293302 546140 328746 546376
rect 328982 546140 329066 546376
rect 329302 546140 364746 546376
rect 364982 546140 365066 546376
rect 365302 546140 400746 546376
rect 400982 546140 401066 546376
rect 401302 546140 436746 546376
rect 436982 546140 437066 546376
rect 437302 546140 472746 546376
rect 472982 546140 473066 546376
rect 473302 546140 508746 546376
rect 508982 546140 509066 546376
rect 509302 546140 544746 546376
rect 544982 546140 545066 546376
rect 545302 546140 580746 546376
rect 580982 546140 581066 546376
rect 581302 546140 588222 546376
rect 588458 546140 588542 546376
rect 588778 546140 592650 546376
rect -8726 546056 592650 546140
rect -8726 545820 -4854 546056
rect -4618 545820 -4534 546056
rect -4298 545820 4746 546056
rect 4982 545820 5066 546056
rect 5302 545820 40746 546056
rect 40982 545820 41066 546056
rect 41302 545820 76746 546056
rect 76982 545820 77066 546056
rect 77302 545820 112746 546056
rect 112982 545820 113066 546056
rect 113302 545820 148746 546056
rect 148982 545820 149066 546056
rect 149302 545820 184746 546056
rect 184982 545820 185066 546056
rect 185302 545820 220746 546056
rect 220982 545820 221066 546056
rect 221302 545820 256746 546056
rect 256982 545820 257066 546056
rect 257302 545820 292746 546056
rect 292982 545820 293066 546056
rect 293302 545820 328746 546056
rect 328982 545820 329066 546056
rect 329302 545820 364746 546056
rect 364982 545820 365066 546056
rect 365302 545820 400746 546056
rect 400982 545820 401066 546056
rect 401302 545820 436746 546056
rect 436982 545820 437066 546056
rect 437302 545820 472746 546056
rect 472982 545820 473066 546056
rect 473302 545820 508746 546056
rect 508982 545820 509066 546056
rect 509302 545820 544746 546056
rect 544982 545820 545066 546056
rect 545302 545820 580746 546056
rect 580982 545820 581066 546056
rect 581302 545820 588222 546056
rect 588458 545820 588542 546056
rect 588778 545820 592650 546056
rect -8726 545788 592650 545820
rect -8726 545136 592650 545168
rect -8726 544900 -3894 545136
rect -3658 544900 -3574 545136
rect -3338 544900 3506 545136
rect 3742 544900 3826 545136
rect 4062 544900 39506 545136
rect 39742 544900 39826 545136
rect 40062 544900 75506 545136
rect 75742 544900 75826 545136
rect 76062 544900 111506 545136
rect 111742 544900 111826 545136
rect 112062 544900 147506 545136
rect 147742 544900 147826 545136
rect 148062 544900 183506 545136
rect 183742 544900 183826 545136
rect 184062 544900 219506 545136
rect 219742 544900 219826 545136
rect 220062 544900 255506 545136
rect 255742 544900 255826 545136
rect 256062 544900 291506 545136
rect 291742 544900 291826 545136
rect 292062 544900 327506 545136
rect 327742 544900 327826 545136
rect 328062 544900 363506 545136
rect 363742 544900 363826 545136
rect 364062 544900 399506 545136
rect 399742 544900 399826 545136
rect 400062 544900 435506 545136
rect 435742 544900 435826 545136
rect 436062 544900 471506 545136
rect 471742 544900 471826 545136
rect 472062 544900 507506 545136
rect 507742 544900 507826 545136
rect 508062 544900 543506 545136
rect 543742 544900 543826 545136
rect 544062 544900 579506 545136
rect 579742 544900 579826 545136
rect 580062 544900 587262 545136
rect 587498 544900 587582 545136
rect 587818 544900 592650 545136
rect -8726 544816 592650 544900
rect -8726 544580 -3894 544816
rect -3658 544580 -3574 544816
rect -3338 544580 3506 544816
rect 3742 544580 3826 544816
rect 4062 544580 39506 544816
rect 39742 544580 39826 544816
rect 40062 544580 75506 544816
rect 75742 544580 75826 544816
rect 76062 544580 111506 544816
rect 111742 544580 111826 544816
rect 112062 544580 147506 544816
rect 147742 544580 147826 544816
rect 148062 544580 183506 544816
rect 183742 544580 183826 544816
rect 184062 544580 219506 544816
rect 219742 544580 219826 544816
rect 220062 544580 255506 544816
rect 255742 544580 255826 544816
rect 256062 544580 291506 544816
rect 291742 544580 291826 544816
rect 292062 544580 327506 544816
rect 327742 544580 327826 544816
rect 328062 544580 363506 544816
rect 363742 544580 363826 544816
rect 364062 544580 399506 544816
rect 399742 544580 399826 544816
rect 400062 544580 435506 544816
rect 435742 544580 435826 544816
rect 436062 544580 471506 544816
rect 471742 544580 471826 544816
rect 472062 544580 507506 544816
rect 507742 544580 507826 544816
rect 508062 544580 543506 544816
rect 543742 544580 543826 544816
rect 544062 544580 579506 544816
rect 579742 544580 579826 544816
rect 580062 544580 587262 544816
rect 587498 544580 587582 544816
rect 587818 544580 592650 544816
rect -8726 544548 592650 544580
rect -8726 543896 592650 543928
rect -8726 543660 -2934 543896
rect -2698 543660 -2614 543896
rect -2378 543660 2266 543896
rect 2502 543660 2586 543896
rect 2822 543660 38266 543896
rect 38502 543660 38586 543896
rect 38822 543660 74266 543896
rect 74502 543660 74586 543896
rect 74822 543660 110266 543896
rect 110502 543660 110586 543896
rect 110822 543660 146266 543896
rect 146502 543660 146586 543896
rect 146822 543660 182266 543896
rect 182502 543660 182586 543896
rect 182822 543660 218266 543896
rect 218502 543660 218586 543896
rect 218822 543660 254266 543896
rect 254502 543660 254586 543896
rect 254822 543660 290266 543896
rect 290502 543660 290586 543896
rect 290822 543660 326266 543896
rect 326502 543660 326586 543896
rect 326822 543660 362266 543896
rect 362502 543660 362586 543896
rect 362822 543660 398266 543896
rect 398502 543660 398586 543896
rect 398822 543660 434266 543896
rect 434502 543660 434586 543896
rect 434822 543660 470266 543896
rect 470502 543660 470586 543896
rect 470822 543660 506266 543896
rect 506502 543660 506586 543896
rect 506822 543660 542266 543896
rect 542502 543660 542586 543896
rect 542822 543660 578266 543896
rect 578502 543660 578586 543896
rect 578822 543660 586302 543896
rect 586538 543660 586622 543896
rect 586858 543660 592650 543896
rect -8726 543576 592650 543660
rect -8726 543340 -2934 543576
rect -2698 543340 -2614 543576
rect -2378 543340 2266 543576
rect 2502 543340 2586 543576
rect 2822 543340 38266 543576
rect 38502 543340 38586 543576
rect 38822 543340 74266 543576
rect 74502 543340 74586 543576
rect 74822 543340 110266 543576
rect 110502 543340 110586 543576
rect 110822 543340 146266 543576
rect 146502 543340 146586 543576
rect 146822 543340 182266 543576
rect 182502 543340 182586 543576
rect 182822 543340 218266 543576
rect 218502 543340 218586 543576
rect 218822 543340 254266 543576
rect 254502 543340 254586 543576
rect 254822 543340 290266 543576
rect 290502 543340 290586 543576
rect 290822 543340 326266 543576
rect 326502 543340 326586 543576
rect 326822 543340 362266 543576
rect 362502 543340 362586 543576
rect 362822 543340 398266 543576
rect 398502 543340 398586 543576
rect 398822 543340 434266 543576
rect 434502 543340 434586 543576
rect 434822 543340 470266 543576
rect 470502 543340 470586 543576
rect 470822 543340 506266 543576
rect 506502 543340 506586 543576
rect 506822 543340 542266 543576
rect 542502 543340 542586 543576
rect 542822 543340 578266 543576
rect 578502 543340 578586 543576
rect 578822 543340 586302 543576
rect 586538 543340 586622 543576
rect 586858 543340 592650 543576
rect -8726 543308 592650 543340
rect -8726 542656 592650 542688
rect -8726 542420 -1974 542656
rect -1738 542420 -1654 542656
rect -1418 542420 1026 542656
rect 1262 542420 1346 542656
rect 1582 542420 37026 542656
rect 37262 542420 37346 542656
rect 37582 542420 73026 542656
rect 73262 542420 73346 542656
rect 73582 542420 109026 542656
rect 109262 542420 109346 542656
rect 109582 542420 145026 542656
rect 145262 542420 145346 542656
rect 145582 542420 181026 542656
rect 181262 542420 181346 542656
rect 181582 542420 217026 542656
rect 217262 542420 217346 542656
rect 217582 542420 253026 542656
rect 253262 542420 253346 542656
rect 253582 542420 289026 542656
rect 289262 542420 289346 542656
rect 289582 542420 325026 542656
rect 325262 542420 325346 542656
rect 325582 542420 361026 542656
rect 361262 542420 361346 542656
rect 361582 542420 397026 542656
rect 397262 542420 397346 542656
rect 397582 542420 433026 542656
rect 433262 542420 433346 542656
rect 433582 542420 469026 542656
rect 469262 542420 469346 542656
rect 469582 542420 505026 542656
rect 505262 542420 505346 542656
rect 505582 542420 541026 542656
rect 541262 542420 541346 542656
rect 541582 542420 577026 542656
rect 577262 542420 577346 542656
rect 577582 542420 585342 542656
rect 585578 542420 585662 542656
rect 585898 542420 592650 542656
rect -8726 542336 592650 542420
rect -8726 542100 -1974 542336
rect -1738 542100 -1654 542336
rect -1418 542100 1026 542336
rect 1262 542100 1346 542336
rect 1582 542100 37026 542336
rect 37262 542100 37346 542336
rect 37582 542100 73026 542336
rect 73262 542100 73346 542336
rect 73582 542100 109026 542336
rect 109262 542100 109346 542336
rect 109582 542100 145026 542336
rect 145262 542100 145346 542336
rect 145582 542100 181026 542336
rect 181262 542100 181346 542336
rect 181582 542100 217026 542336
rect 217262 542100 217346 542336
rect 217582 542100 253026 542336
rect 253262 542100 253346 542336
rect 253582 542100 289026 542336
rect 289262 542100 289346 542336
rect 289582 542100 325026 542336
rect 325262 542100 325346 542336
rect 325582 542100 361026 542336
rect 361262 542100 361346 542336
rect 361582 542100 397026 542336
rect 397262 542100 397346 542336
rect 397582 542100 433026 542336
rect 433262 542100 433346 542336
rect 433582 542100 469026 542336
rect 469262 542100 469346 542336
rect 469582 542100 505026 542336
rect 505262 542100 505346 542336
rect 505582 542100 541026 542336
rect 541262 542100 541346 542336
rect 541582 542100 577026 542336
rect 577262 542100 577346 542336
rect 577582 542100 585342 542336
rect 585578 542100 585662 542336
rect 585898 542100 592650 542336
rect -8726 542068 592650 542100
rect -8726 515336 592650 515368
rect -8726 515100 -8694 515336
rect -8458 515100 -8374 515336
rect -8138 515100 9706 515336
rect 9942 515100 10026 515336
rect 10262 515100 45706 515336
rect 45942 515100 46026 515336
rect 46262 515100 81706 515336
rect 81942 515100 82026 515336
rect 82262 515100 117706 515336
rect 117942 515100 118026 515336
rect 118262 515100 153706 515336
rect 153942 515100 154026 515336
rect 154262 515100 189706 515336
rect 189942 515100 190026 515336
rect 190262 515100 225706 515336
rect 225942 515100 226026 515336
rect 226262 515100 261706 515336
rect 261942 515100 262026 515336
rect 262262 515100 297706 515336
rect 297942 515100 298026 515336
rect 298262 515100 333706 515336
rect 333942 515100 334026 515336
rect 334262 515100 369706 515336
rect 369942 515100 370026 515336
rect 370262 515100 405706 515336
rect 405942 515100 406026 515336
rect 406262 515100 441706 515336
rect 441942 515100 442026 515336
rect 442262 515100 477706 515336
rect 477942 515100 478026 515336
rect 478262 515100 513706 515336
rect 513942 515100 514026 515336
rect 514262 515100 549706 515336
rect 549942 515100 550026 515336
rect 550262 515100 592062 515336
rect 592298 515100 592382 515336
rect 592618 515100 592650 515336
rect -8726 515016 592650 515100
rect -8726 514780 -8694 515016
rect -8458 514780 -8374 515016
rect -8138 514780 9706 515016
rect 9942 514780 10026 515016
rect 10262 514780 45706 515016
rect 45942 514780 46026 515016
rect 46262 514780 81706 515016
rect 81942 514780 82026 515016
rect 82262 514780 117706 515016
rect 117942 514780 118026 515016
rect 118262 514780 153706 515016
rect 153942 514780 154026 515016
rect 154262 514780 189706 515016
rect 189942 514780 190026 515016
rect 190262 514780 225706 515016
rect 225942 514780 226026 515016
rect 226262 514780 261706 515016
rect 261942 514780 262026 515016
rect 262262 514780 297706 515016
rect 297942 514780 298026 515016
rect 298262 514780 333706 515016
rect 333942 514780 334026 515016
rect 334262 514780 369706 515016
rect 369942 514780 370026 515016
rect 370262 514780 405706 515016
rect 405942 514780 406026 515016
rect 406262 514780 441706 515016
rect 441942 514780 442026 515016
rect 442262 514780 477706 515016
rect 477942 514780 478026 515016
rect 478262 514780 513706 515016
rect 513942 514780 514026 515016
rect 514262 514780 549706 515016
rect 549942 514780 550026 515016
rect 550262 514780 592062 515016
rect 592298 514780 592382 515016
rect 592618 514780 592650 515016
rect -8726 514748 592650 514780
rect -8726 514096 592650 514128
rect -8726 513860 -7734 514096
rect -7498 513860 -7414 514096
rect -7178 513860 8466 514096
rect 8702 513860 8786 514096
rect 9022 513860 44466 514096
rect 44702 513860 44786 514096
rect 45022 513860 80466 514096
rect 80702 513860 80786 514096
rect 81022 513860 116466 514096
rect 116702 513860 116786 514096
rect 117022 513860 152466 514096
rect 152702 513860 152786 514096
rect 153022 513860 188466 514096
rect 188702 513860 188786 514096
rect 189022 513860 224466 514096
rect 224702 513860 224786 514096
rect 225022 513860 260466 514096
rect 260702 513860 260786 514096
rect 261022 513860 296466 514096
rect 296702 513860 296786 514096
rect 297022 513860 332466 514096
rect 332702 513860 332786 514096
rect 333022 513860 368466 514096
rect 368702 513860 368786 514096
rect 369022 513860 404466 514096
rect 404702 513860 404786 514096
rect 405022 513860 440466 514096
rect 440702 513860 440786 514096
rect 441022 513860 476466 514096
rect 476702 513860 476786 514096
rect 477022 513860 512466 514096
rect 512702 513860 512786 514096
rect 513022 513860 548466 514096
rect 548702 513860 548786 514096
rect 549022 513860 591102 514096
rect 591338 513860 591422 514096
rect 591658 513860 592650 514096
rect -8726 513776 592650 513860
rect -8726 513540 -7734 513776
rect -7498 513540 -7414 513776
rect -7178 513540 8466 513776
rect 8702 513540 8786 513776
rect 9022 513540 44466 513776
rect 44702 513540 44786 513776
rect 45022 513540 80466 513776
rect 80702 513540 80786 513776
rect 81022 513540 116466 513776
rect 116702 513540 116786 513776
rect 117022 513540 152466 513776
rect 152702 513540 152786 513776
rect 153022 513540 188466 513776
rect 188702 513540 188786 513776
rect 189022 513540 224466 513776
rect 224702 513540 224786 513776
rect 225022 513540 260466 513776
rect 260702 513540 260786 513776
rect 261022 513540 296466 513776
rect 296702 513540 296786 513776
rect 297022 513540 332466 513776
rect 332702 513540 332786 513776
rect 333022 513540 368466 513776
rect 368702 513540 368786 513776
rect 369022 513540 404466 513776
rect 404702 513540 404786 513776
rect 405022 513540 440466 513776
rect 440702 513540 440786 513776
rect 441022 513540 476466 513776
rect 476702 513540 476786 513776
rect 477022 513540 512466 513776
rect 512702 513540 512786 513776
rect 513022 513540 548466 513776
rect 548702 513540 548786 513776
rect 549022 513540 591102 513776
rect 591338 513540 591422 513776
rect 591658 513540 592650 513776
rect -8726 513508 592650 513540
rect -8726 512856 592650 512888
rect -8726 512620 -6774 512856
rect -6538 512620 -6454 512856
rect -6218 512620 7226 512856
rect 7462 512620 7546 512856
rect 7782 512620 43226 512856
rect 43462 512620 43546 512856
rect 43782 512620 79226 512856
rect 79462 512620 79546 512856
rect 79782 512620 115226 512856
rect 115462 512620 115546 512856
rect 115782 512620 151226 512856
rect 151462 512620 151546 512856
rect 151782 512620 187226 512856
rect 187462 512620 187546 512856
rect 187782 512620 223226 512856
rect 223462 512620 223546 512856
rect 223782 512620 259226 512856
rect 259462 512620 259546 512856
rect 259782 512620 295226 512856
rect 295462 512620 295546 512856
rect 295782 512620 331226 512856
rect 331462 512620 331546 512856
rect 331782 512620 367226 512856
rect 367462 512620 367546 512856
rect 367782 512620 403226 512856
rect 403462 512620 403546 512856
rect 403782 512620 439226 512856
rect 439462 512620 439546 512856
rect 439782 512620 475226 512856
rect 475462 512620 475546 512856
rect 475782 512620 511226 512856
rect 511462 512620 511546 512856
rect 511782 512620 547226 512856
rect 547462 512620 547546 512856
rect 547782 512620 590142 512856
rect 590378 512620 590462 512856
rect 590698 512620 592650 512856
rect -8726 512536 592650 512620
rect -8726 512300 -6774 512536
rect -6538 512300 -6454 512536
rect -6218 512300 7226 512536
rect 7462 512300 7546 512536
rect 7782 512300 43226 512536
rect 43462 512300 43546 512536
rect 43782 512300 79226 512536
rect 79462 512300 79546 512536
rect 79782 512300 115226 512536
rect 115462 512300 115546 512536
rect 115782 512300 151226 512536
rect 151462 512300 151546 512536
rect 151782 512300 187226 512536
rect 187462 512300 187546 512536
rect 187782 512300 223226 512536
rect 223462 512300 223546 512536
rect 223782 512300 259226 512536
rect 259462 512300 259546 512536
rect 259782 512300 295226 512536
rect 295462 512300 295546 512536
rect 295782 512300 331226 512536
rect 331462 512300 331546 512536
rect 331782 512300 367226 512536
rect 367462 512300 367546 512536
rect 367782 512300 403226 512536
rect 403462 512300 403546 512536
rect 403782 512300 439226 512536
rect 439462 512300 439546 512536
rect 439782 512300 475226 512536
rect 475462 512300 475546 512536
rect 475782 512300 511226 512536
rect 511462 512300 511546 512536
rect 511782 512300 547226 512536
rect 547462 512300 547546 512536
rect 547782 512300 590142 512536
rect 590378 512300 590462 512536
rect 590698 512300 592650 512536
rect -8726 512268 592650 512300
rect -8726 511616 592650 511648
rect -8726 511380 -5814 511616
rect -5578 511380 -5494 511616
rect -5258 511380 5986 511616
rect 6222 511380 6306 511616
rect 6542 511380 41986 511616
rect 42222 511380 42306 511616
rect 42542 511380 77986 511616
rect 78222 511380 78306 511616
rect 78542 511380 113986 511616
rect 114222 511380 114306 511616
rect 114542 511380 149986 511616
rect 150222 511380 150306 511616
rect 150542 511380 185986 511616
rect 186222 511380 186306 511616
rect 186542 511380 221986 511616
rect 222222 511380 222306 511616
rect 222542 511380 257986 511616
rect 258222 511380 258306 511616
rect 258542 511380 293986 511616
rect 294222 511380 294306 511616
rect 294542 511380 329986 511616
rect 330222 511380 330306 511616
rect 330542 511380 365986 511616
rect 366222 511380 366306 511616
rect 366542 511380 401986 511616
rect 402222 511380 402306 511616
rect 402542 511380 437986 511616
rect 438222 511380 438306 511616
rect 438542 511380 473986 511616
rect 474222 511380 474306 511616
rect 474542 511380 509986 511616
rect 510222 511380 510306 511616
rect 510542 511380 545986 511616
rect 546222 511380 546306 511616
rect 546542 511380 581986 511616
rect 582222 511380 582306 511616
rect 582542 511380 589182 511616
rect 589418 511380 589502 511616
rect 589738 511380 592650 511616
rect -8726 511296 592650 511380
rect -8726 511060 -5814 511296
rect -5578 511060 -5494 511296
rect -5258 511060 5986 511296
rect 6222 511060 6306 511296
rect 6542 511060 41986 511296
rect 42222 511060 42306 511296
rect 42542 511060 77986 511296
rect 78222 511060 78306 511296
rect 78542 511060 113986 511296
rect 114222 511060 114306 511296
rect 114542 511060 149986 511296
rect 150222 511060 150306 511296
rect 150542 511060 185986 511296
rect 186222 511060 186306 511296
rect 186542 511060 221986 511296
rect 222222 511060 222306 511296
rect 222542 511060 257986 511296
rect 258222 511060 258306 511296
rect 258542 511060 293986 511296
rect 294222 511060 294306 511296
rect 294542 511060 329986 511296
rect 330222 511060 330306 511296
rect 330542 511060 365986 511296
rect 366222 511060 366306 511296
rect 366542 511060 401986 511296
rect 402222 511060 402306 511296
rect 402542 511060 437986 511296
rect 438222 511060 438306 511296
rect 438542 511060 473986 511296
rect 474222 511060 474306 511296
rect 474542 511060 509986 511296
rect 510222 511060 510306 511296
rect 510542 511060 545986 511296
rect 546222 511060 546306 511296
rect 546542 511060 581986 511296
rect 582222 511060 582306 511296
rect 582542 511060 589182 511296
rect 589418 511060 589502 511296
rect 589738 511060 592650 511296
rect -8726 511028 592650 511060
rect -8726 510376 592650 510408
rect -8726 510140 -4854 510376
rect -4618 510140 -4534 510376
rect -4298 510140 4746 510376
rect 4982 510140 5066 510376
rect 5302 510140 40746 510376
rect 40982 510140 41066 510376
rect 41302 510140 76746 510376
rect 76982 510140 77066 510376
rect 77302 510140 112746 510376
rect 112982 510140 113066 510376
rect 113302 510140 148746 510376
rect 148982 510140 149066 510376
rect 149302 510140 184746 510376
rect 184982 510140 185066 510376
rect 185302 510140 220746 510376
rect 220982 510140 221066 510376
rect 221302 510140 256746 510376
rect 256982 510140 257066 510376
rect 257302 510140 292746 510376
rect 292982 510140 293066 510376
rect 293302 510140 328746 510376
rect 328982 510140 329066 510376
rect 329302 510140 364746 510376
rect 364982 510140 365066 510376
rect 365302 510140 400746 510376
rect 400982 510140 401066 510376
rect 401302 510140 436746 510376
rect 436982 510140 437066 510376
rect 437302 510140 472746 510376
rect 472982 510140 473066 510376
rect 473302 510140 508746 510376
rect 508982 510140 509066 510376
rect 509302 510140 544746 510376
rect 544982 510140 545066 510376
rect 545302 510140 580746 510376
rect 580982 510140 581066 510376
rect 581302 510140 588222 510376
rect 588458 510140 588542 510376
rect 588778 510140 592650 510376
rect -8726 510056 592650 510140
rect -8726 509820 -4854 510056
rect -4618 509820 -4534 510056
rect -4298 509820 4746 510056
rect 4982 509820 5066 510056
rect 5302 509820 40746 510056
rect 40982 509820 41066 510056
rect 41302 509820 76746 510056
rect 76982 509820 77066 510056
rect 77302 509820 112746 510056
rect 112982 509820 113066 510056
rect 113302 509820 148746 510056
rect 148982 509820 149066 510056
rect 149302 509820 184746 510056
rect 184982 509820 185066 510056
rect 185302 509820 220746 510056
rect 220982 509820 221066 510056
rect 221302 509820 256746 510056
rect 256982 509820 257066 510056
rect 257302 509820 292746 510056
rect 292982 509820 293066 510056
rect 293302 509820 328746 510056
rect 328982 509820 329066 510056
rect 329302 509820 364746 510056
rect 364982 509820 365066 510056
rect 365302 509820 400746 510056
rect 400982 509820 401066 510056
rect 401302 509820 436746 510056
rect 436982 509820 437066 510056
rect 437302 509820 472746 510056
rect 472982 509820 473066 510056
rect 473302 509820 508746 510056
rect 508982 509820 509066 510056
rect 509302 509820 544746 510056
rect 544982 509820 545066 510056
rect 545302 509820 580746 510056
rect 580982 509820 581066 510056
rect 581302 509820 588222 510056
rect 588458 509820 588542 510056
rect 588778 509820 592650 510056
rect -8726 509788 592650 509820
rect -8726 509136 592650 509168
rect -8726 508900 -3894 509136
rect -3658 508900 -3574 509136
rect -3338 508900 3506 509136
rect 3742 508900 3826 509136
rect 4062 508900 39506 509136
rect 39742 508900 39826 509136
rect 40062 508900 75506 509136
rect 75742 508900 75826 509136
rect 76062 508900 111506 509136
rect 111742 508900 111826 509136
rect 112062 508900 147506 509136
rect 147742 508900 147826 509136
rect 148062 508900 183506 509136
rect 183742 508900 183826 509136
rect 184062 508900 219506 509136
rect 219742 508900 219826 509136
rect 220062 508900 255506 509136
rect 255742 508900 255826 509136
rect 256062 508900 291506 509136
rect 291742 508900 291826 509136
rect 292062 508900 327506 509136
rect 327742 508900 327826 509136
rect 328062 508900 363506 509136
rect 363742 508900 363826 509136
rect 364062 508900 399506 509136
rect 399742 508900 399826 509136
rect 400062 508900 435506 509136
rect 435742 508900 435826 509136
rect 436062 508900 471506 509136
rect 471742 508900 471826 509136
rect 472062 508900 507506 509136
rect 507742 508900 507826 509136
rect 508062 508900 543506 509136
rect 543742 508900 543826 509136
rect 544062 508900 579506 509136
rect 579742 508900 579826 509136
rect 580062 508900 587262 509136
rect 587498 508900 587582 509136
rect 587818 508900 592650 509136
rect -8726 508816 592650 508900
rect -8726 508580 -3894 508816
rect -3658 508580 -3574 508816
rect -3338 508580 3506 508816
rect 3742 508580 3826 508816
rect 4062 508580 39506 508816
rect 39742 508580 39826 508816
rect 40062 508580 75506 508816
rect 75742 508580 75826 508816
rect 76062 508580 111506 508816
rect 111742 508580 111826 508816
rect 112062 508580 147506 508816
rect 147742 508580 147826 508816
rect 148062 508580 183506 508816
rect 183742 508580 183826 508816
rect 184062 508580 219506 508816
rect 219742 508580 219826 508816
rect 220062 508580 255506 508816
rect 255742 508580 255826 508816
rect 256062 508580 291506 508816
rect 291742 508580 291826 508816
rect 292062 508580 327506 508816
rect 327742 508580 327826 508816
rect 328062 508580 363506 508816
rect 363742 508580 363826 508816
rect 364062 508580 399506 508816
rect 399742 508580 399826 508816
rect 400062 508580 435506 508816
rect 435742 508580 435826 508816
rect 436062 508580 471506 508816
rect 471742 508580 471826 508816
rect 472062 508580 507506 508816
rect 507742 508580 507826 508816
rect 508062 508580 543506 508816
rect 543742 508580 543826 508816
rect 544062 508580 579506 508816
rect 579742 508580 579826 508816
rect 580062 508580 587262 508816
rect 587498 508580 587582 508816
rect 587818 508580 592650 508816
rect -8726 508548 592650 508580
rect -8726 507896 592650 507928
rect -8726 507660 -2934 507896
rect -2698 507660 -2614 507896
rect -2378 507660 2266 507896
rect 2502 507660 2586 507896
rect 2822 507660 38266 507896
rect 38502 507660 38586 507896
rect 38822 507660 74266 507896
rect 74502 507660 74586 507896
rect 74822 507660 110266 507896
rect 110502 507660 110586 507896
rect 110822 507660 146266 507896
rect 146502 507660 146586 507896
rect 146822 507660 182266 507896
rect 182502 507660 182586 507896
rect 182822 507660 218266 507896
rect 218502 507660 218586 507896
rect 218822 507660 254266 507896
rect 254502 507660 254586 507896
rect 254822 507660 290266 507896
rect 290502 507660 290586 507896
rect 290822 507660 326266 507896
rect 326502 507660 326586 507896
rect 326822 507660 362266 507896
rect 362502 507660 362586 507896
rect 362822 507660 398266 507896
rect 398502 507660 398586 507896
rect 398822 507660 434266 507896
rect 434502 507660 434586 507896
rect 434822 507660 470266 507896
rect 470502 507660 470586 507896
rect 470822 507660 506266 507896
rect 506502 507660 506586 507896
rect 506822 507660 542266 507896
rect 542502 507660 542586 507896
rect 542822 507660 578266 507896
rect 578502 507660 578586 507896
rect 578822 507660 586302 507896
rect 586538 507660 586622 507896
rect 586858 507660 592650 507896
rect -8726 507576 592650 507660
rect -8726 507340 -2934 507576
rect -2698 507340 -2614 507576
rect -2378 507340 2266 507576
rect 2502 507340 2586 507576
rect 2822 507340 38266 507576
rect 38502 507340 38586 507576
rect 38822 507340 74266 507576
rect 74502 507340 74586 507576
rect 74822 507340 110266 507576
rect 110502 507340 110586 507576
rect 110822 507340 146266 507576
rect 146502 507340 146586 507576
rect 146822 507340 182266 507576
rect 182502 507340 182586 507576
rect 182822 507340 218266 507576
rect 218502 507340 218586 507576
rect 218822 507340 254266 507576
rect 254502 507340 254586 507576
rect 254822 507340 290266 507576
rect 290502 507340 290586 507576
rect 290822 507340 326266 507576
rect 326502 507340 326586 507576
rect 326822 507340 362266 507576
rect 362502 507340 362586 507576
rect 362822 507340 398266 507576
rect 398502 507340 398586 507576
rect 398822 507340 434266 507576
rect 434502 507340 434586 507576
rect 434822 507340 470266 507576
rect 470502 507340 470586 507576
rect 470822 507340 506266 507576
rect 506502 507340 506586 507576
rect 506822 507340 542266 507576
rect 542502 507340 542586 507576
rect 542822 507340 578266 507576
rect 578502 507340 578586 507576
rect 578822 507340 586302 507576
rect 586538 507340 586622 507576
rect 586858 507340 592650 507576
rect -8726 507308 592650 507340
rect -8726 506656 592650 506688
rect -8726 506420 -1974 506656
rect -1738 506420 -1654 506656
rect -1418 506420 1026 506656
rect 1262 506420 1346 506656
rect 1582 506420 37026 506656
rect 37262 506420 37346 506656
rect 37582 506420 73026 506656
rect 73262 506420 73346 506656
rect 73582 506420 109026 506656
rect 109262 506420 109346 506656
rect 109582 506420 145026 506656
rect 145262 506420 145346 506656
rect 145582 506420 181026 506656
rect 181262 506420 181346 506656
rect 181582 506420 217026 506656
rect 217262 506420 217346 506656
rect 217582 506420 253026 506656
rect 253262 506420 253346 506656
rect 253582 506420 289026 506656
rect 289262 506420 289346 506656
rect 289582 506420 325026 506656
rect 325262 506420 325346 506656
rect 325582 506420 361026 506656
rect 361262 506420 361346 506656
rect 361582 506420 397026 506656
rect 397262 506420 397346 506656
rect 397582 506420 433026 506656
rect 433262 506420 433346 506656
rect 433582 506420 469026 506656
rect 469262 506420 469346 506656
rect 469582 506420 505026 506656
rect 505262 506420 505346 506656
rect 505582 506420 541026 506656
rect 541262 506420 541346 506656
rect 541582 506420 577026 506656
rect 577262 506420 577346 506656
rect 577582 506420 585342 506656
rect 585578 506420 585662 506656
rect 585898 506420 592650 506656
rect -8726 506336 592650 506420
rect -8726 506100 -1974 506336
rect -1738 506100 -1654 506336
rect -1418 506100 1026 506336
rect 1262 506100 1346 506336
rect 1582 506100 37026 506336
rect 37262 506100 37346 506336
rect 37582 506100 73026 506336
rect 73262 506100 73346 506336
rect 73582 506100 109026 506336
rect 109262 506100 109346 506336
rect 109582 506100 145026 506336
rect 145262 506100 145346 506336
rect 145582 506100 181026 506336
rect 181262 506100 181346 506336
rect 181582 506100 217026 506336
rect 217262 506100 217346 506336
rect 217582 506100 253026 506336
rect 253262 506100 253346 506336
rect 253582 506100 289026 506336
rect 289262 506100 289346 506336
rect 289582 506100 325026 506336
rect 325262 506100 325346 506336
rect 325582 506100 361026 506336
rect 361262 506100 361346 506336
rect 361582 506100 397026 506336
rect 397262 506100 397346 506336
rect 397582 506100 433026 506336
rect 433262 506100 433346 506336
rect 433582 506100 469026 506336
rect 469262 506100 469346 506336
rect 469582 506100 505026 506336
rect 505262 506100 505346 506336
rect 505582 506100 541026 506336
rect 541262 506100 541346 506336
rect 541582 506100 577026 506336
rect 577262 506100 577346 506336
rect 577582 506100 585342 506336
rect 585578 506100 585662 506336
rect 585898 506100 592650 506336
rect -8726 506068 592650 506100
rect -8726 479336 592650 479368
rect -8726 479100 -8694 479336
rect -8458 479100 -8374 479336
rect -8138 479100 9706 479336
rect 9942 479100 10026 479336
rect 10262 479100 45706 479336
rect 45942 479100 46026 479336
rect 46262 479100 81706 479336
rect 81942 479100 82026 479336
rect 82262 479100 117706 479336
rect 117942 479100 118026 479336
rect 118262 479100 153706 479336
rect 153942 479100 154026 479336
rect 154262 479100 189706 479336
rect 189942 479100 190026 479336
rect 190262 479100 225706 479336
rect 225942 479100 226026 479336
rect 226262 479100 261706 479336
rect 261942 479100 262026 479336
rect 262262 479100 297706 479336
rect 297942 479100 298026 479336
rect 298262 479100 333706 479336
rect 333942 479100 334026 479336
rect 334262 479100 369706 479336
rect 369942 479100 370026 479336
rect 370262 479100 405706 479336
rect 405942 479100 406026 479336
rect 406262 479100 441706 479336
rect 441942 479100 442026 479336
rect 442262 479100 477706 479336
rect 477942 479100 478026 479336
rect 478262 479100 513706 479336
rect 513942 479100 514026 479336
rect 514262 479100 549706 479336
rect 549942 479100 550026 479336
rect 550262 479100 592062 479336
rect 592298 479100 592382 479336
rect 592618 479100 592650 479336
rect -8726 479016 592650 479100
rect -8726 478780 -8694 479016
rect -8458 478780 -8374 479016
rect -8138 478780 9706 479016
rect 9942 478780 10026 479016
rect 10262 478780 45706 479016
rect 45942 478780 46026 479016
rect 46262 478780 81706 479016
rect 81942 478780 82026 479016
rect 82262 478780 117706 479016
rect 117942 478780 118026 479016
rect 118262 478780 153706 479016
rect 153942 478780 154026 479016
rect 154262 478780 189706 479016
rect 189942 478780 190026 479016
rect 190262 478780 225706 479016
rect 225942 478780 226026 479016
rect 226262 478780 261706 479016
rect 261942 478780 262026 479016
rect 262262 478780 297706 479016
rect 297942 478780 298026 479016
rect 298262 478780 333706 479016
rect 333942 478780 334026 479016
rect 334262 478780 369706 479016
rect 369942 478780 370026 479016
rect 370262 478780 405706 479016
rect 405942 478780 406026 479016
rect 406262 478780 441706 479016
rect 441942 478780 442026 479016
rect 442262 478780 477706 479016
rect 477942 478780 478026 479016
rect 478262 478780 513706 479016
rect 513942 478780 514026 479016
rect 514262 478780 549706 479016
rect 549942 478780 550026 479016
rect 550262 478780 592062 479016
rect 592298 478780 592382 479016
rect 592618 478780 592650 479016
rect -8726 478748 592650 478780
rect -8726 478096 592650 478128
rect -8726 477860 -7734 478096
rect -7498 477860 -7414 478096
rect -7178 477860 8466 478096
rect 8702 477860 8786 478096
rect 9022 477860 44466 478096
rect 44702 477860 44786 478096
rect 45022 477860 80466 478096
rect 80702 477860 80786 478096
rect 81022 477860 116466 478096
rect 116702 477860 116786 478096
rect 117022 477860 152466 478096
rect 152702 477860 152786 478096
rect 153022 477860 188466 478096
rect 188702 477860 188786 478096
rect 189022 477860 224466 478096
rect 224702 477860 224786 478096
rect 225022 477860 260466 478096
rect 260702 477860 260786 478096
rect 261022 477860 296466 478096
rect 296702 477860 296786 478096
rect 297022 477860 332466 478096
rect 332702 477860 332786 478096
rect 333022 477860 368466 478096
rect 368702 477860 368786 478096
rect 369022 477860 404466 478096
rect 404702 477860 404786 478096
rect 405022 477860 440466 478096
rect 440702 477860 440786 478096
rect 441022 477860 476466 478096
rect 476702 477860 476786 478096
rect 477022 477860 512466 478096
rect 512702 477860 512786 478096
rect 513022 477860 548466 478096
rect 548702 477860 548786 478096
rect 549022 477860 591102 478096
rect 591338 477860 591422 478096
rect 591658 477860 592650 478096
rect -8726 477776 592650 477860
rect -8726 477540 -7734 477776
rect -7498 477540 -7414 477776
rect -7178 477540 8466 477776
rect 8702 477540 8786 477776
rect 9022 477540 44466 477776
rect 44702 477540 44786 477776
rect 45022 477540 80466 477776
rect 80702 477540 80786 477776
rect 81022 477540 116466 477776
rect 116702 477540 116786 477776
rect 117022 477540 152466 477776
rect 152702 477540 152786 477776
rect 153022 477540 188466 477776
rect 188702 477540 188786 477776
rect 189022 477540 224466 477776
rect 224702 477540 224786 477776
rect 225022 477540 260466 477776
rect 260702 477540 260786 477776
rect 261022 477540 296466 477776
rect 296702 477540 296786 477776
rect 297022 477540 332466 477776
rect 332702 477540 332786 477776
rect 333022 477540 368466 477776
rect 368702 477540 368786 477776
rect 369022 477540 404466 477776
rect 404702 477540 404786 477776
rect 405022 477540 440466 477776
rect 440702 477540 440786 477776
rect 441022 477540 476466 477776
rect 476702 477540 476786 477776
rect 477022 477540 512466 477776
rect 512702 477540 512786 477776
rect 513022 477540 548466 477776
rect 548702 477540 548786 477776
rect 549022 477540 591102 477776
rect 591338 477540 591422 477776
rect 591658 477540 592650 477776
rect -8726 477508 592650 477540
rect -8726 476856 592650 476888
rect -8726 476620 -6774 476856
rect -6538 476620 -6454 476856
rect -6218 476620 7226 476856
rect 7462 476620 7546 476856
rect 7782 476620 43226 476856
rect 43462 476620 43546 476856
rect 43782 476620 79226 476856
rect 79462 476620 79546 476856
rect 79782 476620 115226 476856
rect 115462 476620 115546 476856
rect 115782 476620 151226 476856
rect 151462 476620 151546 476856
rect 151782 476620 187226 476856
rect 187462 476620 187546 476856
rect 187782 476620 223226 476856
rect 223462 476620 223546 476856
rect 223782 476620 259226 476856
rect 259462 476620 259546 476856
rect 259782 476620 295226 476856
rect 295462 476620 295546 476856
rect 295782 476620 331226 476856
rect 331462 476620 331546 476856
rect 331782 476620 367226 476856
rect 367462 476620 367546 476856
rect 367782 476620 403226 476856
rect 403462 476620 403546 476856
rect 403782 476620 439226 476856
rect 439462 476620 439546 476856
rect 439782 476620 475226 476856
rect 475462 476620 475546 476856
rect 475782 476620 511226 476856
rect 511462 476620 511546 476856
rect 511782 476620 547226 476856
rect 547462 476620 547546 476856
rect 547782 476620 590142 476856
rect 590378 476620 590462 476856
rect 590698 476620 592650 476856
rect -8726 476536 592650 476620
rect -8726 476300 -6774 476536
rect -6538 476300 -6454 476536
rect -6218 476300 7226 476536
rect 7462 476300 7546 476536
rect 7782 476300 43226 476536
rect 43462 476300 43546 476536
rect 43782 476300 79226 476536
rect 79462 476300 79546 476536
rect 79782 476300 115226 476536
rect 115462 476300 115546 476536
rect 115782 476300 151226 476536
rect 151462 476300 151546 476536
rect 151782 476300 187226 476536
rect 187462 476300 187546 476536
rect 187782 476300 223226 476536
rect 223462 476300 223546 476536
rect 223782 476300 259226 476536
rect 259462 476300 259546 476536
rect 259782 476300 295226 476536
rect 295462 476300 295546 476536
rect 295782 476300 331226 476536
rect 331462 476300 331546 476536
rect 331782 476300 367226 476536
rect 367462 476300 367546 476536
rect 367782 476300 403226 476536
rect 403462 476300 403546 476536
rect 403782 476300 439226 476536
rect 439462 476300 439546 476536
rect 439782 476300 475226 476536
rect 475462 476300 475546 476536
rect 475782 476300 511226 476536
rect 511462 476300 511546 476536
rect 511782 476300 547226 476536
rect 547462 476300 547546 476536
rect 547782 476300 590142 476536
rect 590378 476300 590462 476536
rect 590698 476300 592650 476536
rect -8726 476268 592650 476300
rect -8726 475616 592650 475648
rect -8726 475380 -5814 475616
rect -5578 475380 -5494 475616
rect -5258 475380 5986 475616
rect 6222 475380 6306 475616
rect 6542 475380 41986 475616
rect 42222 475380 42306 475616
rect 42542 475380 77986 475616
rect 78222 475380 78306 475616
rect 78542 475380 113986 475616
rect 114222 475380 114306 475616
rect 114542 475380 149986 475616
rect 150222 475380 150306 475616
rect 150542 475380 185986 475616
rect 186222 475380 186306 475616
rect 186542 475380 221986 475616
rect 222222 475380 222306 475616
rect 222542 475380 257986 475616
rect 258222 475380 258306 475616
rect 258542 475380 293986 475616
rect 294222 475380 294306 475616
rect 294542 475380 329986 475616
rect 330222 475380 330306 475616
rect 330542 475380 365986 475616
rect 366222 475380 366306 475616
rect 366542 475380 401986 475616
rect 402222 475380 402306 475616
rect 402542 475380 437986 475616
rect 438222 475380 438306 475616
rect 438542 475380 473986 475616
rect 474222 475380 474306 475616
rect 474542 475380 509986 475616
rect 510222 475380 510306 475616
rect 510542 475380 545986 475616
rect 546222 475380 546306 475616
rect 546542 475380 581986 475616
rect 582222 475380 582306 475616
rect 582542 475380 589182 475616
rect 589418 475380 589502 475616
rect 589738 475380 592650 475616
rect -8726 475296 592650 475380
rect -8726 475060 -5814 475296
rect -5578 475060 -5494 475296
rect -5258 475060 5986 475296
rect 6222 475060 6306 475296
rect 6542 475060 41986 475296
rect 42222 475060 42306 475296
rect 42542 475060 77986 475296
rect 78222 475060 78306 475296
rect 78542 475060 113986 475296
rect 114222 475060 114306 475296
rect 114542 475060 149986 475296
rect 150222 475060 150306 475296
rect 150542 475060 185986 475296
rect 186222 475060 186306 475296
rect 186542 475060 221986 475296
rect 222222 475060 222306 475296
rect 222542 475060 257986 475296
rect 258222 475060 258306 475296
rect 258542 475060 293986 475296
rect 294222 475060 294306 475296
rect 294542 475060 329986 475296
rect 330222 475060 330306 475296
rect 330542 475060 365986 475296
rect 366222 475060 366306 475296
rect 366542 475060 401986 475296
rect 402222 475060 402306 475296
rect 402542 475060 437986 475296
rect 438222 475060 438306 475296
rect 438542 475060 473986 475296
rect 474222 475060 474306 475296
rect 474542 475060 509986 475296
rect 510222 475060 510306 475296
rect 510542 475060 545986 475296
rect 546222 475060 546306 475296
rect 546542 475060 581986 475296
rect 582222 475060 582306 475296
rect 582542 475060 589182 475296
rect 589418 475060 589502 475296
rect 589738 475060 592650 475296
rect -8726 475028 592650 475060
rect -8726 474376 592650 474408
rect -8726 474140 -4854 474376
rect -4618 474140 -4534 474376
rect -4298 474140 4746 474376
rect 4982 474140 5066 474376
rect 5302 474140 40746 474376
rect 40982 474140 41066 474376
rect 41302 474140 76746 474376
rect 76982 474140 77066 474376
rect 77302 474140 112746 474376
rect 112982 474140 113066 474376
rect 113302 474140 148746 474376
rect 148982 474140 149066 474376
rect 149302 474140 184746 474376
rect 184982 474140 185066 474376
rect 185302 474140 220746 474376
rect 220982 474140 221066 474376
rect 221302 474140 256746 474376
rect 256982 474140 257066 474376
rect 257302 474140 292746 474376
rect 292982 474140 293066 474376
rect 293302 474140 328746 474376
rect 328982 474140 329066 474376
rect 329302 474140 364746 474376
rect 364982 474140 365066 474376
rect 365302 474140 400746 474376
rect 400982 474140 401066 474376
rect 401302 474140 436746 474376
rect 436982 474140 437066 474376
rect 437302 474140 472746 474376
rect 472982 474140 473066 474376
rect 473302 474140 508746 474376
rect 508982 474140 509066 474376
rect 509302 474140 544746 474376
rect 544982 474140 545066 474376
rect 545302 474140 580746 474376
rect 580982 474140 581066 474376
rect 581302 474140 588222 474376
rect 588458 474140 588542 474376
rect 588778 474140 592650 474376
rect -8726 474056 592650 474140
rect -8726 473820 -4854 474056
rect -4618 473820 -4534 474056
rect -4298 473820 4746 474056
rect 4982 473820 5066 474056
rect 5302 473820 40746 474056
rect 40982 473820 41066 474056
rect 41302 473820 76746 474056
rect 76982 473820 77066 474056
rect 77302 473820 112746 474056
rect 112982 473820 113066 474056
rect 113302 473820 148746 474056
rect 148982 473820 149066 474056
rect 149302 473820 184746 474056
rect 184982 473820 185066 474056
rect 185302 473820 220746 474056
rect 220982 473820 221066 474056
rect 221302 473820 256746 474056
rect 256982 473820 257066 474056
rect 257302 473820 292746 474056
rect 292982 473820 293066 474056
rect 293302 473820 328746 474056
rect 328982 473820 329066 474056
rect 329302 473820 364746 474056
rect 364982 473820 365066 474056
rect 365302 473820 400746 474056
rect 400982 473820 401066 474056
rect 401302 473820 436746 474056
rect 436982 473820 437066 474056
rect 437302 473820 472746 474056
rect 472982 473820 473066 474056
rect 473302 473820 508746 474056
rect 508982 473820 509066 474056
rect 509302 473820 544746 474056
rect 544982 473820 545066 474056
rect 545302 473820 580746 474056
rect 580982 473820 581066 474056
rect 581302 473820 588222 474056
rect 588458 473820 588542 474056
rect 588778 473820 592650 474056
rect -8726 473788 592650 473820
rect -8726 473136 592650 473168
rect -8726 472900 -3894 473136
rect -3658 472900 -3574 473136
rect -3338 472900 3506 473136
rect 3742 472900 3826 473136
rect 4062 472900 39506 473136
rect 39742 472900 39826 473136
rect 40062 472900 75506 473136
rect 75742 472900 75826 473136
rect 76062 472900 111506 473136
rect 111742 472900 111826 473136
rect 112062 472900 147506 473136
rect 147742 472900 147826 473136
rect 148062 472900 183506 473136
rect 183742 472900 183826 473136
rect 184062 472900 219506 473136
rect 219742 472900 219826 473136
rect 220062 472900 255506 473136
rect 255742 472900 255826 473136
rect 256062 472900 291506 473136
rect 291742 472900 291826 473136
rect 292062 472900 327506 473136
rect 327742 472900 327826 473136
rect 328062 472900 363506 473136
rect 363742 472900 363826 473136
rect 364062 472900 399506 473136
rect 399742 472900 399826 473136
rect 400062 472900 435506 473136
rect 435742 472900 435826 473136
rect 436062 472900 471506 473136
rect 471742 472900 471826 473136
rect 472062 472900 507506 473136
rect 507742 472900 507826 473136
rect 508062 472900 543506 473136
rect 543742 472900 543826 473136
rect 544062 472900 579506 473136
rect 579742 472900 579826 473136
rect 580062 472900 587262 473136
rect 587498 472900 587582 473136
rect 587818 472900 592650 473136
rect -8726 472816 592650 472900
rect -8726 472580 -3894 472816
rect -3658 472580 -3574 472816
rect -3338 472580 3506 472816
rect 3742 472580 3826 472816
rect 4062 472580 39506 472816
rect 39742 472580 39826 472816
rect 40062 472580 75506 472816
rect 75742 472580 75826 472816
rect 76062 472580 111506 472816
rect 111742 472580 111826 472816
rect 112062 472580 147506 472816
rect 147742 472580 147826 472816
rect 148062 472580 183506 472816
rect 183742 472580 183826 472816
rect 184062 472580 219506 472816
rect 219742 472580 219826 472816
rect 220062 472580 255506 472816
rect 255742 472580 255826 472816
rect 256062 472580 291506 472816
rect 291742 472580 291826 472816
rect 292062 472580 327506 472816
rect 327742 472580 327826 472816
rect 328062 472580 363506 472816
rect 363742 472580 363826 472816
rect 364062 472580 399506 472816
rect 399742 472580 399826 472816
rect 400062 472580 435506 472816
rect 435742 472580 435826 472816
rect 436062 472580 471506 472816
rect 471742 472580 471826 472816
rect 472062 472580 507506 472816
rect 507742 472580 507826 472816
rect 508062 472580 543506 472816
rect 543742 472580 543826 472816
rect 544062 472580 579506 472816
rect 579742 472580 579826 472816
rect 580062 472580 587262 472816
rect 587498 472580 587582 472816
rect 587818 472580 592650 472816
rect -8726 472548 592650 472580
rect -8726 471896 592650 471928
rect -8726 471660 -2934 471896
rect -2698 471660 -2614 471896
rect -2378 471660 2266 471896
rect 2502 471660 2586 471896
rect 2822 471660 38266 471896
rect 38502 471660 38586 471896
rect 38822 471660 74266 471896
rect 74502 471660 74586 471896
rect 74822 471660 110266 471896
rect 110502 471660 110586 471896
rect 110822 471660 146266 471896
rect 146502 471660 146586 471896
rect 146822 471660 182266 471896
rect 182502 471660 182586 471896
rect 182822 471660 218266 471896
rect 218502 471660 218586 471896
rect 218822 471660 254266 471896
rect 254502 471660 254586 471896
rect 254822 471660 290266 471896
rect 290502 471660 290586 471896
rect 290822 471660 326266 471896
rect 326502 471660 326586 471896
rect 326822 471660 362266 471896
rect 362502 471660 362586 471896
rect 362822 471660 398266 471896
rect 398502 471660 398586 471896
rect 398822 471660 434266 471896
rect 434502 471660 434586 471896
rect 434822 471660 470266 471896
rect 470502 471660 470586 471896
rect 470822 471660 506266 471896
rect 506502 471660 506586 471896
rect 506822 471660 542266 471896
rect 542502 471660 542586 471896
rect 542822 471660 578266 471896
rect 578502 471660 578586 471896
rect 578822 471660 586302 471896
rect 586538 471660 586622 471896
rect 586858 471660 592650 471896
rect -8726 471576 592650 471660
rect -8726 471340 -2934 471576
rect -2698 471340 -2614 471576
rect -2378 471340 2266 471576
rect 2502 471340 2586 471576
rect 2822 471340 38266 471576
rect 38502 471340 38586 471576
rect 38822 471340 74266 471576
rect 74502 471340 74586 471576
rect 74822 471340 110266 471576
rect 110502 471340 110586 471576
rect 110822 471340 146266 471576
rect 146502 471340 146586 471576
rect 146822 471340 182266 471576
rect 182502 471340 182586 471576
rect 182822 471340 218266 471576
rect 218502 471340 218586 471576
rect 218822 471340 254266 471576
rect 254502 471340 254586 471576
rect 254822 471340 290266 471576
rect 290502 471340 290586 471576
rect 290822 471340 326266 471576
rect 326502 471340 326586 471576
rect 326822 471340 362266 471576
rect 362502 471340 362586 471576
rect 362822 471340 398266 471576
rect 398502 471340 398586 471576
rect 398822 471340 434266 471576
rect 434502 471340 434586 471576
rect 434822 471340 470266 471576
rect 470502 471340 470586 471576
rect 470822 471340 506266 471576
rect 506502 471340 506586 471576
rect 506822 471340 542266 471576
rect 542502 471340 542586 471576
rect 542822 471340 578266 471576
rect 578502 471340 578586 471576
rect 578822 471340 586302 471576
rect 586538 471340 586622 471576
rect 586858 471340 592650 471576
rect -8726 471308 592650 471340
rect -8726 470656 592650 470688
rect -8726 470420 -1974 470656
rect -1738 470420 -1654 470656
rect -1418 470420 1026 470656
rect 1262 470420 1346 470656
rect 1582 470420 37026 470656
rect 37262 470420 37346 470656
rect 37582 470420 73026 470656
rect 73262 470420 73346 470656
rect 73582 470420 109026 470656
rect 109262 470420 109346 470656
rect 109582 470420 145026 470656
rect 145262 470420 145346 470656
rect 145582 470420 181026 470656
rect 181262 470420 181346 470656
rect 181582 470420 217026 470656
rect 217262 470420 217346 470656
rect 217582 470420 253026 470656
rect 253262 470420 253346 470656
rect 253582 470420 289026 470656
rect 289262 470420 289346 470656
rect 289582 470420 325026 470656
rect 325262 470420 325346 470656
rect 325582 470420 361026 470656
rect 361262 470420 361346 470656
rect 361582 470420 397026 470656
rect 397262 470420 397346 470656
rect 397582 470420 433026 470656
rect 433262 470420 433346 470656
rect 433582 470420 469026 470656
rect 469262 470420 469346 470656
rect 469582 470420 505026 470656
rect 505262 470420 505346 470656
rect 505582 470420 541026 470656
rect 541262 470420 541346 470656
rect 541582 470420 577026 470656
rect 577262 470420 577346 470656
rect 577582 470420 585342 470656
rect 585578 470420 585662 470656
rect 585898 470420 592650 470656
rect -8726 470336 592650 470420
rect -8726 470100 -1974 470336
rect -1738 470100 -1654 470336
rect -1418 470100 1026 470336
rect 1262 470100 1346 470336
rect 1582 470100 37026 470336
rect 37262 470100 37346 470336
rect 37582 470100 73026 470336
rect 73262 470100 73346 470336
rect 73582 470100 109026 470336
rect 109262 470100 109346 470336
rect 109582 470100 145026 470336
rect 145262 470100 145346 470336
rect 145582 470100 181026 470336
rect 181262 470100 181346 470336
rect 181582 470100 217026 470336
rect 217262 470100 217346 470336
rect 217582 470100 253026 470336
rect 253262 470100 253346 470336
rect 253582 470100 289026 470336
rect 289262 470100 289346 470336
rect 289582 470100 325026 470336
rect 325262 470100 325346 470336
rect 325582 470100 361026 470336
rect 361262 470100 361346 470336
rect 361582 470100 397026 470336
rect 397262 470100 397346 470336
rect 397582 470100 433026 470336
rect 433262 470100 433346 470336
rect 433582 470100 469026 470336
rect 469262 470100 469346 470336
rect 469582 470100 505026 470336
rect 505262 470100 505346 470336
rect 505582 470100 541026 470336
rect 541262 470100 541346 470336
rect 541582 470100 577026 470336
rect 577262 470100 577346 470336
rect 577582 470100 585342 470336
rect 585578 470100 585662 470336
rect 585898 470100 592650 470336
rect -8726 470068 592650 470100
rect -8726 443336 592650 443368
rect -8726 443100 -8694 443336
rect -8458 443100 -8374 443336
rect -8138 443100 9706 443336
rect 9942 443100 10026 443336
rect 10262 443100 45706 443336
rect 45942 443100 46026 443336
rect 46262 443100 81706 443336
rect 81942 443100 82026 443336
rect 82262 443100 117706 443336
rect 117942 443100 118026 443336
rect 118262 443100 153706 443336
rect 153942 443100 154026 443336
rect 154262 443100 189706 443336
rect 189942 443100 190026 443336
rect 190262 443100 225706 443336
rect 225942 443100 226026 443336
rect 226262 443100 261706 443336
rect 261942 443100 262026 443336
rect 262262 443100 297706 443336
rect 297942 443100 298026 443336
rect 298262 443100 333706 443336
rect 333942 443100 334026 443336
rect 334262 443100 369706 443336
rect 369942 443100 370026 443336
rect 370262 443100 405706 443336
rect 405942 443100 406026 443336
rect 406262 443100 441706 443336
rect 441942 443100 442026 443336
rect 442262 443100 477706 443336
rect 477942 443100 478026 443336
rect 478262 443100 513706 443336
rect 513942 443100 514026 443336
rect 514262 443100 549706 443336
rect 549942 443100 550026 443336
rect 550262 443100 592062 443336
rect 592298 443100 592382 443336
rect 592618 443100 592650 443336
rect -8726 443016 592650 443100
rect -8726 442780 -8694 443016
rect -8458 442780 -8374 443016
rect -8138 442780 9706 443016
rect 9942 442780 10026 443016
rect 10262 442780 45706 443016
rect 45942 442780 46026 443016
rect 46262 442780 81706 443016
rect 81942 442780 82026 443016
rect 82262 442780 117706 443016
rect 117942 442780 118026 443016
rect 118262 442780 153706 443016
rect 153942 442780 154026 443016
rect 154262 442780 189706 443016
rect 189942 442780 190026 443016
rect 190262 442780 225706 443016
rect 225942 442780 226026 443016
rect 226262 442780 261706 443016
rect 261942 442780 262026 443016
rect 262262 442780 297706 443016
rect 297942 442780 298026 443016
rect 298262 442780 333706 443016
rect 333942 442780 334026 443016
rect 334262 442780 369706 443016
rect 369942 442780 370026 443016
rect 370262 442780 405706 443016
rect 405942 442780 406026 443016
rect 406262 442780 441706 443016
rect 441942 442780 442026 443016
rect 442262 442780 477706 443016
rect 477942 442780 478026 443016
rect 478262 442780 513706 443016
rect 513942 442780 514026 443016
rect 514262 442780 549706 443016
rect 549942 442780 550026 443016
rect 550262 442780 592062 443016
rect 592298 442780 592382 443016
rect 592618 442780 592650 443016
rect -8726 442748 592650 442780
rect -8726 442096 592650 442128
rect -8726 441860 -7734 442096
rect -7498 441860 -7414 442096
rect -7178 441860 8466 442096
rect 8702 441860 8786 442096
rect 9022 441860 44466 442096
rect 44702 441860 44786 442096
rect 45022 441860 80466 442096
rect 80702 441860 80786 442096
rect 81022 441860 116466 442096
rect 116702 441860 116786 442096
rect 117022 441860 152466 442096
rect 152702 441860 152786 442096
rect 153022 441860 188466 442096
rect 188702 441860 188786 442096
rect 189022 441860 224466 442096
rect 224702 441860 224786 442096
rect 225022 441860 260466 442096
rect 260702 441860 260786 442096
rect 261022 441860 296466 442096
rect 296702 441860 296786 442096
rect 297022 441860 332466 442096
rect 332702 441860 332786 442096
rect 333022 441860 368466 442096
rect 368702 441860 368786 442096
rect 369022 441860 404466 442096
rect 404702 441860 404786 442096
rect 405022 441860 440466 442096
rect 440702 441860 440786 442096
rect 441022 441860 476466 442096
rect 476702 441860 476786 442096
rect 477022 441860 512466 442096
rect 512702 441860 512786 442096
rect 513022 441860 548466 442096
rect 548702 441860 548786 442096
rect 549022 441860 591102 442096
rect 591338 441860 591422 442096
rect 591658 441860 592650 442096
rect -8726 441776 592650 441860
rect -8726 441540 -7734 441776
rect -7498 441540 -7414 441776
rect -7178 441540 8466 441776
rect 8702 441540 8786 441776
rect 9022 441540 44466 441776
rect 44702 441540 44786 441776
rect 45022 441540 80466 441776
rect 80702 441540 80786 441776
rect 81022 441540 116466 441776
rect 116702 441540 116786 441776
rect 117022 441540 152466 441776
rect 152702 441540 152786 441776
rect 153022 441540 188466 441776
rect 188702 441540 188786 441776
rect 189022 441540 224466 441776
rect 224702 441540 224786 441776
rect 225022 441540 260466 441776
rect 260702 441540 260786 441776
rect 261022 441540 296466 441776
rect 296702 441540 296786 441776
rect 297022 441540 332466 441776
rect 332702 441540 332786 441776
rect 333022 441540 368466 441776
rect 368702 441540 368786 441776
rect 369022 441540 404466 441776
rect 404702 441540 404786 441776
rect 405022 441540 440466 441776
rect 440702 441540 440786 441776
rect 441022 441540 476466 441776
rect 476702 441540 476786 441776
rect 477022 441540 512466 441776
rect 512702 441540 512786 441776
rect 513022 441540 548466 441776
rect 548702 441540 548786 441776
rect 549022 441540 591102 441776
rect 591338 441540 591422 441776
rect 591658 441540 592650 441776
rect -8726 441508 592650 441540
rect -8726 440856 592650 440888
rect -8726 440620 -6774 440856
rect -6538 440620 -6454 440856
rect -6218 440620 7226 440856
rect 7462 440620 7546 440856
rect 7782 440620 43226 440856
rect 43462 440620 43546 440856
rect 43782 440620 79226 440856
rect 79462 440620 79546 440856
rect 79782 440620 115226 440856
rect 115462 440620 115546 440856
rect 115782 440620 151226 440856
rect 151462 440620 151546 440856
rect 151782 440620 187226 440856
rect 187462 440620 187546 440856
rect 187782 440620 223226 440856
rect 223462 440620 223546 440856
rect 223782 440620 259226 440856
rect 259462 440620 259546 440856
rect 259782 440620 295226 440856
rect 295462 440620 295546 440856
rect 295782 440620 331226 440856
rect 331462 440620 331546 440856
rect 331782 440620 367226 440856
rect 367462 440620 367546 440856
rect 367782 440620 403226 440856
rect 403462 440620 403546 440856
rect 403782 440620 439226 440856
rect 439462 440620 439546 440856
rect 439782 440620 475226 440856
rect 475462 440620 475546 440856
rect 475782 440620 511226 440856
rect 511462 440620 511546 440856
rect 511782 440620 547226 440856
rect 547462 440620 547546 440856
rect 547782 440620 590142 440856
rect 590378 440620 590462 440856
rect 590698 440620 592650 440856
rect -8726 440536 592650 440620
rect -8726 440300 -6774 440536
rect -6538 440300 -6454 440536
rect -6218 440300 7226 440536
rect 7462 440300 7546 440536
rect 7782 440300 43226 440536
rect 43462 440300 43546 440536
rect 43782 440300 79226 440536
rect 79462 440300 79546 440536
rect 79782 440300 115226 440536
rect 115462 440300 115546 440536
rect 115782 440300 151226 440536
rect 151462 440300 151546 440536
rect 151782 440300 187226 440536
rect 187462 440300 187546 440536
rect 187782 440300 223226 440536
rect 223462 440300 223546 440536
rect 223782 440300 259226 440536
rect 259462 440300 259546 440536
rect 259782 440300 295226 440536
rect 295462 440300 295546 440536
rect 295782 440300 331226 440536
rect 331462 440300 331546 440536
rect 331782 440300 367226 440536
rect 367462 440300 367546 440536
rect 367782 440300 403226 440536
rect 403462 440300 403546 440536
rect 403782 440300 439226 440536
rect 439462 440300 439546 440536
rect 439782 440300 475226 440536
rect 475462 440300 475546 440536
rect 475782 440300 511226 440536
rect 511462 440300 511546 440536
rect 511782 440300 547226 440536
rect 547462 440300 547546 440536
rect 547782 440300 590142 440536
rect 590378 440300 590462 440536
rect 590698 440300 592650 440536
rect -8726 440268 592650 440300
rect -8726 439616 592650 439648
rect -8726 439380 -5814 439616
rect -5578 439380 -5494 439616
rect -5258 439380 5986 439616
rect 6222 439380 6306 439616
rect 6542 439380 41986 439616
rect 42222 439380 42306 439616
rect 42542 439380 77986 439616
rect 78222 439380 78306 439616
rect 78542 439380 113986 439616
rect 114222 439380 114306 439616
rect 114542 439380 149986 439616
rect 150222 439380 150306 439616
rect 150542 439380 185986 439616
rect 186222 439380 186306 439616
rect 186542 439380 221986 439616
rect 222222 439380 222306 439616
rect 222542 439380 257986 439616
rect 258222 439380 258306 439616
rect 258542 439380 293986 439616
rect 294222 439380 294306 439616
rect 294542 439380 329986 439616
rect 330222 439380 330306 439616
rect 330542 439380 365986 439616
rect 366222 439380 366306 439616
rect 366542 439380 401986 439616
rect 402222 439380 402306 439616
rect 402542 439380 437986 439616
rect 438222 439380 438306 439616
rect 438542 439380 473986 439616
rect 474222 439380 474306 439616
rect 474542 439380 509986 439616
rect 510222 439380 510306 439616
rect 510542 439380 581986 439616
rect 582222 439380 582306 439616
rect 582542 439380 589182 439616
rect 589418 439380 589502 439616
rect 589738 439380 592650 439616
rect -8726 439296 592650 439380
rect -8726 439060 -5814 439296
rect -5578 439060 -5494 439296
rect -5258 439060 5986 439296
rect 6222 439060 6306 439296
rect 6542 439060 41986 439296
rect 42222 439060 42306 439296
rect 42542 439060 77986 439296
rect 78222 439060 78306 439296
rect 78542 439060 113986 439296
rect 114222 439060 114306 439296
rect 114542 439060 149986 439296
rect 150222 439060 150306 439296
rect 150542 439060 185986 439296
rect 186222 439060 186306 439296
rect 186542 439060 221986 439296
rect 222222 439060 222306 439296
rect 222542 439060 257986 439296
rect 258222 439060 258306 439296
rect 258542 439060 293986 439296
rect 294222 439060 294306 439296
rect 294542 439060 329986 439296
rect 330222 439060 330306 439296
rect 330542 439060 365986 439296
rect 366222 439060 366306 439296
rect 366542 439060 401986 439296
rect 402222 439060 402306 439296
rect 402542 439060 437986 439296
rect 438222 439060 438306 439296
rect 438542 439060 473986 439296
rect 474222 439060 474306 439296
rect 474542 439060 509986 439296
rect 510222 439060 510306 439296
rect 510542 439060 581986 439296
rect 582222 439060 582306 439296
rect 582542 439060 589182 439296
rect 589418 439060 589502 439296
rect 589738 439060 592650 439296
rect -8726 439028 592650 439060
rect -8726 438376 592650 438408
rect -8726 438140 -4854 438376
rect -4618 438140 -4534 438376
rect -4298 438140 4746 438376
rect 4982 438140 5066 438376
rect 5302 438140 40746 438376
rect 40982 438140 41066 438376
rect 41302 438140 76746 438376
rect 76982 438140 77066 438376
rect 77302 438140 112746 438376
rect 112982 438140 113066 438376
rect 113302 438140 148746 438376
rect 148982 438140 149066 438376
rect 149302 438140 184746 438376
rect 184982 438140 185066 438376
rect 185302 438140 220746 438376
rect 220982 438140 221066 438376
rect 221302 438140 256746 438376
rect 256982 438140 257066 438376
rect 257302 438140 292746 438376
rect 292982 438140 293066 438376
rect 293302 438140 328746 438376
rect 328982 438140 329066 438376
rect 329302 438140 364746 438376
rect 364982 438140 365066 438376
rect 365302 438140 400746 438376
rect 400982 438140 401066 438376
rect 401302 438140 436746 438376
rect 436982 438140 437066 438376
rect 437302 438140 472746 438376
rect 472982 438140 473066 438376
rect 473302 438140 508746 438376
rect 508982 438140 509066 438376
rect 509302 438140 580746 438376
rect 580982 438140 581066 438376
rect 581302 438140 588222 438376
rect 588458 438140 588542 438376
rect 588778 438140 592650 438376
rect -8726 438056 592650 438140
rect -8726 437820 -4854 438056
rect -4618 437820 -4534 438056
rect -4298 437820 4746 438056
rect 4982 437820 5066 438056
rect 5302 437820 40746 438056
rect 40982 437820 41066 438056
rect 41302 437820 76746 438056
rect 76982 437820 77066 438056
rect 77302 437820 112746 438056
rect 112982 437820 113066 438056
rect 113302 437820 148746 438056
rect 148982 437820 149066 438056
rect 149302 437820 184746 438056
rect 184982 437820 185066 438056
rect 185302 437820 220746 438056
rect 220982 437820 221066 438056
rect 221302 437820 256746 438056
rect 256982 437820 257066 438056
rect 257302 437820 292746 438056
rect 292982 437820 293066 438056
rect 293302 437820 328746 438056
rect 328982 437820 329066 438056
rect 329302 437820 364746 438056
rect 364982 437820 365066 438056
rect 365302 437820 400746 438056
rect 400982 437820 401066 438056
rect 401302 437820 436746 438056
rect 436982 437820 437066 438056
rect 437302 437820 472746 438056
rect 472982 437820 473066 438056
rect 473302 437820 508746 438056
rect 508982 437820 509066 438056
rect 509302 437820 580746 438056
rect 580982 437820 581066 438056
rect 581302 437820 588222 438056
rect 588458 437820 588542 438056
rect 588778 437820 592650 438056
rect -8726 437788 592650 437820
rect -8726 437136 592650 437168
rect -8726 436900 -3894 437136
rect -3658 436900 -3574 437136
rect -3338 436900 3506 437136
rect 3742 436900 3826 437136
rect 4062 436900 39506 437136
rect 39742 436900 39826 437136
rect 40062 436900 75506 437136
rect 75742 436900 75826 437136
rect 76062 436900 111506 437136
rect 111742 436900 111826 437136
rect 112062 436900 147506 437136
rect 147742 436900 147826 437136
rect 148062 436900 183506 437136
rect 183742 436900 183826 437136
rect 184062 436900 219506 437136
rect 219742 436900 219826 437136
rect 220062 436900 255506 437136
rect 255742 436900 255826 437136
rect 256062 436900 291506 437136
rect 291742 436900 291826 437136
rect 292062 436900 327506 437136
rect 327742 436900 327826 437136
rect 328062 436900 363506 437136
rect 363742 436900 363826 437136
rect 364062 436900 399506 437136
rect 399742 436900 399826 437136
rect 400062 436900 435506 437136
rect 435742 436900 435826 437136
rect 436062 436900 471506 437136
rect 471742 436900 471826 437136
rect 472062 436900 507506 437136
rect 507742 436900 507826 437136
rect 508062 436900 579506 437136
rect 579742 436900 579826 437136
rect 580062 436900 587262 437136
rect 587498 436900 587582 437136
rect 587818 436900 592650 437136
rect -8726 436816 592650 436900
rect -8726 436580 -3894 436816
rect -3658 436580 -3574 436816
rect -3338 436580 3506 436816
rect 3742 436580 3826 436816
rect 4062 436580 39506 436816
rect 39742 436580 39826 436816
rect 40062 436580 75506 436816
rect 75742 436580 75826 436816
rect 76062 436580 111506 436816
rect 111742 436580 111826 436816
rect 112062 436580 147506 436816
rect 147742 436580 147826 436816
rect 148062 436580 183506 436816
rect 183742 436580 183826 436816
rect 184062 436580 219506 436816
rect 219742 436580 219826 436816
rect 220062 436580 255506 436816
rect 255742 436580 255826 436816
rect 256062 436580 291506 436816
rect 291742 436580 291826 436816
rect 292062 436580 327506 436816
rect 327742 436580 327826 436816
rect 328062 436580 363506 436816
rect 363742 436580 363826 436816
rect 364062 436580 399506 436816
rect 399742 436580 399826 436816
rect 400062 436580 435506 436816
rect 435742 436580 435826 436816
rect 436062 436580 471506 436816
rect 471742 436580 471826 436816
rect 472062 436580 507506 436816
rect 507742 436580 507826 436816
rect 508062 436580 579506 436816
rect 579742 436580 579826 436816
rect 580062 436580 587262 436816
rect 587498 436580 587582 436816
rect 587818 436580 592650 436816
rect -8726 436548 592650 436580
rect -8726 435896 592650 435928
rect -8726 435660 -2934 435896
rect -2698 435660 -2614 435896
rect -2378 435660 2266 435896
rect 2502 435660 2586 435896
rect 2822 435660 38266 435896
rect 38502 435660 38586 435896
rect 38822 435660 74266 435896
rect 74502 435660 74586 435896
rect 74822 435660 110266 435896
rect 110502 435660 110586 435896
rect 110822 435660 146266 435896
rect 146502 435660 146586 435896
rect 146822 435660 182266 435896
rect 182502 435660 182586 435896
rect 182822 435660 218266 435896
rect 218502 435660 218586 435896
rect 218822 435660 254266 435896
rect 254502 435660 254586 435896
rect 254822 435660 290266 435896
rect 290502 435660 290586 435896
rect 290822 435660 326266 435896
rect 326502 435660 326586 435896
rect 326822 435660 362266 435896
rect 362502 435660 362586 435896
rect 362822 435660 398266 435896
rect 398502 435660 398586 435896
rect 398822 435660 434266 435896
rect 434502 435660 434586 435896
rect 434822 435660 470266 435896
rect 470502 435660 470586 435896
rect 470822 435660 506266 435896
rect 506502 435660 506586 435896
rect 506822 435660 540918 435896
rect 541154 435660 542850 435896
rect 543086 435660 544782 435896
rect 545018 435660 546714 435896
rect 546950 435660 578266 435896
rect 578502 435660 578586 435896
rect 578822 435660 586302 435896
rect 586538 435660 586622 435896
rect 586858 435660 592650 435896
rect -8726 435576 592650 435660
rect -8726 435340 -2934 435576
rect -2698 435340 -2614 435576
rect -2378 435340 2266 435576
rect 2502 435340 2586 435576
rect 2822 435340 38266 435576
rect 38502 435340 38586 435576
rect 38822 435340 74266 435576
rect 74502 435340 74586 435576
rect 74822 435340 110266 435576
rect 110502 435340 110586 435576
rect 110822 435340 146266 435576
rect 146502 435340 146586 435576
rect 146822 435340 182266 435576
rect 182502 435340 182586 435576
rect 182822 435340 218266 435576
rect 218502 435340 218586 435576
rect 218822 435340 254266 435576
rect 254502 435340 254586 435576
rect 254822 435340 290266 435576
rect 290502 435340 290586 435576
rect 290822 435340 326266 435576
rect 326502 435340 326586 435576
rect 326822 435340 362266 435576
rect 362502 435340 362586 435576
rect 362822 435340 398266 435576
rect 398502 435340 398586 435576
rect 398822 435340 434266 435576
rect 434502 435340 434586 435576
rect 434822 435340 470266 435576
rect 470502 435340 470586 435576
rect 470822 435340 506266 435576
rect 506502 435340 506586 435576
rect 506822 435340 540918 435576
rect 541154 435340 542850 435576
rect 543086 435340 544782 435576
rect 545018 435340 546714 435576
rect 546950 435340 578266 435576
rect 578502 435340 578586 435576
rect 578822 435340 586302 435576
rect 586538 435340 586622 435576
rect 586858 435340 592650 435576
rect -8726 435308 592650 435340
rect -8726 434656 592650 434688
rect -8726 434420 -1974 434656
rect -1738 434420 -1654 434656
rect -1418 434420 1026 434656
rect 1262 434420 1346 434656
rect 1582 434420 37026 434656
rect 37262 434420 37346 434656
rect 37582 434420 73026 434656
rect 73262 434420 73346 434656
rect 73582 434420 109026 434656
rect 109262 434420 109346 434656
rect 109582 434420 145026 434656
rect 145262 434420 145346 434656
rect 145582 434420 181026 434656
rect 181262 434420 181346 434656
rect 181582 434420 217026 434656
rect 217262 434420 217346 434656
rect 217582 434420 253026 434656
rect 253262 434420 253346 434656
rect 253582 434420 289026 434656
rect 289262 434420 289346 434656
rect 289582 434420 325026 434656
rect 325262 434420 325346 434656
rect 325582 434420 361026 434656
rect 361262 434420 361346 434656
rect 361582 434420 397026 434656
rect 397262 434420 397346 434656
rect 397582 434420 433026 434656
rect 433262 434420 433346 434656
rect 433582 434420 469026 434656
rect 469262 434420 469346 434656
rect 469582 434420 505026 434656
rect 505262 434420 505346 434656
rect 505582 434420 539952 434656
rect 540188 434420 541884 434656
rect 542120 434420 543816 434656
rect 544052 434420 545748 434656
rect 545984 434420 577026 434656
rect 577262 434420 577346 434656
rect 577582 434420 585342 434656
rect 585578 434420 585662 434656
rect 585898 434420 592650 434656
rect -8726 434336 592650 434420
rect -8726 434100 -1974 434336
rect -1738 434100 -1654 434336
rect -1418 434100 1026 434336
rect 1262 434100 1346 434336
rect 1582 434100 37026 434336
rect 37262 434100 37346 434336
rect 37582 434100 73026 434336
rect 73262 434100 73346 434336
rect 73582 434100 109026 434336
rect 109262 434100 109346 434336
rect 109582 434100 145026 434336
rect 145262 434100 145346 434336
rect 145582 434100 181026 434336
rect 181262 434100 181346 434336
rect 181582 434100 217026 434336
rect 217262 434100 217346 434336
rect 217582 434100 253026 434336
rect 253262 434100 253346 434336
rect 253582 434100 289026 434336
rect 289262 434100 289346 434336
rect 289582 434100 325026 434336
rect 325262 434100 325346 434336
rect 325582 434100 361026 434336
rect 361262 434100 361346 434336
rect 361582 434100 397026 434336
rect 397262 434100 397346 434336
rect 397582 434100 433026 434336
rect 433262 434100 433346 434336
rect 433582 434100 469026 434336
rect 469262 434100 469346 434336
rect 469582 434100 505026 434336
rect 505262 434100 505346 434336
rect 505582 434100 539952 434336
rect 540188 434100 541884 434336
rect 542120 434100 543816 434336
rect 544052 434100 545748 434336
rect 545984 434100 577026 434336
rect 577262 434100 577346 434336
rect 577582 434100 585342 434336
rect 585578 434100 585662 434336
rect 585898 434100 592650 434336
rect -8726 434068 592650 434100
rect -8726 407336 592650 407368
rect -8726 407100 -8694 407336
rect -8458 407100 -8374 407336
rect -8138 407100 9706 407336
rect 9942 407100 10026 407336
rect 10262 407100 45706 407336
rect 45942 407100 46026 407336
rect 46262 407100 81706 407336
rect 81942 407100 82026 407336
rect 82262 407100 117706 407336
rect 117942 407100 118026 407336
rect 118262 407100 153706 407336
rect 153942 407100 154026 407336
rect 154262 407100 189706 407336
rect 189942 407100 190026 407336
rect 190262 407100 225706 407336
rect 225942 407100 226026 407336
rect 226262 407100 261706 407336
rect 261942 407100 262026 407336
rect 262262 407100 297706 407336
rect 297942 407100 298026 407336
rect 298262 407100 333706 407336
rect 333942 407100 334026 407336
rect 334262 407100 369706 407336
rect 369942 407100 370026 407336
rect 370262 407100 405706 407336
rect 405942 407100 406026 407336
rect 406262 407100 441706 407336
rect 441942 407100 442026 407336
rect 442262 407100 477706 407336
rect 477942 407100 478026 407336
rect 478262 407100 513706 407336
rect 513942 407100 514026 407336
rect 514262 407100 549706 407336
rect 549942 407100 550026 407336
rect 550262 407100 592062 407336
rect 592298 407100 592382 407336
rect 592618 407100 592650 407336
rect -8726 407016 592650 407100
rect -8726 406780 -8694 407016
rect -8458 406780 -8374 407016
rect -8138 406780 9706 407016
rect 9942 406780 10026 407016
rect 10262 406780 45706 407016
rect 45942 406780 46026 407016
rect 46262 406780 81706 407016
rect 81942 406780 82026 407016
rect 82262 406780 117706 407016
rect 117942 406780 118026 407016
rect 118262 406780 153706 407016
rect 153942 406780 154026 407016
rect 154262 406780 189706 407016
rect 189942 406780 190026 407016
rect 190262 406780 225706 407016
rect 225942 406780 226026 407016
rect 226262 406780 261706 407016
rect 261942 406780 262026 407016
rect 262262 406780 297706 407016
rect 297942 406780 298026 407016
rect 298262 406780 333706 407016
rect 333942 406780 334026 407016
rect 334262 406780 369706 407016
rect 369942 406780 370026 407016
rect 370262 406780 405706 407016
rect 405942 406780 406026 407016
rect 406262 406780 441706 407016
rect 441942 406780 442026 407016
rect 442262 406780 477706 407016
rect 477942 406780 478026 407016
rect 478262 406780 513706 407016
rect 513942 406780 514026 407016
rect 514262 406780 549706 407016
rect 549942 406780 550026 407016
rect 550262 406780 592062 407016
rect 592298 406780 592382 407016
rect 592618 406780 592650 407016
rect -8726 406748 592650 406780
rect -8726 406096 592650 406128
rect -8726 405860 -7734 406096
rect -7498 405860 -7414 406096
rect -7178 405860 8466 406096
rect 8702 405860 8786 406096
rect 9022 405860 44466 406096
rect 44702 405860 44786 406096
rect 45022 405860 80466 406096
rect 80702 405860 80786 406096
rect 81022 405860 116466 406096
rect 116702 405860 116786 406096
rect 117022 405860 152466 406096
rect 152702 405860 152786 406096
rect 153022 405860 188466 406096
rect 188702 405860 188786 406096
rect 189022 405860 224466 406096
rect 224702 405860 224786 406096
rect 225022 405860 260466 406096
rect 260702 405860 260786 406096
rect 261022 405860 296466 406096
rect 296702 405860 296786 406096
rect 297022 405860 332466 406096
rect 332702 405860 332786 406096
rect 333022 405860 368466 406096
rect 368702 405860 368786 406096
rect 369022 405860 404466 406096
rect 404702 405860 404786 406096
rect 405022 405860 440466 406096
rect 440702 405860 440786 406096
rect 441022 405860 476466 406096
rect 476702 405860 476786 406096
rect 477022 405860 512466 406096
rect 512702 405860 512786 406096
rect 513022 405860 548466 406096
rect 548702 405860 548786 406096
rect 549022 405860 591102 406096
rect 591338 405860 591422 406096
rect 591658 405860 592650 406096
rect -8726 405776 592650 405860
rect -8726 405540 -7734 405776
rect -7498 405540 -7414 405776
rect -7178 405540 8466 405776
rect 8702 405540 8786 405776
rect 9022 405540 44466 405776
rect 44702 405540 44786 405776
rect 45022 405540 80466 405776
rect 80702 405540 80786 405776
rect 81022 405540 116466 405776
rect 116702 405540 116786 405776
rect 117022 405540 152466 405776
rect 152702 405540 152786 405776
rect 153022 405540 188466 405776
rect 188702 405540 188786 405776
rect 189022 405540 224466 405776
rect 224702 405540 224786 405776
rect 225022 405540 260466 405776
rect 260702 405540 260786 405776
rect 261022 405540 296466 405776
rect 296702 405540 296786 405776
rect 297022 405540 332466 405776
rect 332702 405540 332786 405776
rect 333022 405540 368466 405776
rect 368702 405540 368786 405776
rect 369022 405540 404466 405776
rect 404702 405540 404786 405776
rect 405022 405540 440466 405776
rect 440702 405540 440786 405776
rect 441022 405540 476466 405776
rect 476702 405540 476786 405776
rect 477022 405540 512466 405776
rect 512702 405540 512786 405776
rect 513022 405540 548466 405776
rect 548702 405540 548786 405776
rect 549022 405540 591102 405776
rect 591338 405540 591422 405776
rect 591658 405540 592650 405776
rect -8726 405508 592650 405540
rect -8726 404856 592650 404888
rect -8726 404620 -6774 404856
rect -6538 404620 -6454 404856
rect -6218 404620 7226 404856
rect 7462 404620 7546 404856
rect 7782 404620 43226 404856
rect 43462 404620 43546 404856
rect 43782 404620 79226 404856
rect 79462 404620 79546 404856
rect 79782 404620 115226 404856
rect 115462 404620 115546 404856
rect 115782 404620 151226 404856
rect 151462 404620 151546 404856
rect 151782 404620 187226 404856
rect 187462 404620 187546 404856
rect 187782 404620 223226 404856
rect 223462 404620 223546 404856
rect 223782 404620 259226 404856
rect 259462 404620 259546 404856
rect 259782 404620 295226 404856
rect 295462 404620 295546 404856
rect 295782 404620 331226 404856
rect 331462 404620 331546 404856
rect 331782 404620 367226 404856
rect 367462 404620 367546 404856
rect 367782 404620 403226 404856
rect 403462 404620 403546 404856
rect 403782 404620 439226 404856
rect 439462 404620 439546 404856
rect 439782 404620 475226 404856
rect 475462 404620 475546 404856
rect 475782 404620 511226 404856
rect 511462 404620 511546 404856
rect 511782 404620 547226 404856
rect 547462 404620 547546 404856
rect 547782 404620 590142 404856
rect 590378 404620 590462 404856
rect 590698 404620 592650 404856
rect -8726 404536 592650 404620
rect -8726 404300 -6774 404536
rect -6538 404300 -6454 404536
rect -6218 404300 7226 404536
rect 7462 404300 7546 404536
rect 7782 404300 43226 404536
rect 43462 404300 43546 404536
rect 43782 404300 79226 404536
rect 79462 404300 79546 404536
rect 79782 404300 115226 404536
rect 115462 404300 115546 404536
rect 115782 404300 151226 404536
rect 151462 404300 151546 404536
rect 151782 404300 187226 404536
rect 187462 404300 187546 404536
rect 187782 404300 223226 404536
rect 223462 404300 223546 404536
rect 223782 404300 259226 404536
rect 259462 404300 259546 404536
rect 259782 404300 295226 404536
rect 295462 404300 295546 404536
rect 295782 404300 331226 404536
rect 331462 404300 331546 404536
rect 331782 404300 367226 404536
rect 367462 404300 367546 404536
rect 367782 404300 403226 404536
rect 403462 404300 403546 404536
rect 403782 404300 439226 404536
rect 439462 404300 439546 404536
rect 439782 404300 475226 404536
rect 475462 404300 475546 404536
rect 475782 404300 511226 404536
rect 511462 404300 511546 404536
rect 511782 404300 547226 404536
rect 547462 404300 547546 404536
rect 547782 404300 590142 404536
rect 590378 404300 590462 404536
rect 590698 404300 592650 404536
rect -8726 404268 592650 404300
rect -8726 403616 592650 403648
rect -8726 403380 -5814 403616
rect -5578 403380 -5494 403616
rect -5258 403380 5986 403616
rect 6222 403380 6306 403616
rect 6542 403380 41986 403616
rect 42222 403380 42306 403616
rect 42542 403380 77986 403616
rect 78222 403380 78306 403616
rect 78542 403380 113986 403616
rect 114222 403380 114306 403616
rect 114542 403380 149986 403616
rect 150222 403380 150306 403616
rect 150542 403380 185986 403616
rect 186222 403380 186306 403616
rect 186542 403380 221986 403616
rect 222222 403380 222306 403616
rect 222542 403380 257986 403616
rect 258222 403380 258306 403616
rect 258542 403380 293986 403616
rect 294222 403380 294306 403616
rect 294542 403380 329986 403616
rect 330222 403380 330306 403616
rect 330542 403380 365986 403616
rect 366222 403380 366306 403616
rect 366542 403380 401986 403616
rect 402222 403380 402306 403616
rect 402542 403380 437986 403616
rect 438222 403380 438306 403616
rect 438542 403380 473986 403616
rect 474222 403380 474306 403616
rect 474542 403380 509986 403616
rect 510222 403380 510306 403616
rect 510542 403380 581986 403616
rect 582222 403380 582306 403616
rect 582542 403380 589182 403616
rect 589418 403380 589502 403616
rect 589738 403380 592650 403616
rect -8726 403296 592650 403380
rect -8726 403060 -5814 403296
rect -5578 403060 -5494 403296
rect -5258 403060 5986 403296
rect 6222 403060 6306 403296
rect 6542 403060 41986 403296
rect 42222 403060 42306 403296
rect 42542 403060 77986 403296
rect 78222 403060 78306 403296
rect 78542 403060 113986 403296
rect 114222 403060 114306 403296
rect 114542 403060 149986 403296
rect 150222 403060 150306 403296
rect 150542 403060 185986 403296
rect 186222 403060 186306 403296
rect 186542 403060 221986 403296
rect 222222 403060 222306 403296
rect 222542 403060 257986 403296
rect 258222 403060 258306 403296
rect 258542 403060 293986 403296
rect 294222 403060 294306 403296
rect 294542 403060 329986 403296
rect 330222 403060 330306 403296
rect 330542 403060 365986 403296
rect 366222 403060 366306 403296
rect 366542 403060 401986 403296
rect 402222 403060 402306 403296
rect 402542 403060 437986 403296
rect 438222 403060 438306 403296
rect 438542 403060 473986 403296
rect 474222 403060 474306 403296
rect 474542 403060 509986 403296
rect 510222 403060 510306 403296
rect 510542 403060 581986 403296
rect 582222 403060 582306 403296
rect 582542 403060 589182 403296
rect 589418 403060 589502 403296
rect 589738 403060 592650 403296
rect -8726 403028 592650 403060
rect -8726 402376 592650 402408
rect -8726 402140 -4854 402376
rect -4618 402140 -4534 402376
rect -4298 402140 4746 402376
rect 4982 402140 5066 402376
rect 5302 402140 40746 402376
rect 40982 402140 41066 402376
rect 41302 402140 76746 402376
rect 76982 402140 77066 402376
rect 77302 402140 112746 402376
rect 112982 402140 113066 402376
rect 113302 402140 148746 402376
rect 148982 402140 149066 402376
rect 149302 402140 184746 402376
rect 184982 402140 185066 402376
rect 185302 402140 220746 402376
rect 220982 402140 221066 402376
rect 221302 402140 256746 402376
rect 256982 402140 257066 402376
rect 257302 402140 292746 402376
rect 292982 402140 293066 402376
rect 293302 402140 328746 402376
rect 328982 402140 329066 402376
rect 329302 402140 364746 402376
rect 364982 402140 365066 402376
rect 365302 402140 400746 402376
rect 400982 402140 401066 402376
rect 401302 402140 436746 402376
rect 436982 402140 437066 402376
rect 437302 402140 472746 402376
rect 472982 402140 473066 402376
rect 473302 402140 508746 402376
rect 508982 402140 509066 402376
rect 509302 402140 580746 402376
rect 580982 402140 581066 402376
rect 581302 402140 588222 402376
rect 588458 402140 588542 402376
rect 588778 402140 592650 402376
rect -8726 402056 592650 402140
rect -8726 401820 -4854 402056
rect -4618 401820 -4534 402056
rect -4298 401820 4746 402056
rect 4982 401820 5066 402056
rect 5302 401820 40746 402056
rect 40982 401820 41066 402056
rect 41302 401820 76746 402056
rect 76982 401820 77066 402056
rect 77302 401820 112746 402056
rect 112982 401820 113066 402056
rect 113302 401820 148746 402056
rect 148982 401820 149066 402056
rect 149302 401820 184746 402056
rect 184982 401820 185066 402056
rect 185302 401820 220746 402056
rect 220982 401820 221066 402056
rect 221302 401820 256746 402056
rect 256982 401820 257066 402056
rect 257302 401820 292746 402056
rect 292982 401820 293066 402056
rect 293302 401820 328746 402056
rect 328982 401820 329066 402056
rect 329302 401820 364746 402056
rect 364982 401820 365066 402056
rect 365302 401820 400746 402056
rect 400982 401820 401066 402056
rect 401302 401820 436746 402056
rect 436982 401820 437066 402056
rect 437302 401820 472746 402056
rect 472982 401820 473066 402056
rect 473302 401820 508746 402056
rect 508982 401820 509066 402056
rect 509302 401820 580746 402056
rect 580982 401820 581066 402056
rect 581302 401820 588222 402056
rect 588458 401820 588542 402056
rect 588778 401820 592650 402056
rect -8726 401788 592650 401820
rect -8726 401136 592650 401168
rect -8726 400900 -3894 401136
rect -3658 400900 -3574 401136
rect -3338 400900 3506 401136
rect 3742 400900 3826 401136
rect 4062 400900 39506 401136
rect 39742 400900 39826 401136
rect 40062 400900 75506 401136
rect 75742 400900 75826 401136
rect 76062 400900 111506 401136
rect 111742 400900 111826 401136
rect 112062 400900 147506 401136
rect 147742 400900 147826 401136
rect 148062 400900 183506 401136
rect 183742 400900 183826 401136
rect 184062 400900 219506 401136
rect 219742 400900 219826 401136
rect 220062 400900 255506 401136
rect 255742 400900 255826 401136
rect 256062 400900 291506 401136
rect 291742 400900 291826 401136
rect 292062 400900 327506 401136
rect 327742 400900 327826 401136
rect 328062 400900 363506 401136
rect 363742 400900 363826 401136
rect 364062 400900 399506 401136
rect 399742 400900 399826 401136
rect 400062 400900 435506 401136
rect 435742 400900 435826 401136
rect 436062 400900 471506 401136
rect 471742 400900 471826 401136
rect 472062 400900 507506 401136
rect 507742 400900 507826 401136
rect 508062 400900 579506 401136
rect 579742 400900 579826 401136
rect 580062 400900 587262 401136
rect 587498 400900 587582 401136
rect 587818 400900 592650 401136
rect -8726 400816 592650 400900
rect -8726 400580 -3894 400816
rect -3658 400580 -3574 400816
rect -3338 400580 3506 400816
rect 3742 400580 3826 400816
rect 4062 400580 39506 400816
rect 39742 400580 39826 400816
rect 40062 400580 75506 400816
rect 75742 400580 75826 400816
rect 76062 400580 111506 400816
rect 111742 400580 111826 400816
rect 112062 400580 147506 400816
rect 147742 400580 147826 400816
rect 148062 400580 183506 400816
rect 183742 400580 183826 400816
rect 184062 400580 219506 400816
rect 219742 400580 219826 400816
rect 220062 400580 255506 400816
rect 255742 400580 255826 400816
rect 256062 400580 291506 400816
rect 291742 400580 291826 400816
rect 292062 400580 327506 400816
rect 327742 400580 327826 400816
rect 328062 400580 363506 400816
rect 363742 400580 363826 400816
rect 364062 400580 399506 400816
rect 399742 400580 399826 400816
rect 400062 400580 435506 400816
rect 435742 400580 435826 400816
rect 436062 400580 471506 400816
rect 471742 400580 471826 400816
rect 472062 400580 507506 400816
rect 507742 400580 507826 400816
rect 508062 400580 579506 400816
rect 579742 400580 579826 400816
rect 580062 400580 587262 400816
rect 587498 400580 587582 400816
rect 587818 400580 592650 400816
rect -8726 400548 592650 400580
rect -8726 399896 592650 399928
rect -8726 399660 -2934 399896
rect -2698 399660 -2614 399896
rect -2378 399660 2266 399896
rect 2502 399660 2586 399896
rect 2822 399660 38266 399896
rect 38502 399660 38586 399896
rect 38822 399660 74266 399896
rect 74502 399660 74586 399896
rect 74822 399660 110266 399896
rect 110502 399660 110586 399896
rect 110822 399660 146266 399896
rect 146502 399660 146586 399896
rect 146822 399660 182266 399896
rect 182502 399660 182586 399896
rect 182822 399660 218266 399896
rect 218502 399660 218586 399896
rect 218822 399660 254266 399896
rect 254502 399660 254586 399896
rect 254822 399660 290266 399896
rect 290502 399660 290586 399896
rect 290822 399660 326266 399896
rect 326502 399660 326586 399896
rect 326822 399660 362266 399896
rect 362502 399660 362586 399896
rect 362822 399660 398266 399896
rect 398502 399660 398586 399896
rect 398822 399660 434266 399896
rect 434502 399660 434586 399896
rect 434822 399660 470266 399896
rect 470502 399660 470586 399896
rect 470822 399660 506266 399896
rect 506502 399660 506586 399896
rect 506822 399660 540918 399896
rect 541154 399660 542850 399896
rect 543086 399660 544782 399896
rect 545018 399660 546714 399896
rect 546950 399660 578266 399896
rect 578502 399660 578586 399896
rect 578822 399660 586302 399896
rect 586538 399660 586622 399896
rect 586858 399660 592650 399896
rect -8726 399576 592650 399660
rect -8726 399340 -2934 399576
rect -2698 399340 -2614 399576
rect -2378 399340 2266 399576
rect 2502 399340 2586 399576
rect 2822 399340 38266 399576
rect 38502 399340 38586 399576
rect 38822 399340 74266 399576
rect 74502 399340 74586 399576
rect 74822 399340 110266 399576
rect 110502 399340 110586 399576
rect 110822 399340 146266 399576
rect 146502 399340 146586 399576
rect 146822 399340 182266 399576
rect 182502 399340 182586 399576
rect 182822 399340 218266 399576
rect 218502 399340 218586 399576
rect 218822 399340 254266 399576
rect 254502 399340 254586 399576
rect 254822 399340 290266 399576
rect 290502 399340 290586 399576
rect 290822 399340 326266 399576
rect 326502 399340 326586 399576
rect 326822 399340 362266 399576
rect 362502 399340 362586 399576
rect 362822 399340 398266 399576
rect 398502 399340 398586 399576
rect 398822 399340 434266 399576
rect 434502 399340 434586 399576
rect 434822 399340 470266 399576
rect 470502 399340 470586 399576
rect 470822 399340 506266 399576
rect 506502 399340 506586 399576
rect 506822 399340 540918 399576
rect 541154 399340 542850 399576
rect 543086 399340 544782 399576
rect 545018 399340 546714 399576
rect 546950 399340 578266 399576
rect 578502 399340 578586 399576
rect 578822 399340 586302 399576
rect 586538 399340 586622 399576
rect 586858 399340 592650 399576
rect -8726 399308 592650 399340
rect -8726 398656 592650 398688
rect -8726 398420 -1974 398656
rect -1738 398420 -1654 398656
rect -1418 398420 1026 398656
rect 1262 398420 1346 398656
rect 1582 398420 37026 398656
rect 37262 398420 37346 398656
rect 37582 398420 73026 398656
rect 73262 398420 73346 398656
rect 73582 398420 109026 398656
rect 109262 398420 109346 398656
rect 109582 398420 145026 398656
rect 145262 398420 145346 398656
rect 145582 398420 181026 398656
rect 181262 398420 181346 398656
rect 181582 398420 217026 398656
rect 217262 398420 217346 398656
rect 217582 398420 253026 398656
rect 253262 398420 253346 398656
rect 253582 398420 289026 398656
rect 289262 398420 289346 398656
rect 289582 398420 325026 398656
rect 325262 398420 325346 398656
rect 325582 398420 361026 398656
rect 361262 398420 361346 398656
rect 361582 398420 397026 398656
rect 397262 398420 397346 398656
rect 397582 398420 433026 398656
rect 433262 398420 433346 398656
rect 433582 398420 469026 398656
rect 469262 398420 469346 398656
rect 469582 398420 505026 398656
rect 505262 398420 505346 398656
rect 505582 398420 539952 398656
rect 540188 398420 541884 398656
rect 542120 398420 543816 398656
rect 544052 398420 545748 398656
rect 545984 398420 577026 398656
rect 577262 398420 577346 398656
rect 577582 398420 585342 398656
rect 585578 398420 585662 398656
rect 585898 398420 592650 398656
rect -8726 398336 592650 398420
rect -8726 398100 -1974 398336
rect -1738 398100 -1654 398336
rect -1418 398100 1026 398336
rect 1262 398100 1346 398336
rect 1582 398100 37026 398336
rect 37262 398100 37346 398336
rect 37582 398100 73026 398336
rect 73262 398100 73346 398336
rect 73582 398100 109026 398336
rect 109262 398100 109346 398336
rect 109582 398100 145026 398336
rect 145262 398100 145346 398336
rect 145582 398100 181026 398336
rect 181262 398100 181346 398336
rect 181582 398100 217026 398336
rect 217262 398100 217346 398336
rect 217582 398100 253026 398336
rect 253262 398100 253346 398336
rect 253582 398100 289026 398336
rect 289262 398100 289346 398336
rect 289582 398100 325026 398336
rect 325262 398100 325346 398336
rect 325582 398100 361026 398336
rect 361262 398100 361346 398336
rect 361582 398100 397026 398336
rect 397262 398100 397346 398336
rect 397582 398100 433026 398336
rect 433262 398100 433346 398336
rect 433582 398100 469026 398336
rect 469262 398100 469346 398336
rect 469582 398100 505026 398336
rect 505262 398100 505346 398336
rect 505582 398100 539952 398336
rect 540188 398100 541884 398336
rect 542120 398100 543816 398336
rect 544052 398100 545748 398336
rect 545984 398100 577026 398336
rect 577262 398100 577346 398336
rect 577582 398100 585342 398336
rect 585578 398100 585662 398336
rect 585898 398100 592650 398336
rect -8726 398068 592650 398100
rect -8726 371336 592650 371368
rect -8726 371100 -8694 371336
rect -8458 371100 -8374 371336
rect -8138 371100 9706 371336
rect 9942 371100 10026 371336
rect 10262 371100 45706 371336
rect 45942 371100 46026 371336
rect 46262 371100 81706 371336
rect 81942 371100 82026 371336
rect 82262 371100 117706 371336
rect 117942 371100 118026 371336
rect 118262 371100 153706 371336
rect 153942 371100 154026 371336
rect 154262 371100 189706 371336
rect 189942 371100 190026 371336
rect 190262 371100 225706 371336
rect 225942 371100 226026 371336
rect 226262 371100 261706 371336
rect 261942 371100 262026 371336
rect 262262 371100 297706 371336
rect 297942 371100 298026 371336
rect 298262 371100 333706 371336
rect 333942 371100 334026 371336
rect 334262 371100 369706 371336
rect 369942 371100 370026 371336
rect 370262 371100 405706 371336
rect 405942 371100 406026 371336
rect 406262 371100 441706 371336
rect 441942 371100 442026 371336
rect 442262 371100 477706 371336
rect 477942 371100 478026 371336
rect 478262 371100 513706 371336
rect 513942 371100 514026 371336
rect 514262 371100 549706 371336
rect 549942 371100 550026 371336
rect 550262 371100 592062 371336
rect 592298 371100 592382 371336
rect 592618 371100 592650 371336
rect -8726 371016 592650 371100
rect -8726 370780 -8694 371016
rect -8458 370780 -8374 371016
rect -8138 370780 9706 371016
rect 9942 370780 10026 371016
rect 10262 370780 45706 371016
rect 45942 370780 46026 371016
rect 46262 370780 81706 371016
rect 81942 370780 82026 371016
rect 82262 370780 117706 371016
rect 117942 370780 118026 371016
rect 118262 370780 153706 371016
rect 153942 370780 154026 371016
rect 154262 370780 189706 371016
rect 189942 370780 190026 371016
rect 190262 370780 225706 371016
rect 225942 370780 226026 371016
rect 226262 370780 261706 371016
rect 261942 370780 262026 371016
rect 262262 370780 297706 371016
rect 297942 370780 298026 371016
rect 298262 370780 333706 371016
rect 333942 370780 334026 371016
rect 334262 370780 369706 371016
rect 369942 370780 370026 371016
rect 370262 370780 405706 371016
rect 405942 370780 406026 371016
rect 406262 370780 441706 371016
rect 441942 370780 442026 371016
rect 442262 370780 477706 371016
rect 477942 370780 478026 371016
rect 478262 370780 513706 371016
rect 513942 370780 514026 371016
rect 514262 370780 549706 371016
rect 549942 370780 550026 371016
rect 550262 370780 592062 371016
rect 592298 370780 592382 371016
rect 592618 370780 592650 371016
rect -8726 370748 592650 370780
rect -8726 370096 592650 370128
rect -8726 369860 -7734 370096
rect -7498 369860 -7414 370096
rect -7178 369860 8466 370096
rect 8702 369860 8786 370096
rect 9022 369860 44466 370096
rect 44702 369860 44786 370096
rect 45022 369860 80466 370096
rect 80702 369860 80786 370096
rect 81022 369860 116466 370096
rect 116702 369860 116786 370096
rect 117022 369860 152466 370096
rect 152702 369860 152786 370096
rect 153022 369860 188466 370096
rect 188702 369860 188786 370096
rect 189022 369860 224466 370096
rect 224702 369860 224786 370096
rect 225022 369860 260466 370096
rect 260702 369860 260786 370096
rect 261022 369860 296466 370096
rect 296702 369860 296786 370096
rect 297022 369860 332466 370096
rect 332702 369860 332786 370096
rect 333022 369860 368466 370096
rect 368702 369860 368786 370096
rect 369022 369860 404466 370096
rect 404702 369860 404786 370096
rect 405022 369860 440466 370096
rect 440702 369860 440786 370096
rect 441022 369860 476466 370096
rect 476702 369860 476786 370096
rect 477022 369860 512466 370096
rect 512702 369860 512786 370096
rect 513022 369860 548466 370096
rect 548702 369860 548786 370096
rect 549022 369860 591102 370096
rect 591338 369860 591422 370096
rect 591658 369860 592650 370096
rect -8726 369776 592650 369860
rect -8726 369540 -7734 369776
rect -7498 369540 -7414 369776
rect -7178 369540 8466 369776
rect 8702 369540 8786 369776
rect 9022 369540 44466 369776
rect 44702 369540 44786 369776
rect 45022 369540 80466 369776
rect 80702 369540 80786 369776
rect 81022 369540 116466 369776
rect 116702 369540 116786 369776
rect 117022 369540 152466 369776
rect 152702 369540 152786 369776
rect 153022 369540 188466 369776
rect 188702 369540 188786 369776
rect 189022 369540 224466 369776
rect 224702 369540 224786 369776
rect 225022 369540 260466 369776
rect 260702 369540 260786 369776
rect 261022 369540 296466 369776
rect 296702 369540 296786 369776
rect 297022 369540 332466 369776
rect 332702 369540 332786 369776
rect 333022 369540 368466 369776
rect 368702 369540 368786 369776
rect 369022 369540 404466 369776
rect 404702 369540 404786 369776
rect 405022 369540 440466 369776
rect 440702 369540 440786 369776
rect 441022 369540 476466 369776
rect 476702 369540 476786 369776
rect 477022 369540 512466 369776
rect 512702 369540 512786 369776
rect 513022 369540 548466 369776
rect 548702 369540 548786 369776
rect 549022 369540 591102 369776
rect 591338 369540 591422 369776
rect 591658 369540 592650 369776
rect -8726 369508 592650 369540
rect -8726 368856 592650 368888
rect -8726 368620 -6774 368856
rect -6538 368620 -6454 368856
rect -6218 368620 7226 368856
rect 7462 368620 7546 368856
rect 7782 368620 43226 368856
rect 43462 368620 43546 368856
rect 43782 368620 79226 368856
rect 79462 368620 79546 368856
rect 79782 368620 115226 368856
rect 115462 368620 115546 368856
rect 115782 368620 151226 368856
rect 151462 368620 151546 368856
rect 151782 368620 187226 368856
rect 187462 368620 187546 368856
rect 187782 368620 223226 368856
rect 223462 368620 223546 368856
rect 223782 368620 259226 368856
rect 259462 368620 259546 368856
rect 259782 368620 295226 368856
rect 295462 368620 295546 368856
rect 295782 368620 331226 368856
rect 331462 368620 331546 368856
rect 331782 368620 367226 368856
rect 367462 368620 367546 368856
rect 367782 368620 403226 368856
rect 403462 368620 403546 368856
rect 403782 368620 439226 368856
rect 439462 368620 439546 368856
rect 439782 368620 475226 368856
rect 475462 368620 475546 368856
rect 475782 368620 511226 368856
rect 511462 368620 511546 368856
rect 511782 368620 547226 368856
rect 547462 368620 547546 368856
rect 547782 368620 590142 368856
rect 590378 368620 590462 368856
rect 590698 368620 592650 368856
rect -8726 368536 592650 368620
rect -8726 368300 -6774 368536
rect -6538 368300 -6454 368536
rect -6218 368300 7226 368536
rect 7462 368300 7546 368536
rect 7782 368300 43226 368536
rect 43462 368300 43546 368536
rect 43782 368300 79226 368536
rect 79462 368300 79546 368536
rect 79782 368300 115226 368536
rect 115462 368300 115546 368536
rect 115782 368300 151226 368536
rect 151462 368300 151546 368536
rect 151782 368300 187226 368536
rect 187462 368300 187546 368536
rect 187782 368300 223226 368536
rect 223462 368300 223546 368536
rect 223782 368300 259226 368536
rect 259462 368300 259546 368536
rect 259782 368300 295226 368536
rect 295462 368300 295546 368536
rect 295782 368300 331226 368536
rect 331462 368300 331546 368536
rect 331782 368300 367226 368536
rect 367462 368300 367546 368536
rect 367782 368300 403226 368536
rect 403462 368300 403546 368536
rect 403782 368300 439226 368536
rect 439462 368300 439546 368536
rect 439782 368300 475226 368536
rect 475462 368300 475546 368536
rect 475782 368300 511226 368536
rect 511462 368300 511546 368536
rect 511782 368300 547226 368536
rect 547462 368300 547546 368536
rect 547782 368300 590142 368536
rect 590378 368300 590462 368536
rect 590698 368300 592650 368536
rect -8726 368268 592650 368300
rect -8726 367616 592650 367648
rect -8726 367380 -5814 367616
rect -5578 367380 -5494 367616
rect -5258 367380 5986 367616
rect 6222 367380 6306 367616
rect 6542 367380 41986 367616
rect 42222 367380 42306 367616
rect 42542 367380 77986 367616
rect 78222 367380 78306 367616
rect 78542 367380 113986 367616
rect 114222 367380 114306 367616
rect 114542 367380 149986 367616
rect 150222 367380 150306 367616
rect 150542 367380 185986 367616
rect 186222 367380 186306 367616
rect 186542 367380 221986 367616
rect 222222 367380 222306 367616
rect 222542 367380 257986 367616
rect 258222 367380 258306 367616
rect 258542 367380 293986 367616
rect 294222 367380 294306 367616
rect 294542 367380 329986 367616
rect 330222 367380 330306 367616
rect 330542 367380 365986 367616
rect 366222 367380 366306 367616
rect 366542 367380 401986 367616
rect 402222 367380 402306 367616
rect 402542 367380 437986 367616
rect 438222 367380 438306 367616
rect 438542 367380 473986 367616
rect 474222 367380 474306 367616
rect 474542 367380 509986 367616
rect 510222 367380 510306 367616
rect 510542 367380 581986 367616
rect 582222 367380 582306 367616
rect 582542 367380 589182 367616
rect 589418 367380 589502 367616
rect 589738 367380 592650 367616
rect -8726 367296 592650 367380
rect -8726 367060 -5814 367296
rect -5578 367060 -5494 367296
rect -5258 367060 5986 367296
rect 6222 367060 6306 367296
rect 6542 367060 41986 367296
rect 42222 367060 42306 367296
rect 42542 367060 77986 367296
rect 78222 367060 78306 367296
rect 78542 367060 113986 367296
rect 114222 367060 114306 367296
rect 114542 367060 149986 367296
rect 150222 367060 150306 367296
rect 150542 367060 185986 367296
rect 186222 367060 186306 367296
rect 186542 367060 221986 367296
rect 222222 367060 222306 367296
rect 222542 367060 257986 367296
rect 258222 367060 258306 367296
rect 258542 367060 293986 367296
rect 294222 367060 294306 367296
rect 294542 367060 329986 367296
rect 330222 367060 330306 367296
rect 330542 367060 365986 367296
rect 366222 367060 366306 367296
rect 366542 367060 401986 367296
rect 402222 367060 402306 367296
rect 402542 367060 437986 367296
rect 438222 367060 438306 367296
rect 438542 367060 473986 367296
rect 474222 367060 474306 367296
rect 474542 367060 509986 367296
rect 510222 367060 510306 367296
rect 510542 367060 581986 367296
rect 582222 367060 582306 367296
rect 582542 367060 589182 367296
rect 589418 367060 589502 367296
rect 589738 367060 592650 367296
rect -8726 367028 592650 367060
rect -8726 366376 592650 366408
rect -8726 366140 -4854 366376
rect -4618 366140 -4534 366376
rect -4298 366140 4746 366376
rect 4982 366140 5066 366376
rect 5302 366140 40746 366376
rect 40982 366140 41066 366376
rect 41302 366140 76746 366376
rect 76982 366140 77066 366376
rect 77302 366140 112746 366376
rect 112982 366140 113066 366376
rect 113302 366140 148746 366376
rect 148982 366140 149066 366376
rect 149302 366140 184746 366376
rect 184982 366140 185066 366376
rect 185302 366140 220746 366376
rect 220982 366140 221066 366376
rect 221302 366140 256746 366376
rect 256982 366140 257066 366376
rect 257302 366140 292746 366376
rect 292982 366140 293066 366376
rect 293302 366140 328746 366376
rect 328982 366140 329066 366376
rect 329302 366140 364746 366376
rect 364982 366140 365066 366376
rect 365302 366140 400746 366376
rect 400982 366140 401066 366376
rect 401302 366140 436746 366376
rect 436982 366140 437066 366376
rect 437302 366140 472746 366376
rect 472982 366140 473066 366376
rect 473302 366140 508746 366376
rect 508982 366140 509066 366376
rect 509302 366140 580746 366376
rect 580982 366140 581066 366376
rect 581302 366140 588222 366376
rect 588458 366140 588542 366376
rect 588778 366140 592650 366376
rect -8726 366056 592650 366140
rect -8726 365820 -4854 366056
rect -4618 365820 -4534 366056
rect -4298 365820 4746 366056
rect 4982 365820 5066 366056
rect 5302 365820 40746 366056
rect 40982 365820 41066 366056
rect 41302 365820 76746 366056
rect 76982 365820 77066 366056
rect 77302 365820 112746 366056
rect 112982 365820 113066 366056
rect 113302 365820 148746 366056
rect 148982 365820 149066 366056
rect 149302 365820 184746 366056
rect 184982 365820 185066 366056
rect 185302 365820 220746 366056
rect 220982 365820 221066 366056
rect 221302 365820 256746 366056
rect 256982 365820 257066 366056
rect 257302 365820 292746 366056
rect 292982 365820 293066 366056
rect 293302 365820 328746 366056
rect 328982 365820 329066 366056
rect 329302 365820 364746 366056
rect 364982 365820 365066 366056
rect 365302 365820 400746 366056
rect 400982 365820 401066 366056
rect 401302 365820 436746 366056
rect 436982 365820 437066 366056
rect 437302 365820 472746 366056
rect 472982 365820 473066 366056
rect 473302 365820 508746 366056
rect 508982 365820 509066 366056
rect 509302 365820 580746 366056
rect 580982 365820 581066 366056
rect 581302 365820 588222 366056
rect 588458 365820 588542 366056
rect 588778 365820 592650 366056
rect -8726 365788 592650 365820
rect -8726 365136 592650 365168
rect -8726 364900 -3894 365136
rect -3658 364900 -3574 365136
rect -3338 364900 3506 365136
rect 3742 364900 3826 365136
rect 4062 364900 39506 365136
rect 39742 364900 39826 365136
rect 40062 364900 75506 365136
rect 75742 364900 75826 365136
rect 76062 364900 111506 365136
rect 111742 364900 111826 365136
rect 112062 364900 147506 365136
rect 147742 364900 147826 365136
rect 148062 364900 183506 365136
rect 183742 364900 183826 365136
rect 184062 364900 219506 365136
rect 219742 364900 219826 365136
rect 220062 364900 255506 365136
rect 255742 364900 255826 365136
rect 256062 364900 291506 365136
rect 291742 364900 291826 365136
rect 292062 364900 327506 365136
rect 327742 364900 327826 365136
rect 328062 364900 363506 365136
rect 363742 364900 363826 365136
rect 364062 364900 399506 365136
rect 399742 364900 399826 365136
rect 400062 364900 435506 365136
rect 435742 364900 435826 365136
rect 436062 364900 471506 365136
rect 471742 364900 471826 365136
rect 472062 364900 507506 365136
rect 507742 364900 507826 365136
rect 508062 364900 579506 365136
rect 579742 364900 579826 365136
rect 580062 364900 587262 365136
rect 587498 364900 587582 365136
rect 587818 364900 592650 365136
rect -8726 364816 592650 364900
rect -8726 364580 -3894 364816
rect -3658 364580 -3574 364816
rect -3338 364580 3506 364816
rect 3742 364580 3826 364816
rect 4062 364580 39506 364816
rect 39742 364580 39826 364816
rect 40062 364580 75506 364816
rect 75742 364580 75826 364816
rect 76062 364580 111506 364816
rect 111742 364580 111826 364816
rect 112062 364580 147506 364816
rect 147742 364580 147826 364816
rect 148062 364580 183506 364816
rect 183742 364580 183826 364816
rect 184062 364580 219506 364816
rect 219742 364580 219826 364816
rect 220062 364580 255506 364816
rect 255742 364580 255826 364816
rect 256062 364580 291506 364816
rect 291742 364580 291826 364816
rect 292062 364580 327506 364816
rect 327742 364580 327826 364816
rect 328062 364580 363506 364816
rect 363742 364580 363826 364816
rect 364062 364580 399506 364816
rect 399742 364580 399826 364816
rect 400062 364580 435506 364816
rect 435742 364580 435826 364816
rect 436062 364580 471506 364816
rect 471742 364580 471826 364816
rect 472062 364580 507506 364816
rect 507742 364580 507826 364816
rect 508062 364580 579506 364816
rect 579742 364580 579826 364816
rect 580062 364580 587262 364816
rect 587498 364580 587582 364816
rect 587818 364580 592650 364816
rect -8726 364548 592650 364580
rect -8726 363896 592650 363928
rect -8726 363660 -2934 363896
rect -2698 363660 -2614 363896
rect -2378 363660 2266 363896
rect 2502 363660 2586 363896
rect 2822 363660 38266 363896
rect 38502 363660 38586 363896
rect 38822 363660 74266 363896
rect 74502 363660 74586 363896
rect 74822 363660 110266 363896
rect 110502 363660 110586 363896
rect 110822 363660 146266 363896
rect 146502 363660 146586 363896
rect 146822 363660 182266 363896
rect 182502 363660 182586 363896
rect 182822 363660 218266 363896
rect 218502 363660 218586 363896
rect 218822 363660 254266 363896
rect 254502 363660 254586 363896
rect 254822 363660 290266 363896
rect 290502 363660 290586 363896
rect 290822 363660 326266 363896
rect 326502 363660 326586 363896
rect 326822 363660 362266 363896
rect 362502 363660 362586 363896
rect 362822 363660 398266 363896
rect 398502 363660 398586 363896
rect 398822 363660 434266 363896
rect 434502 363660 434586 363896
rect 434822 363660 470266 363896
rect 470502 363660 470586 363896
rect 470822 363660 506266 363896
rect 506502 363660 506586 363896
rect 506822 363660 540918 363896
rect 541154 363660 542850 363896
rect 543086 363660 544782 363896
rect 545018 363660 546714 363896
rect 546950 363660 578266 363896
rect 578502 363660 578586 363896
rect 578822 363660 586302 363896
rect 586538 363660 586622 363896
rect 586858 363660 592650 363896
rect -8726 363576 592650 363660
rect -8726 363340 -2934 363576
rect -2698 363340 -2614 363576
rect -2378 363340 2266 363576
rect 2502 363340 2586 363576
rect 2822 363340 38266 363576
rect 38502 363340 38586 363576
rect 38822 363340 74266 363576
rect 74502 363340 74586 363576
rect 74822 363340 110266 363576
rect 110502 363340 110586 363576
rect 110822 363340 146266 363576
rect 146502 363340 146586 363576
rect 146822 363340 182266 363576
rect 182502 363340 182586 363576
rect 182822 363340 218266 363576
rect 218502 363340 218586 363576
rect 218822 363340 254266 363576
rect 254502 363340 254586 363576
rect 254822 363340 290266 363576
rect 290502 363340 290586 363576
rect 290822 363340 326266 363576
rect 326502 363340 326586 363576
rect 326822 363340 362266 363576
rect 362502 363340 362586 363576
rect 362822 363340 398266 363576
rect 398502 363340 398586 363576
rect 398822 363340 434266 363576
rect 434502 363340 434586 363576
rect 434822 363340 470266 363576
rect 470502 363340 470586 363576
rect 470822 363340 506266 363576
rect 506502 363340 506586 363576
rect 506822 363340 540918 363576
rect 541154 363340 542850 363576
rect 543086 363340 544782 363576
rect 545018 363340 546714 363576
rect 546950 363340 578266 363576
rect 578502 363340 578586 363576
rect 578822 363340 586302 363576
rect 586538 363340 586622 363576
rect 586858 363340 592650 363576
rect -8726 363308 592650 363340
rect -8726 362656 592650 362688
rect -8726 362420 -1974 362656
rect -1738 362420 -1654 362656
rect -1418 362420 1026 362656
rect 1262 362420 1346 362656
rect 1582 362420 37026 362656
rect 37262 362420 37346 362656
rect 37582 362420 73026 362656
rect 73262 362420 73346 362656
rect 73582 362420 109026 362656
rect 109262 362420 109346 362656
rect 109582 362420 145026 362656
rect 145262 362420 145346 362656
rect 145582 362420 181026 362656
rect 181262 362420 181346 362656
rect 181582 362420 217026 362656
rect 217262 362420 217346 362656
rect 217582 362420 253026 362656
rect 253262 362420 253346 362656
rect 253582 362420 289026 362656
rect 289262 362420 289346 362656
rect 289582 362420 325026 362656
rect 325262 362420 325346 362656
rect 325582 362420 361026 362656
rect 361262 362420 361346 362656
rect 361582 362420 397026 362656
rect 397262 362420 397346 362656
rect 397582 362420 433026 362656
rect 433262 362420 433346 362656
rect 433582 362420 469026 362656
rect 469262 362420 469346 362656
rect 469582 362420 505026 362656
rect 505262 362420 505346 362656
rect 505582 362420 539952 362656
rect 540188 362420 541884 362656
rect 542120 362420 543816 362656
rect 544052 362420 545748 362656
rect 545984 362420 577026 362656
rect 577262 362420 577346 362656
rect 577582 362420 585342 362656
rect 585578 362420 585662 362656
rect 585898 362420 592650 362656
rect -8726 362336 592650 362420
rect -8726 362100 -1974 362336
rect -1738 362100 -1654 362336
rect -1418 362100 1026 362336
rect 1262 362100 1346 362336
rect 1582 362100 37026 362336
rect 37262 362100 37346 362336
rect 37582 362100 73026 362336
rect 73262 362100 73346 362336
rect 73582 362100 109026 362336
rect 109262 362100 109346 362336
rect 109582 362100 145026 362336
rect 145262 362100 145346 362336
rect 145582 362100 181026 362336
rect 181262 362100 181346 362336
rect 181582 362100 217026 362336
rect 217262 362100 217346 362336
rect 217582 362100 253026 362336
rect 253262 362100 253346 362336
rect 253582 362100 289026 362336
rect 289262 362100 289346 362336
rect 289582 362100 325026 362336
rect 325262 362100 325346 362336
rect 325582 362100 361026 362336
rect 361262 362100 361346 362336
rect 361582 362100 397026 362336
rect 397262 362100 397346 362336
rect 397582 362100 433026 362336
rect 433262 362100 433346 362336
rect 433582 362100 469026 362336
rect 469262 362100 469346 362336
rect 469582 362100 505026 362336
rect 505262 362100 505346 362336
rect 505582 362100 539952 362336
rect 540188 362100 541884 362336
rect 542120 362100 543816 362336
rect 544052 362100 545748 362336
rect 545984 362100 577026 362336
rect 577262 362100 577346 362336
rect 577582 362100 585342 362336
rect 585578 362100 585662 362336
rect 585898 362100 592650 362336
rect -8726 362068 592650 362100
rect -8726 335336 592650 335368
rect -8726 335100 -8694 335336
rect -8458 335100 -8374 335336
rect -8138 335100 9706 335336
rect 9942 335100 10026 335336
rect 10262 335100 45706 335336
rect 45942 335100 46026 335336
rect 46262 335100 81706 335336
rect 81942 335100 82026 335336
rect 82262 335100 117706 335336
rect 117942 335100 118026 335336
rect 118262 335100 153706 335336
rect 153942 335100 154026 335336
rect 154262 335100 189706 335336
rect 189942 335100 190026 335336
rect 190262 335100 225706 335336
rect 225942 335100 226026 335336
rect 226262 335100 261706 335336
rect 261942 335100 262026 335336
rect 262262 335100 297706 335336
rect 297942 335100 298026 335336
rect 298262 335100 333706 335336
rect 333942 335100 334026 335336
rect 334262 335100 369706 335336
rect 369942 335100 370026 335336
rect 370262 335100 405706 335336
rect 405942 335100 406026 335336
rect 406262 335100 441706 335336
rect 441942 335100 442026 335336
rect 442262 335100 477706 335336
rect 477942 335100 478026 335336
rect 478262 335100 513706 335336
rect 513942 335100 514026 335336
rect 514262 335100 549706 335336
rect 549942 335100 550026 335336
rect 550262 335100 592062 335336
rect 592298 335100 592382 335336
rect 592618 335100 592650 335336
rect -8726 335016 592650 335100
rect -8726 334780 -8694 335016
rect -8458 334780 -8374 335016
rect -8138 334780 9706 335016
rect 9942 334780 10026 335016
rect 10262 334780 45706 335016
rect 45942 334780 46026 335016
rect 46262 334780 81706 335016
rect 81942 334780 82026 335016
rect 82262 334780 117706 335016
rect 117942 334780 118026 335016
rect 118262 334780 153706 335016
rect 153942 334780 154026 335016
rect 154262 334780 189706 335016
rect 189942 334780 190026 335016
rect 190262 334780 225706 335016
rect 225942 334780 226026 335016
rect 226262 334780 261706 335016
rect 261942 334780 262026 335016
rect 262262 334780 297706 335016
rect 297942 334780 298026 335016
rect 298262 334780 333706 335016
rect 333942 334780 334026 335016
rect 334262 334780 369706 335016
rect 369942 334780 370026 335016
rect 370262 334780 405706 335016
rect 405942 334780 406026 335016
rect 406262 334780 441706 335016
rect 441942 334780 442026 335016
rect 442262 334780 477706 335016
rect 477942 334780 478026 335016
rect 478262 334780 513706 335016
rect 513942 334780 514026 335016
rect 514262 334780 549706 335016
rect 549942 334780 550026 335016
rect 550262 334780 592062 335016
rect 592298 334780 592382 335016
rect 592618 334780 592650 335016
rect -8726 334748 592650 334780
rect -8726 334096 592650 334128
rect -8726 333860 -7734 334096
rect -7498 333860 -7414 334096
rect -7178 333860 8466 334096
rect 8702 333860 8786 334096
rect 9022 333860 44466 334096
rect 44702 333860 44786 334096
rect 45022 333860 80466 334096
rect 80702 333860 80786 334096
rect 81022 333860 116466 334096
rect 116702 333860 116786 334096
rect 117022 333860 152466 334096
rect 152702 333860 152786 334096
rect 153022 333860 188466 334096
rect 188702 333860 188786 334096
rect 189022 333860 224466 334096
rect 224702 333860 224786 334096
rect 225022 333860 260466 334096
rect 260702 333860 260786 334096
rect 261022 333860 296466 334096
rect 296702 333860 296786 334096
rect 297022 333860 332466 334096
rect 332702 333860 332786 334096
rect 333022 333860 368466 334096
rect 368702 333860 368786 334096
rect 369022 333860 404466 334096
rect 404702 333860 404786 334096
rect 405022 333860 440466 334096
rect 440702 333860 440786 334096
rect 441022 333860 476466 334096
rect 476702 333860 476786 334096
rect 477022 333860 512466 334096
rect 512702 333860 512786 334096
rect 513022 333860 548466 334096
rect 548702 333860 548786 334096
rect 549022 333860 591102 334096
rect 591338 333860 591422 334096
rect 591658 333860 592650 334096
rect -8726 333776 592650 333860
rect -8726 333540 -7734 333776
rect -7498 333540 -7414 333776
rect -7178 333540 8466 333776
rect 8702 333540 8786 333776
rect 9022 333540 44466 333776
rect 44702 333540 44786 333776
rect 45022 333540 80466 333776
rect 80702 333540 80786 333776
rect 81022 333540 116466 333776
rect 116702 333540 116786 333776
rect 117022 333540 152466 333776
rect 152702 333540 152786 333776
rect 153022 333540 188466 333776
rect 188702 333540 188786 333776
rect 189022 333540 224466 333776
rect 224702 333540 224786 333776
rect 225022 333540 260466 333776
rect 260702 333540 260786 333776
rect 261022 333540 296466 333776
rect 296702 333540 296786 333776
rect 297022 333540 332466 333776
rect 332702 333540 332786 333776
rect 333022 333540 368466 333776
rect 368702 333540 368786 333776
rect 369022 333540 404466 333776
rect 404702 333540 404786 333776
rect 405022 333540 440466 333776
rect 440702 333540 440786 333776
rect 441022 333540 476466 333776
rect 476702 333540 476786 333776
rect 477022 333540 512466 333776
rect 512702 333540 512786 333776
rect 513022 333540 548466 333776
rect 548702 333540 548786 333776
rect 549022 333540 591102 333776
rect 591338 333540 591422 333776
rect 591658 333540 592650 333776
rect -8726 333508 592650 333540
rect -8726 332856 592650 332888
rect -8726 332620 -6774 332856
rect -6538 332620 -6454 332856
rect -6218 332620 7226 332856
rect 7462 332620 7546 332856
rect 7782 332620 43226 332856
rect 43462 332620 43546 332856
rect 43782 332620 79226 332856
rect 79462 332620 79546 332856
rect 79782 332620 115226 332856
rect 115462 332620 115546 332856
rect 115782 332620 151226 332856
rect 151462 332620 151546 332856
rect 151782 332620 187226 332856
rect 187462 332620 187546 332856
rect 187782 332620 223226 332856
rect 223462 332620 223546 332856
rect 223782 332620 259226 332856
rect 259462 332620 259546 332856
rect 259782 332620 295226 332856
rect 295462 332620 295546 332856
rect 295782 332620 331226 332856
rect 331462 332620 331546 332856
rect 331782 332620 367226 332856
rect 367462 332620 367546 332856
rect 367782 332620 403226 332856
rect 403462 332620 403546 332856
rect 403782 332620 439226 332856
rect 439462 332620 439546 332856
rect 439782 332620 475226 332856
rect 475462 332620 475546 332856
rect 475782 332620 511226 332856
rect 511462 332620 511546 332856
rect 511782 332620 547226 332856
rect 547462 332620 547546 332856
rect 547782 332620 590142 332856
rect 590378 332620 590462 332856
rect 590698 332620 592650 332856
rect -8726 332536 592650 332620
rect -8726 332300 -6774 332536
rect -6538 332300 -6454 332536
rect -6218 332300 7226 332536
rect 7462 332300 7546 332536
rect 7782 332300 43226 332536
rect 43462 332300 43546 332536
rect 43782 332300 79226 332536
rect 79462 332300 79546 332536
rect 79782 332300 115226 332536
rect 115462 332300 115546 332536
rect 115782 332300 151226 332536
rect 151462 332300 151546 332536
rect 151782 332300 187226 332536
rect 187462 332300 187546 332536
rect 187782 332300 223226 332536
rect 223462 332300 223546 332536
rect 223782 332300 259226 332536
rect 259462 332300 259546 332536
rect 259782 332300 295226 332536
rect 295462 332300 295546 332536
rect 295782 332300 331226 332536
rect 331462 332300 331546 332536
rect 331782 332300 367226 332536
rect 367462 332300 367546 332536
rect 367782 332300 403226 332536
rect 403462 332300 403546 332536
rect 403782 332300 439226 332536
rect 439462 332300 439546 332536
rect 439782 332300 475226 332536
rect 475462 332300 475546 332536
rect 475782 332300 511226 332536
rect 511462 332300 511546 332536
rect 511782 332300 547226 332536
rect 547462 332300 547546 332536
rect 547782 332300 590142 332536
rect 590378 332300 590462 332536
rect 590698 332300 592650 332536
rect -8726 332268 592650 332300
rect -8726 331616 592650 331648
rect -8726 331380 -5814 331616
rect -5578 331380 -5494 331616
rect -5258 331380 5986 331616
rect 6222 331380 6306 331616
rect 6542 331380 41986 331616
rect 42222 331380 42306 331616
rect 42542 331380 77986 331616
rect 78222 331380 78306 331616
rect 78542 331380 113986 331616
rect 114222 331380 114306 331616
rect 114542 331380 149986 331616
rect 150222 331380 150306 331616
rect 150542 331380 185986 331616
rect 186222 331380 186306 331616
rect 186542 331380 221986 331616
rect 222222 331380 222306 331616
rect 222542 331380 257986 331616
rect 258222 331380 258306 331616
rect 258542 331380 293986 331616
rect 294222 331380 294306 331616
rect 294542 331380 329986 331616
rect 330222 331380 330306 331616
rect 330542 331380 365986 331616
rect 366222 331380 366306 331616
rect 366542 331380 401986 331616
rect 402222 331380 402306 331616
rect 402542 331380 437986 331616
rect 438222 331380 438306 331616
rect 438542 331380 473986 331616
rect 474222 331380 474306 331616
rect 474542 331380 509986 331616
rect 510222 331380 510306 331616
rect 510542 331380 581986 331616
rect 582222 331380 582306 331616
rect 582542 331380 589182 331616
rect 589418 331380 589502 331616
rect 589738 331380 592650 331616
rect -8726 331296 592650 331380
rect -8726 331060 -5814 331296
rect -5578 331060 -5494 331296
rect -5258 331060 5986 331296
rect 6222 331060 6306 331296
rect 6542 331060 41986 331296
rect 42222 331060 42306 331296
rect 42542 331060 77986 331296
rect 78222 331060 78306 331296
rect 78542 331060 113986 331296
rect 114222 331060 114306 331296
rect 114542 331060 149986 331296
rect 150222 331060 150306 331296
rect 150542 331060 185986 331296
rect 186222 331060 186306 331296
rect 186542 331060 221986 331296
rect 222222 331060 222306 331296
rect 222542 331060 257986 331296
rect 258222 331060 258306 331296
rect 258542 331060 293986 331296
rect 294222 331060 294306 331296
rect 294542 331060 329986 331296
rect 330222 331060 330306 331296
rect 330542 331060 365986 331296
rect 366222 331060 366306 331296
rect 366542 331060 401986 331296
rect 402222 331060 402306 331296
rect 402542 331060 437986 331296
rect 438222 331060 438306 331296
rect 438542 331060 473986 331296
rect 474222 331060 474306 331296
rect 474542 331060 509986 331296
rect 510222 331060 510306 331296
rect 510542 331060 581986 331296
rect 582222 331060 582306 331296
rect 582542 331060 589182 331296
rect 589418 331060 589502 331296
rect 589738 331060 592650 331296
rect -8726 331028 592650 331060
rect -8726 330376 592650 330408
rect -8726 330140 -4854 330376
rect -4618 330140 -4534 330376
rect -4298 330140 4746 330376
rect 4982 330140 5066 330376
rect 5302 330140 40746 330376
rect 40982 330140 41066 330376
rect 41302 330140 76746 330376
rect 76982 330140 77066 330376
rect 77302 330140 112746 330376
rect 112982 330140 113066 330376
rect 113302 330140 148746 330376
rect 148982 330140 149066 330376
rect 149302 330140 184746 330376
rect 184982 330140 185066 330376
rect 185302 330140 220746 330376
rect 220982 330140 221066 330376
rect 221302 330140 256746 330376
rect 256982 330140 257066 330376
rect 257302 330140 292746 330376
rect 292982 330140 293066 330376
rect 293302 330140 328746 330376
rect 328982 330140 329066 330376
rect 329302 330140 364746 330376
rect 364982 330140 365066 330376
rect 365302 330140 400746 330376
rect 400982 330140 401066 330376
rect 401302 330140 436746 330376
rect 436982 330140 437066 330376
rect 437302 330140 472746 330376
rect 472982 330140 473066 330376
rect 473302 330140 508746 330376
rect 508982 330140 509066 330376
rect 509302 330140 580746 330376
rect 580982 330140 581066 330376
rect 581302 330140 588222 330376
rect 588458 330140 588542 330376
rect 588778 330140 592650 330376
rect -8726 330056 592650 330140
rect -8726 329820 -4854 330056
rect -4618 329820 -4534 330056
rect -4298 329820 4746 330056
rect 4982 329820 5066 330056
rect 5302 329820 40746 330056
rect 40982 329820 41066 330056
rect 41302 329820 76746 330056
rect 76982 329820 77066 330056
rect 77302 329820 112746 330056
rect 112982 329820 113066 330056
rect 113302 329820 148746 330056
rect 148982 329820 149066 330056
rect 149302 329820 184746 330056
rect 184982 329820 185066 330056
rect 185302 329820 220746 330056
rect 220982 329820 221066 330056
rect 221302 329820 256746 330056
rect 256982 329820 257066 330056
rect 257302 329820 292746 330056
rect 292982 329820 293066 330056
rect 293302 329820 328746 330056
rect 328982 329820 329066 330056
rect 329302 329820 364746 330056
rect 364982 329820 365066 330056
rect 365302 329820 400746 330056
rect 400982 329820 401066 330056
rect 401302 329820 436746 330056
rect 436982 329820 437066 330056
rect 437302 329820 472746 330056
rect 472982 329820 473066 330056
rect 473302 329820 508746 330056
rect 508982 329820 509066 330056
rect 509302 329820 580746 330056
rect 580982 329820 581066 330056
rect 581302 329820 588222 330056
rect 588458 329820 588542 330056
rect 588778 329820 592650 330056
rect -8726 329788 592650 329820
rect -8726 329136 592650 329168
rect -8726 328900 -3894 329136
rect -3658 328900 -3574 329136
rect -3338 328900 3506 329136
rect 3742 328900 3826 329136
rect 4062 328900 39506 329136
rect 39742 328900 39826 329136
rect 40062 328900 75506 329136
rect 75742 328900 75826 329136
rect 76062 328900 111506 329136
rect 111742 328900 111826 329136
rect 112062 328900 147506 329136
rect 147742 328900 147826 329136
rect 148062 328900 183506 329136
rect 183742 328900 183826 329136
rect 184062 328900 219506 329136
rect 219742 328900 219826 329136
rect 220062 328900 255506 329136
rect 255742 328900 255826 329136
rect 256062 328900 291506 329136
rect 291742 328900 291826 329136
rect 292062 328900 327506 329136
rect 327742 328900 327826 329136
rect 328062 328900 363506 329136
rect 363742 328900 363826 329136
rect 364062 328900 399506 329136
rect 399742 328900 399826 329136
rect 400062 328900 435506 329136
rect 435742 328900 435826 329136
rect 436062 328900 471506 329136
rect 471742 328900 471826 329136
rect 472062 328900 507506 329136
rect 507742 328900 507826 329136
rect 508062 328900 579506 329136
rect 579742 328900 579826 329136
rect 580062 328900 587262 329136
rect 587498 328900 587582 329136
rect 587818 328900 592650 329136
rect -8726 328816 592650 328900
rect -8726 328580 -3894 328816
rect -3658 328580 -3574 328816
rect -3338 328580 3506 328816
rect 3742 328580 3826 328816
rect 4062 328580 39506 328816
rect 39742 328580 39826 328816
rect 40062 328580 75506 328816
rect 75742 328580 75826 328816
rect 76062 328580 111506 328816
rect 111742 328580 111826 328816
rect 112062 328580 147506 328816
rect 147742 328580 147826 328816
rect 148062 328580 183506 328816
rect 183742 328580 183826 328816
rect 184062 328580 219506 328816
rect 219742 328580 219826 328816
rect 220062 328580 255506 328816
rect 255742 328580 255826 328816
rect 256062 328580 291506 328816
rect 291742 328580 291826 328816
rect 292062 328580 327506 328816
rect 327742 328580 327826 328816
rect 328062 328580 363506 328816
rect 363742 328580 363826 328816
rect 364062 328580 399506 328816
rect 399742 328580 399826 328816
rect 400062 328580 435506 328816
rect 435742 328580 435826 328816
rect 436062 328580 471506 328816
rect 471742 328580 471826 328816
rect 472062 328580 507506 328816
rect 507742 328580 507826 328816
rect 508062 328580 579506 328816
rect 579742 328580 579826 328816
rect 580062 328580 587262 328816
rect 587498 328580 587582 328816
rect 587818 328580 592650 328816
rect -8726 328548 592650 328580
rect -8726 327896 592650 327928
rect -8726 327660 -2934 327896
rect -2698 327660 -2614 327896
rect -2378 327660 2266 327896
rect 2502 327660 2586 327896
rect 2822 327660 38266 327896
rect 38502 327660 38586 327896
rect 38822 327660 74266 327896
rect 74502 327660 74586 327896
rect 74822 327660 110266 327896
rect 110502 327660 110586 327896
rect 110822 327660 146266 327896
rect 146502 327660 146586 327896
rect 146822 327660 182266 327896
rect 182502 327660 182586 327896
rect 182822 327660 218266 327896
rect 218502 327660 218586 327896
rect 218822 327660 254266 327896
rect 254502 327660 254586 327896
rect 254822 327660 290266 327896
rect 290502 327660 290586 327896
rect 290822 327660 326266 327896
rect 326502 327660 326586 327896
rect 326822 327660 362266 327896
rect 362502 327660 362586 327896
rect 362822 327660 398266 327896
rect 398502 327660 398586 327896
rect 398822 327660 434266 327896
rect 434502 327660 434586 327896
rect 434822 327660 470266 327896
rect 470502 327660 470586 327896
rect 470822 327660 506266 327896
rect 506502 327660 506586 327896
rect 506822 327660 540918 327896
rect 541154 327660 542850 327896
rect 543086 327660 544782 327896
rect 545018 327660 546714 327896
rect 546950 327660 578266 327896
rect 578502 327660 578586 327896
rect 578822 327660 586302 327896
rect 586538 327660 586622 327896
rect 586858 327660 592650 327896
rect -8726 327576 592650 327660
rect -8726 327340 -2934 327576
rect -2698 327340 -2614 327576
rect -2378 327340 2266 327576
rect 2502 327340 2586 327576
rect 2822 327340 38266 327576
rect 38502 327340 38586 327576
rect 38822 327340 74266 327576
rect 74502 327340 74586 327576
rect 74822 327340 110266 327576
rect 110502 327340 110586 327576
rect 110822 327340 146266 327576
rect 146502 327340 146586 327576
rect 146822 327340 182266 327576
rect 182502 327340 182586 327576
rect 182822 327340 218266 327576
rect 218502 327340 218586 327576
rect 218822 327340 254266 327576
rect 254502 327340 254586 327576
rect 254822 327340 290266 327576
rect 290502 327340 290586 327576
rect 290822 327340 326266 327576
rect 326502 327340 326586 327576
rect 326822 327340 362266 327576
rect 362502 327340 362586 327576
rect 362822 327340 398266 327576
rect 398502 327340 398586 327576
rect 398822 327340 434266 327576
rect 434502 327340 434586 327576
rect 434822 327340 470266 327576
rect 470502 327340 470586 327576
rect 470822 327340 506266 327576
rect 506502 327340 506586 327576
rect 506822 327340 540918 327576
rect 541154 327340 542850 327576
rect 543086 327340 544782 327576
rect 545018 327340 546714 327576
rect 546950 327340 578266 327576
rect 578502 327340 578586 327576
rect 578822 327340 586302 327576
rect 586538 327340 586622 327576
rect 586858 327340 592650 327576
rect -8726 327308 592650 327340
rect -8726 326656 592650 326688
rect -8726 326420 -1974 326656
rect -1738 326420 -1654 326656
rect -1418 326420 1026 326656
rect 1262 326420 1346 326656
rect 1582 326420 37026 326656
rect 37262 326420 37346 326656
rect 37582 326420 73026 326656
rect 73262 326420 73346 326656
rect 73582 326420 109026 326656
rect 109262 326420 109346 326656
rect 109582 326420 145026 326656
rect 145262 326420 145346 326656
rect 145582 326420 181026 326656
rect 181262 326420 181346 326656
rect 181582 326420 217026 326656
rect 217262 326420 217346 326656
rect 217582 326420 253026 326656
rect 253262 326420 253346 326656
rect 253582 326420 289026 326656
rect 289262 326420 289346 326656
rect 289582 326420 325026 326656
rect 325262 326420 325346 326656
rect 325582 326420 361026 326656
rect 361262 326420 361346 326656
rect 361582 326420 397026 326656
rect 397262 326420 397346 326656
rect 397582 326420 433026 326656
rect 433262 326420 433346 326656
rect 433582 326420 469026 326656
rect 469262 326420 469346 326656
rect 469582 326420 505026 326656
rect 505262 326420 505346 326656
rect 505582 326420 539952 326656
rect 540188 326420 541884 326656
rect 542120 326420 543816 326656
rect 544052 326420 545748 326656
rect 545984 326420 577026 326656
rect 577262 326420 577346 326656
rect 577582 326420 585342 326656
rect 585578 326420 585662 326656
rect 585898 326420 592650 326656
rect -8726 326336 592650 326420
rect -8726 326100 -1974 326336
rect -1738 326100 -1654 326336
rect -1418 326100 1026 326336
rect 1262 326100 1346 326336
rect 1582 326100 37026 326336
rect 37262 326100 37346 326336
rect 37582 326100 73026 326336
rect 73262 326100 73346 326336
rect 73582 326100 109026 326336
rect 109262 326100 109346 326336
rect 109582 326100 145026 326336
rect 145262 326100 145346 326336
rect 145582 326100 181026 326336
rect 181262 326100 181346 326336
rect 181582 326100 217026 326336
rect 217262 326100 217346 326336
rect 217582 326100 253026 326336
rect 253262 326100 253346 326336
rect 253582 326100 289026 326336
rect 289262 326100 289346 326336
rect 289582 326100 325026 326336
rect 325262 326100 325346 326336
rect 325582 326100 361026 326336
rect 361262 326100 361346 326336
rect 361582 326100 397026 326336
rect 397262 326100 397346 326336
rect 397582 326100 433026 326336
rect 433262 326100 433346 326336
rect 433582 326100 469026 326336
rect 469262 326100 469346 326336
rect 469582 326100 505026 326336
rect 505262 326100 505346 326336
rect 505582 326100 539952 326336
rect 540188 326100 541884 326336
rect 542120 326100 543816 326336
rect 544052 326100 545748 326336
rect 545984 326100 577026 326336
rect 577262 326100 577346 326336
rect 577582 326100 585342 326336
rect 585578 326100 585662 326336
rect 585898 326100 592650 326336
rect -8726 326068 592650 326100
rect -8726 299336 592650 299368
rect -8726 299100 -8694 299336
rect -8458 299100 -8374 299336
rect -8138 299100 9706 299336
rect 9942 299100 10026 299336
rect 10262 299100 45706 299336
rect 45942 299100 46026 299336
rect 46262 299100 81706 299336
rect 81942 299100 82026 299336
rect 82262 299100 117706 299336
rect 117942 299100 118026 299336
rect 118262 299100 153706 299336
rect 153942 299100 154026 299336
rect 154262 299100 189706 299336
rect 189942 299100 190026 299336
rect 190262 299100 225706 299336
rect 225942 299100 226026 299336
rect 226262 299100 261706 299336
rect 261942 299100 262026 299336
rect 262262 299100 297706 299336
rect 297942 299100 298026 299336
rect 298262 299100 333706 299336
rect 333942 299100 334026 299336
rect 334262 299100 369706 299336
rect 369942 299100 370026 299336
rect 370262 299100 405706 299336
rect 405942 299100 406026 299336
rect 406262 299100 441706 299336
rect 441942 299100 442026 299336
rect 442262 299100 477706 299336
rect 477942 299100 478026 299336
rect 478262 299100 513706 299336
rect 513942 299100 514026 299336
rect 514262 299100 549706 299336
rect 549942 299100 550026 299336
rect 550262 299100 592062 299336
rect 592298 299100 592382 299336
rect 592618 299100 592650 299336
rect -8726 299016 592650 299100
rect -8726 298780 -8694 299016
rect -8458 298780 -8374 299016
rect -8138 298780 9706 299016
rect 9942 298780 10026 299016
rect 10262 298780 45706 299016
rect 45942 298780 46026 299016
rect 46262 298780 81706 299016
rect 81942 298780 82026 299016
rect 82262 298780 117706 299016
rect 117942 298780 118026 299016
rect 118262 298780 153706 299016
rect 153942 298780 154026 299016
rect 154262 298780 189706 299016
rect 189942 298780 190026 299016
rect 190262 298780 225706 299016
rect 225942 298780 226026 299016
rect 226262 298780 261706 299016
rect 261942 298780 262026 299016
rect 262262 298780 297706 299016
rect 297942 298780 298026 299016
rect 298262 298780 333706 299016
rect 333942 298780 334026 299016
rect 334262 298780 369706 299016
rect 369942 298780 370026 299016
rect 370262 298780 405706 299016
rect 405942 298780 406026 299016
rect 406262 298780 441706 299016
rect 441942 298780 442026 299016
rect 442262 298780 477706 299016
rect 477942 298780 478026 299016
rect 478262 298780 513706 299016
rect 513942 298780 514026 299016
rect 514262 298780 549706 299016
rect 549942 298780 550026 299016
rect 550262 298780 592062 299016
rect 592298 298780 592382 299016
rect 592618 298780 592650 299016
rect -8726 298748 592650 298780
rect -8726 298096 592650 298128
rect -8726 297860 -7734 298096
rect -7498 297860 -7414 298096
rect -7178 297860 8466 298096
rect 8702 297860 8786 298096
rect 9022 297860 44466 298096
rect 44702 297860 44786 298096
rect 45022 297860 80466 298096
rect 80702 297860 80786 298096
rect 81022 297860 116466 298096
rect 116702 297860 116786 298096
rect 117022 297860 152466 298096
rect 152702 297860 152786 298096
rect 153022 297860 188466 298096
rect 188702 297860 188786 298096
rect 189022 297860 224466 298096
rect 224702 297860 224786 298096
rect 225022 297860 260466 298096
rect 260702 297860 260786 298096
rect 261022 297860 296466 298096
rect 296702 297860 296786 298096
rect 297022 297860 332466 298096
rect 332702 297860 332786 298096
rect 333022 297860 368466 298096
rect 368702 297860 368786 298096
rect 369022 297860 404466 298096
rect 404702 297860 404786 298096
rect 405022 297860 440466 298096
rect 440702 297860 440786 298096
rect 441022 297860 476466 298096
rect 476702 297860 476786 298096
rect 477022 297860 512466 298096
rect 512702 297860 512786 298096
rect 513022 297860 548466 298096
rect 548702 297860 548786 298096
rect 549022 297860 591102 298096
rect 591338 297860 591422 298096
rect 591658 297860 592650 298096
rect -8726 297776 592650 297860
rect -8726 297540 -7734 297776
rect -7498 297540 -7414 297776
rect -7178 297540 8466 297776
rect 8702 297540 8786 297776
rect 9022 297540 44466 297776
rect 44702 297540 44786 297776
rect 45022 297540 80466 297776
rect 80702 297540 80786 297776
rect 81022 297540 116466 297776
rect 116702 297540 116786 297776
rect 117022 297540 152466 297776
rect 152702 297540 152786 297776
rect 153022 297540 188466 297776
rect 188702 297540 188786 297776
rect 189022 297540 224466 297776
rect 224702 297540 224786 297776
rect 225022 297540 260466 297776
rect 260702 297540 260786 297776
rect 261022 297540 296466 297776
rect 296702 297540 296786 297776
rect 297022 297540 332466 297776
rect 332702 297540 332786 297776
rect 333022 297540 368466 297776
rect 368702 297540 368786 297776
rect 369022 297540 404466 297776
rect 404702 297540 404786 297776
rect 405022 297540 440466 297776
rect 440702 297540 440786 297776
rect 441022 297540 476466 297776
rect 476702 297540 476786 297776
rect 477022 297540 512466 297776
rect 512702 297540 512786 297776
rect 513022 297540 548466 297776
rect 548702 297540 548786 297776
rect 549022 297540 591102 297776
rect 591338 297540 591422 297776
rect 591658 297540 592650 297776
rect -8726 297508 592650 297540
rect -8726 296856 592650 296888
rect -8726 296620 -6774 296856
rect -6538 296620 -6454 296856
rect -6218 296620 7226 296856
rect 7462 296620 7546 296856
rect 7782 296620 43226 296856
rect 43462 296620 43546 296856
rect 43782 296620 79226 296856
rect 79462 296620 79546 296856
rect 79782 296620 115226 296856
rect 115462 296620 115546 296856
rect 115782 296620 151226 296856
rect 151462 296620 151546 296856
rect 151782 296620 187226 296856
rect 187462 296620 187546 296856
rect 187782 296620 223226 296856
rect 223462 296620 223546 296856
rect 223782 296620 259226 296856
rect 259462 296620 259546 296856
rect 259782 296620 295226 296856
rect 295462 296620 295546 296856
rect 295782 296620 331226 296856
rect 331462 296620 331546 296856
rect 331782 296620 367226 296856
rect 367462 296620 367546 296856
rect 367782 296620 403226 296856
rect 403462 296620 403546 296856
rect 403782 296620 439226 296856
rect 439462 296620 439546 296856
rect 439782 296620 475226 296856
rect 475462 296620 475546 296856
rect 475782 296620 511226 296856
rect 511462 296620 511546 296856
rect 511782 296620 547226 296856
rect 547462 296620 547546 296856
rect 547782 296620 590142 296856
rect 590378 296620 590462 296856
rect 590698 296620 592650 296856
rect -8726 296536 592650 296620
rect -8726 296300 -6774 296536
rect -6538 296300 -6454 296536
rect -6218 296300 7226 296536
rect 7462 296300 7546 296536
rect 7782 296300 43226 296536
rect 43462 296300 43546 296536
rect 43782 296300 79226 296536
rect 79462 296300 79546 296536
rect 79782 296300 115226 296536
rect 115462 296300 115546 296536
rect 115782 296300 151226 296536
rect 151462 296300 151546 296536
rect 151782 296300 187226 296536
rect 187462 296300 187546 296536
rect 187782 296300 223226 296536
rect 223462 296300 223546 296536
rect 223782 296300 259226 296536
rect 259462 296300 259546 296536
rect 259782 296300 295226 296536
rect 295462 296300 295546 296536
rect 295782 296300 331226 296536
rect 331462 296300 331546 296536
rect 331782 296300 367226 296536
rect 367462 296300 367546 296536
rect 367782 296300 403226 296536
rect 403462 296300 403546 296536
rect 403782 296300 439226 296536
rect 439462 296300 439546 296536
rect 439782 296300 475226 296536
rect 475462 296300 475546 296536
rect 475782 296300 511226 296536
rect 511462 296300 511546 296536
rect 511782 296300 547226 296536
rect 547462 296300 547546 296536
rect 547782 296300 590142 296536
rect 590378 296300 590462 296536
rect 590698 296300 592650 296536
rect -8726 296268 592650 296300
rect -8726 295616 592650 295648
rect -8726 295380 -5814 295616
rect -5578 295380 -5494 295616
rect -5258 295380 5986 295616
rect 6222 295380 6306 295616
rect 6542 295380 41986 295616
rect 42222 295380 42306 295616
rect 42542 295380 77986 295616
rect 78222 295380 78306 295616
rect 78542 295380 113986 295616
rect 114222 295380 114306 295616
rect 114542 295380 149986 295616
rect 150222 295380 150306 295616
rect 150542 295380 185986 295616
rect 186222 295380 186306 295616
rect 186542 295380 221986 295616
rect 222222 295380 222306 295616
rect 222542 295380 257986 295616
rect 258222 295380 258306 295616
rect 258542 295380 293986 295616
rect 294222 295380 294306 295616
rect 294542 295380 329986 295616
rect 330222 295380 330306 295616
rect 330542 295380 365986 295616
rect 366222 295380 366306 295616
rect 366542 295380 401986 295616
rect 402222 295380 402306 295616
rect 402542 295380 437986 295616
rect 438222 295380 438306 295616
rect 438542 295380 473986 295616
rect 474222 295380 474306 295616
rect 474542 295380 509986 295616
rect 510222 295380 510306 295616
rect 510542 295380 581986 295616
rect 582222 295380 582306 295616
rect 582542 295380 589182 295616
rect 589418 295380 589502 295616
rect 589738 295380 592650 295616
rect -8726 295296 592650 295380
rect -8726 295060 -5814 295296
rect -5578 295060 -5494 295296
rect -5258 295060 5986 295296
rect 6222 295060 6306 295296
rect 6542 295060 41986 295296
rect 42222 295060 42306 295296
rect 42542 295060 77986 295296
rect 78222 295060 78306 295296
rect 78542 295060 113986 295296
rect 114222 295060 114306 295296
rect 114542 295060 149986 295296
rect 150222 295060 150306 295296
rect 150542 295060 185986 295296
rect 186222 295060 186306 295296
rect 186542 295060 221986 295296
rect 222222 295060 222306 295296
rect 222542 295060 257986 295296
rect 258222 295060 258306 295296
rect 258542 295060 293986 295296
rect 294222 295060 294306 295296
rect 294542 295060 329986 295296
rect 330222 295060 330306 295296
rect 330542 295060 365986 295296
rect 366222 295060 366306 295296
rect 366542 295060 401986 295296
rect 402222 295060 402306 295296
rect 402542 295060 437986 295296
rect 438222 295060 438306 295296
rect 438542 295060 473986 295296
rect 474222 295060 474306 295296
rect 474542 295060 509986 295296
rect 510222 295060 510306 295296
rect 510542 295060 581986 295296
rect 582222 295060 582306 295296
rect 582542 295060 589182 295296
rect 589418 295060 589502 295296
rect 589738 295060 592650 295296
rect -8726 295028 592650 295060
rect -8726 294376 592650 294408
rect -8726 294140 -4854 294376
rect -4618 294140 -4534 294376
rect -4298 294140 4746 294376
rect 4982 294140 5066 294376
rect 5302 294140 40746 294376
rect 40982 294140 41066 294376
rect 41302 294140 76746 294376
rect 76982 294140 77066 294376
rect 77302 294140 112746 294376
rect 112982 294140 113066 294376
rect 113302 294140 148746 294376
rect 148982 294140 149066 294376
rect 149302 294140 184746 294376
rect 184982 294140 185066 294376
rect 185302 294140 220746 294376
rect 220982 294140 221066 294376
rect 221302 294140 256746 294376
rect 256982 294140 257066 294376
rect 257302 294140 292746 294376
rect 292982 294140 293066 294376
rect 293302 294140 328746 294376
rect 328982 294140 329066 294376
rect 329302 294140 364746 294376
rect 364982 294140 365066 294376
rect 365302 294140 400746 294376
rect 400982 294140 401066 294376
rect 401302 294140 436746 294376
rect 436982 294140 437066 294376
rect 437302 294140 472746 294376
rect 472982 294140 473066 294376
rect 473302 294140 508746 294376
rect 508982 294140 509066 294376
rect 509302 294140 580746 294376
rect 580982 294140 581066 294376
rect 581302 294140 588222 294376
rect 588458 294140 588542 294376
rect 588778 294140 592650 294376
rect -8726 294056 592650 294140
rect -8726 293820 -4854 294056
rect -4618 293820 -4534 294056
rect -4298 293820 4746 294056
rect 4982 293820 5066 294056
rect 5302 293820 40746 294056
rect 40982 293820 41066 294056
rect 41302 293820 76746 294056
rect 76982 293820 77066 294056
rect 77302 293820 112746 294056
rect 112982 293820 113066 294056
rect 113302 293820 148746 294056
rect 148982 293820 149066 294056
rect 149302 293820 184746 294056
rect 184982 293820 185066 294056
rect 185302 293820 220746 294056
rect 220982 293820 221066 294056
rect 221302 293820 256746 294056
rect 256982 293820 257066 294056
rect 257302 293820 292746 294056
rect 292982 293820 293066 294056
rect 293302 293820 328746 294056
rect 328982 293820 329066 294056
rect 329302 293820 364746 294056
rect 364982 293820 365066 294056
rect 365302 293820 400746 294056
rect 400982 293820 401066 294056
rect 401302 293820 436746 294056
rect 436982 293820 437066 294056
rect 437302 293820 472746 294056
rect 472982 293820 473066 294056
rect 473302 293820 508746 294056
rect 508982 293820 509066 294056
rect 509302 293820 580746 294056
rect 580982 293820 581066 294056
rect 581302 293820 588222 294056
rect 588458 293820 588542 294056
rect 588778 293820 592650 294056
rect -8726 293788 592650 293820
rect -8726 293136 592650 293168
rect -8726 292900 -3894 293136
rect -3658 292900 -3574 293136
rect -3338 292900 3506 293136
rect 3742 292900 3826 293136
rect 4062 292900 39506 293136
rect 39742 292900 39826 293136
rect 40062 292900 75506 293136
rect 75742 292900 75826 293136
rect 76062 292900 111506 293136
rect 111742 292900 111826 293136
rect 112062 292900 147506 293136
rect 147742 292900 147826 293136
rect 148062 292900 183506 293136
rect 183742 292900 183826 293136
rect 184062 292900 219506 293136
rect 219742 292900 219826 293136
rect 220062 292900 255506 293136
rect 255742 292900 255826 293136
rect 256062 292900 291506 293136
rect 291742 292900 291826 293136
rect 292062 292900 327506 293136
rect 327742 292900 327826 293136
rect 328062 292900 363506 293136
rect 363742 292900 363826 293136
rect 364062 292900 399506 293136
rect 399742 292900 399826 293136
rect 400062 292900 435506 293136
rect 435742 292900 435826 293136
rect 436062 292900 471506 293136
rect 471742 292900 471826 293136
rect 472062 292900 507506 293136
rect 507742 292900 507826 293136
rect 508062 292900 579506 293136
rect 579742 292900 579826 293136
rect 580062 292900 587262 293136
rect 587498 292900 587582 293136
rect 587818 292900 592650 293136
rect -8726 292816 592650 292900
rect -8726 292580 -3894 292816
rect -3658 292580 -3574 292816
rect -3338 292580 3506 292816
rect 3742 292580 3826 292816
rect 4062 292580 39506 292816
rect 39742 292580 39826 292816
rect 40062 292580 75506 292816
rect 75742 292580 75826 292816
rect 76062 292580 111506 292816
rect 111742 292580 111826 292816
rect 112062 292580 147506 292816
rect 147742 292580 147826 292816
rect 148062 292580 183506 292816
rect 183742 292580 183826 292816
rect 184062 292580 219506 292816
rect 219742 292580 219826 292816
rect 220062 292580 255506 292816
rect 255742 292580 255826 292816
rect 256062 292580 291506 292816
rect 291742 292580 291826 292816
rect 292062 292580 327506 292816
rect 327742 292580 327826 292816
rect 328062 292580 363506 292816
rect 363742 292580 363826 292816
rect 364062 292580 399506 292816
rect 399742 292580 399826 292816
rect 400062 292580 435506 292816
rect 435742 292580 435826 292816
rect 436062 292580 471506 292816
rect 471742 292580 471826 292816
rect 472062 292580 507506 292816
rect 507742 292580 507826 292816
rect 508062 292580 579506 292816
rect 579742 292580 579826 292816
rect 580062 292580 587262 292816
rect 587498 292580 587582 292816
rect 587818 292580 592650 292816
rect -8726 292548 592650 292580
rect -8726 291896 592650 291928
rect -8726 291660 -2934 291896
rect -2698 291660 -2614 291896
rect -2378 291660 2266 291896
rect 2502 291660 2586 291896
rect 2822 291660 38266 291896
rect 38502 291660 38586 291896
rect 38822 291660 74266 291896
rect 74502 291660 74586 291896
rect 74822 291660 110266 291896
rect 110502 291660 110586 291896
rect 110822 291660 146266 291896
rect 146502 291660 146586 291896
rect 146822 291660 182266 291896
rect 182502 291660 182586 291896
rect 182822 291660 218266 291896
rect 218502 291660 218586 291896
rect 218822 291660 254266 291896
rect 254502 291660 254586 291896
rect 254822 291660 290266 291896
rect 290502 291660 290586 291896
rect 290822 291660 326266 291896
rect 326502 291660 326586 291896
rect 326822 291660 362266 291896
rect 362502 291660 362586 291896
rect 362822 291660 398266 291896
rect 398502 291660 398586 291896
rect 398822 291660 434266 291896
rect 434502 291660 434586 291896
rect 434822 291660 470266 291896
rect 470502 291660 470586 291896
rect 470822 291660 506266 291896
rect 506502 291660 506586 291896
rect 506822 291660 540918 291896
rect 541154 291660 542850 291896
rect 543086 291660 544782 291896
rect 545018 291660 546714 291896
rect 546950 291660 578266 291896
rect 578502 291660 578586 291896
rect 578822 291660 586302 291896
rect 586538 291660 586622 291896
rect 586858 291660 592650 291896
rect -8726 291576 592650 291660
rect -8726 291340 -2934 291576
rect -2698 291340 -2614 291576
rect -2378 291340 2266 291576
rect 2502 291340 2586 291576
rect 2822 291340 38266 291576
rect 38502 291340 38586 291576
rect 38822 291340 74266 291576
rect 74502 291340 74586 291576
rect 74822 291340 110266 291576
rect 110502 291340 110586 291576
rect 110822 291340 146266 291576
rect 146502 291340 146586 291576
rect 146822 291340 182266 291576
rect 182502 291340 182586 291576
rect 182822 291340 218266 291576
rect 218502 291340 218586 291576
rect 218822 291340 254266 291576
rect 254502 291340 254586 291576
rect 254822 291340 290266 291576
rect 290502 291340 290586 291576
rect 290822 291340 326266 291576
rect 326502 291340 326586 291576
rect 326822 291340 362266 291576
rect 362502 291340 362586 291576
rect 362822 291340 398266 291576
rect 398502 291340 398586 291576
rect 398822 291340 434266 291576
rect 434502 291340 434586 291576
rect 434822 291340 470266 291576
rect 470502 291340 470586 291576
rect 470822 291340 506266 291576
rect 506502 291340 506586 291576
rect 506822 291340 540918 291576
rect 541154 291340 542850 291576
rect 543086 291340 544782 291576
rect 545018 291340 546714 291576
rect 546950 291340 578266 291576
rect 578502 291340 578586 291576
rect 578822 291340 586302 291576
rect 586538 291340 586622 291576
rect 586858 291340 592650 291576
rect -8726 291308 592650 291340
rect -8726 290656 592650 290688
rect -8726 290420 -1974 290656
rect -1738 290420 -1654 290656
rect -1418 290420 1026 290656
rect 1262 290420 1346 290656
rect 1582 290420 37026 290656
rect 37262 290420 37346 290656
rect 37582 290420 73026 290656
rect 73262 290420 73346 290656
rect 73582 290420 109026 290656
rect 109262 290420 109346 290656
rect 109582 290420 145026 290656
rect 145262 290420 145346 290656
rect 145582 290420 181026 290656
rect 181262 290420 181346 290656
rect 181582 290420 217026 290656
rect 217262 290420 217346 290656
rect 217582 290420 253026 290656
rect 253262 290420 253346 290656
rect 253582 290420 289026 290656
rect 289262 290420 289346 290656
rect 289582 290420 325026 290656
rect 325262 290420 325346 290656
rect 325582 290420 361026 290656
rect 361262 290420 361346 290656
rect 361582 290420 397026 290656
rect 397262 290420 397346 290656
rect 397582 290420 433026 290656
rect 433262 290420 433346 290656
rect 433582 290420 469026 290656
rect 469262 290420 469346 290656
rect 469582 290420 505026 290656
rect 505262 290420 505346 290656
rect 505582 290420 539952 290656
rect 540188 290420 541884 290656
rect 542120 290420 543816 290656
rect 544052 290420 545748 290656
rect 545984 290420 577026 290656
rect 577262 290420 577346 290656
rect 577582 290420 585342 290656
rect 585578 290420 585662 290656
rect 585898 290420 592650 290656
rect -8726 290336 592650 290420
rect -8726 290100 -1974 290336
rect -1738 290100 -1654 290336
rect -1418 290100 1026 290336
rect 1262 290100 1346 290336
rect 1582 290100 37026 290336
rect 37262 290100 37346 290336
rect 37582 290100 73026 290336
rect 73262 290100 73346 290336
rect 73582 290100 109026 290336
rect 109262 290100 109346 290336
rect 109582 290100 145026 290336
rect 145262 290100 145346 290336
rect 145582 290100 181026 290336
rect 181262 290100 181346 290336
rect 181582 290100 217026 290336
rect 217262 290100 217346 290336
rect 217582 290100 253026 290336
rect 253262 290100 253346 290336
rect 253582 290100 289026 290336
rect 289262 290100 289346 290336
rect 289582 290100 325026 290336
rect 325262 290100 325346 290336
rect 325582 290100 361026 290336
rect 361262 290100 361346 290336
rect 361582 290100 397026 290336
rect 397262 290100 397346 290336
rect 397582 290100 433026 290336
rect 433262 290100 433346 290336
rect 433582 290100 469026 290336
rect 469262 290100 469346 290336
rect 469582 290100 505026 290336
rect 505262 290100 505346 290336
rect 505582 290100 539952 290336
rect 540188 290100 541884 290336
rect 542120 290100 543816 290336
rect 544052 290100 545748 290336
rect 545984 290100 577026 290336
rect 577262 290100 577346 290336
rect 577582 290100 585342 290336
rect 585578 290100 585662 290336
rect 585898 290100 592650 290336
rect -8726 290068 592650 290100
rect -8726 263336 592650 263368
rect -8726 263100 -8694 263336
rect -8458 263100 -8374 263336
rect -8138 263100 9706 263336
rect 9942 263100 10026 263336
rect 10262 263100 45706 263336
rect 45942 263100 46026 263336
rect 46262 263100 81706 263336
rect 81942 263100 82026 263336
rect 82262 263100 117706 263336
rect 117942 263100 118026 263336
rect 118262 263100 153706 263336
rect 153942 263100 154026 263336
rect 154262 263100 189706 263336
rect 189942 263100 190026 263336
rect 190262 263100 225706 263336
rect 225942 263100 226026 263336
rect 226262 263100 261706 263336
rect 261942 263100 262026 263336
rect 262262 263100 297706 263336
rect 297942 263100 298026 263336
rect 298262 263100 333706 263336
rect 333942 263100 334026 263336
rect 334262 263100 369706 263336
rect 369942 263100 370026 263336
rect 370262 263100 405706 263336
rect 405942 263100 406026 263336
rect 406262 263100 441706 263336
rect 441942 263100 442026 263336
rect 442262 263100 477706 263336
rect 477942 263100 478026 263336
rect 478262 263100 513706 263336
rect 513942 263100 514026 263336
rect 514262 263100 549706 263336
rect 549942 263100 550026 263336
rect 550262 263100 592062 263336
rect 592298 263100 592382 263336
rect 592618 263100 592650 263336
rect -8726 263016 592650 263100
rect -8726 262780 -8694 263016
rect -8458 262780 -8374 263016
rect -8138 262780 9706 263016
rect 9942 262780 10026 263016
rect 10262 262780 45706 263016
rect 45942 262780 46026 263016
rect 46262 262780 81706 263016
rect 81942 262780 82026 263016
rect 82262 262780 117706 263016
rect 117942 262780 118026 263016
rect 118262 262780 153706 263016
rect 153942 262780 154026 263016
rect 154262 262780 189706 263016
rect 189942 262780 190026 263016
rect 190262 262780 225706 263016
rect 225942 262780 226026 263016
rect 226262 262780 261706 263016
rect 261942 262780 262026 263016
rect 262262 262780 297706 263016
rect 297942 262780 298026 263016
rect 298262 262780 333706 263016
rect 333942 262780 334026 263016
rect 334262 262780 369706 263016
rect 369942 262780 370026 263016
rect 370262 262780 405706 263016
rect 405942 262780 406026 263016
rect 406262 262780 441706 263016
rect 441942 262780 442026 263016
rect 442262 262780 477706 263016
rect 477942 262780 478026 263016
rect 478262 262780 513706 263016
rect 513942 262780 514026 263016
rect 514262 262780 549706 263016
rect 549942 262780 550026 263016
rect 550262 262780 592062 263016
rect 592298 262780 592382 263016
rect 592618 262780 592650 263016
rect -8726 262748 592650 262780
rect -8726 262096 592650 262128
rect -8726 261860 -7734 262096
rect -7498 261860 -7414 262096
rect -7178 261860 8466 262096
rect 8702 261860 8786 262096
rect 9022 261860 44466 262096
rect 44702 261860 44786 262096
rect 45022 261860 80466 262096
rect 80702 261860 80786 262096
rect 81022 261860 116466 262096
rect 116702 261860 116786 262096
rect 117022 261860 152466 262096
rect 152702 261860 152786 262096
rect 153022 261860 188466 262096
rect 188702 261860 188786 262096
rect 189022 261860 224466 262096
rect 224702 261860 224786 262096
rect 225022 261860 260466 262096
rect 260702 261860 260786 262096
rect 261022 261860 296466 262096
rect 296702 261860 296786 262096
rect 297022 261860 332466 262096
rect 332702 261860 332786 262096
rect 333022 261860 368466 262096
rect 368702 261860 368786 262096
rect 369022 261860 404466 262096
rect 404702 261860 404786 262096
rect 405022 261860 440466 262096
rect 440702 261860 440786 262096
rect 441022 261860 476466 262096
rect 476702 261860 476786 262096
rect 477022 261860 512466 262096
rect 512702 261860 512786 262096
rect 513022 261860 548466 262096
rect 548702 261860 548786 262096
rect 549022 261860 591102 262096
rect 591338 261860 591422 262096
rect 591658 261860 592650 262096
rect -8726 261776 592650 261860
rect -8726 261540 -7734 261776
rect -7498 261540 -7414 261776
rect -7178 261540 8466 261776
rect 8702 261540 8786 261776
rect 9022 261540 44466 261776
rect 44702 261540 44786 261776
rect 45022 261540 80466 261776
rect 80702 261540 80786 261776
rect 81022 261540 116466 261776
rect 116702 261540 116786 261776
rect 117022 261540 152466 261776
rect 152702 261540 152786 261776
rect 153022 261540 188466 261776
rect 188702 261540 188786 261776
rect 189022 261540 224466 261776
rect 224702 261540 224786 261776
rect 225022 261540 260466 261776
rect 260702 261540 260786 261776
rect 261022 261540 296466 261776
rect 296702 261540 296786 261776
rect 297022 261540 332466 261776
rect 332702 261540 332786 261776
rect 333022 261540 368466 261776
rect 368702 261540 368786 261776
rect 369022 261540 404466 261776
rect 404702 261540 404786 261776
rect 405022 261540 440466 261776
rect 440702 261540 440786 261776
rect 441022 261540 476466 261776
rect 476702 261540 476786 261776
rect 477022 261540 512466 261776
rect 512702 261540 512786 261776
rect 513022 261540 548466 261776
rect 548702 261540 548786 261776
rect 549022 261540 591102 261776
rect 591338 261540 591422 261776
rect 591658 261540 592650 261776
rect -8726 261508 592650 261540
rect -8726 260856 592650 260888
rect -8726 260620 -6774 260856
rect -6538 260620 -6454 260856
rect -6218 260620 7226 260856
rect 7462 260620 7546 260856
rect 7782 260620 43226 260856
rect 43462 260620 43546 260856
rect 43782 260620 79226 260856
rect 79462 260620 79546 260856
rect 79782 260620 115226 260856
rect 115462 260620 115546 260856
rect 115782 260620 151226 260856
rect 151462 260620 151546 260856
rect 151782 260620 187226 260856
rect 187462 260620 187546 260856
rect 187782 260620 223226 260856
rect 223462 260620 223546 260856
rect 223782 260620 259226 260856
rect 259462 260620 259546 260856
rect 259782 260620 295226 260856
rect 295462 260620 295546 260856
rect 295782 260620 331226 260856
rect 331462 260620 331546 260856
rect 331782 260620 367226 260856
rect 367462 260620 367546 260856
rect 367782 260620 403226 260856
rect 403462 260620 403546 260856
rect 403782 260620 439226 260856
rect 439462 260620 439546 260856
rect 439782 260620 475226 260856
rect 475462 260620 475546 260856
rect 475782 260620 511226 260856
rect 511462 260620 511546 260856
rect 511782 260620 547226 260856
rect 547462 260620 547546 260856
rect 547782 260620 590142 260856
rect 590378 260620 590462 260856
rect 590698 260620 592650 260856
rect -8726 260536 592650 260620
rect -8726 260300 -6774 260536
rect -6538 260300 -6454 260536
rect -6218 260300 7226 260536
rect 7462 260300 7546 260536
rect 7782 260300 43226 260536
rect 43462 260300 43546 260536
rect 43782 260300 79226 260536
rect 79462 260300 79546 260536
rect 79782 260300 115226 260536
rect 115462 260300 115546 260536
rect 115782 260300 151226 260536
rect 151462 260300 151546 260536
rect 151782 260300 187226 260536
rect 187462 260300 187546 260536
rect 187782 260300 223226 260536
rect 223462 260300 223546 260536
rect 223782 260300 259226 260536
rect 259462 260300 259546 260536
rect 259782 260300 295226 260536
rect 295462 260300 295546 260536
rect 295782 260300 331226 260536
rect 331462 260300 331546 260536
rect 331782 260300 367226 260536
rect 367462 260300 367546 260536
rect 367782 260300 403226 260536
rect 403462 260300 403546 260536
rect 403782 260300 439226 260536
rect 439462 260300 439546 260536
rect 439782 260300 475226 260536
rect 475462 260300 475546 260536
rect 475782 260300 511226 260536
rect 511462 260300 511546 260536
rect 511782 260300 547226 260536
rect 547462 260300 547546 260536
rect 547782 260300 590142 260536
rect 590378 260300 590462 260536
rect 590698 260300 592650 260536
rect -8726 260268 592650 260300
rect -8726 259616 592650 259648
rect -8726 259380 -5814 259616
rect -5578 259380 -5494 259616
rect -5258 259380 5986 259616
rect 6222 259380 6306 259616
rect 6542 259380 41986 259616
rect 42222 259380 42306 259616
rect 42542 259380 77986 259616
rect 78222 259380 78306 259616
rect 78542 259380 113986 259616
rect 114222 259380 114306 259616
rect 114542 259380 149986 259616
rect 150222 259380 150306 259616
rect 150542 259380 185986 259616
rect 186222 259380 186306 259616
rect 186542 259380 221986 259616
rect 222222 259380 222306 259616
rect 222542 259380 257986 259616
rect 258222 259380 258306 259616
rect 258542 259380 293986 259616
rect 294222 259380 294306 259616
rect 294542 259380 329986 259616
rect 330222 259380 330306 259616
rect 330542 259380 365986 259616
rect 366222 259380 366306 259616
rect 366542 259380 401986 259616
rect 402222 259380 402306 259616
rect 402542 259380 437986 259616
rect 438222 259380 438306 259616
rect 438542 259380 473986 259616
rect 474222 259380 474306 259616
rect 474542 259380 509986 259616
rect 510222 259380 510306 259616
rect 510542 259380 545986 259616
rect 546222 259380 546306 259616
rect 546542 259380 581986 259616
rect 582222 259380 582306 259616
rect 582542 259380 589182 259616
rect 589418 259380 589502 259616
rect 589738 259380 592650 259616
rect -8726 259296 592650 259380
rect -8726 259060 -5814 259296
rect -5578 259060 -5494 259296
rect -5258 259060 5986 259296
rect 6222 259060 6306 259296
rect 6542 259060 41986 259296
rect 42222 259060 42306 259296
rect 42542 259060 77986 259296
rect 78222 259060 78306 259296
rect 78542 259060 113986 259296
rect 114222 259060 114306 259296
rect 114542 259060 149986 259296
rect 150222 259060 150306 259296
rect 150542 259060 185986 259296
rect 186222 259060 186306 259296
rect 186542 259060 221986 259296
rect 222222 259060 222306 259296
rect 222542 259060 257986 259296
rect 258222 259060 258306 259296
rect 258542 259060 293986 259296
rect 294222 259060 294306 259296
rect 294542 259060 329986 259296
rect 330222 259060 330306 259296
rect 330542 259060 365986 259296
rect 366222 259060 366306 259296
rect 366542 259060 401986 259296
rect 402222 259060 402306 259296
rect 402542 259060 437986 259296
rect 438222 259060 438306 259296
rect 438542 259060 473986 259296
rect 474222 259060 474306 259296
rect 474542 259060 509986 259296
rect 510222 259060 510306 259296
rect 510542 259060 545986 259296
rect 546222 259060 546306 259296
rect 546542 259060 581986 259296
rect 582222 259060 582306 259296
rect 582542 259060 589182 259296
rect 589418 259060 589502 259296
rect 589738 259060 592650 259296
rect -8726 259028 592650 259060
rect -8726 258376 592650 258408
rect -8726 258140 -4854 258376
rect -4618 258140 -4534 258376
rect -4298 258140 4746 258376
rect 4982 258140 5066 258376
rect 5302 258140 40746 258376
rect 40982 258140 41066 258376
rect 41302 258140 76746 258376
rect 76982 258140 77066 258376
rect 77302 258140 112746 258376
rect 112982 258140 113066 258376
rect 113302 258140 148746 258376
rect 148982 258140 149066 258376
rect 149302 258140 184746 258376
rect 184982 258140 185066 258376
rect 185302 258140 220746 258376
rect 220982 258140 221066 258376
rect 221302 258140 256746 258376
rect 256982 258140 257066 258376
rect 257302 258140 292746 258376
rect 292982 258140 293066 258376
rect 293302 258140 328746 258376
rect 328982 258140 329066 258376
rect 329302 258140 364746 258376
rect 364982 258140 365066 258376
rect 365302 258140 400746 258376
rect 400982 258140 401066 258376
rect 401302 258140 436746 258376
rect 436982 258140 437066 258376
rect 437302 258140 472746 258376
rect 472982 258140 473066 258376
rect 473302 258140 508746 258376
rect 508982 258140 509066 258376
rect 509302 258140 544746 258376
rect 544982 258140 545066 258376
rect 545302 258140 580746 258376
rect 580982 258140 581066 258376
rect 581302 258140 588222 258376
rect 588458 258140 588542 258376
rect 588778 258140 592650 258376
rect -8726 258056 592650 258140
rect -8726 257820 -4854 258056
rect -4618 257820 -4534 258056
rect -4298 257820 4746 258056
rect 4982 257820 5066 258056
rect 5302 257820 40746 258056
rect 40982 257820 41066 258056
rect 41302 257820 76746 258056
rect 76982 257820 77066 258056
rect 77302 257820 112746 258056
rect 112982 257820 113066 258056
rect 113302 257820 148746 258056
rect 148982 257820 149066 258056
rect 149302 257820 184746 258056
rect 184982 257820 185066 258056
rect 185302 257820 220746 258056
rect 220982 257820 221066 258056
rect 221302 257820 256746 258056
rect 256982 257820 257066 258056
rect 257302 257820 292746 258056
rect 292982 257820 293066 258056
rect 293302 257820 328746 258056
rect 328982 257820 329066 258056
rect 329302 257820 364746 258056
rect 364982 257820 365066 258056
rect 365302 257820 400746 258056
rect 400982 257820 401066 258056
rect 401302 257820 436746 258056
rect 436982 257820 437066 258056
rect 437302 257820 472746 258056
rect 472982 257820 473066 258056
rect 473302 257820 508746 258056
rect 508982 257820 509066 258056
rect 509302 257820 544746 258056
rect 544982 257820 545066 258056
rect 545302 257820 580746 258056
rect 580982 257820 581066 258056
rect 581302 257820 588222 258056
rect 588458 257820 588542 258056
rect 588778 257820 592650 258056
rect -8726 257788 592650 257820
rect -8726 257136 592650 257168
rect -8726 256900 -3894 257136
rect -3658 256900 -3574 257136
rect -3338 256900 3506 257136
rect 3742 256900 3826 257136
rect 4062 256900 39506 257136
rect 39742 256900 39826 257136
rect 40062 256900 75506 257136
rect 75742 256900 75826 257136
rect 76062 256900 111506 257136
rect 111742 256900 111826 257136
rect 112062 256900 147506 257136
rect 147742 256900 147826 257136
rect 148062 256900 183506 257136
rect 183742 256900 183826 257136
rect 184062 256900 219506 257136
rect 219742 256900 219826 257136
rect 220062 256900 255506 257136
rect 255742 256900 255826 257136
rect 256062 256900 291506 257136
rect 291742 256900 291826 257136
rect 292062 256900 327506 257136
rect 327742 256900 327826 257136
rect 328062 256900 363506 257136
rect 363742 256900 363826 257136
rect 364062 256900 399506 257136
rect 399742 256900 399826 257136
rect 400062 256900 435506 257136
rect 435742 256900 435826 257136
rect 436062 256900 471506 257136
rect 471742 256900 471826 257136
rect 472062 256900 507506 257136
rect 507742 256900 507826 257136
rect 508062 256900 543506 257136
rect 543742 256900 543826 257136
rect 544062 256900 579506 257136
rect 579742 256900 579826 257136
rect 580062 256900 587262 257136
rect 587498 256900 587582 257136
rect 587818 256900 592650 257136
rect -8726 256816 592650 256900
rect -8726 256580 -3894 256816
rect -3658 256580 -3574 256816
rect -3338 256580 3506 256816
rect 3742 256580 3826 256816
rect 4062 256580 39506 256816
rect 39742 256580 39826 256816
rect 40062 256580 75506 256816
rect 75742 256580 75826 256816
rect 76062 256580 111506 256816
rect 111742 256580 111826 256816
rect 112062 256580 147506 256816
rect 147742 256580 147826 256816
rect 148062 256580 183506 256816
rect 183742 256580 183826 256816
rect 184062 256580 219506 256816
rect 219742 256580 219826 256816
rect 220062 256580 255506 256816
rect 255742 256580 255826 256816
rect 256062 256580 291506 256816
rect 291742 256580 291826 256816
rect 292062 256580 327506 256816
rect 327742 256580 327826 256816
rect 328062 256580 363506 256816
rect 363742 256580 363826 256816
rect 364062 256580 399506 256816
rect 399742 256580 399826 256816
rect 400062 256580 435506 256816
rect 435742 256580 435826 256816
rect 436062 256580 471506 256816
rect 471742 256580 471826 256816
rect 472062 256580 507506 256816
rect 507742 256580 507826 256816
rect 508062 256580 543506 256816
rect 543742 256580 543826 256816
rect 544062 256580 579506 256816
rect 579742 256580 579826 256816
rect 580062 256580 587262 256816
rect 587498 256580 587582 256816
rect 587818 256580 592650 256816
rect -8726 256548 592650 256580
rect -8726 255896 592650 255928
rect -8726 255660 -2934 255896
rect -2698 255660 -2614 255896
rect -2378 255660 2266 255896
rect 2502 255660 2586 255896
rect 2822 255660 38266 255896
rect 38502 255660 38586 255896
rect 38822 255660 74266 255896
rect 74502 255660 74586 255896
rect 74822 255660 110266 255896
rect 110502 255660 110586 255896
rect 110822 255660 146266 255896
rect 146502 255660 146586 255896
rect 146822 255660 182266 255896
rect 182502 255660 182586 255896
rect 182822 255660 218266 255896
rect 218502 255660 218586 255896
rect 218822 255660 254266 255896
rect 254502 255660 254586 255896
rect 254822 255660 290266 255896
rect 290502 255660 290586 255896
rect 290822 255660 326266 255896
rect 326502 255660 326586 255896
rect 326822 255660 362266 255896
rect 362502 255660 362586 255896
rect 362822 255660 398266 255896
rect 398502 255660 398586 255896
rect 398822 255660 434266 255896
rect 434502 255660 434586 255896
rect 434822 255660 470266 255896
rect 470502 255660 470586 255896
rect 470822 255660 506266 255896
rect 506502 255660 506586 255896
rect 506822 255660 542266 255896
rect 542502 255660 542586 255896
rect 542822 255660 578266 255896
rect 578502 255660 578586 255896
rect 578822 255660 586302 255896
rect 586538 255660 586622 255896
rect 586858 255660 592650 255896
rect -8726 255576 592650 255660
rect -8726 255340 -2934 255576
rect -2698 255340 -2614 255576
rect -2378 255340 2266 255576
rect 2502 255340 2586 255576
rect 2822 255340 38266 255576
rect 38502 255340 38586 255576
rect 38822 255340 74266 255576
rect 74502 255340 74586 255576
rect 74822 255340 110266 255576
rect 110502 255340 110586 255576
rect 110822 255340 146266 255576
rect 146502 255340 146586 255576
rect 146822 255340 182266 255576
rect 182502 255340 182586 255576
rect 182822 255340 218266 255576
rect 218502 255340 218586 255576
rect 218822 255340 254266 255576
rect 254502 255340 254586 255576
rect 254822 255340 290266 255576
rect 290502 255340 290586 255576
rect 290822 255340 326266 255576
rect 326502 255340 326586 255576
rect 326822 255340 362266 255576
rect 362502 255340 362586 255576
rect 362822 255340 398266 255576
rect 398502 255340 398586 255576
rect 398822 255340 434266 255576
rect 434502 255340 434586 255576
rect 434822 255340 470266 255576
rect 470502 255340 470586 255576
rect 470822 255340 506266 255576
rect 506502 255340 506586 255576
rect 506822 255340 542266 255576
rect 542502 255340 542586 255576
rect 542822 255340 578266 255576
rect 578502 255340 578586 255576
rect 578822 255340 586302 255576
rect 586538 255340 586622 255576
rect 586858 255340 592650 255576
rect -8726 255308 592650 255340
rect -8726 254656 592650 254688
rect -8726 254420 -1974 254656
rect -1738 254420 -1654 254656
rect -1418 254420 1026 254656
rect 1262 254420 1346 254656
rect 1582 254420 37026 254656
rect 37262 254420 37346 254656
rect 37582 254420 73026 254656
rect 73262 254420 73346 254656
rect 73582 254420 109026 254656
rect 109262 254420 109346 254656
rect 109582 254420 145026 254656
rect 145262 254420 145346 254656
rect 145582 254420 181026 254656
rect 181262 254420 181346 254656
rect 181582 254420 217026 254656
rect 217262 254420 217346 254656
rect 217582 254420 253026 254656
rect 253262 254420 253346 254656
rect 253582 254420 289026 254656
rect 289262 254420 289346 254656
rect 289582 254420 325026 254656
rect 325262 254420 325346 254656
rect 325582 254420 361026 254656
rect 361262 254420 361346 254656
rect 361582 254420 397026 254656
rect 397262 254420 397346 254656
rect 397582 254420 433026 254656
rect 433262 254420 433346 254656
rect 433582 254420 469026 254656
rect 469262 254420 469346 254656
rect 469582 254420 505026 254656
rect 505262 254420 505346 254656
rect 505582 254420 541026 254656
rect 541262 254420 541346 254656
rect 541582 254420 577026 254656
rect 577262 254420 577346 254656
rect 577582 254420 585342 254656
rect 585578 254420 585662 254656
rect 585898 254420 592650 254656
rect -8726 254336 592650 254420
rect -8726 254100 -1974 254336
rect -1738 254100 -1654 254336
rect -1418 254100 1026 254336
rect 1262 254100 1346 254336
rect 1582 254100 37026 254336
rect 37262 254100 37346 254336
rect 37582 254100 73026 254336
rect 73262 254100 73346 254336
rect 73582 254100 109026 254336
rect 109262 254100 109346 254336
rect 109582 254100 145026 254336
rect 145262 254100 145346 254336
rect 145582 254100 181026 254336
rect 181262 254100 181346 254336
rect 181582 254100 217026 254336
rect 217262 254100 217346 254336
rect 217582 254100 253026 254336
rect 253262 254100 253346 254336
rect 253582 254100 289026 254336
rect 289262 254100 289346 254336
rect 289582 254100 325026 254336
rect 325262 254100 325346 254336
rect 325582 254100 361026 254336
rect 361262 254100 361346 254336
rect 361582 254100 397026 254336
rect 397262 254100 397346 254336
rect 397582 254100 433026 254336
rect 433262 254100 433346 254336
rect 433582 254100 469026 254336
rect 469262 254100 469346 254336
rect 469582 254100 505026 254336
rect 505262 254100 505346 254336
rect 505582 254100 541026 254336
rect 541262 254100 541346 254336
rect 541582 254100 577026 254336
rect 577262 254100 577346 254336
rect 577582 254100 585342 254336
rect 585578 254100 585662 254336
rect 585898 254100 592650 254336
rect -8726 254068 592650 254100
rect -8726 227336 592650 227368
rect -8726 227100 -8694 227336
rect -8458 227100 -8374 227336
rect -8138 227100 9706 227336
rect 9942 227100 10026 227336
rect 10262 227100 45706 227336
rect 45942 227100 46026 227336
rect 46262 227100 81706 227336
rect 81942 227100 82026 227336
rect 82262 227100 117706 227336
rect 117942 227100 118026 227336
rect 118262 227100 153706 227336
rect 153942 227100 154026 227336
rect 154262 227100 189706 227336
rect 189942 227100 190026 227336
rect 190262 227100 225706 227336
rect 225942 227100 226026 227336
rect 226262 227100 261706 227336
rect 261942 227100 262026 227336
rect 262262 227100 297706 227336
rect 297942 227100 298026 227336
rect 298262 227100 333706 227336
rect 333942 227100 334026 227336
rect 334262 227100 369706 227336
rect 369942 227100 370026 227336
rect 370262 227100 405706 227336
rect 405942 227100 406026 227336
rect 406262 227100 441706 227336
rect 441942 227100 442026 227336
rect 442262 227100 477706 227336
rect 477942 227100 478026 227336
rect 478262 227100 513706 227336
rect 513942 227100 514026 227336
rect 514262 227100 549706 227336
rect 549942 227100 550026 227336
rect 550262 227100 592062 227336
rect 592298 227100 592382 227336
rect 592618 227100 592650 227336
rect -8726 227016 592650 227100
rect -8726 226780 -8694 227016
rect -8458 226780 -8374 227016
rect -8138 226780 9706 227016
rect 9942 226780 10026 227016
rect 10262 226780 45706 227016
rect 45942 226780 46026 227016
rect 46262 226780 81706 227016
rect 81942 226780 82026 227016
rect 82262 226780 117706 227016
rect 117942 226780 118026 227016
rect 118262 226780 153706 227016
rect 153942 226780 154026 227016
rect 154262 226780 189706 227016
rect 189942 226780 190026 227016
rect 190262 226780 225706 227016
rect 225942 226780 226026 227016
rect 226262 226780 261706 227016
rect 261942 226780 262026 227016
rect 262262 226780 297706 227016
rect 297942 226780 298026 227016
rect 298262 226780 333706 227016
rect 333942 226780 334026 227016
rect 334262 226780 369706 227016
rect 369942 226780 370026 227016
rect 370262 226780 405706 227016
rect 405942 226780 406026 227016
rect 406262 226780 441706 227016
rect 441942 226780 442026 227016
rect 442262 226780 477706 227016
rect 477942 226780 478026 227016
rect 478262 226780 513706 227016
rect 513942 226780 514026 227016
rect 514262 226780 549706 227016
rect 549942 226780 550026 227016
rect 550262 226780 592062 227016
rect 592298 226780 592382 227016
rect 592618 226780 592650 227016
rect -8726 226748 592650 226780
rect -8726 226096 592650 226128
rect -8726 225860 -7734 226096
rect -7498 225860 -7414 226096
rect -7178 225860 8466 226096
rect 8702 225860 8786 226096
rect 9022 225860 44466 226096
rect 44702 225860 44786 226096
rect 45022 225860 80466 226096
rect 80702 225860 80786 226096
rect 81022 225860 116466 226096
rect 116702 225860 116786 226096
rect 117022 225860 152466 226096
rect 152702 225860 152786 226096
rect 153022 225860 188466 226096
rect 188702 225860 188786 226096
rect 189022 225860 224466 226096
rect 224702 225860 224786 226096
rect 225022 225860 260466 226096
rect 260702 225860 260786 226096
rect 261022 225860 296466 226096
rect 296702 225860 296786 226096
rect 297022 225860 332466 226096
rect 332702 225860 332786 226096
rect 333022 225860 368466 226096
rect 368702 225860 368786 226096
rect 369022 225860 404466 226096
rect 404702 225860 404786 226096
rect 405022 225860 440466 226096
rect 440702 225860 440786 226096
rect 441022 225860 476466 226096
rect 476702 225860 476786 226096
rect 477022 225860 512466 226096
rect 512702 225860 512786 226096
rect 513022 225860 548466 226096
rect 548702 225860 548786 226096
rect 549022 225860 591102 226096
rect 591338 225860 591422 226096
rect 591658 225860 592650 226096
rect -8726 225776 592650 225860
rect -8726 225540 -7734 225776
rect -7498 225540 -7414 225776
rect -7178 225540 8466 225776
rect 8702 225540 8786 225776
rect 9022 225540 44466 225776
rect 44702 225540 44786 225776
rect 45022 225540 80466 225776
rect 80702 225540 80786 225776
rect 81022 225540 116466 225776
rect 116702 225540 116786 225776
rect 117022 225540 152466 225776
rect 152702 225540 152786 225776
rect 153022 225540 188466 225776
rect 188702 225540 188786 225776
rect 189022 225540 224466 225776
rect 224702 225540 224786 225776
rect 225022 225540 260466 225776
rect 260702 225540 260786 225776
rect 261022 225540 296466 225776
rect 296702 225540 296786 225776
rect 297022 225540 332466 225776
rect 332702 225540 332786 225776
rect 333022 225540 368466 225776
rect 368702 225540 368786 225776
rect 369022 225540 404466 225776
rect 404702 225540 404786 225776
rect 405022 225540 440466 225776
rect 440702 225540 440786 225776
rect 441022 225540 476466 225776
rect 476702 225540 476786 225776
rect 477022 225540 512466 225776
rect 512702 225540 512786 225776
rect 513022 225540 548466 225776
rect 548702 225540 548786 225776
rect 549022 225540 591102 225776
rect 591338 225540 591422 225776
rect 591658 225540 592650 225776
rect -8726 225508 592650 225540
rect -8726 224856 592650 224888
rect -8726 224620 -6774 224856
rect -6538 224620 -6454 224856
rect -6218 224620 7226 224856
rect 7462 224620 7546 224856
rect 7782 224620 43226 224856
rect 43462 224620 43546 224856
rect 43782 224620 79226 224856
rect 79462 224620 79546 224856
rect 79782 224620 115226 224856
rect 115462 224620 115546 224856
rect 115782 224620 151226 224856
rect 151462 224620 151546 224856
rect 151782 224620 187226 224856
rect 187462 224620 187546 224856
rect 187782 224620 223226 224856
rect 223462 224620 223546 224856
rect 223782 224620 259226 224856
rect 259462 224620 259546 224856
rect 259782 224620 295226 224856
rect 295462 224620 295546 224856
rect 295782 224620 331226 224856
rect 331462 224620 331546 224856
rect 331782 224620 367226 224856
rect 367462 224620 367546 224856
rect 367782 224620 403226 224856
rect 403462 224620 403546 224856
rect 403782 224620 439226 224856
rect 439462 224620 439546 224856
rect 439782 224620 475226 224856
rect 475462 224620 475546 224856
rect 475782 224620 511226 224856
rect 511462 224620 511546 224856
rect 511782 224620 547226 224856
rect 547462 224620 547546 224856
rect 547782 224620 590142 224856
rect 590378 224620 590462 224856
rect 590698 224620 592650 224856
rect -8726 224536 592650 224620
rect -8726 224300 -6774 224536
rect -6538 224300 -6454 224536
rect -6218 224300 7226 224536
rect 7462 224300 7546 224536
rect 7782 224300 43226 224536
rect 43462 224300 43546 224536
rect 43782 224300 79226 224536
rect 79462 224300 79546 224536
rect 79782 224300 115226 224536
rect 115462 224300 115546 224536
rect 115782 224300 151226 224536
rect 151462 224300 151546 224536
rect 151782 224300 187226 224536
rect 187462 224300 187546 224536
rect 187782 224300 223226 224536
rect 223462 224300 223546 224536
rect 223782 224300 259226 224536
rect 259462 224300 259546 224536
rect 259782 224300 295226 224536
rect 295462 224300 295546 224536
rect 295782 224300 331226 224536
rect 331462 224300 331546 224536
rect 331782 224300 367226 224536
rect 367462 224300 367546 224536
rect 367782 224300 403226 224536
rect 403462 224300 403546 224536
rect 403782 224300 439226 224536
rect 439462 224300 439546 224536
rect 439782 224300 475226 224536
rect 475462 224300 475546 224536
rect 475782 224300 511226 224536
rect 511462 224300 511546 224536
rect 511782 224300 547226 224536
rect 547462 224300 547546 224536
rect 547782 224300 590142 224536
rect 590378 224300 590462 224536
rect 590698 224300 592650 224536
rect -8726 224268 592650 224300
rect -8726 223616 592650 223648
rect -8726 223380 -5814 223616
rect -5578 223380 -5494 223616
rect -5258 223380 5986 223616
rect 6222 223380 6306 223616
rect 6542 223380 41986 223616
rect 42222 223380 42306 223616
rect 42542 223380 77986 223616
rect 78222 223380 78306 223616
rect 78542 223380 113986 223616
rect 114222 223380 114306 223616
rect 114542 223380 149986 223616
rect 150222 223380 150306 223616
rect 150542 223380 185986 223616
rect 186222 223380 186306 223616
rect 186542 223380 221986 223616
rect 222222 223380 222306 223616
rect 222542 223380 257986 223616
rect 258222 223380 258306 223616
rect 258542 223380 293986 223616
rect 294222 223380 294306 223616
rect 294542 223380 329986 223616
rect 330222 223380 330306 223616
rect 330542 223380 365986 223616
rect 366222 223380 366306 223616
rect 366542 223380 401986 223616
rect 402222 223380 402306 223616
rect 402542 223380 437986 223616
rect 438222 223380 438306 223616
rect 438542 223380 473986 223616
rect 474222 223380 474306 223616
rect 474542 223380 509986 223616
rect 510222 223380 510306 223616
rect 510542 223380 545986 223616
rect 546222 223380 546306 223616
rect 546542 223380 581986 223616
rect 582222 223380 582306 223616
rect 582542 223380 589182 223616
rect 589418 223380 589502 223616
rect 589738 223380 592650 223616
rect -8726 223296 592650 223380
rect -8726 223060 -5814 223296
rect -5578 223060 -5494 223296
rect -5258 223060 5986 223296
rect 6222 223060 6306 223296
rect 6542 223060 41986 223296
rect 42222 223060 42306 223296
rect 42542 223060 77986 223296
rect 78222 223060 78306 223296
rect 78542 223060 113986 223296
rect 114222 223060 114306 223296
rect 114542 223060 149986 223296
rect 150222 223060 150306 223296
rect 150542 223060 185986 223296
rect 186222 223060 186306 223296
rect 186542 223060 221986 223296
rect 222222 223060 222306 223296
rect 222542 223060 257986 223296
rect 258222 223060 258306 223296
rect 258542 223060 293986 223296
rect 294222 223060 294306 223296
rect 294542 223060 329986 223296
rect 330222 223060 330306 223296
rect 330542 223060 365986 223296
rect 366222 223060 366306 223296
rect 366542 223060 401986 223296
rect 402222 223060 402306 223296
rect 402542 223060 437986 223296
rect 438222 223060 438306 223296
rect 438542 223060 473986 223296
rect 474222 223060 474306 223296
rect 474542 223060 509986 223296
rect 510222 223060 510306 223296
rect 510542 223060 545986 223296
rect 546222 223060 546306 223296
rect 546542 223060 581986 223296
rect 582222 223060 582306 223296
rect 582542 223060 589182 223296
rect 589418 223060 589502 223296
rect 589738 223060 592650 223296
rect -8726 223028 592650 223060
rect -8726 222376 592650 222408
rect -8726 222140 -4854 222376
rect -4618 222140 -4534 222376
rect -4298 222140 4746 222376
rect 4982 222140 5066 222376
rect 5302 222140 40746 222376
rect 40982 222140 41066 222376
rect 41302 222140 76746 222376
rect 76982 222140 77066 222376
rect 77302 222140 112746 222376
rect 112982 222140 113066 222376
rect 113302 222140 148746 222376
rect 148982 222140 149066 222376
rect 149302 222140 184746 222376
rect 184982 222140 185066 222376
rect 185302 222140 220746 222376
rect 220982 222140 221066 222376
rect 221302 222140 256746 222376
rect 256982 222140 257066 222376
rect 257302 222140 292746 222376
rect 292982 222140 293066 222376
rect 293302 222140 328746 222376
rect 328982 222140 329066 222376
rect 329302 222140 364746 222376
rect 364982 222140 365066 222376
rect 365302 222140 400746 222376
rect 400982 222140 401066 222376
rect 401302 222140 436746 222376
rect 436982 222140 437066 222376
rect 437302 222140 472746 222376
rect 472982 222140 473066 222376
rect 473302 222140 508746 222376
rect 508982 222140 509066 222376
rect 509302 222140 544746 222376
rect 544982 222140 545066 222376
rect 545302 222140 580746 222376
rect 580982 222140 581066 222376
rect 581302 222140 588222 222376
rect 588458 222140 588542 222376
rect 588778 222140 592650 222376
rect -8726 222056 592650 222140
rect -8726 221820 -4854 222056
rect -4618 221820 -4534 222056
rect -4298 221820 4746 222056
rect 4982 221820 5066 222056
rect 5302 221820 40746 222056
rect 40982 221820 41066 222056
rect 41302 221820 76746 222056
rect 76982 221820 77066 222056
rect 77302 221820 112746 222056
rect 112982 221820 113066 222056
rect 113302 221820 148746 222056
rect 148982 221820 149066 222056
rect 149302 221820 184746 222056
rect 184982 221820 185066 222056
rect 185302 221820 220746 222056
rect 220982 221820 221066 222056
rect 221302 221820 256746 222056
rect 256982 221820 257066 222056
rect 257302 221820 292746 222056
rect 292982 221820 293066 222056
rect 293302 221820 328746 222056
rect 328982 221820 329066 222056
rect 329302 221820 364746 222056
rect 364982 221820 365066 222056
rect 365302 221820 400746 222056
rect 400982 221820 401066 222056
rect 401302 221820 436746 222056
rect 436982 221820 437066 222056
rect 437302 221820 472746 222056
rect 472982 221820 473066 222056
rect 473302 221820 508746 222056
rect 508982 221820 509066 222056
rect 509302 221820 544746 222056
rect 544982 221820 545066 222056
rect 545302 221820 580746 222056
rect 580982 221820 581066 222056
rect 581302 221820 588222 222056
rect 588458 221820 588542 222056
rect 588778 221820 592650 222056
rect -8726 221788 592650 221820
rect -8726 221136 592650 221168
rect -8726 220900 -3894 221136
rect -3658 220900 -3574 221136
rect -3338 220900 3506 221136
rect 3742 220900 3826 221136
rect 4062 220900 39506 221136
rect 39742 220900 39826 221136
rect 40062 220900 75506 221136
rect 75742 220900 75826 221136
rect 76062 220900 111506 221136
rect 111742 220900 111826 221136
rect 112062 220900 147506 221136
rect 147742 220900 147826 221136
rect 148062 220900 183506 221136
rect 183742 220900 183826 221136
rect 184062 220900 219506 221136
rect 219742 220900 219826 221136
rect 220062 220900 255506 221136
rect 255742 220900 255826 221136
rect 256062 220900 291506 221136
rect 291742 220900 291826 221136
rect 292062 220900 327506 221136
rect 327742 220900 327826 221136
rect 328062 220900 363506 221136
rect 363742 220900 363826 221136
rect 364062 220900 399506 221136
rect 399742 220900 399826 221136
rect 400062 220900 435506 221136
rect 435742 220900 435826 221136
rect 436062 220900 471506 221136
rect 471742 220900 471826 221136
rect 472062 220900 507506 221136
rect 507742 220900 507826 221136
rect 508062 220900 543506 221136
rect 543742 220900 543826 221136
rect 544062 220900 579506 221136
rect 579742 220900 579826 221136
rect 580062 220900 587262 221136
rect 587498 220900 587582 221136
rect 587818 220900 592650 221136
rect -8726 220816 592650 220900
rect -8726 220580 -3894 220816
rect -3658 220580 -3574 220816
rect -3338 220580 3506 220816
rect 3742 220580 3826 220816
rect 4062 220580 39506 220816
rect 39742 220580 39826 220816
rect 40062 220580 75506 220816
rect 75742 220580 75826 220816
rect 76062 220580 111506 220816
rect 111742 220580 111826 220816
rect 112062 220580 147506 220816
rect 147742 220580 147826 220816
rect 148062 220580 183506 220816
rect 183742 220580 183826 220816
rect 184062 220580 219506 220816
rect 219742 220580 219826 220816
rect 220062 220580 255506 220816
rect 255742 220580 255826 220816
rect 256062 220580 291506 220816
rect 291742 220580 291826 220816
rect 292062 220580 327506 220816
rect 327742 220580 327826 220816
rect 328062 220580 363506 220816
rect 363742 220580 363826 220816
rect 364062 220580 399506 220816
rect 399742 220580 399826 220816
rect 400062 220580 435506 220816
rect 435742 220580 435826 220816
rect 436062 220580 471506 220816
rect 471742 220580 471826 220816
rect 472062 220580 507506 220816
rect 507742 220580 507826 220816
rect 508062 220580 543506 220816
rect 543742 220580 543826 220816
rect 544062 220580 579506 220816
rect 579742 220580 579826 220816
rect 580062 220580 587262 220816
rect 587498 220580 587582 220816
rect 587818 220580 592650 220816
rect -8726 220548 592650 220580
rect -8726 219896 592650 219928
rect -8726 219660 -2934 219896
rect -2698 219660 -2614 219896
rect -2378 219660 2266 219896
rect 2502 219660 2586 219896
rect 2822 219660 38266 219896
rect 38502 219660 38586 219896
rect 38822 219660 74266 219896
rect 74502 219660 74586 219896
rect 74822 219660 110266 219896
rect 110502 219660 110586 219896
rect 110822 219660 146266 219896
rect 146502 219660 146586 219896
rect 146822 219660 182266 219896
rect 182502 219660 182586 219896
rect 182822 219660 218266 219896
rect 218502 219660 218586 219896
rect 218822 219660 254266 219896
rect 254502 219660 254586 219896
rect 254822 219660 290266 219896
rect 290502 219660 290586 219896
rect 290822 219660 326266 219896
rect 326502 219660 326586 219896
rect 326822 219660 362266 219896
rect 362502 219660 362586 219896
rect 362822 219660 398266 219896
rect 398502 219660 398586 219896
rect 398822 219660 434266 219896
rect 434502 219660 434586 219896
rect 434822 219660 470266 219896
rect 470502 219660 470586 219896
rect 470822 219660 506266 219896
rect 506502 219660 506586 219896
rect 506822 219660 542266 219896
rect 542502 219660 542586 219896
rect 542822 219660 578266 219896
rect 578502 219660 578586 219896
rect 578822 219660 586302 219896
rect 586538 219660 586622 219896
rect 586858 219660 592650 219896
rect -8726 219576 592650 219660
rect -8726 219340 -2934 219576
rect -2698 219340 -2614 219576
rect -2378 219340 2266 219576
rect 2502 219340 2586 219576
rect 2822 219340 38266 219576
rect 38502 219340 38586 219576
rect 38822 219340 74266 219576
rect 74502 219340 74586 219576
rect 74822 219340 110266 219576
rect 110502 219340 110586 219576
rect 110822 219340 146266 219576
rect 146502 219340 146586 219576
rect 146822 219340 182266 219576
rect 182502 219340 182586 219576
rect 182822 219340 218266 219576
rect 218502 219340 218586 219576
rect 218822 219340 254266 219576
rect 254502 219340 254586 219576
rect 254822 219340 290266 219576
rect 290502 219340 290586 219576
rect 290822 219340 326266 219576
rect 326502 219340 326586 219576
rect 326822 219340 362266 219576
rect 362502 219340 362586 219576
rect 362822 219340 398266 219576
rect 398502 219340 398586 219576
rect 398822 219340 434266 219576
rect 434502 219340 434586 219576
rect 434822 219340 470266 219576
rect 470502 219340 470586 219576
rect 470822 219340 506266 219576
rect 506502 219340 506586 219576
rect 506822 219340 542266 219576
rect 542502 219340 542586 219576
rect 542822 219340 578266 219576
rect 578502 219340 578586 219576
rect 578822 219340 586302 219576
rect 586538 219340 586622 219576
rect 586858 219340 592650 219576
rect -8726 219308 592650 219340
rect -8726 218656 592650 218688
rect -8726 218420 -1974 218656
rect -1738 218420 -1654 218656
rect -1418 218420 1026 218656
rect 1262 218420 1346 218656
rect 1582 218420 37026 218656
rect 37262 218420 37346 218656
rect 37582 218420 73026 218656
rect 73262 218420 73346 218656
rect 73582 218420 109026 218656
rect 109262 218420 109346 218656
rect 109582 218420 145026 218656
rect 145262 218420 145346 218656
rect 145582 218420 181026 218656
rect 181262 218420 181346 218656
rect 181582 218420 217026 218656
rect 217262 218420 217346 218656
rect 217582 218420 253026 218656
rect 253262 218420 253346 218656
rect 253582 218420 289026 218656
rect 289262 218420 289346 218656
rect 289582 218420 325026 218656
rect 325262 218420 325346 218656
rect 325582 218420 361026 218656
rect 361262 218420 361346 218656
rect 361582 218420 397026 218656
rect 397262 218420 397346 218656
rect 397582 218420 433026 218656
rect 433262 218420 433346 218656
rect 433582 218420 469026 218656
rect 469262 218420 469346 218656
rect 469582 218420 505026 218656
rect 505262 218420 505346 218656
rect 505582 218420 541026 218656
rect 541262 218420 541346 218656
rect 541582 218420 577026 218656
rect 577262 218420 577346 218656
rect 577582 218420 585342 218656
rect 585578 218420 585662 218656
rect 585898 218420 592650 218656
rect -8726 218336 592650 218420
rect -8726 218100 -1974 218336
rect -1738 218100 -1654 218336
rect -1418 218100 1026 218336
rect 1262 218100 1346 218336
rect 1582 218100 37026 218336
rect 37262 218100 37346 218336
rect 37582 218100 73026 218336
rect 73262 218100 73346 218336
rect 73582 218100 109026 218336
rect 109262 218100 109346 218336
rect 109582 218100 145026 218336
rect 145262 218100 145346 218336
rect 145582 218100 181026 218336
rect 181262 218100 181346 218336
rect 181582 218100 217026 218336
rect 217262 218100 217346 218336
rect 217582 218100 253026 218336
rect 253262 218100 253346 218336
rect 253582 218100 289026 218336
rect 289262 218100 289346 218336
rect 289582 218100 325026 218336
rect 325262 218100 325346 218336
rect 325582 218100 361026 218336
rect 361262 218100 361346 218336
rect 361582 218100 397026 218336
rect 397262 218100 397346 218336
rect 397582 218100 433026 218336
rect 433262 218100 433346 218336
rect 433582 218100 469026 218336
rect 469262 218100 469346 218336
rect 469582 218100 505026 218336
rect 505262 218100 505346 218336
rect 505582 218100 541026 218336
rect 541262 218100 541346 218336
rect 541582 218100 577026 218336
rect 577262 218100 577346 218336
rect 577582 218100 585342 218336
rect 585578 218100 585662 218336
rect 585898 218100 592650 218336
rect -8726 218068 592650 218100
rect -8726 191336 592650 191368
rect -8726 191100 -8694 191336
rect -8458 191100 -8374 191336
rect -8138 191100 9706 191336
rect 9942 191100 10026 191336
rect 10262 191100 45706 191336
rect 45942 191100 46026 191336
rect 46262 191100 81706 191336
rect 81942 191100 82026 191336
rect 82262 191100 117706 191336
rect 117942 191100 118026 191336
rect 118262 191100 153706 191336
rect 153942 191100 154026 191336
rect 154262 191100 189706 191336
rect 189942 191100 190026 191336
rect 190262 191100 225706 191336
rect 225942 191100 226026 191336
rect 226262 191100 261706 191336
rect 261942 191100 262026 191336
rect 262262 191100 297706 191336
rect 297942 191100 298026 191336
rect 298262 191100 333706 191336
rect 333942 191100 334026 191336
rect 334262 191100 369706 191336
rect 369942 191100 370026 191336
rect 370262 191100 405706 191336
rect 405942 191100 406026 191336
rect 406262 191100 441706 191336
rect 441942 191100 442026 191336
rect 442262 191100 477706 191336
rect 477942 191100 478026 191336
rect 478262 191100 513706 191336
rect 513942 191100 514026 191336
rect 514262 191100 549706 191336
rect 549942 191100 550026 191336
rect 550262 191100 592062 191336
rect 592298 191100 592382 191336
rect 592618 191100 592650 191336
rect -8726 191016 592650 191100
rect -8726 190780 -8694 191016
rect -8458 190780 -8374 191016
rect -8138 190780 9706 191016
rect 9942 190780 10026 191016
rect 10262 190780 45706 191016
rect 45942 190780 46026 191016
rect 46262 190780 81706 191016
rect 81942 190780 82026 191016
rect 82262 190780 117706 191016
rect 117942 190780 118026 191016
rect 118262 190780 153706 191016
rect 153942 190780 154026 191016
rect 154262 190780 189706 191016
rect 189942 190780 190026 191016
rect 190262 190780 225706 191016
rect 225942 190780 226026 191016
rect 226262 190780 261706 191016
rect 261942 190780 262026 191016
rect 262262 190780 297706 191016
rect 297942 190780 298026 191016
rect 298262 190780 333706 191016
rect 333942 190780 334026 191016
rect 334262 190780 369706 191016
rect 369942 190780 370026 191016
rect 370262 190780 405706 191016
rect 405942 190780 406026 191016
rect 406262 190780 441706 191016
rect 441942 190780 442026 191016
rect 442262 190780 477706 191016
rect 477942 190780 478026 191016
rect 478262 190780 513706 191016
rect 513942 190780 514026 191016
rect 514262 190780 549706 191016
rect 549942 190780 550026 191016
rect 550262 190780 592062 191016
rect 592298 190780 592382 191016
rect 592618 190780 592650 191016
rect -8726 190748 592650 190780
rect -8726 190096 592650 190128
rect -8726 189860 -7734 190096
rect -7498 189860 -7414 190096
rect -7178 189860 8466 190096
rect 8702 189860 8786 190096
rect 9022 189860 44466 190096
rect 44702 189860 44786 190096
rect 45022 189860 80466 190096
rect 80702 189860 80786 190096
rect 81022 189860 116466 190096
rect 116702 189860 116786 190096
rect 117022 189860 152466 190096
rect 152702 189860 152786 190096
rect 153022 189860 188466 190096
rect 188702 189860 188786 190096
rect 189022 189860 224466 190096
rect 224702 189860 224786 190096
rect 225022 189860 260466 190096
rect 260702 189860 260786 190096
rect 261022 189860 296466 190096
rect 296702 189860 296786 190096
rect 297022 189860 332466 190096
rect 332702 189860 332786 190096
rect 333022 189860 368466 190096
rect 368702 189860 368786 190096
rect 369022 189860 404466 190096
rect 404702 189860 404786 190096
rect 405022 189860 440466 190096
rect 440702 189860 440786 190096
rect 441022 189860 476466 190096
rect 476702 189860 476786 190096
rect 477022 189860 512466 190096
rect 512702 189860 512786 190096
rect 513022 189860 548466 190096
rect 548702 189860 548786 190096
rect 549022 189860 591102 190096
rect 591338 189860 591422 190096
rect 591658 189860 592650 190096
rect -8726 189776 592650 189860
rect -8726 189540 -7734 189776
rect -7498 189540 -7414 189776
rect -7178 189540 8466 189776
rect 8702 189540 8786 189776
rect 9022 189540 44466 189776
rect 44702 189540 44786 189776
rect 45022 189540 80466 189776
rect 80702 189540 80786 189776
rect 81022 189540 116466 189776
rect 116702 189540 116786 189776
rect 117022 189540 152466 189776
rect 152702 189540 152786 189776
rect 153022 189540 188466 189776
rect 188702 189540 188786 189776
rect 189022 189540 224466 189776
rect 224702 189540 224786 189776
rect 225022 189540 260466 189776
rect 260702 189540 260786 189776
rect 261022 189540 296466 189776
rect 296702 189540 296786 189776
rect 297022 189540 332466 189776
rect 332702 189540 332786 189776
rect 333022 189540 368466 189776
rect 368702 189540 368786 189776
rect 369022 189540 404466 189776
rect 404702 189540 404786 189776
rect 405022 189540 440466 189776
rect 440702 189540 440786 189776
rect 441022 189540 476466 189776
rect 476702 189540 476786 189776
rect 477022 189540 512466 189776
rect 512702 189540 512786 189776
rect 513022 189540 548466 189776
rect 548702 189540 548786 189776
rect 549022 189540 591102 189776
rect 591338 189540 591422 189776
rect 591658 189540 592650 189776
rect -8726 189508 592650 189540
rect -8726 188856 592650 188888
rect -8726 188620 -6774 188856
rect -6538 188620 -6454 188856
rect -6218 188620 7226 188856
rect 7462 188620 7546 188856
rect 7782 188620 43226 188856
rect 43462 188620 43546 188856
rect 43782 188620 79226 188856
rect 79462 188620 79546 188856
rect 79782 188620 115226 188856
rect 115462 188620 115546 188856
rect 115782 188620 151226 188856
rect 151462 188620 151546 188856
rect 151782 188620 187226 188856
rect 187462 188620 187546 188856
rect 187782 188620 223226 188856
rect 223462 188620 223546 188856
rect 223782 188620 259226 188856
rect 259462 188620 259546 188856
rect 259782 188620 295226 188856
rect 295462 188620 295546 188856
rect 295782 188620 331226 188856
rect 331462 188620 331546 188856
rect 331782 188620 367226 188856
rect 367462 188620 367546 188856
rect 367782 188620 403226 188856
rect 403462 188620 403546 188856
rect 403782 188620 439226 188856
rect 439462 188620 439546 188856
rect 439782 188620 475226 188856
rect 475462 188620 475546 188856
rect 475782 188620 511226 188856
rect 511462 188620 511546 188856
rect 511782 188620 547226 188856
rect 547462 188620 547546 188856
rect 547782 188620 590142 188856
rect 590378 188620 590462 188856
rect 590698 188620 592650 188856
rect -8726 188536 592650 188620
rect -8726 188300 -6774 188536
rect -6538 188300 -6454 188536
rect -6218 188300 7226 188536
rect 7462 188300 7546 188536
rect 7782 188300 43226 188536
rect 43462 188300 43546 188536
rect 43782 188300 79226 188536
rect 79462 188300 79546 188536
rect 79782 188300 115226 188536
rect 115462 188300 115546 188536
rect 115782 188300 151226 188536
rect 151462 188300 151546 188536
rect 151782 188300 187226 188536
rect 187462 188300 187546 188536
rect 187782 188300 223226 188536
rect 223462 188300 223546 188536
rect 223782 188300 259226 188536
rect 259462 188300 259546 188536
rect 259782 188300 295226 188536
rect 295462 188300 295546 188536
rect 295782 188300 331226 188536
rect 331462 188300 331546 188536
rect 331782 188300 367226 188536
rect 367462 188300 367546 188536
rect 367782 188300 403226 188536
rect 403462 188300 403546 188536
rect 403782 188300 439226 188536
rect 439462 188300 439546 188536
rect 439782 188300 475226 188536
rect 475462 188300 475546 188536
rect 475782 188300 511226 188536
rect 511462 188300 511546 188536
rect 511782 188300 547226 188536
rect 547462 188300 547546 188536
rect 547782 188300 590142 188536
rect 590378 188300 590462 188536
rect 590698 188300 592650 188536
rect -8726 188268 592650 188300
rect -8726 187616 592650 187648
rect -8726 187380 -5814 187616
rect -5578 187380 -5494 187616
rect -5258 187380 5986 187616
rect 6222 187380 6306 187616
rect 6542 187380 41986 187616
rect 42222 187380 42306 187616
rect 42542 187380 77986 187616
rect 78222 187380 78306 187616
rect 78542 187380 113986 187616
rect 114222 187380 114306 187616
rect 114542 187380 149986 187616
rect 150222 187380 150306 187616
rect 150542 187380 185986 187616
rect 186222 187380 186306 187616
rect 186542 187380 221986 187616
rect 222222 187380 222306 187616
rect 222542 187380 257986 187616
rect 258222 187380 258306 187616
rect 258542 187380 293986 187616
rect 294222 187380 294306 187616
rect 294542 187380 329986 187616
rect 330222 187380 330306 187616
rect 330542 187380 365986 187616
rect 366222 187380 366306 187616
rect 366542 187380 401986 187616
rect 402222 187380 402306 187616
rect 402542 187380 437986 187616
rect 438222 187380 438306 187616
rect 438542 187380 473986 187616
rect 474222 187380 474306 187616
rect 474542 187380 509986 187616
rect 510222 187380 510306 187616
rect 510542 187380 545986 187616
rect 546222 187380 546306 187616
rect 546542 187380 581986 187616
rect 582222 187380 582306 187616
rect 582542 187380 589182 187616
rect 589418 187380 589502 187616
rect 589738 187380 592650 187616
rect -8726 187296 592650 187380
rect -8726 187060 -5814 187296
rect -5578 187060 -5494 187296
rect -5258 187060 5986 187296
rect 6222 187060 6306 187296
rect 6542 187060 41986 187296
rect 42222 187060 42306 187296
rect 42542 187060 77986 187296
rect 78222 187060 78306 187296
rect 78542 187060 113986 187296
rect 114222 187060 114306 187296
rect 114542 187060 149986 187296
rect 150222 187060 150306 187296
rect 150542 187060 185986 187296
rect 186222 187060 186306 187296
rect 186542 187060 221986 187296
rect 222222 187060 222306 187296
rect 222542 187060 257986 187296
rect 258222 187060 258306 187296
rect 258542 187060 293986 187296
rect 294222 187060 294306 187296
rect 294542 187060 329986 187296
rect 330222 187060 330306 187296
rect 330542 187060 365986 187296
rect 366222 187060 366306 187296
rect 366542 187060 401986 187296
rect 402222 187060 402306 187296
rect 402542 187060 437986 187296
rect 438222 187060 438306 187296
rect 438542 187060 473986 187296
rect 474222 187060 474306 187296
rect 474542 187060 509986 187296
rect 510222 187060 510306 187296
rect 510542 187060 545986 187296
rect 546222 187060 546306 187296
rect 546542 187060 581986 187296
rect 582222 187060 582306 187296
rect 582542 187060 589182 187296
rect 589418 187060 589502 187296
rect 589738 187060 592650 187296
rect -8726 187028 592650 187060
rect -8726 186376 592650 186408
rect -8726 186140 -4854 186376
rect -4618 186140 -4534 186376
rect -4298 186140 4746 186376
rect 4982 186140 5066 186376
rect 5302 186140 40746 186376
rect 40982 186140 41066 186376
rect 41302 186140 76746 186376
rect 76982 186140 77066 186376
rect 77302 186140 112746 186376
rect 112982 186140 113066 186376
rect 113302 186140 148746 186376
rect 148982 186140 149066 186376
rect 149302 186140 184746 186376
rect 184982 186140 185066 186376
rect 185302 186140 220746 186376
rect 220982 186140 221066 186376
rect 221302 186140 256746 186376
rect 256982 186140 257066 186376
rect 257302 186140 292746 186376
rect 292982 186140 293066 186376
rect 293302 186140 328746 186376
rect 328982 186140 329066 186376
rect 329302 186140 364746 186376
rect 364982 186140 365066 186376
rect 365302 186140 400746 186376
rect 400982 186140 401066 186376
rect 401302 186140 436746 186376
rect 436982 186140 437066 186376
rect 437302 186140 472746 186376
rect 472982 186140 473066 186376
rect 473302 186140 508746 186376
rect 508982 186140 509066 186376
rect 509302 186140 544746 186376
rect 544982 186140 545066 186376
rect 545302 186140 580746 186376
rect 580982 186140 581066 186376
rect 581302 186140 588222 186376
rect 588458 186140 588542 186376
rect 588778 186140 592650 186376
rect -8726 186056 592650 186140
rect -8726 185820 -4854 186056
rect -4618 185820 -4534 186056
rect -4298 185820 4746 186056
rect 4982 185820 5066 186056
rect 5302 185820 40746 186056
rect 40982 185820 41066 186056
rect 41302 185820 76746 186056
rect 76982 185820 77066 186056
rect 77302 185820 112746 186056
rect 112982 185820 113066 186056
rect 113302 185820 148746 186056
rect 148982 185820 149066 186056
rect 149302 185820 184746 186056
rect 184982 185820 185066 186056
rect 185302 185820 220746 186056
rect 220982 185820 221066 186056
rect 221302 185820 256746 186056
rect 256982 185820 257066 186056
rect 257302 185820 292746 186056
rect 292982 185820 293066 186056
rect 293302 185820 328746 186056
rect 328982 185820 329066 186056
rect 329302 185820 364746 186056
rect 364982 185820 365066 186056
rect 365302 185820 400746 186056
rect 400982 185820 401066 186056
rect 401302 185820 436746 186056
rect 436982 185820 437066 186056
rect 437302 185820 472746 186056
rect 472982 185820 473066 186056
rect 473302 185820 508746 186056
rect 508982 185820 509066 186056
rect 509302 185820 544746 186056
rect 544982 185820 545066 186056
rect 545302 185820 580746 186056
rect 580982 185820 581066 186056
rect 581302 185820 588222 186056
rect 588458 185820 588542 186056
rect 588778 185820 592650 186056
rect -8726 185788 592650 185820
rect -8726 185136 592650 185168
rect -8726 184900 -3894 185136
rect -3658 184900 -3574 185136
rect -3338 184900 3506 185136
rect 3742 184900 3826 185136
rect 4062 184900 39506 185136
rect 39742 184900 39826 185136
rect 40062 184900 75506 185136
rect 75742 184900 75826 185136
rect 76062 184900 111506 185136
rect 111742 184900 111826 185136
rect 112062 184900 147506 185136
rect 147742 184900 147826 185136
rect 148062 184900 183506 185136
rect 183742 184900 183826 185136
rect 184062 184900 219506 185136
rect 219742 184900 219826 185136
rect 220062 184900 255506 185136
rect 255742 184900 255826 185136
rect 256062 184900 291506 185136
rect 291742 184900 291826 185136
rect 292062 184900 327506 185136
rect 327742 184900 327826 185136
rect 328062 184900 363506 185136
rect 363742 184900 363826 185136
rect 364062 184900 399506 185136
rect 399742 184900 399826 185136
rect 400062 184900 435506 185136
rect 435742 184900 435826 185136
rect 436062 184900 471506 185136
rect 471742 184900 471826 185136
rect 472062 184900 507506 185136
rect 507742 184900 507826 185136
rect 508062 184900 543506 185136
rect 543742 184900 543826 185136
rect 544062 184900 579506 185136
rect 579742 184900 579826 185136
rect 580062 184900 587262 185136
rect 587498 184900 587582 185136
rect 587818 184900 592650 185136
rect -8726 184816 592650 184900
rect -8726 184580 -3894 184816
rect -3658 184580 -3574 184816
rect -3338 184580 3506 184816
rect 3742 184580 3826 184816
rect 4062 184580 39506 184816
rect 39742 184580 39826 184816
rect 40062 184580 75506 184816
rect 75742 184580 75826 184816
rect 76062 184580 111506 184816
rect 111742 184580 111826 184816
rect 112062 184580 147506 184816
rect 147742 184580 147826 184816
rect 148062 184580 183506 184816
rect 183742 184580 183826 184816
rect 184062 184580 219506 184816
rect 219742 184580 219826 184816
rect 220062 184580 255506 184816
rect 255742 184580 255826 184816
rect 256062 184580 291506 184816
rect 291742 184580 291826 184816
rect 292062 184580 327506 184816
rect 327742 184580 327826 184816
rect 328062 184580 363506 184816
rect 363742 184580 363826 184816
rect 364062 184580 399506 184816
rect 399742 184580 399826 184816
rect 400062 184580 435506 184816
rect 435742 184580 435826 184816
rect 436062 184580 471506 184816
rect 471742 184580 471826 184816
rect 472062 184580 507506 184816
rect 507742 184580 507826 184816
rect 508062 184580 543506 184816
rect 543742 184580 543826 184816
rect 544062 184580 579506 184816
rect 579742 184580 579826 184816
rect 580062 184580 587262 184816
rect 587498 184580 587582 184816
rect 587818 184580 592650 184816
rect -8726 184548 592650 184580
rect -8726 183896 592650 183928
rect -8726 183660 -2934 183896
rect -2698 183660 -2614 183896
rect -2378 183660 2266 183896
rect 2502 183660 2586 183896
rect 2822 183660 38266 183896
rect 38502 183660 38586 183896
rect 38822 183660 74266 183896
rect 74502 183660 74586 183896
rect 74822 183660 110266 183896
rect 110502 183660 110586 183896
rect 110822 183660 146266 183896
rect 146502 183660 146586 183896
rect 146822 183660 182266 183896
rect 182502 183660 182586 183896
rect 182822 183660 218266 183896
rect 218502 183660 218586 183896
rect 218822 183660 254266 183896
rect 254502 183660 254586 183896
rect 254822 183660 290266 183896
rect 290502 183660 290586 183896
rect 290822 183660 326266 183896
rect 326502 183660 326586 183896
rect 326822 183660 362266 183896
rect 362502 183660 362586 183896
rect 362822 183660 398266 183896
rect 398502 183660 398586 183896
rect 398822 183660 434266 183896
rect 434502 183660 434586 183896
rect 434822 183660 470266 183896
rect 470502 183660 470586 183896
rect 470822 183660 506266 183896
rect 506502 183660 506586 183896
rect 506822 183660 542266 183896
rect 542502 183660 542586 183896
rect 542822 183660 578266 183896
rect 578502 183660 578586 183896
rect 578822 183660 586302 183896
rect 586538 183660 586622 183896
rect 586858 183660 592650 183896
rect -8726 183576 592650 183660
rect -8726 183340 -2934 183576
rect -2698 183340 -2614 183576
rect -2378 183340 2266 183576
rect 2502 183340 2586 183576
rect 2822 183340 38266 183576
rect 38502 183340 38586 183576
rect 38822 183340 74266 183576
rect 74502 183340 74586 183576
rect 74822 183340 110266 183576
rect 110502 183340 110586 183576
rect 110822 183340 146266 183576
rect 146502 183340 146586 183576
rect 146822 183340 182266 183576
rect 182502 183340 182586 183576
rect 182822 183340 218266 183576
rect 218502 183340 218586 183576
rect 218822 183340 254266 183576
rect 254502 183340 254586 183576
rect 254822 183340 290266 183576
rect 290502 183340 290586 183576
rect 290822 183340 326266 183576
rect 326502 183340 326586 183576
rect 326822 183340 362266 183576
rect 362502 183340 362586 183576
rect 362822 183340 398266 183576
rect 398502 183340 398586 183576
rect 398822 183340 434266 183576
rect 434502 183340 434586 183576
rect 434822 183340 470266 183576
rect 470502 183340 470586 183576
rect 470822 183340 506266 183576
rect 506502 183340 506586 183576
rect 506822 183340 542266 183576
rect 542502 183340 542586 183576
rect 542822 183340 578266 183576
rect 578502 183340 578586 183576
rect 578822 183340 586302 183576
rect 586538 183340 586622 183576
rect 586858 183340 592650 183576
rect -8726 183308 592650 183340
rect -8726 182656 592650 182688
rect -8726 182420 -1974 182656
rect -1738 182420 -1654 182656
rect -1418 182420 1026 182656
rect 1262 182420 1346 182656
rect 1582 182420 37026 182656
rect 37262 182420 37346 182656
rect 37582 182420 73026 182656
rect 73262 182420 73346 182656
rect 73582 182420 109026 182656
rect 109262 182420 109346 182656
rect 109582 182420 145026 182656
rect 145262 182420 145346 182656
rect 145582 182420 181026 182656
rect 181262 182420 181346 182656
rect 181582 182420 217026 182656
rect 217262 182420 217346 182656
rect 217582 182420 253026 182656
rect 253262 182420 253346 182656
rect 253582 182420 289026 182656
rect 289262 182420 289346 182656
rect 289582 182420 325026 182656
rect 325262 182420 325346 182656
rect 325582 182420 361026 182656
rect 361262 182420 361346 182656
rect 361582 182420 397026 182656
rect 397262 182420 397346 182656
rect 397582 182420 433026 182656
rect 433262 182420 433346 182656
rect 433582 182420 469026 182656
rect 469262 182420 469346 182656
rect 469582 182420 505026 182656
rect 505262 182420 505346 182656
rect 505582 182420 541026 182656
rect 541262 182420 541346 182656
rect 541582 182420 577026 182656
rect 577262 182420 577346 182656
rect 577582 182420 585342 182656
rect 585578 182420 585662 182656
rect 585898 182420 592650 182656
rect -8726 182336 592650 182420
rect -8726 182100 -1974 182336
rect -1738 182100 -1654 182336
rect -1418 182100 1026 182336
rect 1262 182100 1346 182336
rect 1582 182100 37026 182336
rect 37262 182100 37346 182336
rect 37582 182100 73026 182336
rect 73262 182100 73346 182336
rect 73582 182100 109026 182336
rect 109262 182100 109346 182336
rect 109582 182100 145026 182336
rect 145262 182100 145346 182336
rect 145582 182100 181026 182336
rect 181262 182100 181346 182336
rect 181582 182100 217026 182336
rect 217262 182100 217346 182336
rect 217582 182100 253026 182336
rect 253262 182100 253346 182336
rect 253582 182100 289026 182336
rect 289262 182100 289346 182336
rect 289582 182100 325026 182336
rect 325262 182100 325346 182336
rect 325582 182100 361026 182336
rect 361262 182100 361346 182336
rect 361582 182100 397026 182336
rect 397262 182100 397346 182336
rect 397582 182100 433026 182336
rect 433262 182100 433346 182336
rect 433582 182100 469026 182336
rect 469262 182100 469346 182336
rect 469582 182100 505026 182336
rect 505262 182100 505346 182336
rect 505582 182100 541026 182336
rect 541262 182100 541346 182336
rect 541582 182100 577026 182336
rect 577262 182100 577346 182336
rect 577582 182100 585342 182336
rect 585578 182100 585662 182336
rect 585898 182100 592650 182336
rect -8726 182068 592650 182100
rect -8726 155336 592650 155368
rect -8726 155100 -8694 155336
rect -8458 155100 -8374 155336
rect -8138 155100 9706 155336
rect 9942 155100 10026 155336
rect 10262 155100 45706 155336
rect 45942 155100 46026 155336
rect 46262 155100 81706 155336
rect 81942 155100 82026 155336
rect 82262 155100 117706 155336
rect 117942 155100 118026 155336
rect 118262 155100 153706 155336
rect 153942 155100 154026 155336
rect 154262 155100 189706 155336
rect 189942 155100 190026 155336
rect 190262 155100 225706 155336
rect 225942 155100 226026 155336
rect 226262 155100 261706 155336
rect 261942 155100 262026 155336
rect 262262 155100 297706 155336
rect 297942 155100 298026 155336
rect 298262 155100 333706 155336
rect 333942 155100 334026 155336
rect 334262 155100 369706 155336
rect 369942 155100 370026 155336
rect 370262 155100 405706 155336
rect 405942 155100 406026 155336
rect 406262 155100 441706 155336
rect 441942 155100 442026 155336
rect 442262 155100 477706 155336
rect 477942 155100 478026 155336
rect 478262 155100 513706 155336
rect 513942 155100 514026 155336
rect 514262 155100 549706 155336
rect 549942 155100 550026 155336
rect 550262 155100 592062 155336
rect 592298 155100 592382 155336
rect 592618 155100 592650 155336
rect -8726 155016 592650 155100
rect -8726 154780 -8694 155016
rect -8458 154780 -8374 155016
rect -8138 154780 9706 155016
rect 9942 154780 10026 155016
rect 10262 154780 45706 155016
rect 45942 154780 46026 155016
rect 46262 154780 81706 155016
rect 81942 154780 82026 155016
rect 82262 154780 117706 155016
rect 117942 154780 118026 155016
rect 118262 154780 153706 155016
rect 153942 154780 154026 155016
rect 154262 154780 189706 155016
rect 189942 154780 190026 155016
rect 190262 154780 225706 155016
rect 225942 154780 226026 155016
rect 226262 154780 261706 155016
rect 261942 154780 262026 155016
rect 262262 154780 297706 155016
rect 297942 154780 298026 155016
rect 298262 154780 333706 155016
rect 333942 154780 334026 155016
rect 334262 154780 369706 155016
rect 369942 154780 370026 155016
rect 370262 154780 405706 155016
rect 405942 154780 406026 155016
rect 406262 154780 441706 155016
rect 441942 154780 442026 155016
rect 442262 154780 477706 155016
rect 477942 154780 478026 155016
rect 478262 154780 513706 155016
rect 513942 154780 514026 155016
rect 514262 154780 549706 155016
rect 549942 154780 550026 155016
rect 550262 154780 592062 155016
rect 592298 154780 592382 155016
rect 592618 154780 592650 155016
rect -8726 154748 592650 154780
rect -8726 154096 592650 154128
rect -8726 153860 -7734 154096
rect -7498 153860 -7414 154096
rect -7178 153860 8466 154096
rect 8702 153860 8786 154096
rect 9022 153860 44466 154096
rect 44702 153860 44786 154096
rect 45022 153860 80466 154096
rect 80702 153860 80786 154096
rect 81022 153860 116466 154096
rect 116702 153860 116786 154096
rect 117022 153860 152466 154096
rect 152702 153860 152786 154096
rect 153022 153860 188466 154096
rect 188702 153860 188786 154096
rect 189022 153860 224466 154096
rect 224702 153860 224786 154096
rect 225022 153860 260466 154096
rect 260702 153860 260786 154096
rect 261022 153860 296466 154096
rect 296702 153860 296786 154096
rect 297022 153860 332466 154096
rect 332702 153860 332786 154096
rect 333022 153860 368466 154096
rect 368702 153860 368786 154096
rect 369022 153860 404466 154096
rect 404702 153860 404786 154096
rect 405022 153860 440466 154096
rect 440702 153860 440786 154096
rect 441022 153860 476466 154096
rect 476702 153860 476786 154096
rect 477022 153860 512466 154096
rect 512702 153860 512786 154096
rect 513022 153860 548466 154096
rect 548702 153860 548786 154096
rect 549022 153860 591102 154096
rect 591338 153860 591422 154096
rect 591658 153860 592650 154096
rect -8726 153776 592650 153860
rect -8726 153540 -7734 153776
rect -7498 153540 -7414 153776
rect -7178 153540 8466 153776
rect 8702 153540 8786 153776
rect 9022 153540 44466 153776
rect 44702 153540 44786 153776
rect 45022 153540 80466 153776
rect 80702 153540 80786 153776
rect 81022 153540 116466 153776
rect 116702 153540 116786 153776
rect 117022 153540 152466 153776
rect 152702 153540 152786 153776
rect 153022 153540 188466 153776
rect 188702 153540 188786 153776
rect 189022 153540 224466 153776
rect 224702 153540 224786 153776
rect 225022 153540 260466 153776
rect 260702 153540 260786 153776
rect 261022 153540 296466 153776
rect 296702 153540 296786 153776
rect 297022 153540 332466 153776
rect 332702 153540 332786 153776
rect 333022 153540 368466 153776
rect 368702 153540 368786 153776
rect 369022 153540 404466 153776
rect 404702 153540 404786 153776
rect 405022 153540 440466 153776
rect 440702 153540 440786 153776
rect 441022 153540 476466 153776
rect 476702 153540 476786 153776
rect 477022 153540 512466 153776
rect 512702 153540 512786 153776
rect 513022 153540 548466 153776
rect 548702 153540 548786 153776
rect 549022 153540 591102 153776
rect 591338 153540 591422 153776
rect 591658 153540 592650 153776
rect -8726 153508 592650 153540
rect -8726 152856 592650 152888
rect -8726 152620 -6774 152856
rect -6538 152620 -6454 152856
rect -6218 152620 7226 152856
rect 7462 152620 7546 152856
rect 7782 152620 43226 152856
rect 43462 152620 43546 152856
rect 43782 152620 79226 152856
rect 79462 152620 79546 152856
rect 79782 152620 115226 152856
rect 115462 152620 115546 152856
rect 115782 152620 151226 152856
rect 151462 152620 151546 152856
rect 151782 152620 187226 152856
rect 187462 152620 187546 152856
rect 187782 152620 223226 152856
rect 223462 152620 223546 152856
rect 223782 152620 259226 152856
rect 259462 152620 259546 152856
rect 259782 152620 295226 152856
rect 295462 152620 295546 152856
rect 295782 152620 331226 152856
rect 331462 152620 331546 152856
rect 331782 152620 367226 152856
rect 367462 152620 367546 152856
rect 367782 152620 403226 152856
rect 403462 152620 403546 152856
rect 403782 152620 439226 152856
rect 439462 152620 439546 152856
rect 439782 152620 475226 152856
rect 475462 152620 475546 152856
rect 475782 152620 511226 152856
rect 511462 152620 511546 152856
rect 511782 152620 547226 152856
rect 547462 152620 547546 152856
rect 547782 152620 590142 152856
rect 590378 152620 590462 152856
rect 590698 152620 592650 152856
rect -8726 152536 592650 152620
rect -8726 152300 -6774 152536
rect -6538 152300 -6454 152536
rect -6218 152300 7226 152536
rect 7462 152300 7546 152536
rect 7782 152300 43226 152536
rect 43462 152300 43546 152536
rect 43782 152300 79226 152536
rect 79462 152300 79546 152536
rect 79782 152300 115226 152536
rect 115462 152300 115546 152536
rect 115782 152300 151226 152536
rect 151462 152300 151546 152536
rect 151782 152300 187226 152536
rect 187462 152300 187546 152536
rect 187782 152300 223226 152536
rect 223462 152300 223546 152536
rect 223782 152300 259226 152536
rect 259462 152300 259546 152536
rect 259782 152300 295226 152536
rect 295462 152300 295546 152536
rect 295782 152300 331226 152536
rect 331462 152300 331546 152536
rect 331782 152300 367226 152536
rect 367462 152300 367546 152536
rect 367782 152300 403226 152536
rect 403462 152300 403546 152536
rect 403782 152300 439226 152536
rect 439462 152300 439546 152536
rect 439782 152300 475226 152536
rect 475462 152300 475546 152536
rect 475782 152300 511226 152536
rect 511462 152300 511546 152536
rect 511782 152300 547226 152536
rect 547462 152300 547546 152536
rect 547782 152300 590142 152536
rect 590378 152300 590462 152536
rect 590698 152300 592650 152536
rect -8726 152268 592650 152300
rect -8726 151616 592650 151648
rect -8726 151380 -5814 151616
rect -5578 151380 -5494 151616
rect -5258 151380 5986 151616
rect 6222 151380 6306 151616
rect 6542 151380 41986 151616
rect 42222 151380 42306 151616
rect 42542 151380 77986 151616
rect 78222 151380 78306 151616
rect 78542 151380 113986 151616
rect 114222 151380 114306 151616
rect 114542 151380 149986 151616
rect 150222 151380 150306 151616
rect 150542 151380 185986 151616
rect 186222 151380 186306 151616
rect 186542 151380 221986 151616
rect 222222 151380 222306 151616
rect 222542 151380 257986 151616
rect 258222 151380 258306 151616
rect 258542 151380 293986 151616
rect 294222 151380 294306 151616
rect 294542 151380 329986 151616
rect 330222 151380 330306 151616
rect 330542 151380 365986 151616
rect 366222 151380 366306 151616
rect 366542 151380 401986 151616
rect 402222 151380 402306 151616
rect 402542 151380 437986 151616
rect 438222 151380 438306 151616
rect 438542 151380 473986 151616
rect 474222 151380 474306 151616
rect 474542 151380 509986 151616
rect 510222 151380 510306 151616
rect 510542 151380 545986 151616
rect 546222 151380 546306 151616
rect 546542 151380 581986 151616
rect 582222 151380 582306 151616
rect 582542 151380 589182 151616
rect 589418 151380 589502 151616
rect 589738 151380 592650 151616
rect -8726 151296 592650 151380
rect -8726 151060 -5814 151296
rect -5578 151060 -5494 151296
rect -5258 151060 5986 151296
rect 6222 151060 6306 151296
rect 6542 151060 41986 151296
rect 42222 151060 42306 151296
rect 42542 151060 77986 151296
rect 78222 151060 78306 151296
rect 78542 151060 113986 151296
rect 114222 151060 114306 151296
rect 114542 151060 149986 151296
rect 150222 151060 150306 151296
rect 150542 151060 185986 151296
rect 186222 151060 186306 151296
rect 186542 151060 221986 151296
rect 222222 151060 222306 151296
rect 222542 151060 257986 151296
rect 258222 151060 258306 151296
rect 258542 151060 293986 151296
rect 294222 151060 294306 151296
rect 294542 151060 329986 151296
rect 330222 151060 330306 151296
rect 330542 151060 365986 151296
rect 366222 151060 366306 151296
rect 366542 151060 401986 151296
rect 402222 151060 402306 151296
rect 402542 151060 437986 151296
rect 438222 151060 438306 151296
rect 438542 151060 473986 151296
rect 474222 151060 474306 151296
rect 474542 151060 509986 151296
rect 510222 151060 510306 151296
rect 510542 151060 545986 151296
rect 546222 151060 546306 151296
rect 546542 151060 581986 151296
rect 582222 151060 582306 151296
rect 582542 151060 589182 151296
rect 589418 151060 589502 151296
rect 589738 151060 592650 151296
rect -8726 151028 592650 151060
rect -8726 150376 592650 150408
rect -8726 150140 -4854 150376
rect -4618 150140 -4534 150376
rect -4298 150140 4746 150376
rect 4982 150140 5066 150376
rect 5302 150140 40746 150376
rect 40982 150140 41066 150376
rect 41302 150140 76746 150376
rect 76982 150140 77066 150376
rect 77302 150140 112746 150376
rect 112982 150140 113066 150376
rect 113302 150140 148746 150376
rect 148982 150140 149066 150376
rect 149302 150140 184746 150376
rect 184982 150140 185066 150376
rect 185302 150140 220746 150376
rect 220982 150140 221066 150376
rect 221302 150140 256746 150376
rect 256982 150140 257066 150376
rect 257302 150140 292746 150376
rect 292982 150140 293066 150376
rect 293302 150140 328746 150376
rect 328982 150140 329066 150376
rect 329302 150140 364746 150376
rect 364982 150140 365066 150376
rect 365302 150140 400746 150376
rect 400982 150140 401066 150376
rect 401302 150140 436746 150376
rect 436982 150140 437066 150376
rect 437302 150140 472746 150376
rect 472982 150140 473066 150376
rect 473302 150140 508746 150376
rect 508982 150140 509066 150376
rect 509302 150140 544746 150376
rect 544982 150140 545066 150376
rect 545302 150140 580746 150376
rect 580982 150140 581066 150376
rect 581302 150140 588222 150376
rect 588458 150140 588542 150376
rect 588778 150140 592650 150376
rect -8726 150056 592650 150140
rect -8726 149820 -4854 150056
rect -4618 149820 -4534 150056
rect -4298 149820 4746 150056
rect 4982 149820 5066 150056
rect 5302 149820 40746 150056
rect 40982 149820 41066 150056
rect 41302 149820 76746 150056
rect 76982 149820 77066 150056
rect 77302 149820 112746 150056
rect 112982 149820 113066 150056
rect 113302 149820 148746 150056
rect 148982 149820 149066 150056
rect 149302 149820 184746 150056
rect 184982 149820 185066 150056
rect 185302 149820 220746 150056
rect 220982 149820 221066 150056
rect 221302 149820 256746 150056
rect 256982 149820 257066 150056
rect 257302 149820 292746 150056
rect 292982 149820 293066 150056
rect 293302 149820 328746 150056
rect 328982 149820 329066 150056
rect 329302 149820 364746 150056
rect 364982 149820 365066 150056
rect 365302 149820 400746 150056
rect 400982 149820 401066 150056
rect 401302 149820 436746 150056
rect 436982 149820 437066 150056
rect 437302 149820 472746 150056
rect 472982 149820 473066 150056
rect 473302 149820 508746 150056
rect 508982 149820 509066 150056
rect 509302 149820 544746 150056
rect 544982 149820 545066 150056
rect 545302 149820 580746 150056
rect 580982 149820 581066 150056
rect 581302 149820 588222 150056
rect 588458 149820 588542 150056
rect 588778 149820 592650 150056
rect -8726 149788 592650 149820
rect -8726 149136 592650 149168
rect -8726 148900 -3894 149136
rect -3658 148900 -3574 149136
rect -3338 148900 3506 149136
rect 3742 148900 3826 149136
rect 4062 148900 39506 149136
rect 39742 148900 39826 149136
rect 40062 148900 75506 149136
rect 75742 148900 75826 149136
rect 76062 148900 111506 149136
rect 111742 148900 111826 149136
rect 112062 148900 147506 149136
rect 147742 148900 147826 149136
rect 148062 148900 183506 149136
rect 183742 148900 183826 149136
rect 184062 148900 219506 149136
rect 219742 148900 219826 149136
rect 220062 148900 255506 149136
rect 255742 148900 255826 149136
rect 256062 148900 291506 149136
rect 291742 148900 291826 149136
rect 292062 148900 327506 149136
rect 327742 148900 327826 149136
rect 328062 148900 363506 149136
rect 363742 148900 363826 149136
rect 364062 148900 399506 149136
rect 399742 148900 399826 149136
rect 400062 148900 435506 149136
rect 435742 148900 435826 149136
rect 436062 148900 471506 149136
rect 471742 148900 471826 149136
rect 472062 148900 507506 149136
rect 507742 148900 507826 149136
rect 508062 148900 543506 149136
rect 543742 148900 543826 149136
rect 544062 148900 579506 149136
rect 579742 148900 579826 149136
rect 580062 148900 587262 149136
rect 587498 148900 587582 149136
rect 587818 148900 592650 149136
rect -8726 148816 592650 148900
rect -8726 148580 -3894 148816
rect -3658 148580 -3574 148816
rect -3338 148580 3506 148816
rect 3742 148580 3826 148816
rect 4062 148580 39506 148816
rect 39742 148580 39826 148816
rect 40062 148580 75506 148816
rect 75742 148580 75826 148816
rect 76062 148580 111506 148816
rect 111742 148580 111826 148816
rect 112062 148580 147506 148816
rect 147742 148580 147826 148816
rect 148062 148580 183506 148816
rect 183742 148580 183826 148816
rect 184062 148580 219506 148816
rect 219742 148580 219826 148816
rect 220062 148580 255506 148816
rect 255742 148580 255826 148816
rect 256062 148580 291506 148816
rect 291742 148580 291826 148816
rect 292062 148580 327506 148816
rect 327742 148580 327826 148816
rect 328062 148580 363506 148816
rect 363742 148580 363826 148816
rect 364062 148580 399506 148816
rect 399742 148580 399826 148816
rect 400062 148580 435506 148816
rect 435742 148580 435826 148816
rect 436062 148580 471506 148816
rect 471742 148580 471826 148816
rect 472062 148580 507506 148816
rect 507742 148580 507826 148816
rect 508062 148580 543506 148816
rect 543742 148580 543826 148816
rect 544062 148580 579506 148816
rect 579742 148580 579826 148816
rect 580062 148580 587262 148816
rect 587498 148580 587582 148816
rect 587818 148580 592650 148816
rect -8726 148548 592650 148580
rect -8726 147896 592650 147928
rect -8726 147660 -2934 147896
rect -2698 147660 -2614 147896
rect -2378 147660 2266 147896
rect 2502 147660 2586 147896
rect 2822 147660 38266 147896
rect 38502 147660 38586 147896
rect 38822 147660 74266 147896
rect 74502 147660 74586 147896
rect 74822 147660 110266 147896
rect 110502 147660 110586 147896
rect 110822 147660 146266 147896
rect 146502 147660 146586 147896
rect 146822 147660 182266 147896
rect 182502 147660 182586 147896
rect 182822 147660 218266 147896
rect 218502 147660 218586 147896
rect 218822 147660 254266 147896
rect 254502 147660 254586 147896
rect 254822 147660 290266 147896
rect 290502 147660 290586 147896
rect 290822 147660 326266 147896
rect 326502 147660 326586 147896
rect 326822 147660 362266 147896
rect 362502 147660 362586 147896
rect 362822 147660 398266 147896
rect 398502 147660 398586 147896
rect 398822 147660 434266 147896
rect 434502 147660 434586 147896
rect 434822 147660 470266 147896
rect 470502 147660 470586 147896
rect 470822 147660 506266 147896
rect 506502 147660 506586 147896
rect 506822 147660 542266 147896
rect 542502 147660 542586 147896
rect 542822 147660 578266 147896
rect 578502 147660 578586 147896
rect 578822 147660 586302 147896
rect 586538 147660 586622 147896
rect 586858 147660 592650 147896
rect -8726 147576 592650 147660
rect -8726 147340 -2934 147576
rect -2698 147340 -2614 147576
rect -2378 147340 2266 147576
rect 2502 147340 2586 147576
rect 2822 147340 38266 147576
rect 38502 147340 38586 147576
rect 38822 147340 74266 147576
rect 74502 147340 74586 147576
rect 74822 147340 110266 147576
rect 110502 147340 110586 147576
rect 110822 147340 146266 147576
rect 146502 147340 146586 147576
rect 146822 147340 182266 147576
rect 182502 147340 182586 147576
rect 182822 147340 218266 147576
rect 218502 147340 218586 147576
rect 218822 147340 254266 147576
rect 254502 147340 254586 147576
rect 254822 147340 290266 147576
rect 290502 147340 290586 147576
rect 290822 147340 326266 147576
rect 326502 147340 326586 147576
rect 326822 147340 362266 147576
rect 362502 147340 362586 147576
rect 362822 147340 398266 147576
rect 398502 147340 398586 147576
rect 398822 147340 434266 147576
rect 434502 147340 434586 147576
rect 434822 147340 470266 147576
rect 470502 147340 470586 147576
rect 470822 147340 506266 147576
rect 506502 147340 506586 147576
rect 506822 147340 542266 147576
rect 542502 147340 542586 147576
rect 542822 147340 578266 147576
rect 578502 147340 578586 147576
rect 578822 147340 586302 147576
rect 586538 147340 586622 147576
rect 586858 147340 592650 147576
rect -8726 147308 592650 147340
rect -8726 146656 592650 146688
rect -8726 146420 -1974 146656
rect -1738 146420 -1654 146656
rect -1418 146420 1026 146656
rect 1262 146420 1346 146656
rect 1582 146420 37026 146656
rect 37262 146420 37346 146656
rect 37582 146420 73026 146656
rect 73262 146420 73346 146656
rect 73582 146420 109026 146656
rect 109262 146420 109346 146656
rect 109582 146420 145026 146656
rect 145262 146420 145346 146656
rect 145582 146420 181026 146656
rect 181262 146420 181346 146656
rect 181582 146420 217026 146656
rect 217262 146420 217346 146656
rect 217582 146420 253026 146656
rect 253262 146420 253346 146656
rect 253582 146420 289026 146656
rect 289262 146420 289346 146656
rect 289582 146420 325026 146656
rect 325262 146420 325346 146656
rect 325582 146420 361026 146656
rect 361262 146420 361346 146656
rect 361582 146420 397026 146656
rect 397262 146420 397346 146656
rect 397582 146420 433026 146656
rect 433262 146420 433346 146656
rect 433582 146420 469026 146656
rect 469262 146420 469346 146656
rect 469582 146420 505026 146656
rect 505262 146420 505346 146656
rect 505582 146420 541026 146656
rect 541262 146420 541346 146656
rect 541582 146420 577026 146656
rect 577262 146420 577346 146656
rect 577582 146420 585342 146656
rect 585578 146420 585662 146656
rect 585898 146420 592650 146656
rect -8726 146336 592650 146420
rect -8726 146100 -1974 146336
rect -1738 146100 -1654 146336
rect -1418 146100 1026 146336
rect 1262 146100 1346 146336
rect 1582 146100 37026 146336
rect 37262 146100 37346 146336
rect 37582 146100 73026 146336
rect 73262 146100 73346 146336
rect 73582 146100 109026 146336
rect 109262 146100 109346 146336
rect 109582 146100 145026 146336
rect 145262 146100 145346 146336
rect 145582 146100 181026 146336
rect 181262 146100 181346 146336
rect 181582 146100 217026 146336
rect 217262 146100 217346 146336
rect 217582 146100 253026 146336
rect 253262 146100 253346 146336
rect 253582 146100 289026 146336
rect 289262 146100 289346 146336
rect 289582 146100 325026 146336
rect 325262 146100 325346 146336
rect 325582 146100 361026 146336
rect 361262 146100 361346 146336
rect 361582 146100 397026 146336
rect 397262 146100 397346 146336
rect 397582 146100 433026 146336
rect 433262 146100 433346 146336
rect 433582 146100 469026 146336
rect 469262 146100 469346 146336
rect 469582 146100 505026 146336
rect 505262 146100 505346 146336
rect 505582 146100 541026 146336
rect 541262 146100 541346 146336
rect 541582 146100 577026 146336
rect 577262 146100 577346 146336
rect 577582 146100 585342 146336
rect 585578 146100 585662 146336
rect 585898 146100 592650 146336
rect -8726 146068 592650 146100
rect -8726 119336 592650 119368
rect -8726 119100 -8694 119336
rect -8458 119100 -8374 119336
rect -8138 119100 9706 119336
rect 9942 119100 10026 119336
rect 10262 119100 45706 119336
rect 45942 119100 46026 119336
rect 46262 119100 81706 119336
rect 81942 119100 82026 119336
rect 82262 119100 117706 119336
rect 117942 119100 118026 119336
rect 118262 119100 153706 119336
rect 153942 119100 154026 119336
rect 154262 119100 189706 119336
rect 189942 119100 190026 119336
rect 190262 119100 225706 119336
rect 225942 119100 226026 119336
rect 226262 119100 261706 119336
rect 261942 119100 262026 119336
rect 262262 119100 297706 119336
rect 297942 119100 298026 119336
rect 298262 119100 333706 119336
rect 333942 119100 334026 119336
rect 334262 119100 369706 119336
rect 369942 119100 370026 119336
rect 370262 119100 405706 119336
rect 405942 119100 406026 119336
rect 406262 119100 441706 119336
rect 441942 119100 442026 119336
rect 442262 119100 477706 119336
rect 477942 119100 478026 119336
rect 478262 119100 513706 119336
rect 513942 119100 514026 119336
rect 514262 119100 549706 119336
rect 549942 119100 550026 119336
rect 550262 119100 592062 119336
rect 592298 119100 592382 119336
rect 592618 119100 592650 119336
rect -8726 119016 592650 119100
rect -8726 118780 -8694 119016
rect -8458 118780 -8374 119016
rect -8138 118780 9706 119016
rect 9942 118780 10026 119016
rect 10262 118780 45706 119016
rect 45942 118780 46026 119016
rect 46262 118780 81706 119016
rect 81942 118780 82026 119016
rect 82262 118780 117706 119016
rect 117942 118780 118026 119016
rect 118262 118780 153706 119016
rect 153942 118780 154026 119016
rect 154262 118780 189706 119016
rect 189942 118780 190026 119016
rect 190262 118780 225706 119016
rect 225942 118780 226026 119016
rect 226262 118780 261706 119016
rect 261942 118780 262026 119016
rect 262262 118780 297706 119016
rect 297942 118780 298026 119016
rect 298262 118780 333706 119016
rect 333942 118780 334026 119016
rect 334262 118780 369706 119016
rect 369942 118780 370026 119016
rect 370262 118780 405706 119016
rect 405942 118780 406026 119016
rect 406262 118780 441706 119016
rect 441942 118780 442026 119016
rect 442262 118780 477706 119016
rect 477942 118780 478026 119016
rect 478262 118780 513706 119016
rect 513942 118780 514026 119016
rect 514262 118780 549706 119016
rect 549942 118780 550026 119016
rect 550262 118780 592062 119016
rect 592298 118780 592382 119016
rect 592618 118780 592650 119016
rect -8726 118748 592650 118780
rect -8726 118096 592650 118128
rect -8726 117860 -7734 118096
rect -7498 117860 -7414 118096
rect -7178 117860 8466 118096
rect 8702 117860 8786 118096
rect 9022 117860 44466 118096
rect 44702 117860 44786 118096
rect 45022 117860 80466 118096
rect 80702 117860 80786 118096
rect 81022 117860 116466 118096
rect 116702 117860 116786 118096
rect 117022 117860 152466 118096
rect 152702 117860 152786 118096
rect 153022 117860 188466 118096
rect 188702 117860 188786 118096
rect 189022 117860 224466 118096
rect 224702 117860 224786 118096
rect 225022 117860 260466 118096
rect 260702 117860 260786 118096
rect 261022 117860 296466 118096
rect 296702 117860 296786 118096
rect 297022 117860 332466 118096
rect 332702 117860 332786 118096
rect 333022 117860 368466 118096
rect 368702 117860 368786 118096
rect 369022 117860 404466 118096
rect 404702 117860 404786 118096
rect 405022 117860 440466 118096
rect 440702 117860 440786 118096
rect 441022 117860 476466 118096
rect 476702 117860 476786 118096
rect 477022 117860 512466 118096
rect 512702 117860 512786 118096
rect 513022 117860 548466 118096
rect 548702 117860 548786 118096
rect 549022 117860 591102 118096
rect 591338 117860 591422 118096
rect 591658 117860 592650 118096
rect -8726 117776 592650 117860
rect -8726 117540 -7734 117776
rect -7498 117540 -7414 117776
rect -7178 117540 8466 117776
rect 8702 117540 8786 117776
rect 9022 117540 44466 117776
rect 44702 117540 44786 117776
rect 45022 117540 80466 117776
rect 80702 117540 80786 117776
rect 81022 117540 116466 117776
rect 116702 117540 116786 117776
rect 117022 117540 152466 117776
rect 152702 117540 152786 117776
rect 153022 117540 188466 117776
rect 188702 117540 188786 117776
rect 189022 117540 224466 117776
rect 224702 117540 224786 117776
rect 225022 117540 260466 117776
rect 260702 117540 260786 117776
rect 261022 117540 296466 117776
rect 296702 117540 296786 117776
rect 297022 117540 332466 117776
rect 332702 117540 332786 117776
rect 333022 117540 368466 117776
rect 368702 117540 368786 117776
rect 369022 117540 404466 117776
rect 404702 117540 404786 117776
rect 405022 117540 440466 117776
rect 440702 117540 440786 117776
rect 441022 117540 476466 117776
rect 476702 117540 476786 117776
rect 477022 117540 512466 117776
rect 512702 117540 512786 117776
rect 513022 117540 548466 117776
rect 548702 117540 548786 117776
rect 549022 117540 591102 117776
rect 591338 117540 591422 117776
rect 591658 117540 592650 117776
rect -8726 117508 592650 117540
rect -8726 116856 592650 116888
rect -8726 116620 -6774 116856
rect -6538 116620 -6454 116856
rect -6218 116620 7226 116856
rect 7462 116620 7546 116856
rect 7782 116620 43226 116856
rect 43462 116620 43546 116856
rect 43782 116620 79226 116856
rect 79462 116620 79546 116856
rect 79782 116620 115226 116856
rect 115462 116620 115546 116856
rect 115782 116620 151226 116856
rect 151462 116620 151546 116856
rect 151782 116620 187226 116856
rect 187462 116620 187546 116856
rect 187782 116620 223226 116856
rect 223462 116620 223546 116856
rect 223782 116620 259226 116856
rect 259462 116620 259546 116856
rect 259782 116620 295226 116856
rect 295462 116620 295546 116856
rect 295782 116620 331226 116856
rect 331462 116620 331546 116856
rect 331782 116620 367226 116856
rect 367462 116620 367546 116856
rect 367782 116620 403226 116856
rect 403462 116620 403546 116856
rect 403782 116620 439226 116856
rect 439462 116620 439546 116856
rect 439782 116620 475226 116856
rect 475462 116620 475546 116856
rect 475782 116620 511226 116856
rect 511462 116620 511546 116856
rect 511782 116620 547226 116856
rect 547462 116620 547546 116856
rect 547782 116620 590142 116856
rect 590378 116620 590462 116856
rect 590698 116620 592650 116856
rect -8726 116536 592650 116620
rect -8726 116300 -6774 116536
rect -6538 116300 -6454 116536
rect -6218 116300 7226 116536
rect 7462 116300 7546 116536
rect 7782 116300 43226 116536
rect 43462 116300 43546 116536
rect 43782 116300 79226 116536
rect 79462 116300 79546 116536
rect 79782 116300 115226 116536
rect 115462 116300 115546 116536
rect 115782 116300 151226 116536
rect 151462 116300 151546 116536
rect 151782 116300 187226 116536
rect 187462 116300 187546 116536
rect 187782 116300 223226 116536
rect 223462 116300 223546 116536
rect 223782 116300 259226 116536
rect 259462 116300 259546 116536
rect 259782 116300 295226 116536
rect 295462 116300 295546 116536
rect 295782 116300 331226 116536
rect 331462 116300 331546 116536
rect 331782 116300 367226 116536
rect 367462 116300 367546 116536
rect 367782 116300 403226 116536
rect 403462 116300 403546 116536
rect 403782 116300 439226 116536
rect 439462 116300 439546 116536
rect 439782 116300 475226 116536
rect 475462 116300 475546 116536
rect 475782 116300 511226 116536
rect 511462 116300 511546 116536
rect 511782 116300 547226 116536
rect 547462 116300 547546 116536
rect 547782 116300 590142 116536
rect 590378 116300 590462 116536
rect 590698 116300 592650 116536
rect -8726 116268 592650 116300
rect -8726 115616 592650 115648
rect -8726 115380 -5814 115616
rect -5578 115380 -5494 115616
rect -5258 115380 5986 115616
rect 6222 115380 6306 115616
rect 6542 115380 41986 115616
rect 42222 115380 42306 115616
rect 42542 115380 77986 115616
rect 78222 115380 78306 115616
rect 78542 115380 113986 115616
rect 114222 115380 114306 115616
rect 114542 115380 149986 115616
rect 150222 115380 150306 115616
rect 150542 115380 185986 115616
rect 186222 115380 186306 115616
rect 186542 115380 221986 115616
rect 222222 115380 222306 115616
rect 222542 115380 257986 115616
rect 258222 115380 258306 115616
rect 258542 115380 293986 115616
rect 294222 115380 294306 115616
rect 294542 115380 329986 115616
rect 330222 115380 330306 115616
rect 330542 115380 365986 115616
rect 366222 115380 366306 115616
rect 366542 115380 401986 115616
rect 402222 115380 402306 115616
rect 402542 115380 437986 115616
rect 438222 115380 438306 115616
rect 438542 115380 473986 115616
rect 474222 115380 474306 115616
rect 474542 115380 509986 115616
rect 510222 115380 510306 115616
rect 510542 115380 545986 115616
rect 546222 115380 546306 115616
rect 546542 115380 581986 115616
rect 582222 115380 582306 115616
rect 582542 115380 589182 115616
rect 589418 115380 589502 115616
rect 589738 115380 592650 115616
rect -8726 115296 592650 115380
rect -8726 115060 -5814 115296
rect -5578 115060 -5494 115296
rect -5258 115060 5986 115296
rect 6222 115060 6306 115296
rect 6542 115060 41986 115296
rect 42222 115060 42306 115296
rect 42542 115060 77986 115296
rect 78222 115060 78306 115296
rect 78542 115060 113986 115296
rect 114222 115060 114306 115296
rect 114542 115060 149986 115296
rect 150222 115060 150306 115296
rect 150542 115060 185986 115296
rect 186222 115060 186306 115296
rect 186542 115060 221986 115296
rect 222222 115060 222306 115296
rect 222542 115060 257986 115296
rect 258222 115060 258306 115296
rect 258542 115060 293986 115296
rect 294222 115060 294306 115296
rect 294542 115060 329986 115296
rect 330222 115060 330306 115296
rect 330542 115060 365986 115296
rect 366222 115060 366306 115296
rect 366542 115060 401986 115296
rect 402222 115060 402306 115296
rect 402542 115060 437986 115296
rect 438222 115060 438306 115296
rect 438542 115060 473986 115296
rect 474222 115060 474306 115296
rect 474542 115060 509986 115296
rect 510222 115060 510306 115296
rect 510542 115060 545986 115296
rect 546222 115060 546306 115296
rect 546542 115060 581986 115296
rect 582222 115060 582306 115296
rect 582542 115060 589182 115296
rect 589418 115060 589502 115296
rect 589738 115060 592650 115296
rect -8726 115028 592650 115060
rect -8726 114376 592650 114408
rect -8726 114140 -4854 114376
rect -4618 114140 -4534 114376
rect -4298 114140 4746 114376
rect 4982 114140 5066 114376
rect 5302 114140 40746 114376
rect 40982 114140 41066 114376
rect 41302 114140 76746 114376
rect 76982 114140 77066 114376
rect 77302 114140 112746 114376
rect 112982 114140 113066 114376
rect 113302 114140 148746 114376
rect 148982 114140 149066 114376
rect 149302 114140 184746 114376
rect 184982 114140 185066 114376
rect 185302 114140 220746 114376
rect 220982 114140 221066 114376
rect 221302 114140 256746 114376
rect 256982 114140 257066 114376
rect 257302 114140 292746 114376
rect 292982 114140 293066 114376
rect 293302 114140 328746 114376
rect 328982 114140 329066 114376
rect 329302 114140 364746 114376
rect 364982 114140 365066 114376
rect 365302 114140 400746 114376
rect 400982 114140 401066 114376
rect 401302 114140 436746 114376
rect 436982 114140 437066 114376
rect 437302 114140 472746 114376
rect 472982 114140 473066 114376
rect 473302 114140 508746 114376
rect 508982 114140 509066 114376
rect 509302 114140 544746 114376
rect 544982 114140 545066 114376
rect 545302 114140 580746 114376
rect 580982 114140 581066 114376
rect 581302 114140 588222 114376
rect 588458 114140 588542 114376
rect 588778 114140 592650 114376
rect -8726 114056 592650 114140
rect -8726 113820 -4854 114056
rect -4618 113820 -4534 114056
rect -4298 113820 4746 114056
rect 4982 113820 5066 114056
rect 5302 113820 40746 114056
rect 40982 113820 41066 114056
rect 41302 113820 76746 114056
rect 76982 113820 77066 114056
rect 77302 113820 112746 114056
rect 112982 113820 113066 114056
rect 113302 113820 148746 114056
rect 148982 113820 149066 114056
rect 149302 113820 184746 114056
rect 184982 113820 185066 114056
rect 185302 113820 220746 114056
rect 220982 113820 221066 114056
rect 221302 113820 256746 114056
rect 256982 113820 257066 114056
rect 257302 113820 292746 114056
rect 292982 113820 293066 114056
rect 293302 113820 328746 114056
rect 328982 113820 329066 114056
rect 329302 113820 364746 114056
rect 364982 113820 365066 114056
rect 365302 113820 400746 114056
rect 400982 113820 401066 114056
rect 401302 113820 436746 114056
rect 436982 113820 437066 114056
rect 437302 113820 472746 114056
rect 472982 113820 473066 114056
rect 473302 113820 508746 114056
rect 508982 113820 509066 114056
rect 509302 113820 544746 114056
rect 544982 113820 545066 114056
rect 545302 113820 580746 114056
rect 580982 113820 581066 114056
rect 581302 113820 588222 114056
rect 588458 113820 588542 114056
rect 588778 113820 592650 114056
rect -8726 113788 592650 113820
rect -8726 113136 592650 113168
rect -8726 112900 -3894 113136
rect -3658 112900 -3574 113136
rect -3338 112900 3506 113136
rect 3742 112900 3826 113136
rect 4062 112900 39506 113136
rect 39742 112900 39826 113136
rect 40062 112900 75506 113136
rect 75742 112900 75826 113136
rect 76062 112900 111506 113136
rect 111742 112900 111826 113136
rect 112062 112900 147506 113136
rect 147742 112900 147826 113136
rect 148062 112900 183506 113136
rect 183742 112900 183826 113136
rect 184062 112900 219506 113136
rect 219742 112900 219826 113136
rect 220062 112900 255506 113136
rect 255742 112900 255826 113136
rect 256062 112900 291506 113136
rect 291742 112900 291826 113136
rect 292062 112900 327506 113136
rect 327742 112900 327826 113136
rect 328062 112900 363506 113136
rect 363742 112900 363826 113136
rect 364062 112900 399506 113136
rect 399742 112900 399826 113136
rect 400062 112900 435506 113136
rect 435742 112900 435826 113136
rect 436062 112900 471506 113136
rect 471742 112900 471826 113136
rect 472062 112900 507506 113136
rect 507742 112900 507826 113136
rect 508062 112900 543506 113136
rect 543742 112900 543826 113136
rect 544062 112900 579506 113136
rect 579742 112900 579826 113136
rect 580062 112900 587262 113136
rect 587498 112900 587582 113136
rect 587818 112900 592650 113136
rect -8726 112816 592650 112900
rect -8726 112580 -3894 112816
rect -3658 112580 -3574 112816
rect -3338 112580 3506 112816
rect 3742 112580 3826 112816
rect 4062 112580 39506 112816
rect 39742 112580 39826 112816
rect 40062 112580 75506 112816
rect 75742 112580 75826 112816
rect 76062 112580 111506 112816
rect 111742 112580 111826 112816
rect 112062 112580 147506 112816
rect 147742 112580 147826 112816
rect 148062 112580 183506 112816
rect 183742 112580 183826 112816
rect 184062 112580 219506 112816
rect 219742 112580 219826 112816
rect 220062 112580 255506 112816
rect 255742 112580 255826 112816
rect 256062 112580 291506 112816
rect 291742 112580 291826 112816
rect 292062 112580 327506 112816
rect 327742 112580 327826 112816
rect 328062 112580 363506 112816
rect 363742 112580 363826 112816
rect 364062 112580 399506 112816
rect 399742 112580 399826 112816
rect 400062 112580 435506 112816
rect 435742 112580 435826 112816
rect 436062 112580 471506 112816
rect 471742 112580 471826 112816
rect 472062 112580 507506 112816
rect 507742 112580 507826 112816
rect 508062 112580 543506 112816
rect 543742 112580 543826 112816
rect 544062 112580 579506 112816
rect 579742 112580 579826 112816
rect 580062 112580 587262 112816
rect 587498 112580 587582 112816
rect 587818 112580 592650 112816
rect -8726 112548 592650 112580
rect -8726 111896 592650 111928
rect -8726 111660 -2934 111896
rect -2698 111660 -2614 111896
rect -2378 111660 2266 111896
rect 2502 111660 2586 111896
rect 2822 111660 38266 111896
rect 38502 111660 38586 111896
rect 38822 111660 74266 111896
rect 74502 111660 74586 111896
rect 74822 111660 110266 111896
rect 110502 111660 110586 111896
rect 110822 111660 146266 111896
rect 146502 111660 146586 111896
rect 146822 111660 182266 111896
rect 182502 111660 182586 111896
rect 182822 111660 218266 111896
rect 218502 111660 218586 111896
rect 218822 111660 254266 111896
rect 254502 111660 254586 111896
rect 254822 111660 290266 111896
rect 290502 111660 290586 111896
rect 290822 111660 326266 111896
rect 326502 111660 326586 111896
rect 326822 111660 362266 111896
rect 362502 111660 362586 111896
rect 362822 111660 398266 111896
rect 398502 111660 398586 111896
rect 398822 111660 434266 111896
rect 434502 111660 434586 111896
rect 434822 111660 470266 111896
rect 470502 111660 470586 111896
rect 470822 111660 506266 111896
rect 506502 111660 506586 111896
rect 506822 111660 542266 111896
rect 542502 111660 542586 111896
rect 542822 111660 578266 111896
rect 578502 111660 578586 111896
rect 578822 111660 586302 111896
rect 586538 111660 586622 111896
rect 586858 111660 592650 111896
rect -8726 111576 592650 111660
rect -8726 111340 -2934 111576
rect -2698 111340 -2614 111576
rect -2378 111340 2266 111576
rect 2502 111340 2586 111576
rect 2822 111340 38266 111576
rect 38502 111340 38586 111576
rect 38822 111340 74266 111576
rect 74502 111340 74586 111576
rect 74822 111340 110266 111576
rect 110502 111340 110586 111576
rect 110822 111340 146266 111576
rect 146502 111340 146586 111576
rect 146822 111340 182266 111576
rect 182502 111340 182586 111576
rect 182822 111340 218266 111576
rect 218502 111340 218586 111576
rect 218822 111340 254266 111576
rect 254502 111340 254586 111576
rect 254822 111340 290266 111576
rect 290502 111340 290586 111576
rect 290822 111340 326266 111576
rect 326502 111340 326586 111576
rect 326822 111340 362266 111576
rect 362502 111340 362586 111576
rect 362822 111340 398266 111576
rect 398502 111340 398586 111576
rect 398822 111340 434266 111576
rect 434502 111340 434586 111576
rect 434822 111340 470266 111576
rect 470502 111340 470586 111576
rect 470822 111340 506266 111576
rect 506502 111340 506586 111576
rect 506822 111340 542266 111576
rect 542502 111340 542586 111576
rect 542822 111340 578266 111576
rect 578502 111340 578586 111576
rect 578822 111340 586302 111576
rect 586538 111340 586622 111576
rect 586858 111340 592650 111576
rect -8726 111308 592650 111340
rect -8726 110656 592650 110688
rect -8726 110420 -1974 110656
rect -1738 110420 -1654 110656
rect -1418 110420 1026 110656
rect 1262 110420 1346 110656
rect 1582 110420 37026 110656
rect 37262 110420 37346 110656
rect 37582 110420 73026 110656
rect 73262 110420 73346 110656
rect 73582 110420 109026 110656
rect 109262 110420 109346 110656
rect 109582 110420 145026 110656
rect 145262 110420 145346 110656
rect 145582 110420 181026 110656
rect 181262 110420 181346 110656
rect 181582 110420 217026 110656
rect 217262 110420 217346 110656
rect 217582 110420 253026 110656
rect 253262 110420 253346 110656
rect 253582 110420 289026 110656
rect 289262 110420 289346 110656
rect 289582 110420 325026 110656
rect 325262 110420 325346 110656
rect 325582 110420 361026 110656
rect 361262 110420 361346 110656
rect 361582 110420 397026 110656
rect 397262 110420 397346 110656
rect 397582 110420 433026 110656
rect 433262 110420 433346 110656
rect 433582 110420 469026 110656
rect 469262 110420 469346 110656
rect 469582 110420 505026 110656
rect 505262 110420 505346 110656
rect 505582 110420 541026 110656
rect 541262 110420 541346 110656
rect 541582 110420 577026 110656
rect 577262 110420 577346 110656
rect 577582 110420 585342 110656
rect 585578 110420 585662 110656
rect 585898 110420 592650 110656
rect -8726 110336 592650 110420
rect -8726 110100 -1974 110336
rect -1738 110100 -1654 110336
rect -1418 110100 1026 110336
rect 1262 110100 1346 110336
rect 1582 110100 37026 110336
rect 37262 110100 37346 110336
rect 37582 110100 73026 110336
rect 73262 110100 73346 110336
rect 73582 110100 109026 110336
rect 109262 110100 109346 110336
rect 109582 110100 145026 110336
rect 145262 110100 145346 110336
rect 145582 110100 181026 110336
rect 181262 110100 181346 110336
rect 181582 110100 217026 110336
rect 217262 110100 217346 110336
rect 217582 110100 253026 110336
rect 253262 110100 253346 110336
rect 253582 110100 289026 110336
rect 289262 110100 289346 110336
rect 289582 110100 325026 110336
rect 325262 110100 325346 110336
rect 325582 110100 361026 110336
rect 361262 110100 361346 110336
rect 361582 110100 397026 110336
rect 397262 110100 397346 110336
rect 397582 110100 433026 110336
rect 433262 110100 433346 110336
rect 433582 110100 469026 110336
rect 469262 110100 469346 110336
rect 469582 110100 505026 110336
rect 505262 110100 505346 110336
rect 505582 110100 541026 110336
rect 541262 110100 541346 110336
rect 541582 110100 577026 110336
rect 577262 110100 577346 110336
rect 577582 110100 585342 110336
rect 585578 110100 585662 110336
rect 585898 110100 592650 110336
rect -8726 110068 592650 110100
rect -8726 83336 592650 83368
rect -8726 83100 -8694 83336
rect -8458 83100 -8374 83336
rect -8138 83100 9706 83336
rect 9942 83100 10026 83336
rect 10262 83100 45706 83336
rect 45942 83100 46026 83336
rect 46262 83100 81706 83336
rect 81942 83100 82026 83336
rect 82262 83100 117706 83336
rect 117942 83100 118026 83336
rect 118262 83100 153706 83336
rect 153942 83100 154026 83336
rect 154262 83100 189706 83336
rect 189942 83100 190026 83336
rect 190262 83100 225706 83336
rect 225942 83100 226026 83336
rect 226262 83100 261706 83336
rect 261942 83100 262026 83336
rect 262262 83100 297706 83336
rect 297942 83100 298026 83336
rect 298262 83100 333706 83336
rect 333942 83100 334026 83336
rect 334262 83100 369706 83336
rect 369942 83100 370026 83336
rect 370262 83100 405706 83336
rect 405942 83100 406026 83336
rect 406262 83100 441706 83336
rect 441942 83100 442026 83336
rect 442262 83100 477706 83336
rect 477942 83100 478026 83336
rect 478262 83100 513706 83336
rect 513942 83100 514026 83336
rect 514262 83100 549706 83336
rect 549942 83100 550026 83336
rect 550262 83100 592062 83336
rect 592298 83100 592382 83336
rect 592618 83100 592650 83336
rect -8726 83016 592650 83100
rect -8726 82780 -8694 83016
rect -8458 82780 -8374 83016
rect -8138 82780 9706 83016
rect 9942 82780 10026 83016
rect 10262 82780 45706 83016
rect 45942 82780 46026 83016
rect 46262 82780 81706 83016
rect 81942 82780 82026 83016
rect 82262 82780 117706 83016
rect 117942 82780 118026 83016
rect 118262 82780 153706 83016
rect 153942 82780 154026 83016
rect 154262 82780 189706 83016
rect 189942 82780 190026 83016
rect 190262 82780 225706 83016
rect 225942 82780 226026 83016
rect 226262 82780 261706 83016
rect 261942 82780 262026 83016
rect 262262 82780 297706 83016
rect 297942 82780 298026 83016
rect 298262 82780 333706 83016
rect 333942 82780 334026 83016
rect 334262 82780 369706 83016
rect 369942 82780 370026 83016
rect 370262 82780 405706 83016
rect 405942 82780 406026 83016
rect 406262 82780 441706 83016
rect 441942 82780 442026 83016
rect 442262 82780 477706 83016
rect 477942 82780 478026 83016
rect 478262 82780 513706 83016
rect 513942 82780 514026 83016
rect 514262 82780 549706 83016
rect 549942 82780 550026 83016
rect 550262 82780 592062 83016
rect 592298 82780 592382 83016
rect 592618 82780 592650 83016
rect -8726 82748 592650 82780
rect -8726 82096 592650 82128
rect -8726 81860 -7734 82096
rect -7498 81860 -7414 82096
rect -7178 81860 8466 82096
rect 8702 81860 8786 82096
rect 9022 81860 44466 82096
rect 44702 81860 44786 82096
rect 45022 81860 80466 82096
rect 80702 81860 80786 82096
rect 81022 81860 116466 82096
rect 116702 81860 116786 82096
rect 117022 81860 152466 82096
rect 152702 81860 152786 82096
rect 153022 81860 188466 82096
rect 188702 81860 188786 82096
rect 189022 81860 224466 82096
rect 224702 81860 224786 82096
rect 225022 81860 260466 82096
rect 260702 81860 260786 82096
rect 261022 81860 296466 82096
rect 296702 81860 296786 82096
rect 297022 81860 332466 82096
rect 332702 81860 332786 82096
rect 333022 81860 368466 82096
rect 368702 81860 368786 82096
rect 369022 81860 404466 82096
rect 404702 81860 404786 82096
rect 405022 81860 440466 82096
rect 440702 81860 440786 82096
rect 441022 81860 476466 82096
rect 476702 81860 476786 82096
rect 477022 81860 512466 82096
rect 512702 81860 512786 82096
rect 513022 81860 548466 82096
rect 548702 81860 548786 82096
rect 549022 81860 591102 82096
rect 591338 81860 591422 82096
rect 591658 81860 592650 82096
rect -8726 81776 592650 81860
rect -8726 81540 -7734 81776
rect -7498 81540 -7414 81776
rect -7178 81540 8466 81776
rect 8702 81540 8786 81776
rect 9022 81540 44466 81776
rect 44702 81540 44786 81776
rect 45022 81540 80466 81776
rect 80702 81540 80786 81776
rect 81022 81540 116466 81776
rect 116702 81540 116786 81776
rect 117022 81540 152466 81776
rect 152702 81540 152786 81776
rect 153022 81540 188466 81776
rect 188702 81540 188786 81776
rect 189022 81540 224466 81776
rect 224702 81540 224786 81776
rect 225022 81540 260466 81776
rect 260702 81540 260786 81776
rect 261022 81540 296466 81776
rect 296702 81540 296786 81776
rect 297022 81540 332466 81776
rect 332702 81540 332786 81776
rect 333022 81540 368466 81776
rect 368702 81540 368786 81776
rect 369022 81540 404466 81776
rect 404702 81540 404786 81776
rect 405022 81540 440466 81776
rect 440702 81540 440786 81776
rect 441022 81540 476466 81776
rect 476702 81540 476786 81776
rect 477022 81540 512466 81776
rect 512702 81540 512786 81776
rect 513022 81540 548466 81776
rect 548702 81540 548786 81776
rect 549022 81540 591102 81776
rect 591338 81540 591422 81776
rect 591658 81540 592650 81776
rect -8726 81508 592650 81540
rect -8726 80856 592650 80888
rect -8726 80620 -6774 80856
rect -6538 80620 -6454 80856
rect -6218 80620 7226 80856
rect 7462 80620 7546 80856
rect 7782 80620 43226 80856
rect 43462 80620 43546 80856
rect 43782 80620 79226 80856
rect 79462 80620 79546 80856
rect 79782 80620 115226 80856
rect 115462 80620 115546 80856
rect 115782 80620 151226 80856
rect 151462 80620 151546 80856
rect 151782 80620 187226 80856
rect 187462 80620 187546 80856
rect 187782 80620 223226 80856
rect 223462 80620 223546 80856
rect 223782 80620 259226 80856
rect 259462 80620 259546 80856
rect 259782 80620 295226 80856
rect 295462 80620 295546 80856
rect 295782 80620 331226 80856
rect 331462 80620 331546 80856
rect 331782 80620 367226 80856
rect 367462 80620 367546 80856
rect 367782 80620 403226 80856
rect 403462 80620 403546 80856
rect 403782 80620 439226 80856
rect 439462 80620 439546 80856
rect 439782 80620 475226 80856
rect 475462 80620 475546 80856
rect 475782 80620 511226 80856
rect 511462 80620 511546 80856
rect 511782 80620 547226 80856
rect 547462 80620 547546 80856
rect 547782 80620 590142 80856
rect 590378 80620 590462 80856
rect 590698 80620 592650 80856
rect -8726 80536 592650 80620
rect -8726 80300 -6774 80536
rect -6538 80300 -6454 80536
rect -6218 80300 7226 80536
rect 7462 80300 7546 80536
rect 7782 80300 43226 80536
rect 43462 80300 43546 80536
rect 43782 80300 79226 80536
rect 79462 80300 79546 80536
rect 79782 80300 115226 80536
rect 115462 80300 115546 80536
rect 115782 80300 151226 80536
rect 151462 80300 151546 80536
rect 151782 80300 187226 80536
rect 187462 80300 187546 80536
rect 187782 80300 223226 80536
rect 223462 80300 223546 80536
rect 223782 80300 259226 80536
rect 259462 80300 259546 80536
rect 259782 80300 295226 80536
rect 295462 80300 295546 80536
rect 295782 80300 331226 80536
rect 331462 80300 331546 80536
rect 331782 80300 367226 80536
rect 367462 80300 367546 80536
rect 367782 80300 403226 80536
rect 403462 80300 403546 80536
rect 403782 80300 439226 80536
rect 439462 80300 439546 80536
rect 439782 80300 475226 80536
rect 475462 80300 475546 80536
rect 475782 80300 511226 80536
rect 511462 80300 511546 80536
rect 511782 80300 547226 80536
rect 547462 80300 547546 80536
rect 547782 80300 590142 80536
rect 590378 80300 590462 80536
rect 590698 80300 592650 80536
rect -8726 80268 592650 80300
rect -8726 79616 592650 79648
rect -8726 79380 -5814 79616
rect -5578 79380 -5494 79616
rect -5258 79380 5986 79616
rect 6222 79380 6306 79616
rect 6542 79380 41986 79616
rect 42222 79380 42306 79616
rect 42542 79380 77986 79616
rect 78222 79380 78306 79616
rect 78542 79380 113986 79616
rect 114222 79380 114306 79616
rect 114542 79380 149986 79616
rect 150222 79380 150306 79616
rect 150542 79380 185986 79616
rect 186222 79380 186306 79616
rect 186542 79380 221986 79616
rect 222222 79380 222306 79616
rect 222542 79380 257986 79616
rect 258222 79380 258306 79616
rect 258542 79380 293986 79616
rect 294222 79380 294306 79616
rect 294542 79380 329986 79616
rect 330222 79380 330306 79616
rect 330542 79380 365986 79616
rect 366222 79380 366306 79616
rect 366542 79380 401986 79616
rect 402222 79380 402306 79616
rect 402542 79380 437986 79616
rect 438222 79380 438306 79616
rect 438542 79380 473986 79616
rect 474222 79380 474306 79616
rect 474542 79380 509986 79616
rect 510222 79380 510306 79616
rect 510542 79380 545986 79616
rect 546222 79380 546306 79616
rect 546542 79380 581986 79616
rect 582222 79380 582306 79616
rect 582542 79380 589182 79616
rect 589418 79380 589502 79616
rect 589738 79380 592650 79616
rect -8726 79296 592650 79380
rect -8726 79060 -5814 79296
rect -5578 79060 -5494 79296
rect -5258 79060 5986 79296
rect 6222 79060 6306 79296
rect 6542 79060 41986 79296
rect 42222 79060 42306 79296
rect 42542 79060 77986 79296
rect 78222 79060 78306 79296
rect 78542 79060 113986 79296
rect 114222 79060 114306 79296
rect 114542 79060 149986 79296
rect 150222 79060 150306 79296
rect 150542 79060 185986 79296
rect 186222 79060 186306 79296
rect 186542 79060 221986 79296
rect 222222 79060 222306 79296
rect 222542 79060 257986 79296
rect 258222 79060 258306 79296
rect 258542 79060 293986 79296
rect 294222 79060 294306 79296
rect 294542 79060 329986 79296
rect 330222 79060 330306 79296
rect 330542 79060 365986 79296
rect 366222 79060 366306 79296
rect 366542 79060 401986 79296
rect 402222 79060 402306 79296
rect 402542 79060 437986 79296
rect 438222 79060 438306 79296
rect 438542 79060 473986 79296
rect 474222 79060 474306 79296
rect 474542 79060 509986 79296
rect 510222 79060 510306 79296
rect 510542 79060 545986 79296
rect 546222 79060 546306 79296
rect 546542 79060 581986 79296
rect 582222 79060 582306 79296
rect 582542 79060 589182 79296
rect 589418 79060 589502 79296
rect 589738 79060 592650 79296
rect -8726 79028 592650 79060
rect -8726 78376 592650 78408
rect -8726 78140 -4854 78376
rect -4618 78140 -4534 78376
rect -4298 78140 4746 78376
rect 4982 78140 5066 78376
rect 5302 78140 40746 78376
rect 40982 78140 41066 78376
rect 41302 78140 76746 78376
rect 76982 78140 77066 78376
rect 77302 78140 112746 78376
rect 112982 78140 113066 78376
rect 113302 78140 148746 78376
rect 148982 78140 149066 78376
rect 149302 78140 184746 78376
rect 184982 78140 185066 78376
rect 185302 78140 220746 78376
rect 220982 78140 221066 78376
rect 221302 78140 256746 78376
rect 256982 78140 257066 78376
rect 257302 78140 292746 78376
rect 292982 78140 293066 78376
rect 293302 78140 328746 78376
rect 328982 78140 329066 78376
rect 329302 78140 364746 78376
rect 364982 78140 365066 78376
rect 365302 78140 400746 78376
rect 400982 78140 401066 78376
rect 401302 78140 436746 78376
rect 436982 78140 437066 78376
rect 437302 78140 472746 78376
rect 472982 78140 473066 78376
rect 473302 78140 508746 78376
rect 508982 78140 509066 78376
rect 509302 78140 544746 78376
rect 544982 78140 545066 78376
rect 545302 78140 580746 78376
rect 580982 78140 581066 78376
rect 581302 78140 588222 78376
rect 588458 78140 588542 78376
rect 588778 78140 592650 78376
rect -8726 78056 592650 78140
rect -8726 77820 -4854 78056
rect -4618 77820 -4534 78056
rect -4298 77820 4746 78056
rect 4982 77820 5066 78056
rect 5302 77820 40746 78056
rect 40982 77820 41066 78056
rect 41302 77820 76746 78056
rect 76982 77820 77066 78056
rect 77302 77820 112746 78056
rect 112982 77820 113066 78056
rect 113302 77820 148746 78056
rect 148982 77820 149066 78056
rect 149302 77820 184746 78056
rect 184982 77820 185066 78056
rect 185302 77820 220746 78056
rect 220982 77820 221066 78056
rect 221302 77820 256746 78056
rect 256982 77820 257066 78056
rect 257302 77820 292746 78056
rect 292982 77820 293066 78056
rect 293302 77820 328746 78056
rect 328982 77820 329066 78056
rect 329302 77820 364746 78056
rect 364982 77820 365066 78056
rect 365302 77820 400746 78056
rect 400982 77820 401066 78056
rect 401302 77820 436746 78056
rect 436982 77820 437066 78056
rect 437302 77820 472746 78056
rect 472982 77820 473066 78056
rect 473302 77820 508746 78056
rect 508982 77820 509066 78056
rect 509302 77820 544746 78056
rect 544982 77820 545066 78056
rect 545302 77820 580746 78056
rect 580982 77820 581066 78056
rect 581302 77820 588222 78056
rect 588458 77820 588542 78056
rect 588778 77820 592650 78056
rect -8726 77788 592650 77820
rect -8726 77136 592650 77168
rect -8726 76900 -3894 77136
rect -3658 76900 -3574 77136
rect -3338 76900 3506 77136
rect 3742 76900 3826 77136
rect 4062 76900 39506 77136
rect 39742 76900 39826 77136
rect 40062 76900 75506 77136
rect 75742 76900 75826 77136
rect 76062 76900 111506 77136
rect 111742 76900 111826 77136
rect 112062 76900 147506 77136
rect 147742 76900 147826 77136
rect 148062 76900 183506 77136
rect 183742 76900 183826 77136
rect 184062 76900 219506 77136
rect 219742 76900 219826 77136
rect 220062 76900 255506 77136
rect 255742 76900 255826 77136
rect 256062 76900 291506 77136
rect 291742 76900 291826 77136
rect 292062 76900 327506 77136
rect 327742 76900 327826 77136
rect 328062 76900 363506 77136
rect 363742 76900 363826 77136
rect 364062 76900 399506 77136
rect 399742 76900 399826 77136
rect 400062 76900 435506 77136
rect 435742 76900 435826 77136
rect 436062 76900 471506 77136
rect 471742 76900 471826 77136
rect 472062 76900 507506 77136
rect 507742 76900 507826 77136
rect 508062 76900 543506 77136
rect 543742 76900 543826 77136
rect 544062 76900 579506 77136
rect 579742 76900 579826 77136
rect 580062 76900 587262 77136
rect 587498 76900 587582 77136
rect 587818 76900 592650 77136
rect -8726 76816 592650 76900
rect -8726 76580 -3894 76816
rect -3658 76580 -3574 76816
rect -3338 76580 3506 76816
rect 3742 76580 3826 76816
rect 4062 76580 39506 76816
rect 39742 76580 39826 76816
rect 40062 76580 75506 76816
rect 75742 76580 75826 76816
rect 76062 76580 111506 76816
rect 111742 76580 111826 76816
rect 112062 76580 147506 76816
rect 147742 76580 147826 76816
rect 148062 76580 183506 76816
rect 183742 76580 183826 76816
rect 184062 76580 219506 76816
rect 219742 76580 219826 76816
rect 220062 76580 255506 76816
rect 255742 76580 255826 76816
rect 256062 76580 291506 76816
rect 291742 76580 291826 76816
rect 292062 76580 327506 76816
rect 327742 76580 327826 76816
rect 328062 76580 363506 76816
rect 363742 76580 363826 76816
rect 364062 76580 399506 76816
rect 399742 76580 399826 76816
rect 400062 76580 435506 76816
rect 435742 76580 435826 76816
rect 436062 76580 471506 76816
rect 471742 76580 471826 76816
rect 472062 76580 507506 76816
rect 507742 76580 507826 76816
rect 508062 76580 543506 76816
rect 543742 76580 543826 76816
rect 544062 76580 579506 76816
rect 579742 76580 579826 76816
rect 580062 76580 587262 76816
rect 587498 76580 587582 76816
rect 587818 76580 592650 76816
rect -8726 76548 592650 76580
rect -8726 75896 592650 75928
rect -8726 75660 -2934 75896
rect -2698 75660 -2614 75896
rect -2378 75660 2266 75896
rect 2502 75660 2586 75896
rect 2822 75660 38266 75896
rect 38502 75660 38586 75896
rect 38822 75660 74266 75896
rect 74502 75660 74586 75896
rect 74822 75660 110266 75896
rect 110502 75660 110586 75896
rect 110822 75660 146266 75896
rect 146502 75660 146586 75896
rect 146822 75660 182266 75896
rect 182502 75660 182586 75896
rect 182822 75660 218266 75896
rect 218502 75660 218586 75896
rect 218822 75660 254266 75896
rect 254502 75660 254586 75896
rect 254822 75660 290266 75896
rect 290502 75660 290586 75896
rect 290822 75660 326266 75896
rect 326502 75660 326586 75896
rect 326822 75660 362266 75896
rect 362502 75660 362586 75896
rect 362822 75660 398266 75896
rect 398502 75660 398586 75896
rect 398822 75660 434266 75896
rect 434502 75660 434586 75896
rect 434822 75660 470266 75896
rect 470502 75660 470586 75896
rect 470822 75660 506266 75896
rect 506502 75660 506586 75896
rect 506822 75660 542266 75896
rect 542502 75660 542586 75896
rect 542822 75660 578266 75896
rect 578502 75660 578586 75896
rect 578822 75660 586302 75896
rect 586538 75660 586622 75896
rect 586858 75660 592650 75896
rect -8726 75576 592650 75660
rect -8726 75340 -2934 75576
rect -2698 75340 -2614 75576
rect -2378 75340 2266 75576
rect 2502 75340 2586 75576
rect 2822 75340 38266 75576
rect 38502 75340 38586 75576
rect 38822 75340 74266 75576
rect 74502 75340 74586 75576
rect 74822 75340 110266 75576
rect 110502 75340 110586 75576
rect 110822 75340 146266 75576
rect 146502 75340 146586 75576
rect 146822 75340 182266 75576
rect 182502 75340 182586 75576
rect 182822 75340 218266 75576
rect 218502 75340 218586 75576
rect 218822 75340 254266 75576
rect 254502 75340 254586 75576
rect 254822 75340 290266 75576
rect 290502 75340 290586 75576
rect 290822 75340 326266 75576
rect 326502 75340 326586 75576
rect 326822 75340 362266 75576
rect 362502 75340 362586 75576
rect 362822 75340 398266 75576
rect 398502 75340 398586 75576
rect 398822 75340 434266 75576
rect 434502 75340 434586 75576
rect 434822 75340 470266 75576
rect 470502 75340 470586 75576
rect 470822 75340 506266 75576
rect 506502 75340 506586 75576
rect 506822 75340 542266 75576
rect 542502 75340 542586 75576
rect 542822 75340 578266 75576
rect 578502 75340 578586 75576
rect 578822 75340 586302 75576
rect 586538 75340 586622 75576
rect 586858 75340 592650 75576
rect -8726 75308 592650 75340
rect -8726 74656 592650 74688
rect -8726 74420 -1974 74656
rect -1738 74420 -1654 74656
rect -1418 74420 1026 74656
rect 1262 74420 1346 74656
rect 1582 74420 37026 74656
rect 37262 74420 37346 74656
rect 37582 74420 73026 74656
rect 73262 74420 73346 74656
rect 73582 74420 109026 74656
rect 109262 74420 109346 74656
rect 109582 74420 145026 74656
rect 145262 74420 145346 74656
rect 145582 74420 181026 74656
rect 181262 74420 181346 74656
rect 181582 74420 217026 74656
rect 217262 74420 217346 74656
rect 217582 74420 253026 74656
rect 253262 74420 253346 74656
rect 253582 74420 289026 74656
rect 289262 74420 289346 74656
rect 289582 74420 325026 74656
rect 325262 74420 325346 74656
rect 325582 74420 361026 74656
rect 361262 74420 361346 74656
rect 361582 74420 397026 74656
rect 397262 74420 397346 74656
rect 397582 74420 433026 74656
rect 433262 74420 433346 74656
rect 433582 74420 469026 74656
rect 469262 74420 469346 74656
rect 469582 74420 505026 74656
rect 505262 74420 505346 74656
rect 505582 74420 541026 74656
rect 541262 74420 541346 74656
rect 541582 74420 577026 74656
rect 577262 74420 577346 74656
rect 577582 74420 585342 74656
rect 585578 74420 585662 74656
rect 585898 74420 592650 74656
rect -8726 74336 592650 74420
rect -8726 74100 -1974 74336
rect -1738 74100 -1654 74336
rect -1418 74100 1026 74336
rect 1262 74100 1346 74336
rect 1582 74100 37026 74336
rect 37262 74100 37346 74336
rect 37582 74100 73026 74336
rect 73262 74100 73346 74336
rect 73582 74100 109026 74336
rect 109262 74100 109346 74336
rect 109582 74100 145026 74336
rect 145262 74100 145346 74336
rect 145582 74100 181026 74336
rect 181262 74100 181346 74336
rect 181582 74100 217026 74336
rect 217262 74100 217346 74336
rect 217582 74100 253026 74336
rect 253262 74100 253346 74336
rect 253582 74100 289026 74336
rect 289262 74100 289346 74336
rect 289582 74100 325026 74336
rect 325262 74100 325346 74336
rect 325582 74100 361026 74336
rect 361262 74100 361346 74336
rect 361582 74100 397026 74336
rect 397262 74100 397346 74336
rect 397582 74100 433026 74336
rect 433262 74100 433346 74336
rect 433582 74100 469026 74336
rect 469262 74100 469346 74336
rect 469582 74100 505026 74336
rect 505262 74100 505346 74336
rect 505582 74100 541026 74336
rect 541262 74100 541346 74336
rect 541582 74100 577026 74336
rect 577262 74100 577346 74336
rect 577582 74100 585342 74336
rect 585578 74100 585662 74336
rect 585898 74100 592650 74336
rect -8726 74068 592650 74100
rect -8726 47336 592650 47368
rect -8726 47100 -8694 47336
rect -8458 47100 -8374 47336
rect -8138 47100 9706 47336
rect 9942 47100 10026 47336
rect 10262 47100 45706 47336
rect 45942 47100 46026 47336
rect 46262 47100 81706 47336
rect 81942 47100 82026 47336
rect 82262 47100 117706 47336
rect 117942 47100 118026 47336
rect 118262 47100 153706 47336
rect 153942 47100 154026 47336
rect 154262 47100 189706 47336
rect 189942 47100 190026 47336
rect 190262 47100 225706 47336
rect 225942 47100 226026 47336
rect 226262 47100 261706 47336
rect 261942 47100 262026 47336
rect 262262 47100 297706 47336
rect 297942 47100 298026 47336
rect 298262 47100 333706 47336
rect 333942 47100 334026 47336
rect 334262 47100 369706 47336
rect 369942 47100 370026 47336
rect 370262 47100 405706 47336
rect 405942 47100 406026 47336
rect 406262 47100 441706 47336
rect 441942 47100 442026 47336
rect 442262 47100 477706 47336
rect 477942 47100 478026 47336
rect 478262 47100 513706 47336
rect 513942 47100 514026 47336
rect 514262 47100 549706 47336
rect 549942 47100 550026 47336
rect 550262 47100 592062 47336
rect 592298 47100 592382 47336
rect 592618 47100 592650 47336
rect -8726 47016 592650 47100
rect -8726 46780 -8694 47016
rect -8458 46780 -8374 47016
rect -8138 46780 9706 47016
rect 9942 46780 10026 47016
rect 10262 46780 45706 47016
rect 45942 46780 46026 47016
rect 46262 46780 81706 47016
rect 81942 46780 82026 47016
rect 82262 46780 117706 47016
rect 117942 46780 118026 47016
rect 118262 46780 153706 47016
rect 153942 46780 154026 47016
rect 154262 46780 189706 47016
rect 189942 46780 190026 47016
rect 190262 46780 225706 47016
rect 225942 46780 226026 47016
rect 226262 46780 261706 47016
rect 261942 46780 262026 47016
rect 262262 46780 297706 47016
rect 297942 46780 298026 47016
rect 298262 46780 333706 47016
rect 333942 46780 334026 47016
rect 334262 46780 369706 47016
rect 369942 46780 370026 47016
rect 370262 46780 405706 47016
rect 405942 46780 406026 47016
rect 406262 46780 441706 47016
rect 441942 46780 442026 47016
rect 442262 46780 477706 47016
rect 477942 46780 478026 47016
rect 478262 46780 513706 47016
rect 513942 46780 514026 47016
rect 514262 46780 549706 47016
rect 549942 46780 550026 47016
rect 550262 46780 592062 47016
rect 592298 46780 592382 47016
rect 592618 46780 592650 47016
rect -8726 46748 592650 46780
rect -8726 46096 592650 46128
rect -8726 45860 -7734 46096
rect -7498 45860 -7414 46096
rect -7178 45860 8466 46096
rect 8702 45860 8786 46096
rect 9022 45860 44466 46096
rect 44702 45860 44786 46096
rect 45022 45860 80466 46096
rect 80702 45860 80786 46096
rect 81022 45860 116466 46096
rect 116702 45860 116786 46096
rect 117022 45860 152466 46096
rect 152702 45860 152786 46096
rect 153022 45860 188466 46096
rect 188702 45860 188786 46096
rect 189022 45860 224466 46096
rect 224702 45860 224786 46096
rect 225022 45860 260466 46096
rect 260702 45860 260786 46096
rect 261022 45860 296466 46096
rect 296702 45860 296786 46096
rect 297022 45860 332466 46096
rect 332702 45860 332786 46096
rect 333022 45860 368466 46096
rect 368702 45860 368786 46096
rect 369022 45860 404466 46096
rect 404702 45860 404786 46096
rect 405022 45860 440466 46096
rect 440702 45860 440786 46096
rect 441022 45860 476466 46096
rect 476702 45860 476786 46096
rect 477022 45860 512466 46096
rect 512702 45860 512786 46096
rect 513022 45860 548466 46096
rect 548702 45860 548786 46096
rect 549022 45860 591102 46096
rect 591338 45860 591422 46096
rect 591658 45860 592650 46096
rect -8726 45776 592650 45860
rect -8726 45540 -7734 45776
rect -7498 45540 -7414 45776
rect -7178 45540 8466 45776
rect 8702 45540 8786 45776
rect 9022 45540 44466 45776
rect 44702 45540 44786 45776
rect 45022 45540 80466 45776
rect 80702 45540 80786 45776
rect 81022 45540 116466 45776
rect 116702 45540 116786 45776
rect 117022 45540 152466 45776
rect 152702 45540 152786 45776
rect 153022 45540 188466 45776
rect 188702 45540 188786 45776
rect 189022 45540 224466 45776
rect 224702 45540 224786 45776
rect 225022 45540 260466 45776
rect 260702 45540 260786 45776
rect 261022 45540 296466 45776
rect 296702 45540 296786 45776
rect 297022 45540 332466 45776
rect 332702 45540 332786 45776
rect 333022 45540 368466 45776
rect 368702 45540 368786 45776
rect 369022 45540 404466 45776
rect 404702 45540 404786 45776
rect 405022 45540 440466 45776
rect 440702 45540 440786 45776
rect 441022 45540 476466 45776
rect 476702 45540 476786 45776
rect 477022 45540 512466 45776
rect 512702 45540 512786 45776
rect 513022 45540 548466 45776
rect 548702 45540 548786 45776
rect 549022 45540 591102 45776
rect 591338 45540 591422 45776
rect 591658 45540 592650 45776
rect -8726 45508 592650 45540
rect -8726 44856 592650 44888
rect -8726 44620 -6774 44856
rect -6538 44620 -6454 44856
rect -6218 44620 7226 44856
rect 7462 44620 7546 44856
rect 7782 44620 43226 44856
rect 43462 44620 43546 44856
rect 43782 44620 79226 44856
rect 79462 44620 79546 44856
rect 79782 44620 115226 44856
rect 115462 44620 115546 44856
rect 115782 44620 151226 44856
rect 151462 44620 151546 44856
rect 151782 44620 187226 44856
rect 187462 44620 187546 44856
rect 187782 44620 223226 44856
rect 223462 44620 223546 44856
rect 223782 44620 259226 44856
rect 259462 44620 259546 44856
rect 259782 44620 295226 44856
rect 295462 44620 295546 44856
rect 295782 44620 331226 44856
rect 331462 44620 331546 44856
rect 331782 44620 367226 44856
rect 367462 44620 367546 44856
rect 367782 44620 403226 44856
rect 403462 44620 403546 44856
rect 403782 44620 439226 44856
rect 439462 44620 439546 44856
rect 439782 44620 475226 44856
rect 475462 44620 475546 44856
rect 475782 44620 511226 44856
rect 511462 44620 511546 44856
rect 511782 44620 547226 44856
rect 547462 44620 547546 44856
rect 547782 44620 590142 44856
rect 590378 44620 590462 44856
rect 590698 44620 592650 44856
rect -8726 44536 592650 44620
rect -8726 44300 -6774 44536
rect -6538 44300 -6454 44536
rect -6218 44300 7226 44536
rect 7462 44300 7546 44536
rect 7782 44300 43226 44536
rect 43462 44300 43546 44536
rect 43782 44300 79226 44536
rect 79462 44300 79546 44536
rect 79782 44300 115226 44536
rect 115462 44300 115546 44536
rect 115782 44300 151226 44536
rect 151462 44300 151546 44536
rect 151782 44300 187226 44536
rect 187462 44300 187546 44536
rect 187782 44300 223226 44536
rect 223462 44300 223546 44536
rect 223782 44300 259226 44536
rect 259462 44300 259546 44536
rect 259782 44300 295226 44536
rect 295462 44300 295546 44536
rect 295782 44300 331226 44536
rect 331462 44300 331546 44536
rect 331782 44300 367226 44536
rect 367462 44300 367546 44536
rect 367782 44300 403226 44536
rect 403462 44300 403546 44536
rect 403782 44300 439226 44536
rect 439462 44300 439546 44536
rect 439782 44300 475226 44536
rect 475462 44300 475546 44536
rect 475782 44300 511226 44536
rect 511462 44300 511546 44536
rect 511782 44300 547226 44536
rect 547462 44300 547546 44536
rect 547782 44300 590142 44536
rect 590378 44300 590462 44536
rect 590698 44300 592650 44536
rect -8726 44268 592650 44300
rect -8726 43616 592650 43648
rect -8726 43380 -5814 43616
rect -5578 43380 -5494 43616
rect -5258 43380 5986 43616
rect 6222 43380 6306 43616
rect 6542 43380 41986 43616
rect 42222 43380 42306 43616
rect 42542 43380 77986 43616
rect 78222 43380 78306 43616
rect 78542 43380 113986 43616
rect 114222 43380 114306 43616
rect 114542 43380 149986 43616
rect 150222 43380 150306 43616
rect 150542 43380 185986 43616
rect 186222 43380 186306 43616
rect 186542 43380 221986 43616
rect 222222 43380 222306 43616
rect 222542 43380 257986 43616
rect 258222 43380 258306 43616
rect 258542 43380 293986 43616
rect 294222 43380 294306 43616
rect 294542 43380 329986 43616
rect 330222 43380 330306 43616
rect 330542 43380 365986 43616
rect 366222 43380 366306 43616
rect 366542 43380 401986 43616
rect 402222 43380 402306 43616
rect 402542 43380 437986 43616
rect 438222 43380 438306 43616
rect 438542 43380 473986 43616
rect 474222 43380 474306 43616
rect 474542 43380 509986 43616
rect 510222 43380 510306 43616
rect 510542 43380 545986 43616
rect 546222 43380 546306 43616
rect 546542 43380 581986 43616
rect 582222 43380 582306 43616
rect 582542 43380 589182 43616
rect 589418 43380 589502 43616
rect 589738 43380 592650 43616
rect -8726 43296 592650 43380
rect -8726 43060 -5814 43296
rect -5578 43060 -5494 43296
rect -5258 43060 5986 43296
rect 6222 43060 6306 43296
rect 6542 43060 41986 43296
rect 42222 43060 42306 43296
rect 42542 43060 77986 43296
rect 78222 43060 78306 43296
rect 78542 43060 113986 43296
rect 114222 43060 114306 43296
rect 114542 43060 149986 43296
rect 150222 43060 150306 43296
rect 150542 43060 185986 43296
rect 186222 43060 186306 43296
rect 186542 43060 221986 43296
rect 222222 43060 222306 43296
rect 222542 43060 257986 43296
rect 258222 43060 258306 43296
rect 258542 43060 293986 43296
rect 294222 43060 294306 43296
rect 294542 43060 329986 43296
rect 330222 43060 330306 43296
rect 330542 43060 365986 43296
rect 366222 43060 366306 43296
rect 366542 43060 401986 43296
rect 402222 43060 402306 43296
rect 402542 43060 437986 43296
rect 438222 43060 438306 43296
rect 438542 43060 473986 43296
rect 474222 43060 474306 43296
rect 474542 43060 509986 43296
rect 510222 43060 510306 43296
rect 510542 43060 545986 43296
rect 546222 43060 546306 43296
rect 546542 43060 581986 43296
rect 582222 43060 582306 43296
rect 582542 43060 589182 43296
rect 589418 43060 589502 43296
rect 589738 43060 592650 43296
rect -8726 43028 592650 43060
rect -8726 42376 592650 42408
rect -8726 42140 -4854 42376
rect -4618 42140 -4534 42376
rect -4298 42140 4746 42376
rect 4982 42140 5066 42376
rect 5302 42140 40746 42376
rect 40982 42140 41066 42376
rect 41302 42140 76746 42376
rect 76982 42140 77066 42376
rect 77302 42140 112746 42376
rect 112982 42140 113066 42376
rect 113302 42140 148746 42376
rect 148982 42140 149066 42376
rect 149302 42140 184746 42376
rect 184982 42140 185066 42376
rect 185302 42140 220746 42376
rect 220982 42140 221066 42376
rect 221302 42140 256746 42376
rect 256982 42140 257066 42376
rect 257302 42140 292746 42376
rect 292982 42140 293066 42376
rect 293302 42140 328746 42376
rect 328982 42140 329066 42376
rect 329302 42140 364746 42376
rect 364982 42140 365066 42376
rect 365302 42140 400746 42376
rect 400982 42140 401066 42376
rect 401302 42140 436746 42376
rect 436982 42140 437066 42376
rect 437302 42140 472746 42376
rect 472982 42140 473066 42376
rect 473302 42140 508746 42376
rect 508982 42140 509066 42376
rect 509302 42140 544746 42376
rect 544982 42140 545066 42376
rect 545302 42140 580746 42376
rect 580982 42140 581066 42376
rect 581302 42140 588222 42376
rect 588458 42140 588542 42376
rect 588778 42140 592650 42376
rect -8726 42056 592650 42140
rect -8726 41820 -4854 42056
rect -4618 41820 -4534 42056
rect -4298 41820 4746 42056
rect 4982 41820 5066 42056
rect 5302 41820 40746 42056
rect 40982 41820 41066 42056
rect 41302 41820 76746 42056
rect 76982 41820 77066 42056
rect 77302 41820 112746 42056
rect 112982 41820 113066 42056
rect 113302 41820 148746 42056
rect 148982 41820 149066 42056
rect 149302 41820 184746 42056
rect 184982 41820 185066 42056
rect 185302 41820 220746 42056
rect 220982 41820 221066 42056
rect 221302 41820 256746 42056
rect 256982 41820 257066 42056
rect 257302 41820 292746 42056
rect 292982 41820 293066 42056
rect 293302 41820 328746 42056
rect 328982 41820 329066 42056
rect 329302 41820 364746 42056
rect 364982 41820 365066 42056
rect 365302 41820 400746 42056
rect 400982 41820 401066 42056
rect 401302 41820 436746 42056
rect 436982 41820 437066 42056
rect 437302 41820 472746 42056
rect 472982 41820 473066 42056
rect 473302 41820 508746 42056
rect 508982 41820 509066 42056
rect 509302 41820 544746 42056
rect 544982 41820 545066 42056
rect 545302 41820 580746 42056
rect 580982 41820 581066 42056
rect 581302 41820 588222 42056
rect 588458 41820 588542 42056
rect 588778 41820 592650 42056
rect -8726 41788 592650 41820
rect -8726 41136 592650 41168
rect -8726 40900 -3894 41136
rect -3658 40900 -3574 41136
rect -3338 40900 3506 41136
rect 3742 40900 3826 41136
rect 4062 40900 39506 41136
rect 39742 40900 39826 41136
rect 40062 40900 75506 41136
rect 75742 40900 75826 41136
rect 76062 40900 111506 41136
rect 111742 40900 111826 41136
rect 112062 40900 147506 41136
rect 147742 40900 147826 41136
rect 148062 40900 183506 41136
rect 183742 40900 183826 41136
rect 184062 40900 219506 41136
rect 219742 40900 219826 41136
rect 220062 40900 255506 41136
rect 255742 40900 255826 41136
rect 256062 40900 291506 41136
rect 291742 40900 291826 41136
rect 292062 40900 327506 41136
rect 327742 40900 327826 41136
rect 328062 40900 363506 41136
rect 363742 40900 363826 41136
rect 364062 40900 399506 41136
rect 399742 40900 399826 41136
rect 400062 40900 435506 41136
rect 435742 40900 435826 41136
rect 436062 40900 471506 41136
rect 471742 40900 471826 41136
rect 472062 40900 507506 41136
rect 507742 40900 507826 41136
rect 508062 40900 543506 41136
rect 543742 40900 543826 41136
rect 544062 40900 579506 41136
rect 579742 40900 579826 41136
rect 580062 40900 587262 41136
rect 587498 40900 587582 41136
rect 587818 40900 592650 41136
rect -8726 40816 592650 40900
rect -8726 40580 -3894 40816
rect -3658 40580 -3574 40816
rect -3338 40580 3506 40816
rect 3742 40580 3826 40816
rect 4062 40580 39506 40816
rect 39742 40580 39826 40816
rect 40062 40580 75506 40816
rect 75742 40580 75826 40816
rect 76062 40580 111506 40816
rect 111742 40580 111826 40816
rect 112062 40580 147506 40816
rect 147742 40580 147826 40816
rect 148062 40580 183506 40816
rect 183742 40580 183826 40816
rect 184062 40580 219506 40816
rect 219742 40580 219826 40816
rect 220062 40580 255506 40816
rect 255742 40580 255826 40816
rect 256062 40580 291506 40816
rect 291742 40580 291826 40816
rect 292062 40580 327506 40816
rect 327742 40580 327826 40816
rect 328062 40580 363506 40816
rect 363742 40580 363826 40816
rect 364062 40580 399506 40816
rect 399742 40580 399826 40816
rect 400062 40580 435506 40816
rect 435742 40580 435826 40816
rect 436062 40580 471506 40816
rect 471742 40580 471826 40816
rect 472062 40580 507506 40816
rect 507742 40580 507826 40816
rect 508062 40580 543506 40816
rect 543742 40580 543826 40816
rect 544062 40580 579506 40816
rect 579742 40580 579826 40816
rect 580062 40580 587262 40816
rect 587498 40580 587582 40816
rect 587818 40580 592650 40816
rect -8726 40548 592650 40580
rect -8726 39896 592650 39928
rect -8726 39660 -2934 39896
rect -2698 39660 -2614 39896
rect -2378 39660 2266 39896
rect 2502 39660 2586 39896
rect 2822 39660 38266 39896
rect 38502 39660 38586 39896
rect 38822 39660 74266 39896
rect 74502 39660 74586 39896
rect 74822 39660 110266 39896
rect 110502 39660 110586 39896
rect 110822 39660 146266 39896
rect 146502 39660 146586 39896
rect 146822 39660 182266 39896
rect 182502 39660 182586 39896
rect 182822 39660 218266 39896
rect 218502 39660 218586 39896
rect 218822 39660 254266 39896
rect 254502 39660 254586 39896
rect 254822 39660 290266 39896
rect 290502 39660 290586 39896
rect 290822 39660 326266 39896
rect 326502 39660 326586 39896
rect 326822 39660 362266 39896
rect 362502 39660 362586 39896
rect 362822 39660 398266 39896
rect 398502 39660 398586 39896
rect 398822 39660 434266 39896
rect 434502 39660 434586 39896
rect 434822 39660 470266 39896
rect 470502 39660 470586 39896
rect 470822 39660 506266 39896
rect 506502 39660 506586 39896
rect 506822 39660 542266 39896
rect 542502 39660 542586 39896
rect 542822 39660 578266 39896
rect 578502 39660 578586 39896
rect 578822 39660 586302 39896
rect 586538 39660 586622 39896
rect 586858 39660 592650 39896
rect -8726 39576 592650 39660
rect -8726 39340 -2934 39576
rect -2698 39340 -2614 39576
rect -2378 39340 2266 39576
rect 2502 39340 2586 39576
rect 2822 39340 38266 39576
rect 38502 39340 38586 39576
rect 38822 39340 74266 39576
rect 74502 39340 74586 39576
rect 74822 39340 110266 39576
rect 110502 39340 110586 39576
rect 110822 39340 146266 39576
rect 146502 39340 146586 39576
rect 146822 39340 182266 39576
rect 182502 39340 182586 39576
rect 182822 39340 218266 39576
rect 218502 39340 218586 39576
rect 218822 39340 254266 39576
rect 254502 39340 254586 39576
rect 254822 39340 290266 39576
rect 290502 39340 290586 39576
rect 290822 39340 326266 39576
rect 326502 39340 326586 39576
rect 326822 39340 362266 39576
rect 362502 39340 362586 39576
rect 362822 39340 398266 39576
rect 398502 39340 398586 39576
rect 398822 39340 434266 39576
rect 434502 39340 434586 39576
rect 434822 39340 470266 39576
rect 470502 39340 470586 39576
rect 470822 39340 506266 39576
rect 506502 39340 506586 39576
rect 506822 39340 542266 39576
rect 542502 39340 542586 39576
rect 542822 39340 578266 39576
rect 578502 39340 578586 39576
rect 578822 39340 586302 39576
rect 586538 39340 586622 39576
rect 586858 39340 592650 39576
rect -8726 39308 592650 39340
rect -8726 38656 592650 38688
rect -8726 38420 -1974 38656
rect -1738 38420 -1654 38656
rect -1418 38420 1026 38656
rect 1262 38420 1346 38656
rect 1582 38420 37026 38656
rect 37262 38420 37346 38656
rect 37582 38420 73026 38656
rect 73262 38420 73346 38656
rect 73582 38420 109026 38656
rect 109262 38420 109346 38656
rect 109582 38420 145026 38656
rect 145262 38420 145346 38656
rect 145582 38420 181026 38656
rect 181262 38420 181346 38656
rect 181582 38420 217026 38656
rect 217262 38420 217346 38656
rect 217582 38420 253026 38656
rect 253262 38420 253346 38656
rect 253582 38420 289026 38656
rect 289262 38420 289346 38656
rect 289582 38420 325026 38656
rect 325262 38420 325346 38656
rect 325582 38420 361026 38656
rect 361262 38420 361346 38656
rect 361582 38420 397026 38656
rect 397262 38420 397346 38656
rect 397582 38420 433026 38656
rect 433262 38420 433346 38656
rect 433582 38420 469026 38656
rect 469262 38420 469346 38656
rect 469582 38420 505026 38656
rect 505262 38420 505346 38656
rect 505582 38420 541026 38656
rect 541262 38420 541346 38656
rect 541582 38420 577026 38656
rect 577262 38420 577346 38656
rect 577582 38420 585342 38656
rect 585578 38420 585662 38656
rect 585898 38420 592650 38656
rect -8726 38336 592650 38420
rect -8726 38100 -1974 38336
rect -1738 38100 -1654 38336
rect -1418 38100 1026 38336
rect 1262 38100 1346 38336
rect 1582 38100 37026 38336
rect 37262 38100 37346 38336
rect 37582 38100 73026 38336
rect 73262 38100 73346 38336
rect 73582 38100 109026 38336
rect 109262 38100 109346 38336
rect 109582 38100 145026 38336
rect 145262 38100 145346 38336
rect 145582 38100 181026 38336
rect 181262 38100 181346 38336
rect 181582 38100 217026 38336
rect 217262 38100 217346 38336
rect 217582 38100 253026 38336
rect 253262 38100 253346 38336
rect 253582 38100 289026 38336
rect 289262 38100 289346 38336
rect 289582 38100 325026 38336
rect 325262 38100 325346 38336
rect 325582 38100 361026 38336
rect 361262 38100 361346 38336
rect 361582 38100 397026 38336
rect 397262 38100 397346 38336
rect 397582 38100 433026 38336
rect 433262 38100 433346 38336
rect 433582 38100 469026 38336
rect 469262 38100 469346 38336
rect 469582 38100 505026 38336
rect 505262 38100 505346 38336
rect 505582 38100 541026 38336
rect 541262 38100 541346 38336
rect 541582 38100 577026 38336
rect 577262 38100 577346 38336
rect 577582 38100 585342 38336
rect 585578 38100 585662 38336
rect 585898 38100 592650 38336
rect -8726 38068 592650 38100
rect -8726 11336 592650 11368
rect -8726 11100 -8694 11336
rect -8458 11100 -8374 11336
rect -8138 11100 9706 11336
rect 9942 11100 10026 11336
rect 10262 11100 45706 11336
rect 45942 11100 46026 11336
rect 46262 11100 81706 11336
rect 81942 11100 82026 11336
rect 82262 11100 117706 11336
rect 117942 11100 118026 11336
rect 118262 11100 153706 11336
rect 153942 11100 154026 11336
rect 154262 11100 189706 11336
rect 189942 11100 190026 11336
rect 190262 11100 225706 11336
rect 225942 11100 226026 11336
rect 226262 11100 261706 11336
rect 261942 11100 262026 11336
rect 262262 11100 297706 11336
rect 297942 11100 298026 11336
rect 298262 11100 333706 11336
rect 333942 11100 334026 11336
rect 334262 11100 369706 11336
rect 369942 11100 370026 11336
rect 370262 11100 405706 11336
rect 405942 11100 406026 11336
rect 406262 11100 441706 11336
rect 441942 11100 442026 11336
rect 442262 11100 477706 11336
rect 477942 11100 478026 11336
rect 478262 11100 513706 11336
rect 513942 11100 514026 11336
rect 514262 11100 549706 11336
rect 549942 11100 550026 11336
rect 550262 11100 592062 11336
rect 592298 11100 592382 11336
rect 592618 11100 592650 11336
rect -8726 11016 592650 11100
rect -8726 10780 -8694 11016
rect -8458 10780 -8374 11016
rect -8138 10780 9706 11016
rect 9942 10780 10026 11016
rect 10262 10780 45706 11016
rect 45942 10780 46026 11016
rect 46262 10780 81706 11016
rect 81942 10780 82026 11016
rect 82262 10780 117706 11016
rect 117942 10780 118026 11016
rect 118262 10780 153706 11016
rect 153942 10780 154026 11016
rect 154262 10780 189706 11016
rect 189942 10780 190026 11016
rect 190262 10780 225706 11016
rect 225942 10780 226026 11016
rect 226262 10780 261706 11016
rect 261942 10780 262026 11016
rect 262262 10780 297706 11016
rect 297942 10780 298026 11016
rect 298262 10780 333706 11016
rect 333942 10780 334026 11016
rect 334262 10780 369706 11016
rect 369942 10780 370026 11016
rect 370262 10780 405706 11016
rect 405942 10780 406026 11016
rect 406262 10780 441706 11016
rect 441942 10780 442026 11016
rect 442262 10780 477706 11016
rect 477942 10780 478026 11016
rect 478262 10780 513706 11016
rect 513942 10780 514026 11016
rect 514262 10780 549706 11016
rect 549942 10780 550026 11016
rect 550262 10780 592062 11016
rect 592298 10780 592382 11016
rect 592618 10780 592650 11016
rect -8726 10748 592650 10780
rect -8726 10096 592650 10128
rect -8726 9860 -7734 10096
rect -7498 9860 -7414 10096
rect -7178 9860 8466 10096
rect 8702 9860 8786 10096
rect 9022 9860 44466 10096
rect 44702 9860 44786 10096
rect 45022 9860 80466 10096
rect 80702 9860 80786 10096
rect 81022 9860 116466 10096
rect 116702 9860 116786 10096
rect 117022 9860 152466 10096
rect 152702 9860 152786 10096
rect 153022 9860 188466 10096
rect 188702 9860 188786 10096
rect 189022 9860 224466 10096
rect 224702 9860 224786 10096
rect 225022 9860 260466 10096
rect 260702 9860 260786 10096
rect 261022 9860 296466 10096
rect 296702 9860 296786 10096
rect 297022 9860 332466 10096
rect 332702 9860 332786 10096
rect 333022 9860 368466 10096
rect 368702 9860 368786 10096
rect 369022 9860 404466 10096
rect 404702 9860 404786 10096
rect 405022 9860 440466 10096
rect 440702 9860 440786 10096
rect 441022 9860 476466 10096
rect 476702 9860 476786 10096
rect 477022 9860 512466 10096
rect 512702 9860 512786 10096
rect 513022 9860 548466 10096
rect 548702 9860 548786 10096
rect 549022 9860 591102 10096
rect 591338 9860 591422 10096
rect 591658 9860 592650 10096
rect -8726 9776 592650 9860
rect -8726 9540 -7734 9776
rect -7498 9540 -7414 9776
rect -7178 9540 8466 9776
rect 8702 9540 8786 9776
rect 9022 9540 44466 9776
rect 44702 9540 44786 9776
rect 45022 9540 80466 9776
rect 80702 9540 80786 9776
rect 81022 9540 116466 9776
rect 116702 9540 116786 9776
rect 117022 9540 152466 9776
rect 152702 9540 152786 9776
rect 153022 9540 188466 9776
rect 188702 9540 188786 9776
rect 189022 9540 224466 9776
rect 224702 9540 224786 9776
rect 225022 9540 260466 9776
rect 260702 9540 260786 9776
rect 261022 9540 296466 9776
rect 296702 9540 296786 9776
rect 297022 9540 332466 9776
rect 332702 9540 332786 9776
rect 333022 9540 368466 9776
rect 368702 9540 368786 9776
rect 369022 9540 404466 9776
rect 404702 9540 404786 9776
rect 405022 9540 440466 9776
rect 440702 9540 440786 9776
rect 441022 9540 476466 9776
rect 476702 9540 476786 9776
rect 477022 9540 512466 9776
rect 512702 9540 512786 9776
rect 513022 9540 548466 9776
rect 548702 9540 548786 9776
rect 549022 9540 591102 9776
rect 591338 9540 591422 9776
rect 591658 9540 592650 9776
rect -8726 9508 592650 9540
rect -8726 8856 592650 8888
rect -8726 8620 -6774 8856
rect -6538 8620 -6454 8856
rect -6218 8620 7226 8856
rect 7462 8620 7546 8856
rect 7782 8620 43226 8856
rect 43462 8620 43546 8856
rect 43782 8620 79226 8856
rect 79462 8620 79546 8856
rect 79782 8620 115226 8856
rect 115462 8620 115546 8856
rect 115782 8620 151226 8856
rect 151462 8620 151546 8856
rect 151782 8620 187226 8856
rect 187462 8620 187546 8856
rect 187782 8620 223226 8856
rect 223462 8620 223546 8856
rect 223782 8620 259226 8856
rect 259462 8620 259546 8856
rect 259782 8620 295226 8856
rect 295462 8620 295546 8856
rect 295782 8620 331226 8856
rect 331462 8620 331546 8856
rect 331782 8620 367226 8856
rect 367462 8620 367546 8856
rect 367782 8620 403226 8856
rect 403462 8620 403546 8856
rect 403782 8620 439226 8856
rect 439462 8620 439546 8856
rect 439782 8620 475226 8856
rect 475462 8620 475546 8856
rect 475782 8620 511226 8856
rect 511462 8620 511546 8856
rect 511782 8620 547226 8856
rect 547462 8620 547546 8856
rect 547782 8620 590142 8856
rect 590378 8620 590462 8856
rect 590698 8620 592650 8856
rect -8726 8536 592650 8620
rect -8726 8300 -6774 8536
rect -6538 8300 -6454 8536
rect -6218 8300 7226 8536
rect 7462 8300 7546 8536
rect 7782 8300 43226 8536
rect 43462 8300 43546 8536
rect 43782 8300 79226 8536
rect 79462 8300 79546 8536
rect 79782 8300 115226 8536
rect 115462 8300 115546 8536
rect 115782 8300 151226 8536
rect 151462 8300 151546 8536
rect 151782 8300 187226 8536
rect 187462 8300 187546 8536
rect 187782 8300 223226 8536
rect 223462 8300 223546 8536
rect 223782 8300 259226 8536
rect 259462 8300 259546 8536
rect 259782 8300 295226 8536
rect 295462 8300 295546 8536
rect 295782 8300 331226 8536
rect 331462 8300 331546 8536
rect 331782 8300 367226 8536
rect 367462 8300 367546 8536
rect 367782 8300 403226 8536
rect 403462 8300 403546 8536
rect 403782 8300 439226 8536
rect 439462 8300 439546 8536
rect 439782 8300 475226 8536
rect 475462 8300 475546 8536
rect 475782 8300 511226 8536
rect 511462 8300 511546 8536
rect 511782 8300 547226 8536
rect 547462 8300 547546 8536
rect 547782 8300 590142 8536
rect 590378 8300 590462 8536
rect 590698 8300 592650 8536
rect -8726 8268 592650 8300
rect -8726 7616 592650 7648
rect -8726 7380 -5814 7616
rect -5578 7380 -5494 7616
rect -5258 7380 5986 7616
rect 6222 7380 6306 7616
rect 6542 7380 41986 7616
rect 42222 7380 42306 7616
rect 42542 7380 77986 7616
rect 78222 7380 78306 7616
rect 78542 7380 113986 7616
rect 114222 7380 114306 7616
rect 114542 7380 149986 7616
rect 150222 7380 150306 7616
rect 150542 7380 185986 7616
rect 186222 7380 186306 7616
rect 186542 7380 221986 7616
rect 222222 7380 222306 7616
rect 222542 7380 257986 7616
rect 258222 7380 258306 7616
rect 258542 7380 293986 7616
rect 294222 7380 294306 7616
rect 294542 7380 329986 7616
rect 330222 7380 330306 7616
rect 330542 7380 365986 7616
rect 366222 7380 366306 7616
rect 366542 7380 401986 7616
rect 402222 7380 402306 7616
rect 402542 7380 437986 7616
rect 438222 7380 438306 7616
rect 438542 7380 473986 7616
rect 474222 7380 474306 7616
rect 474542 7380 509986 7616
rect 510222 7380 510306 7616
rect 510542 7380 545986 7616
rect 546222 7380 546306 7616
rect 546542 7380 581986 7616
rect 582222 7380 582306 7616
rect 582542 7380 589182 7616
rect 589418 7380 589502 7616
rect 589738 7380 592650 7616
rect -8726 7296 592650 7380
rect -8726 7060 -5814 7296
rect -5578 7060 -5494 7296
rect -5258 7060 5986 7296
rect 6222 7060 6306 7296
rect 6542 7060 41986 7296
rect 42222 7060 42306 7296
rect 42542 7060 77986 7296
rect 78222 7060 78306 7296
rect 78542 7060 113986 7296
rect 114222 7060 114306 7296
rect 114542 7060 149986 7296
rect 150222 7060 150306 7296
rect 150542 7060 185986 7296
rect 186222 7060 186306 7296
rect 186542 7060 221986 7296
rect 222222 7060 222306 7296
rect 222542 7060 257986 7296
rect 258222 7060 258306 7296
rect 258542 7060 293986 7296
rect 294222 7060 294306 7296
rect 294542 7060 329986 7296
rect 330222 7060 330306 7296
rect 330542 7060 365986 7296
rect 366222 7060 366306 7296
rect 366542 7060 401986 7296
rect 402222 7060 402306 7296
rect 402542 7060 437986 7296
rect 438222 7060 438306 7296
rect 438542 7060 473986 7296
rect 474222 7060 474306 7296
rect 474542 7060 509986 7296
rect 510222 7060 510306 7296
rect 510542 7060 545986 7296
rect 546222 7060 546306 7296
rect 546542 7060 581986 7296
rect 582222 7060 582306 7296
rect 582542 7060 589182 7296
rect 589418 7060 589502 7296
rect 589738 7060 592650 7296
rect -8726 7028 592650 7060
rect -8726 6376 592650 6408
rect -8726 6140 -4854 6376
rect -4618 6140 -4534 6376
rect -4298 6140 4746 6376
rect 4982 6140 5066 6376
rect 5302 6140 40746 6376
rect 40982 6140 41066 6376
rect 41302 6140 76746 6376
rect 76982 6140 77066 6376
rect 77302 6140 112746 6376
rect 112982 6140 113066 6376
rect 113302 6140 148746 6376
rect 148982 6140 149066 6376
rect 149302 6140 184746 6376
rect 184982 6140 185066 6376
rect 185302 6140 220746 6376
rect 220982 6140 221066 6376
rect 221302 6140 256746 6376
rect 256982 6140 257066 6376
rect 257302 6140 292746 6376
rect 292982 6140 293066 6376
rect 293302 6140 328746 6376
rect 328982 6140 329066 6376
rect 329302 6140 364746 6376
rect 364982 6140 365066 6376
rect 365302 6140 400746 6376
rect 400982 6140 401066 6376
rect 401302 6140 436746 6376
rect 436982 6140 437066 6376
rect 437302 6140 472746 6376
rect 472982 6140 473066 6376
rect 473302 6140 508746 6376
rect 508982 6140 509066 6376
rect 509302 6140 544746 6376
rect 544982 6140 545066 6376
rect 545302 6140 580746 6376
rect 580982 6140 581066 6376
rect 581302 6140 588222 6376
rect 588458 6140 588542 6376
rect 588778 6140 592650 6376
rect -8726 6056 592650 6140
rect -8726 5820 -4854 6056
rect -4618 5820 -4534 6056
rect -4298 5820 4746 6056
rect 4982 5820 5066 6056
rect 5302 5820 40746 6056
rect 40982 5820 41066 6056
rect 41302 5820 76746 6056
rect 76982 5820 77066 6056
rect 77302 5820 112746 6056
rect 112982 5820 113066 6056
rect 113302 5820 148746 6056
rect 148982 5820 149066 6056
rect 149302 5820 184746 6056
rect 184982 5820 185066 6056
rect 185302 5820 220746 6056
rect 220982 5820 221066 6056
rect 221302 5820 256746 6056
rect 256982 5820 257066 6056
rect 257302 5820 292746 6056
rect 292982 5820 293066 6056
rect 293302 5820 328746 6056
rect 328982 5820 329066 6056
rect 329302 5820 364746 6056
rect 364982 5820 365066 6056
rect 365302 5820 400746 6056
rect 400982 5820 401066 6056
rect 401302 5820 436746 6056
rect 436982 5820 437066 6056
rect 437302 5820 472746 6056
rect 472982 5820 473066 6056
rect 473302 5820 508746 6056
rect 508982 5820 509066 6056
rect 509302 5820 544746 6056
rect 544982 5820 545066 6056
rect 545302 5820 580746 6056
rect 580982 5820 581066 6056
rect 581302 5820 588222 6056
rect 588458 5820 588542 6056
rect 588778 5820 592650 6056
rect -8726 5788 592650 5820
rect -8726 5136 592650 5168
rect -8726 4900 -3894 5136
rect -3658 4900 -3574 5136
rect -3338 4900 3506 5136
rect 3742 4900 3826 5136
rect 4062 4900 39506 5136
rect 39742 4900 39826 5136
rect 40062 4900 75506 5136
rect 75742 4900 75826 5136
rect 76062 4900 111506 5136
rect 111742 4900 111826 5136
rect 112062 4900 147506 5136
rect 147742 4900 147826 5136
rect 148062 4900 183506 5136
rect 183742 4900 183826 5136
rect 184062 4900 219506 5136
rect 219742 4900 219826 5136
rect 220062 4900 255506 5136
rect 255742 4900 255826 5136
rect 256062 4900 291506 5136
rect 291742 4900 291826 5136
rect 292062 4900 327506 5136
rect 327742 4900 327826 5136
rect 328062 4900 363506 5136
rect 363742 4900 363826 5136
rect 364062 4900 399506 5136
rect 399742 4900 399826 5136
rect 400062 4900 435506 5136
rect 435742 4900 435826 5136
rect 436062 4900 471506 5136
rect 471742 4900 471826 5136
rect 472062 4900 507506 5136
rect 507742 4900 507826 5136
rect 508062 4900 543506 5136
rect 543742 4900 543826 5136
rect 544062 4900 579506 5136
rect 579742 4900 579826 5136
rect 580062 4900 587262 5136
rect 587498 4900 587582 5136
rect 587818 4900 592650 5136
rect -8726 4816 592650 4900
rect -8726 4580 -3894 4816
rect -3658 4580 -3574 4816
rect -3338 4580 3506 4816
rect 3742 4580 3826 4816
rect 4062 4580 39506 4816
rect 39742 4580 39826 4816
rect 40062 4580 75506 4816
rect 75742 4580 75826 4816
rect 76062 4580 111506 4816
rect 111742 4580 111826 4816
rect 112062 4580 147506 4816
rect 147742 4580 147826 4816
rect 148062 4580 183506 4816
rect 183742 4580 183826 4816
rect 184062 4580 219506 4816
rect 219742 4580 219826 4816
rect 220062 4580 255506 4816
rect 255742 4580 255826 4816
rect 256062 4580 291506 4816
rect 291742 4580 291826 4816
rect 292062 4580 327506 4816
rect 327742 4580 327826 4816
rect 328062 4580 363506 4816
rect 363742 4580 363826 4816
rect 364062 4580 399506 4816
rect 399742 4580 399826 4816
rect 400062 4580 435506 4816
rect 435742 4580 435826 4816
rect 436062 4580 471506 4816
rect 471742 4580 471826 4816
rect 472062 4580 507506 4816
rect 507742 4580 507826 4816
rect 508062 4580 543506 4816
rect 543742 4580 543826 4816
rect 544062 4580 579506 4816
rect 579742 4580 579826 4816
rect 580062 4580 587262 4816
rect 587498 4580 587582 4816
rect 587818 4580 592650 4816
rect -8726 4548 592650 4580
rect -8726 3896 592650 3928
rect -8726 3660 -2934 3896
rect -2698 3660 -2614 3896
rect -2378 3660 2266 3896
rect 2502 3660 2586 3896
rect 2822 3660 38266 3896
rect 38502 3660 38586 3896
rect 38822 3660 74266 3896
rect 74502 3660 74586 3896
rect 74822 3660 110266 3896
rect 110502 3660 110586 3896
rect 110822 3660 146266 3896
rect 146502 3660 146586 3896
rect 146822 3660 182266 3896
rect 182502 3660 182586 3896
rect 182822 3660 218266 3896
rect 218502 3660 218586 3896
rect 218822 3660 254266 3896
rect 254502 3660 254586 3896
rect 254822 3660 290266 3896
rect 290502 3660 290586 3896
rect 290822 3660 326266 3896
rect 326502 3660 326586 3896
rect 326822 3660 362266 3896
rect 362502 3660 362586 3896
rect 362822 3660 398266 3896
rect 398502 3660 398586 3896
rect 398822 3660 434266 3896
rect 434502 3660 434586 3896
rect 434822 3660 470266 3896
rect 470502 3660 470586 3896
rect 470822 3660 506266 3896
rect 506502 3660 506586 3896
rect 506822 3660 542266 3896
rect 542502 3660 542586 3896
rect 542822 3660 578266 3896
rect 578502 3660 578586 3896
rect 578822 3660 586302 3896
rect 586538 3660 586622 3896
rect 586858 3660 592650 3896
rect -8726 3576 592650 3660
rect -8726 3340 -2934 3576
rect -2698 3340 -2614 3576
rect -2378 3340 2266 3576
rect 2502 3340 2586 3576
rect 2822 3340 38266 3576
rect 38502 3340 38586 3576
rect 38822 3340 74266 3576
rect 74502 3340 74586 3576
rect 74822 3340 110266 3576
rect 110502 3340 110586 3576
rect 110822 3340 146266 3576
rect 146502 3340 146586 3576
rect 146822 3340 182266 3576
rect 182502 3340 182586 3576
rect 182822 3340 218266 3576
rect 218502 3340 218586 3576
rect 218822 3340 254266 3576
rect 254502 3340 254586 3576
rect 254822 3340 290266 3576
rect 290502 3340 290586 3576
rect 290822 3340 326266 3576
rect 326502 3340 326586 3576
rect 326822 3340 362266 3576
rect 362502 3340 362586 3576
rect 362822 3340 398266 3576
rect 398502 3340 398586 3576
rect 398822 3340 434266 3576
rect 434502 3340 434586 3576
rect 434822 3340 470266 3576
rect 470502 3340 470586 3576
rect 470822 3340 506266 3576
rect 506502 3340 506586 3576
rect 506822 3340 542266 3576
rect 542502 3340 542586 3576
rect 542822 3340 578266 3576
rect 578502 3340 578586 3576
rect 578822 3340 586302 3576
rect 586538 3340 586622 3576
rect 586858 3340 592650 3576
rect -8726 3308 592650 3340
rect -8726 2656 592650 2688
rect -8726 2420 -1974 2656
rect -1738 2420 -1654 2656
rect -1418 2420 1026 2656
rect 1262 2420 1346 2656
rect 1582 2420 37026 2656
rect 37262 2420 37346 2656
rect 37582 2420 73026 2656
rect 73262 2420 73346 2656
rect 73582 2420 109026 2656
rect 109262 2420 109346 2656
rect 109582 2420 145026 2656
rect 145262 2420 145346 2656
rect 145582 2420 181026 2656
rect 181262 2420 181346 2656
rect 181582 2420 217026 2656
rect 217262 2420 217346 2656
rect 217582 2420 253026 2656
rect 253262 2420 253346 2656
rect 253582 2420 289026 2656
rect 289262 2420 289346 2656
rect 289582 2420 325026 2656
rect 325262 2420 325346 2656
rect 325582 2420 361026 2656
rect 361262 2420 361346 2656
rect 361582 2420 397026 2656
rect 397262 2420 397346 2656
rect 397582 2420 433026 2656
rect 433262 2420 433346 2656
rect 433582 2420 469026 2656
rect 469262 2420 469346 2656
rect 469582 2420 505026 2656
rect 505262 2420 505346 2656
rect 505582 2420 541026 2656
rect 541262 2420 541346 2656
rect 541582 2420 577026 2656
rect 577262 2420 577346 2656
rect 577582 2420 585342 2656
rect 585578 2420 585662 2656
rect 585898 2420 592650 2656
rect -8726 2336 592650 2420
rect -8726 2100 -1974 2336
rect -1738 2100 -1654 2336
rect -1418 2100 1026 2336
rect 1262 2100 1346 2336
rect 1582 2100 37026 2336
rect 37262 2100 37346 2336
rect 37582 2100 73026 2336
rect 73262 2100 73346 2336
rect 73582 2100 109026 2336
rect 109262 2100 109346 2336
rect 109582 2100 145026 2336
rect 145262 2100 145346 2336
rect 145582 2100 181026 2336
rect 181262 2100 181346 2336
rect 181582 2100 217026 2336
rect 217262 2100 217346 2336
rect 217582 2100 253026 2336
rect 253262 2100 253346 2336
rect 253582 2100 289026 2336
rect 289262 2100 289346 2336
rect 289582 2100 325026 2336
rect 325262 2100 325346 2336
rect 325582 2100 361026 2336
rect 361262 2100 361346 2336
rect 361582 2100 397026 2336
rect 397262 2100 397346 2336
rect 397582 2100 433026 2336
rect 433262 2100 433346 2336
rect 433582 2100 469026 2336
rect 469262 2100 469346 2336
rect 469582 2100 505026 2336
rect 505262 2100 505346 2336
rect 505582 2100 541026 2336
rect 541262 2100 541346 2336
rect 541582 2100 577026 2336
rect 577262 2100 577346 2336
rect 577582 2100 585342 2336
rect 585578 2100 585662 2336
rect 585898 2100 592650 2336
rect -8726 2068 592650 2100
rect -2006 -344 585930 -312
rect -2006 -580 -1974 -344
rect -1738 -580 -1654 -344
rect -1418 -580 1026 -344
rect 1262 -580 1346 -344
rect 1582 -580 37026 -344
rect 37262 -580 37346 -344
rect 37582 -580 73026 -344
rect 73262 -580 73346 -344
rect 73582 -580 109026 -344
rect 109262 -580 109346 -344
rect 109582 -580 145026 -344
rect 145262 -580 145346 -344
rect 145582 -580 181026 -344
rect 181262 -580 181346 -344
rect 181582 -580 217026 -344
rect 217262 -580 217346 -344
rect 217582 -580 253026 -344
rect 253262 -580 253346 -344
rect 253582 -580 289026 -344
rect 289262 -580 289346 -344
rect 289582 -580 325026 -344
rect 325262 -580 325346 -344
rect 325582 -580 361026 -344
rect 361262 -580 361346 -344
rect 361582 -580 397026 -344
rect 397262 -580 397346 -344
rect 397582 -580 433026 -344
rect 433262 -580 433346 -344
rect 433582 -580 469026 -344
rect 469262 -580 469346 -344
rect 469582 -580 505026 -344
rect 505262 -580 505346 -344
rect 505582 -580 541026 -344
rect 541262 -580 541346 -344
rect 541582 -580 577026 -344
rect 577262 -580 577346 -344
rect 577582 -580 585342 -344
rect 585578 -580 585662 -344
rect 585898 -580 585930 -344
rect -2006 -664 585930 -580
rect -2006 -900 -1974 -664
rect -1738 -900 -1654 -664
rect -1418 -900 1026 -664
rect 1262 -900 1346 -664
rect 1582 -900 37026 -664
rect 37262 -900 37346 -664
rect 37582 -900 73026 -664
rect 73262 -900 73346 -664
rect 73582 -900 109026 -664
rect 109262 -900 109346 -664
rect 109582 -900 145026 -664
rect 145262 -900 145346 -664
rect 145582 -900 181026 -664
rect 181262 -900 181346 -664
rect 181582 -900 217026 -664
rect 217262 -900 217346 -664
rect 217582 -900 253026 -664
rect 253262 -900 253346 -664
rect 253582 -900 289026 -664
rect 289262 -900 289346 -664
rect 289582 -900 325026 -664
rect 325262 -900 325346 -664
rect 325582 -900 361026 -664
rect 361262 -900 361346 -664
rect 361582 -900 397026 -664
rect 397262 -900 397346 -664
rect 397582 -900 433026 -664
rect 433262 -900 433346 -664
rect 433582 -900 469026 -664
rect 469262 -900 469346 -664
rect 469582 -900 505026 -664
rect 505262 -900 505346 -664
rect 505582 -900 541026 -664
rect 541262 -900 541346 -664
rect 541582 -900 577026 -664
rect 577262 -900 577346 -664
rect 577582 -900 585342 -664
rect 585578 -900 585662 -664
rect 585898 -900 585930 -664
rect -2006 -932 585930 -900
rect -2966 -1304 586890 -1272
rect -2966 -1540 -2934 -1304
rect -2698 -1540 -2614 -1304
rect -2378 -1540 2266 -1304
rect 2502 -1540 2586 -1304
rect 2822 -1540 38266 -1304
rect 38502 -1540 38586 -1304
rect 38822 -1540 74266 -1304
rect 74502 -1540 74586 -1304
rect 74822 -1540 110266 -1304
rect 110502 -1540 110586 -1304
rect 110822 -1540 146266 -1304
rect 146502 -1540 146586 -1304
rect 146822 -1540 182266 -1304
rect 182502 -1540 182586 -1304
rect 182822 -1540 218266 -1304
rect 218502 -1540 218586 -1304
rect 218822 -1540 254266 -1304
rect 254502 -1540 254586 -1304
rect 254822 -1540 290266 -1304
rect 290502 -1540 290586 -1304
rect 290822 -1540 326266 -1304
rect 326502 -1540 326586 -1304
rect 326822 -1540 362266 -1304
rect 362502 -1540 362586 -1304
rect 362822 -1540 398266 -1304
rect 398502 -1540 398586 -1304
rect 398822 -1540 434266 -1304
rect 434502 -1540 434586 -1304
rect 434822 -1540 470266 -1304
rect 470502 -1540 470586 -1304
rect 470822 -1540 506266 -1304
rect 506502 -1540 506586 -1304
rect 506822 -1540 542266 -1304
rect 542502 -1540 542586 -1304
rect 542822 -1540 578266 -1304
rect 578502 -1540 578586 -1304
rect 578822 -1540 586302 -1304
rect 586538 -1540 586622 -1304
rect 586858 -1540 586890 -1304
rect -2966 -1624 586890 -1540
rect -2966 -1860 -2934 -1624
rect -2698 -1860 -2614 -1624
rect -2378 -1860 2266 -1624
rect 2502 -1860 2586 -1624
rect 2822 -1860 38266 -1624
rect 38502 -1860 38586 -1624
rect 38822 -1860 74266 -1624
rect 74502 -1860 74586 -1624
rect 74822 -1860 110266 -1624
rect 110502 -1860 110586 -1624
rect 110822 -1860 146266 -1624
rect 146502 -1860 146586 -1624
rect 146822 -1860 182266 -1624
rect 182502 -1860 182586 -1624
rect 182822 -1860 218266 -1624
rect 218502 -1860 218586 -1624
rect 218822 -1860 254266 -1624
rect 254502 -1860 254586 -1624
rect 254822 -1860 290266 -1624
rect 290502 -1860 290586 -1624
rect 290822 -1860 326266 -1624
rect 326502 -1860 326586 -1624
rect 326822 -1860 362266 -1624
rect 362502 -1860 362586 -1624
rect 362822 -1860 398266 -1624
rect 398502 -1860 398586 -1624
rect 398822 -1860 434266 -1624
rect 434502 -1860 434586 -1624
rect 434822 -1860 470266 -1624
rect 470502 -1860 470586 -1624
rect 470822 -1860 506266 -1624
rect 506502 -1860 506586 -1624
rect 506822 -1860 542266 -1624
rect 542502 -1860 542586 -1624
rect 542822 -1860 578266 -1624
rect 578502 -1860 578586 -1624
rect 578822 -1860 586302 -1624
rect 586538 -1860 586622 -1624
rect 586858 -1860 586890 -1624
rect -2966 -1892 586890 -1860
rect -3926 -2264 587850 -2232
rect -3926 -2500 -3894 -2264
rect -3658 -2500 -3574 -2264
rect -3338 -2500 3506 -2264
rect 3742 -2500 3826 -2264
rect 4062 -2500 39506 -2264
rect 39742 -2500 39826 -2264
rect 40062 -2500 75506 -2264
rect 75742 -2500 75826 -2264
rect 76062 -2500 111506 -2264
rect 111742 -2500 111826 -2264
rect 112062 -2500 147506 -2264
rect 147742 -2500 147826 -2264
rect 148062 -2500 183506 -2264
rect 183742 -2500 183826 -2264
rect 184062 -2500 219506 -2264
rect 219742 -2500 219826 -2264
rect 220062 -2500 255506 -2264
rect 255742 -2500 255826 -2264
rect 256062 -2500 291506 -2264
rect 291742 -2500 291826 -2264
rect 292062 -2500 327506 -2264
rect 327742 -2500 327826 -2264
rect 328062 -2500 363506 -2264
rect 363742 -2500 363826 -2264
rect 364062 -2500 399506 -2264
rect 399742 -2500 399826 -2264
rect 400062 -2500 435506 -2264
rect 435742 -2500 435826 -2264
rect 436062 -2500 471506 -2264
rect 471742 -2500 471826 -2264
rect 472062 -2500 507506 -2264
rect 507742 -2500 507826 -2264
rect 508062 -2500 543506 -2264
rect 543742 -2500 543826 -2264
rect 544062 -2500 579506 -2264
rect 579742 -2500 579826 -2264
rect 580062 -2500 587262 -2264
rect 587498 -2500 587582 -2264
rect 587818 -2500 587850 -2264
rect -3926 -2584 587850 -2500
rect -3926 -2820 -3894 -2584
rect -3658 -2820 -3574 -2584
rect -3338 -2820 3506 -2584
rect 3742 -2820 3826 -2584
rect 4062 -2820 39506 -2584
rect 39742 -2820 39826 -2584
rect 40062 -2820 75506 -2584
rect 75742 -2820 75826 -2584
rect 76062 -2820 111506 -2584
rect 111742 -2820 111826 -2584
rect 112062 -2820 147506 -2584
rect 147742 -2820 147826 -2584
rect 148062 -2820 183506 -2584
rect 183742 -2820 183826 -2584
rect 184062 -2820 219506 -2584
rect 219742 -2820 219826 -2584
rect 220062 -2820 255506 -2584
rect 255742 -2820 255826 -2584
rect 256062 -2820 291506 -2584
rect 291742 -2820 291826 -2584
rect 292062 -2820 327506 -2584
rect 327742 -2820 327826 -2584
rect 328062 -2820 363506 -2584
rect 363742 -2820 363826 -2584
rect 364062 -2820 399506 -2584
rect 399742 -2820 399826 -2584
rect 400062 -2820 435506 -2584
rect 435742 -2820 435826 -2584
rect 436062 -2820 471506 -2584
rect 471742 -2820 471826 -2584
rect 472062 -2820 507506 -2584
rect 507742 -2820 507826 -2584
rect 508062 -2820 543506 -2584
rect 543742 -2820 543826 -2584
rect 544062 -2820 579506 -2584
rect 579742 -2820 579826 -2584
rect 580062 -2820 587262 -2584
rect 587498 -2820 587582 -2584
rect 587818 -2820 587850 -2584
rect -3926 -2852 587850 -2820
rect -4886 -3224 588810 -3192
rect -4886 -3460 -4854 -3224
rect -4618 -3460 -4534 -3224
rect -4298 -3460 4746 -3224
rect 4982 -3460 5066 -3224
rect 5302 -3460 40746 -3224
rect 40982 -3460 41066 -3224
rect 41302 -3460 76746 -3224
rect 76982 -3460 77066 -3224
rect 77302 -3460 112746 -3224
rect 112982 -3460 113066 -3224
rect 113302 -3460 148746 -3224
rect 148982 -3460 149066 -3224
rect 149302 -3460 184746 -3224
rect 184982 -3460 185066 -3224
rect 185302 -3460 220746 -3224
rect 220982 -3460 221066 -3224
rect 221302 -3460 256746 -3224
rect 256982 -3460 257066 -3224
rect 257302 -3460 292746 -3224
rect 292982 -3460 293066 -3224
rect 293302 -3460 328746 -3224
rect 328982 -3460 329066 -3224
rect 329302 -3460 364746 -3224
rect 364982 -3460 365066 -3224
rect 365302 -3460 400746 -3224
rect 400982 -3460 401066 -3224
rect 401302 -3460 436746 -3224
rect 436982 -3460 437066 -3224
rect 437302 -3460 472746 -3224
rect 472982 -3460 473066 -3224
rect 473302 -3460 508746 -3224
rect 508982 -3460 509066 -3224
rect 509302 -3460 544746 -3224
rect 544982 -3460 545066 -3224
rect 545302 -3460 580746 -3224
rect 580982 -3460 581066 -3224
rect 581302 -3460 588222 -3224
rect 588458 -3460 588542 -3224
rect 588778 -3460 588810 -3224
rect -4886 -3544 588810 -3460
rect -4886 -3780 -4854 -3544
rect -4618 -3780 -4534 -3544
rect -4298 -3780 4746 -3544
rect 4982 -3780 5066 -3544
rect 5302 -3780 40746 -3544
rect 40982 -3780 41066 -3544
rect 41302 -3780 76746 -3544
rect 76982 -3780 77066 -3544
rect 77302 -3780 112746 -3544
rect 112982 -3780 113066 -3544
rect 113302 -3780 148746 -3544
rect 148982 -3780 149066 -3544
rect 149302 -3780 184746 -3544
rect 184982 -3780 185066 -3544
rect 185302 -3780 220746 -3544
rect 220982 -3780 221066 -3544
rect 221302 -3780 256746 -3544
rect 256982 -3780 257066 -3544
rect 257302 -3780 292746 -3544
rect 292982 -3780 293066 -3544
rect 293302 -3780 328746 -3544
rect 328982 -3780 329066 -3544
rect 329302 -3780 364746 -3544
rect 364982 -3780 365066 -3544
rect 365302 -3780 400746 -3544
rect 400982 -3780 401066 -3544
rect 401302 -3780 436746 -3544
rect 436982 -3780 437066 -3544
rect 437302 -3780 472746 -3544
rect 472982 -3780 473066 -3544
rect 473302 -3780 508746 -3544
rect 508982 -3780 509066 -3544
rect 509302 -3780 544746 -3544
rect 544982 -3780 545066 -3544
rect 545302 -3780 580746 -3544
rect 580982 -3780 581066 -3544
rect 581302 -3780 588222 -3544
rect 588458 -3780 588542 -3544
rect 588778 -3780 588810 -3544
rect -4886 -3812 588810 -3780
rect -5846 -4184 589770 -4152
rect -5846 -4420 -5814 -4184
rect -5578 -4420 -5494 -4184
rect -5258 -4420 5986 -4184
rect 6222 -4420 6306 -4184
rect 6542 -4420 41986 -4184
rect 42222 -4420 42306 -4184
rect 42542 -4420 77986 -4184
rect 78222 -4420 78306 -4184
rect 78542 -4420 113986 -4184
rect 114222 -4420 114306 -4184
rect 114542 -4420 149986 -4184
rect 150222 -4420 150306 -4184
rect 150542 -4420 185986 -4184
rect 186222 -4420 186306 -4184
rect 186542 -4420 221986 -4184
rect 222222 -4420 222306 -4184
rect 222542 -4420 257986 -4184
rect 258222 -4420 258306 -4184
rect 258542 -4420 293986 -4184
rect 294222 -4420 294306 -4184
rect 294542 -4420 329986 -4184
rect 330222 -4420 330306 -4184
rect 330542 -4420 365986 -4184
rect 366222 -4420 366306 -4184
rect 366542 -4420 401986 -4184
rect 402222 -4420 402306 -4184
rect 402542 -4420 437986 -4184
rect 438222 -4420 438306 -4184
rect 438542 -4420 473986 -4184
rect 474222 -4420 474306 -4184
rect 474542 -4420 509986 -4184
rect 510222 -4420 510306 -4184
rect 510542 -4420 545986 -4184
rect 546222 -4420 546306 -4184
rect 546542 -4420 581986 -4184
rect 582222 -4420 582306 -4184
rect 582542 -4420 589182 -4184
rect 589418 -4420 589502 -4184
rect 589738 -4420 589770 -4184
rect -5846 -4504 589770 -4420
rect -5846 -4740 -5814 -4504
rect -5578 -4740 -5494 -4504
rect -5258 -4740 5986 -4504
rect 6222 -4740 6306 -4504
rect 6542 -4740 41986 -4504
rect 42222 -4740 42306 -4504
rect 42542 -4740 77986 -4504
rect 78222 -4740 78306 -4504
rect 78542 -4740 113986 -4504
rect 114222 -4740 114306 -4504
rect 114542 -4740 149986 -4504
rect 150222 -4740 150306 -4504
rect 150542 -4740 185986 -4504
rect 186222 -4740 186306 -4504
rect 186542 -4740 221986 -4504
rect 222222 -4740 222306 -4504
rect 222542 -4740 257986 -4504
rect 258222 -4740 258306 -4504
rect 258542 -4740 293986 -4504
rect 294222 -4740 294306 -4504
rect 294542 -4740 329986 -4504
rect 330222 -4740 330306 -4504
rect 330542 -4740 365986 -4504
rect 366222 -4740 366306 -4504
rect 366542 -4740 401986 -4504
rect 402222 -4740 402306 -4504
rect 402542 -4740 437986 -4504
rect 438222 -4740 438306 -4504
rect 438542 -4740 473986 -4504
rect 474222 -4740 474306 -4504
rect 474542 -4740 509986 -4504
rect 510222 -4740 510306 -4504
rect 510542 -4740 545986 -4504
rect 546222 -4740 546306 -4504
rect 546542 -4740 581986 -4504
rect 582222 -4740 582306 -4504
rect 582542 -4740 589182 -4504
rect 589418 -4740 589502 -4504
rect 589738 -4740 589770 -4504
rect -5846 -4772 589770 -4740
rect -6806 -5144 590730 -5112
rect -6806 -5380 -6774 -5144
rect -6538 -5380 -6454 -5144
rect -6218 -5380 7226 -5144
rect 7462 -5380 7546 -5144
rect 7782 -5380 43226 -5144
rect 43462 -5380 43546 -5144
rect 43782 -5380 79226 -5144
rect 79462 -5380 79546 -5144
rect 79782 -5380 115226 -5144
rect 115462 -5380 115546 -5144
rect 115782 -5380 151226 -5144
rect 151462 -5380 151546 -5144
rect 151782 -5380 187226 -5144
rect 187462 -5380 187546 -5144
rect 187782 -5380 223226 -5144
rect 223462 -5380 223546 -5144
rect 223782 -5380 259226 -5144
rect 259462 -5380 259546 -5144
rect 259782 -5380 295226 -5144
rect 295462 -5380 295546 -5144
rect 295782 -5380 331226 -5144
rect 331462 -5380 331546 -5144
rect 331782 -5380 367226 -5144
rect 367462 -5380 367546 -5144
rect 367782 -5380 403226 -5144
rect 403462 -5380 403546 -5144
rect 403782 -5380 439226 -5144
rect 439462 -5380 439546 -5144
rect 439782 -5380 475226 -5144
rect 475462 -5380 475546 -5144
rect 475782 -5380 511226 -5144
rect 511462 -5380 511546 -5144
rect 511782 -5380 547226 -5144
rect 547462 -5380 547546 -5144
rect 547782 -5380 590142 -5144
rect 590378 -5380 590462 -5144
rect 590698 -5380 590730 -5144
rect -6806 -5464 590730 -5380
rect -6806 -5700 -6774 -5464
rect -6538 -5700 -6454 -5464
rect -6218 -5700 7226 -5464
rect 7462 -5700 7546 -5464
rect 7782 -5700 43226 -5464
rect 43462 -5700 43546 -5464
rect 43782 -5700 79226 -5464
rect 79462 -5700 79546 -5464
rect 79782 -5700 115226 -5464
rect 115462 -5700 115546 -5464
rect 115782 -5700 151226 -5464
rect 151462 -5700 151546 -5464
rect 151782 -5700 187226 -5464
rect 187462 -5700 187546 -5464
rect 187782 -5700 223226 -5464
rect 223462 -5700 223546 -5464
rect 223782 -5700 259226 -5464
rect 259462 -5700 259546 -5464
rect 259782 -5700 295226 -5464
rect 295462 -5700 295546 -5464
rect 295782 -5700 331226 -5464
rect 331462 -5700 331546 -5464
rect 331782 -5700 367226 -5464
rect 367462 -5700 367546 -5464
rect 367782 -5700 403226 -5464
rect 403462 -5700 403546 -5464
rect 403782 -5700 439226 -5464
rect 439462 -5700 439546 -5464
rect 439782 -5700 475226 -5464
rect 475462 -5700 475546 -5464
rect 475782 -5700 511226 -5464
rect 511462 -5700 511546 -5464
rect 511782 -5700 547226 -5464
rect 547462 -5700 547546 -5464
rect 547782 -5700 590142 -5464
rect 590378 -5700 590462 -5464
rect 590698 -5700 590730 -5464
rect -6806 -5732 590730 -5700
rect -7766 -6104 591690 -6072
rect -7766 -6340 -7734 -6104
rect -7498 -6340 -7414 -6104
rect -7178 -6340 8466 -6104
rect 8702 -6340 8786 -6104
rect 9022 -6340 44466 -6104
rect 44702 -6340 44786 -6104
rect 45022 -6340 80466 -6104
rect 80702 -6340 80786 -6104
rect 81022 -6340 116466 -6104
rect 116702 -6340 116786 -6104
rect 117022 -6340 152466 -6104
rect 152702 -6340 152786 -6104
rect 153022 -6340 188466 -6104
rect 188702 -6340 188786 -6104
rect 189022 -6340 224466 -6104
rect 224702 -6340 224786 -6104
rect 225022 -6340 260466 -6104
rect 260702 -6340 260786 -6104
rect 261022 -6340 296466 -6104
rect 296702 -6340 296786 -6104
rect 297022 -6340 332466 -6104
rect 332702 -6340 332786 -6104
rect 333022 -6340 368466 -6104
rect 368702 -6340 368786 -6104
rect 369022 -6340 404466 -6104
rect 404702 -6340 404786 -6104
rect 405022 -6340 440466 -6104
rect 440702 -6340 440786 -6104
rect 441022 -6340 476466 -6104
rect 476702 -6340 476786 -6104
rect 477022 -6340 512466 -6104
rect 512702 -6340 512786 -6104
rect 513022 -6340 548466 -6104
rect 548702 -6340 548786 -6104
rect 549022 -6340 591102 -6104
rect 591338 -6340 591422 -6104
rect 591658 -6340 591690 -6104
rect -7766 -6424 591690 -6340
rect -7766 -6660 -7734 -6424
rect -7498 -6660 -7414 -6424
rect -7178 -6660 8466 -6424
rect 8702 -6660 8786 -6424
rect 9022 -6660 44466 -6424
rect 44702 -6660 44786 -6424
rect 45022 -6660 80466 -6424
rect 80702 -6660 80786 -6424
rect 81022 -6660 116466 -6424
rect 116702 -6660 116786 -6424
rect 117022 -6660 152466 -6424
rect 152702 -6660 152786 -6424
rect 153022 -6660 188466 -6424
rect 188702 -6660 188786 -6424
rect 189022 -6660 224466 -6424
rect 224702 -6660 224786 -6424
rect 225022 -6660 260466 -6424
rect 260702 -6660 260786 -6424
rect 261022 -6660 296466 -6424
rect 296702 -6660 296786 -6424
rect 297022 -6660 332466 -6424
rect 332702 -6660 332786 -6424
rect 333022 -6660 368466 -6424
rect 368702 -6660 368786 -6424
rect 369022 -6660 404466 -6424
rect 404702 -6660 404786 -6424
rect 405022 -6660 440466 -6424
rect 440702 -6660 440786 -6424
rect 441022 -6660 476466 -6424
rect 476702 -6660 476786 -6424
rect 477022 -6660 512466 -6424
rect 512702 -6660 512786 -6424
rect 513022 -6660 548466 -6424
rect 548702 -6660 548786 -6424
rect 549022 -6660 591102 -6424
rect 591338 -6660 591422 -6424
rect 591658 -6660 591690 -6424
rect -7766 -6692 591690 -6660
rect -8726 -7064 592650 -7032
rect -8726 -7300 -8694 -7064
rect -8458 -7300 -8374 -7064
rect -8138 -7300 9706 -7064
rect 9942 -7300 10026 -7064
rect 10262 -7300 45706 -7064
rect 45942 -7300 46026 -7064
rect 46262 -7300 81706 -7064
rect 81942 -7300 82026 -7064
rect 82262 -7300 117706 -7064
rect 117942 -7300 118026 -7064
rect 118262 -7300 153706 -7064
rect 153942 -7300 154026 -7064
rect 154262 -7300 189706 -7064
rect 189942 -7300 190026 -7064
rect 190262 -7300 225706 -7064
rect 225942 -7300 226026 -7064
rect 226262 -7300 261706 -7064
rect 261942 -7300 262026 -7064
rect 262262 -7300 297706 -7064
rect 297942 -7300 298026 -7064
rect 298262 -7300 333706 -7064
rect 333942 -7300 334026 -7064
rect 334262 -7300 369706 -7064
rect 369942 -7300 370026 -7064
rect 370262 -7300 405706 -7064
rect 405942 -7300 406026 -7064
rect 406262 -7300 441706 -7064
rect 441942 -7300 442026 -7064
rect 442262 -7300 477706 -7064
rect 477942 -7300 478026 -7064
rect 478262 -7300 513706 -7064
rect 513942 -7300 514026 -7064
rect 514262 -7300 549706 -7064
rect 549942 -7300 550026 -7064
rect 550262 -7300 592062 -7064
rect 592298 -7300 592382 -7064
rect 592618 -7300 592650 -7064
rect -8726 -7384 592650 -7300
rect -8726 -7620 -8694 -7384
rect -8458 -7620 -8374 -7384
rect -8138 -7620 9706 -7384
rect 9942 -7620 10026 -7384
rect 10262 -7620 45706 -7384
rect 45942 -7620 46026 -7384
rect 46262 -7620 81706 -7384
rect 81942 -7620 82026 -7384
rect 82262 -7620 117706 -7384
rect 117942 -7620 118026 -7384
rect 118262 -7620 153706 -7384
rect 153942 -7620 154026 -7384
rect 154262 -7620 189706 -7384
rect 189942 -7620 190026 -7384
rect 190262 -7620 225706 -7384
rect 225942 -7620 226026 -7384
rect 226262 -7620 261706 -7384
rect 261942 -7620 262026 -7384
rect 262262 -7620 297706 -7384
rect 297942 -7620 298026 -7384
rect 298262 -7620 333706 -7384
rect 333942 -7620 334026 -7384
rect 334262 -7620 369706 -7384
rect 369942 -7620 370026 -7384
rect 370262 -7620 405706 -7384
rect 405942 -7620 406026 -7384
rect 406262 -7620 441706 -7384
rect 441942 -7620 442026 -7384
rect 442262 -7620 477706 -7384
rect 477942 -7620 478026 -7384
rect 478262 -7620 513706 -7384
rect 513942 -7620 514026 -7384
rect 514262 -7620 549706 -7384
rect 549942 -7620 550026 -7384
rect 550262 -7620 592062 -7384
rect 592298 -7620 592382 -7384
rect 592618 -7620 592650 -7384
rect -8726 -7652 592650 -7620
use mux16x1_project  mprj1
timestamp 1714498238
transform 1 0 538000 0 1 423802
box 0 552 10000 22000
use mux16x1_project  mprj2
timestamp 1714498238
transform 1 0 538000 0 1 387802
box 0 552 10000 22000
use mux16x1_project  mprj3
timestamp 1714498238
transform 1 0 538000 0 1 351802
box 0 552 10000 22000
use mux16x1_project  mprj4
timestamp 1714498238
transform 1 0 538000 0 1 315802
box 0 552 10000 22000
use mux16x1_project  mprj5
timestamp 1714498238
transform 1 0 538000 0 1 279802
box 0 552 10000 22000
use sky130_osu_ring_oscillator_mpr2ca_8_b0r1  ro1
timestamp 1714079683
transform 1 0 468600 0 1 449002
box 0 0 20145 2491
use sky130_osu_ring_oscillator_mpr2ct_8_b0r1  ro2
timestamp 1714057498
transform 1 0 468600 0 1 430602
box 0 0 20785 2492
use sky130_osu_ring_oscillator_mpr2ea_8_b0r1  ro3
timestamp 1714062703
transform 1 0 468600 0 1 409602
box 0 0 19886 2492
use sky130_osu_ring_oscillator_mpr2et_8_b0r1  ro4
timestamp 1714057805
transform 1 0 468600 0 1 388602
box 0 0 22123 2493
use sky130_osu_ring_oscillator_mpr2xa_8_b0r1  ro5
timestamp 1714057206
transform 1 0 468600 0 1 356002
box 0 0 20809 2493
use sky130_osu_ring_oscillator_mpr2ca_8_b0r2  ro6
timestamp 1714079683
transform 1 0 468600 0 1 340002
box 0 0 20217 2494
use sky130_osu_ring_oscillator_mpr2ct_8_b0r2  ro7
timestamp 1714057574
transform 1 0 468600 0 1 320002
box 0 0 20783 2493
use sky130_osu_ring_oscillator_mpr2ea_8_b0r2  ro8
timestamp 1714057774
transform 1 0 468600 0 1 304602
box 0 0 19885 2492
use sky130_osu_ring_oscillator_mpr2et_8_b0r2  ro9
timestamp 1714057841
transform 1 0 468600 0 1 285002
box 0 0 22120 2493
use sky130_osu_ring_oscillator_mpr2xa_8_b0r2  ro10
timestamp 1714057206
transform 1 0 468600 0 1 265002
box 0 0 20819 2493
use sky130_fd_sc_hd__conb_1  sky130_fd_sc_hd__conb_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform -1 0 576676 0 1 697102
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  sky130_fd_sc_hd__conb_1_1
timestamp 1692646696
transform -1 0 576676 0 1 232255
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  sky130_fd_sc_hd__conb_1_2
timestamp 1692646696
transform -1 0 576676 0 1 272102
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  sky130_fd_sc_hd__conb_1_3
timestamp 1692646696
transform -1 0 576676 0 1 325142
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  sky130_fd_sc_hd__conb_1_4
timestamp 1692646696
transform -1 0 576676 0 1 378318
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  sky130_fd_sc_hd__conb_1_5
timestamp 1692646696
transform -1 0 576676 0 1 431494
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  sky130_fd_sc_hd__conb_1_6
timestamp 1692646696
transform -1 0 576676 0 1 484534
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  sky130_fd_sc_hd__conb_1_7
timestamp 1692646696
transform -1 0 576676 0 1 537710
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  sky130_fd_sc_hd__conb_1_8
timestamp 1692646696
transform -1 0 576676 0 1 590886
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  sky130_fd_sc_hd__conb_1_9
timestamp 1692646696
transform -1 0 576676 0 1 643926
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  sky130_fd_sc_hd__conb_1_10
timestamp 1692646696
transform 1 0 504548 0 -1 702267
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  sky130_fd_sc_hd__conb_1_11
timestamp 1692646696
transform 1 0 252559 0 -1 703079
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  sky130_fd_sc_hd__conb_1_12
timestamp 1692646696
transform 1 0 324561 0 -1 703119
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  sky130_fd_sc_hd__conb_1_13
timestamp 1692646696
transform 1 0 360593 0 -1 702650
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  sky130_fd_sc_hd__conb_1_14
timestamp 1692646696
transform 1 0 432553 0 -1 702513
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  TIE_ZERO_zero_
timestamp 1692646696
transform 1 0 504306 0 1 553794
box -38 -48 314 592
<< labels >>
flabel metal3 s 583520 285278 584960 285518 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703522 446210 704962 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703522 381258 704962 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703522 316398 704962 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703522 251538 704962 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703522 186586 704962 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703522 121726 704962 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703522 56866 704962 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697222 480 697462 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644998 480 645238 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592910 480 593150 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338454 584960 338694 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540686 480 540926 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488598 480 488838 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436510 480 436750 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384286 480 384526 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332198 480 332438 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279974 480 280214 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227886 480 228126 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175798 480 176038 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123574 480 123814 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391630 584960 391870 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444670 584960 444910 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497846 584960 498086 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551022 584960 551262 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604062 584960 604302 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657238 584960 657478 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703522 575930 704962 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703522 511070 704962 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6478 584960 6718 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457998 584960 458238 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511174 584960 511414 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564214 584960 564454 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617390 584960 617630 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670566 584960 670806 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703522 559738 704962 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703522 494878 704962 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703522 429926 704962 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703522 365066 704962 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703522 300206 704962 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46190 584960 46430 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703522 235254 704962 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703522 170394 704962 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703522 105534 704962 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703522 40582 704962 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684166 480 684406 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631942 480 632182 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579854 480 580094 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527766 480 528006 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475542 480 475782 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423454 480 423694 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86038 584960 86278 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371230 480 371470 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319142 480 319382 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267054 480 267294 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214830 480 215070 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162742 480 162982 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110518 480 110758 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71486 480 71726 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32318 480 32558 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125886 584960 126126 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165734 584960 165974 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205582 584960 205822 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245430 584960 245670 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298606 584960 298846 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351782 584960 352022 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404822 584960 405062 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32998 584960 33238 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484518 584960 484758 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537694 584960 537934 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590870 584960 591110 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643910 584960 644150 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697086 584960 697326 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703522 527262 704962 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703522 462402 704962 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703522 397542 704962 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703522 332590 704962 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703522 267730 704962 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72846 584960 73086 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703522 202870 704962 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703522 137918 704962 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703522 73058 704962 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703522 8198 704962 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658054 480 658294 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605966 480 606206 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553742 480 553982 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501654 480 501894 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449430 480 449670 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397342 480 397582 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112694 584960 112934 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345254 480 345494 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293030 480 293270 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240942 480 241182 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188718 480 188958 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136630 480 136870 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84542 480 84782 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45374 480 45614 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6342 480 6582 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152542 584960 152782 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192390 584960 192630 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232238 584960 232478 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272086 584960 272326 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325126 584960 325366 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378302 584960 378542 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431478 584960 431718 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19670 584960 19910 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471326 584960 471566 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524366 584960 524606 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577542 584960 577782 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630718 584960 630958 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683758 584960 683998 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703522 543546 704962 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703522 478594 704962 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703522 413734 704962 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703522 348874 704962 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703522 283922 704962 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59518 584960 59758 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703522 219062 704962 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703522 154202 704962 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703522 89250 704962 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703522 24390 704962 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671110 480 671350 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619022 480 619262 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566798 480 567038 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514710 480 514950 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462486 480 462726 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410398 480 410638 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99366 584960 99606 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358310 480 358550 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306086 480 306326 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253998 480 254238 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201774 480 202014 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149686 480 149926 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97462 480 97702 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58430 480 58670 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19262 480 19502 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139214 584960 139454 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179062 584960 179302 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218910 584960 219150 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258758 584960 258998 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311934 584960 312174 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364974 584960 365214 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418150 584960 418390 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -958 125958 482 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -958 480618 482 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -958 484114 482 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -958 487702 482 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -958 491198 482 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -958 494786 482 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -958 498282 482 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -958 501870 482 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -958 505458 482 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -958 508954 482 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -958 512542 482 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -958 161378 482 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -958 516038 482 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -958 519626 482 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -958 523122 482 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -958 526710 482 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -958 530206 482 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -958 533794 482 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -958 537290 482 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -958 540878 482 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -958 544466 482 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -958 547962 482 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -958 164966 482 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -958 551550 482 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -958 555046 482 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -958 558634 482 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -958 562130 482 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -958 565718 482 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -958 569214 482 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -958 572802 482 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -958 576390 482 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -958 168462 482 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -958 172050 482 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -958 175546 482 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -958 179134 482 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -958 182630 482 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -958 186218 482 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -958 189806 482 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -958 193302 482 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -958 129454 482 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -958 196890 482 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -958 200386 482 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -958 203974 482 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -958 207470 482 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -958 211058 482 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -958 214554 482 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -958 218142 482 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -958 221638 482 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -958 225226 482 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -958 228814 482 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -958 133042 482 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -958 232310 482 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -958 235898 482 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -958 239394 482 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -958 242982 482 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -958 246478 482 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -958 250066 482 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -958 253562 482 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -958 257150 482 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -958 260738 482 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -958 264234 482 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -958 136538 482 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -958 267822 482 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -958 271318 482 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -958 274906 482 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -958 278402 482 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -958 281990 482 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -958 285486 482 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -958 289074 482 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -958 292662 482 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -958 296158 482 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -958 299746 482 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -958 140126 482 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -958 303242 482 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -958 306830 482 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -958 310326 482 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -958 313914 482 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -958 317410 482 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -958 320998 482 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -958 324494 482 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -958 328082 482 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -958 331670 482 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -958 335166 482 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -958 143622 482 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -958 338754 482 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -958 342250 482 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -958 345838 482 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -958 349334 482 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -958 352922 482 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -958 356418 482 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -958 360006 482 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -958 363594 482 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -958 367090 482 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -958 370678 482 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -958 147210 482 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -958 374174 482 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -958 377762 482 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -958 381258 482 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -958 384846 482 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -958 388342 482 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -958 391930 482 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -958 395426 482 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -958 399014 482 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -958 402602 482 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -958 406098 482 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -958 150706 482 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -958 409686 482 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -958 413182 482 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -958 416770 482 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -958 420266 482 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -958 423854 482 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -958 427350 482 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -958 430938 482 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -958 434526 482 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -958 438022 482 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -958 441610 482 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -958 154294 482 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -958 445106 482 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -958 448694 482 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -958 452190 482 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -958 455778 482 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -958 459274 482 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -958 462862 482 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -958 466358 482 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -958 469946 482 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -958 473534 482 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -958 477030 482 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -958 157882 482 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -958 127062 482 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -958 481814 482 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -958 485310 482 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -958 488898 482 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -958 492394 482 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -958 495982 482 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -958 499478 482 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -958 503066 482 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -958 506562 482 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -958 510150 482 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -958 513646 482 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -958 162574 482 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -958 517234 482 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -958 520822 482 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -958 524318 482 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -958 527906 482 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -958 531402 482 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -958 534990 482 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -958 538486 482 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -958 542074 482 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -958 545570 482 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -958 549158 482 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -958 166162 482 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -958 552746 482 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -958 556242 482 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -958 559830 482 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -958 563326 482 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -958 566914 482 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -958 570410 482 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -958 573998 482 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -958 577494 482 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -958 169658 482 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -958 173246 482 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -958 176742 482 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -958 180330 482 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -958 183826 482 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -958 187414 482 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -958 190910 482 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -958 194498 482 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -958 130650 482 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -958 197994 482 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -958 201582 482 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -958 205170 482 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -958 208666 482 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -958 212254 482 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -958 215750 482 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -958 219338 482 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -958 222834 482 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -958 226422 482 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -958 229918 482 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -958 134238 482 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -958 233506 482 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -958 237094 482 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -958 240590 482 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -958 244178 482 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -958 247674 482 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -958 251262 482 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -958 254758 482 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -958 258346 482 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -958 261842 482 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -958 265430 482 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -958 137734 482 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -958 268926 482 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -958 272514 482 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -958 276102 482 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -958 279598 482 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -958 283186 482 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -958 286682 482 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -958 290270 482 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -958 293766 482 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -958 297354 482 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -958 300850 482 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -958 141322 482 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -958 304438 482 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -958 308026 482 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -958 311522 482 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -958 315110 482 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -958 318606 482 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -958 322194 482 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -958 325690 482 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -958 329278 482 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -958 332774 482 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -958 336362 482 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -958 144818 482 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -958 339950 482 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -958 343446 482 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -958 347034 482 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -958 350530 482 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -958 354118 482 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -958 357614 482 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -958 361202 482 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -958 364698 482 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -958 368286 482 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -958 371782 482 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -958 148406 482 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -958 375370 482 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -958 378958 482 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -958 382454 482 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -958 386042 482 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -958 389538 482 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -958 393126 482 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -958 396622 482 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -958 400210 482 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -958 403706 482 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -958 407294 482 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -958 151902 482 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -958 410882 482 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -958 414378 482 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -958 417966 482 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -958 421462 482 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -958 425050 482 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -958 428546 482 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -958 432134 482 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -958 435630 482 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -958 439218 482 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -958 442714 482 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -958 155490 482 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -958 446302 482 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -958 449890 482 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -958 453386 482 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -958 456974 482 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -958 460470 482 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -958 464058 482 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -958 467554 482 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -958 471142 482 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -958 474638 482 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -958 478226 482 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -958 158986 482 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -958 128258 482 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -958 482918 482 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -958 486506 482 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -958 490002 482 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -958 493590 482 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -958 497178 482 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -958 500674 482 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -958 504262 482 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -958 507758 482 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -958 511346 482 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -958 514842 482 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -958 163770 482 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -958 518430 482 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -958 521926 482 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -958 525514 482 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -958 529102 482 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -958 532598 482 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -958 536186 482 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -958 539682 482 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -958 543270 482 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -958 546766 482 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -958 550354 482 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -958 167266 482 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -958 553850 482 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -958 557438 482 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -958 560934 482 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -958 564522 482 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -958 568110 482 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -958 571606 482 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -958 575194 482 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -958 578690 482 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -958 170854 482 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -958 174350 482 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -958 177938 482 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -958 181526 482 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -958 185022 482 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -958 188610 482 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -958 192106 482 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -958 195694 482 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -958 131846 482 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -958 199190 482 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -958 202778 482 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -958 206274 482 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -958 209862 482 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -958 213450 482 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -958 216946 482 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -958 220534 482 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -958 224030 482 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -958 227618 482 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -958 231114 482 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -958 135342 482 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -958 234702 482 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -958 238198 482 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -958 241786 482 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -958 245282 482 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -958 248870 482 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -958 252458 482 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -958 255954 482 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -958 259542 482 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -958 263038 482 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -958 266626 482 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -958 138930 482 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -958 270122 482 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -958 273710 482 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -958 277206 482 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -958 280794 482 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -958 284382 482 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -958 287878 482 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -958 291466 482 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -958 294962 482 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -958 298550 482 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -958 302046 482 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -958 142518 482 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -958 305634 482 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -958 309130 482 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -958 312718 482 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -958 316306 482 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -958 319802 482 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -958 323390 482 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -958 326886 482 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -958 330474 482 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -958 333970 482 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -958 337558 482 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -958 146014 482 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -958 341054 482 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -958 344642 482 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -958 348138 482 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -958 351726 482 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -958 355314 482 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -958 358810 482 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -958 362398 482 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -958 365894 482 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -958 369482 482 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -958 372978 482 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -958 149602 482 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -958 376566 482 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -958 380062 482 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -958 383650 482 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -958 387238 482 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -958 390734 482 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -958 394322 482 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -958 397818 482 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -958 401406 482 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -958 404902 482 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -958 408490 482 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -958 153098 482 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -958 411986 482 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -958 415574 482 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -958 419070 482 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -958 422658 482 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -958 426246 482 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -958 429742 482 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -958 433330 482 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -958 436826 482 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -958 440414 482 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -958 443910 482 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -958 156686 482 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -958 447498 482 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -958 450994 482 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -958 454582 482 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -958 458170 482 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -958 461666 482 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -958 465254 482 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -958 468750 482 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -958 472338 482 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -958 475834 482 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -958 479422 482 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -958 160182 482 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -958 579886 482 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -958 581082 482 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -958 582278 482 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -958 583474 482 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -932 -1386 704872 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -932 585930 -312 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704252 585930 704872 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -932 585930 704872 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 994 -7652 1614 711592 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 36994 -7652 37614 711592 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 72994 -7652 73614 711592 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 108994 -7652 109614 711592 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 144994 -7652 145614 711592 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 180994 -7652 181614 711592 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 216994 -7652 217614 711592 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 252994 -7652 253614 711592 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 288994 -7652 289614 711592 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 324994 -7652 325614 711592 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 360994 -7652 361614 711592 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 396994 -7652 397614 711592 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 432994 -7652 433614 711592 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 468994 -7652 469614 711592 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 504994 -7652 505614 711592 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 540994 -7652 541614 279790 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 540994 445574 541614 711592 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 576994 -7652 577614 711592 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 2068 592650 2688 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 38068 592650 38688 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 74068 592650 74688 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 110068 592650 110688 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 146068 592650 146688 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 182068 592650 182688 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 218068 592650 218688 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 254068 592650 254688 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 290068 592650 290688 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 326068 592650 326688 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 362068 592650 362688 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 398068 592650 398688 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 434068 592650 434688 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 470068 592650 470688 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 506068 592650 506688 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 542068 592650 542688 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 578068 592650 578688 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 614068 592650 614688 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 650068 592650 650688 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 686068 592650 686688 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -3926 -2852 -3306 706792 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 -2852 587850 -2232 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 706172 587850 706792 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 587230 -2852 587850 706792 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 3474 -7652 4094 711592 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 39474 -7652 40094 711592 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 75474 -7652 76094 711592 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 111474 -7652 112094 711592 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 147474 -7652 148094 711592 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 183474 -7652 184094 711592 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 219474 -7652 220094 711592 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 255474 -7652 256094 711592 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 291474 -7652 292094 711592 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 327474 -7652 328094 711592 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 363474 -7652 364094 711592 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 399474 -7652 400094 711592 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 435474 -7652 436094 711592 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 471474 -7652 472094 711592 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 507474 -7652 508094 711592 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 543474 -7652 544094 279790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 543474 445574 544094 711592 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 579474 -7652 580094 711592 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 4548 592650 5168 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 40548 592650 41168 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 76548 592650 77168 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 112548 592650 113168 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 148548 592650 149168 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 184548 592650 185168 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 220548 592650 221168 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 256548 592650 257168 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 292548 592650 293168 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 328548 592650 329168 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 364548 592650 365168 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 400548 592650 401168 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 436548 592650 437168 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 472548 592650 473168 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 508548 592650 509168 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 544548 592650 545168 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 580548 592650 581168 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 616548 592650 617168 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 652548 592650 653168 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 688548 592650 689168 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -5846 -4772 -5226 708712 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 -4772 589770 -4152 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 708092 589770 708712 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 589150 -4772 589770 708712 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 5954 -7652 6574 711592 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 41954 -7652 42574 711592 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 77954 -7652 78574 711592 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 113954 -7652 114574 711592 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 149954 -7652 150574 711592 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 185954 -7652 186574 711592 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 221954 -7652 222574 711592 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 257954 -7652 258574 711592 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 293954 -7652 294574 711592 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 329954 -7652 330574 711592 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 365954 -7652 366574 711592 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 401954 -7652 402574 711592 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 437954 -7652 438574 711592 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 473954 -7652 474574 263617 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 473954 268062 474574 354617 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 473954 359062 474574 711592 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 509954 -7652 510574 711592 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 545954 -7652 546574 279790 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 545954 445574 546574 711592 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 581954 -7652 582574 711592 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 7028 592650 7648 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 43028 592650 43648 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 79028 592650 79648 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 115028 592650 115648 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 151028 592650 151648 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 187028 592650 187648 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 223028 592650 223648 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 259028 592650 259648 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 295028 592650 295648 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 331028 592650 331648 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 367028 592650 367648 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 403028 592650 403648 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 439028 592650 439648 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 475028 592650 475648 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 511028 592650 511648 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 547028 592650 547648 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 583028 592650 583648 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 619028 592650 619648 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 655028 592650 655648 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 691028 592650 691648 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -7766 -6692 -7146 710632 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 -6692 591690 -6072 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 710012 591690 710632 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 591070 -6692 591690 710632 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 8434 -7652 9054 711592 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 44434 -7652 45054 711592 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 80434 -7652 81054 711592 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 116434 -7652 117054 711592 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 152434 -7652 153054 711592 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 188434 -7652 189054 711592 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 224434 -7652 225054 711592 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 260434 -7652 261054 711592 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 296434 -7652 297054 711592 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 332434 -7652 333054 711592 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 368434 -7652 369054 711592 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 404434 -7652 405054 711592 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 440434 -7652 441054 711592 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 476434 -7652 477054 263617 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 476434 268062 477054 354617 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 476434 359062 477054 711592 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 512434 -7652 513054 711592 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 548434 -7652 549054 711592 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 9508 592650 10128 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 45508 592650 46128 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 81508 592650 82128 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 117508 592650 118128 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 153508 592650 154128 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 189508 592650 190128 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 225508 592650 226128 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 261508 592650 262128 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 297508 592650 298128 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 333508 592650 334128 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 369508 592650 370128 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 405508 592650 406128 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 441508 592650 442128 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 477508 592650 478128 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 513508 592650 514128 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 549508 592650 550128 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 585508 592650 586128 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 621508 592650 622128 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 657508 592650 658128 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 693508 592650 694128 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s -6806 -5732 -6186 709672 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 -5732 590730 -5112 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 709052 590730 709672 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 590110 -5732 590730 709672 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 7194 -7652 7814 711592 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 43194 -7652 43814 711592 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 79194 -7652 79814 711592 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 115194 -7652 115814 711592 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 151194 -7652 151814 711592 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 187194 -7652 187814 711592 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 223194 -7652 223814 711592 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 259194 -7652 259814 711592 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 295194 -7652 295814 711592 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 331194 -7652 331814 711592 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 367194 -7652 367814 711592 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 403194 -7652 403814 711592 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 439194 -7652 439814 711592 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 475194 -7652 475814 263617 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 475194 268062 475814 354617 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 475194 359062 475814 711592 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 511194 -7652 511814 711592 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 547194 -7652 547814 711592 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 8268 592650 8888 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 44268 592650 44888 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 80268 592650 80888 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 116268 592650 116888 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 152268 592650 152888 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 188268 592650 188888 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 224268 592650 224888 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 260268 592650 260888 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 296268 592650 296888 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 332268 592650 332888 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 368268 592650 368888 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 404268 592650 404888 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 440268 592650 440888 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 476268 592650 476888 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 512268 592650 512888 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 548268 592650 548888 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 584268 592650 584888 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 620268 592650 620888 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 656268 592650 656888 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 692268 592650 692888 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -8726 -7652 -8106 711592 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 -7652 592650 -7032 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 710972 592650 711592 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 592030 -7652 592650 711592 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 9674 -7652 10294 711592 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 45674 -7652 46294 711592 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 81674 -7652 82294 711592 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 117674 -7652 118294 711592 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 153674 -7652 154294 711592 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 189674 -7652 190294 711592 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 225674 -7652 226294 711592 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 261674 -7652 262294 711592 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 297674 -7652 298294 711592 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 333674 -7652 334294 711592 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 369674 -7652 370294 711592 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 405674 -7652 406294 711592 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 441674 -7652 442294 711592 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 477674 -7652 478294 263617 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 477674 268062 478294 354617 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 477674 359062 478294 711592 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 513674 -7652 514294 711592 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 549674 -7652 550294 711592 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 10748 592650 11368 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 46748 592650 47368 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 82748 592650 83368 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 118748 592650 119368 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 154748 592650 155368 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 190748 592650 191368 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 226748 592650 227368 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 262748 592650 263368 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 298748 592650 299368 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 334748 592650 335368 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 370748 592650 371368 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 406748 592650 407368 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 442748 592650 443368 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 478748 592650 479368 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 514748 592650 515368 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 550748 592650 551368 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 586748 592650 587368 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 622748 592650 623368 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 658748 592650 659368 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 694748 592650 695368 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -2966 -1892 -2346 705832 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 -1892 586890 -1272 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 705212 586890 705832 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 586270 -1892 586890 705832 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 2234 -7652 2854 711592 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 38234 -7652 38854 711592 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 74234 -7652 74854 711592 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 110234 -7652 110854 711592 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 146234 -7652 146854 711592 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 182234 -7652 182854 711592 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 218234 -7652 218854 711592 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 254234 -7652 254854 711592 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 290234 -7652 290854 711592 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 326234 -7652 326854 711592 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 362234 -7652 362854 711592 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 398234 -7652 398854 711592 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 434234 -7652 434854 711592 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 470234 -7652 470854 711592 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 506234 -7652 506854 711592 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 542234 -7652 542854 279790 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 542234 445574 542854 711592 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 578234 -7652 578854 711592 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 3308 592650 3928 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 39308 592650 39928 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 75308 592650 75928 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 111308 592650 111928 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 147308 592650 147928 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 183308 592650 183928 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 219308 592650 219928 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 255308 592650 255928 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 291308 592650 291928 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 327308 592650 327928 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 363308 592650 363928 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 399308 592650 399928 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 435308 592650 435928 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 471308 592650 471928 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 507308 592650 507928 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 543308 592650 543928 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 579308 592650 579928 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 615308 592650 615928 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 651308 592650 651928 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 687308 592650 687928 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -4886 -3812 -4266 707752 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 -3812 588810 -3192 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 707132 588810 707752 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 588190 -3812 588810 707752 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 4714 -7652 5334 711592 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 40714 -7652 41334 711592 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 76714 -7652 77334 711592 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 112714 -7652 113334 711592 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 148714 -7652 149334 711592 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 184714 -7652 185334 711592 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 220714 -7652 221334 711592 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 256714 -7652 257334 711592 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 292714 -7652 293334 711592 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 328714 -7652 329334 711592 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 364714 -7652 365334 711592 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 400714 -7652 401334 711592 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 436714 -7652 437334 711592 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 472714 -7652 473334 263617 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 472714 268062 473334 354617 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 472714 359062 473334 711592 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 508714 -7652 509334 711592 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 544714 -7652 545334 279790 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 544714 445574 545334 711592 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 580714 -7652 581334 711592 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 5788 592650 6408 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 41788 592650 42408 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 77788 592650 78408 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 113788 592650 114408 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 149788 592650 150408 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 185788 592650 186408 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 221788 592650 222408 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 257788 592650 258408 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 293788 592650 294408 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 329788 592650 330408 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 365788 592650 366408 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 401788 592650 402408 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 437788 592650 438408 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 473788 592650 474408 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 509788 592650 510408 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 545788 592650 546408 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 581788 592650 582408 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 617788 592650 618408 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 653788 592650 654408 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 689788 592650 690408 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -958 654 482 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -958 1758 482 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -958 2954 482 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -958 7738 482 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -958 47942 482 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -958 51438 482 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -958 55026 482 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -958 58522 482 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -958 62110 482 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -958 65606 482 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -958 69194 482 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -958 72690 482 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -958 76278 482 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -958 79774 482 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -958 12430 482 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -958 83362 482 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -958 86950 482 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -958 90446 482 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -958 94034 482 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -958 97530 482 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -958 101118 482 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -958 104614 482 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -958 108202 482 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -958 111698 482 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -958 115286 482 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -958 17122 482 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -958 118874 482 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -958 122370 482 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -958 21906 482 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -958 26598 482 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -958 30186 482 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -958 33682 482 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -958 37270 482 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -958 40766 482 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -958 44354 482 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -958 4150 482 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -958 8842 482 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -958 49046 482 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -958 52634 482 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -958 56130 482 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -958 59718 482 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -958 63306 482 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -958 66802 482 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -958 70390 482 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -958 73886 482 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -958 77474 482 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -958 80970 482 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -958 13626 482 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -958 84558 482 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -958 88054 482 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -958 91642 482 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -958 95230 482 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -958 98726 482 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -958 102314 482 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -958 105810 482 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -958 109398 482 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -958 112894 482 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -958 116482 482 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -958 18318 482 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -958 119978 482 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -958 123566 482 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -958 23102 482 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -958 27794 482 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -958 31382 482 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -958 34878 482 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -958 38466 482 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -958 41962 482 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -958 45550 482 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -958 10038 482 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -958 50242 482 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -958 53830 482 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -958 57326 482 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -958 60914 482 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -958 64410 482 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -958 67998 482 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -958 71586 482 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -958 75082 482 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -958 78670 482 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -958 82166 482 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -958 14822 482 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -958 85754 482 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -958 89250 482 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -958 92838 482 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -958 96334 482 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -958 99922 482 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -958 103418 482 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -958 107006 482 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -958 110594 482 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -958 114090 482 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -958 117678 482 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -958 19514 482 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -958 121174 482 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -958 124762 482 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -958 24298 482 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -958 28990 482 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -958 32486 482 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -958 36074 482 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -958 39662 482 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -958 43158 482 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -958 46746 482 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -958 11234 482 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -958 16018 482 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -958 20710 482 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -958 25402 482 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -958 5346 482 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -958 6542 482 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
