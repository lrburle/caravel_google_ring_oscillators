magic
tech sky130A
magscale 1 2
timestamp 1708620019
<< error_s >>
rect 3122 2133 3123 2144
rect 3312 2133 3313 2144
rect 3398 2133 3399 2144
rect 5328 2133 5329 2144
rect 5518 2133 5519 2144
rect 5604 2133 5605 2144
rect 6280 2133 6281 2144
rect 6470 2133 6471 2144
rect 6556 2133 6557 2144
rect 6829 2133 6830 2144
rect 7027 2133 7028 2144
rect 8913 2133 8914 2144
rect 9103 2133 9104 2144
rect 9189 2133 9190 2144
rect 9865 2133 9866 2144
rect 10055 2133 10056 2144
rect 10141 2133 10142 2144
rect 10414 2133 10415 2144
rect 10612 2133 10613 2144
rect 12498 2133 12499 2144
rect 12688 2133 12689 2144
rect 12774 2133 12775 2144
rect 13450 2133 13451 2144
rect 13640 2133 13641 2144
rect 13726 2133 13727 2144
rect 13999 2133 14000 2144
rect 14197 2133 14198 2144
rect 16083 2133 16084 2144
rect 16273 2133 16274 2144
rect 16359 2133 16360 2144
rect 17035 2133 17036 2144
rect 17225 2133 17226 2144
rect 17311 2133 17312 2144
rect 17584 2133 17585 2144
rect 17782 2133 17783 2144
rect 19668 2133 19669 2144
rect 19858 2133 19859 2144
rect 19944 2133 19945 2144
rect 20620 2133 20621 2144
rect 20810 2133 20811 2144
rect 20896 2133 20897 2144
rect 21169 2133 21170 2144
rect 21367 2133 21368 2144
rect 3133 2093 3134 2133
rect 3323 2093 3324 2133
rect 3409 2093 3410 2133
rect 5339 2093 5340 2133
rect 5529 2093 5530 2133
rect 5615 2093 5616 2133
rect 6291 2093 6292 2133
rect 6481 2093 6482 2133
rect 6567 2093 6568 2133
rect 6840 2093 6841 2133
rect 7038 2093 7039 2133
rect 8924 2093 8925 2133
rect 9114 2093 9115 2133
rect 9200 2093 9201 2133
rect 9876 2093 9877 2133
rect 10066 2093 10067 2133
rect 10152 2093 10153 2133
rect 10425 2093 10426 2133
rect 10623 2093 10624 2133
rect 12509 2093 12510 2133
rect 12699 2093 12700 2133
rect 12785 2093 12786 2133
rect 13461 2093 13462 2133
rect 13651 2093 13652 2133
rect 13737 2093 13738 2133
rect 14010 2093 14011 2133
rect 14208 2093 14209 2133
rect 16094 2093 16095 2133
rect 16284 2093 16285 2133
rect 16370 2093 16371 2133
rect 17046 2093 17047 2133
rect 17236 2093 17237 2133
rect 17322 2093 17323 2133
rect 17595 2093 17596 2133
rect 17793 2093 17794 2133
rect 19679 2093 19680 2133
rect 19869 2093 19870 2133
rect 19955 2093 19956 2133
rect 20631 2093 20632 2133
rect 20821 2093 20822 2133
rect 20907 2093 20908 2133
rect 21180 2093 21181 2133
rect 21378 2093 21379 2133
rect 6488 1966 6515 1973
rect 10073 1966 10100 1973
rect 13658 1966 13685 1973
rect 17243 1966 17270 1973
rect 20828 1966 20855 1973
rect 6488 1945 6556 1966
rect 10073 1945 10141 1966
rect 13658 1945 13726 1966
rect 17243 1945 17311 1966
rect 20828 1945 20896 1966
rect 6488 1939 6543 1945
rect 10073 1939 10128 1945
rect 13658 1939 13713 1945
rect 17243 1939 17298 1945
rect 20828 1939 20883 1945
rect 6527 1938 6528 1939
rect 10112 1938 10113 1939
rect 13697 1938 13698 1939
rect 17282 1938 17283 1939
rect 20867 1938 20868 1939
rect 6500 1932 6555 1938
rect 10085 1932 10140 1938
rect 13670 1932 13725 1938
rect 17255 1932 17310 1938
rect 20840 1932 20895 1938
rect 6527 1910 6528 1932
rect 10112 1910 10113 1932
rect 13697 1910 13698 1932
rect 17282 1910 17283 1932
rect 20867 1910 20868 1932
rect 3122 1703 3123 1714
rect 3312 1703 3313 1714
rect 3398 1703 3399 1714
rect 5328 1703 5329 1714
rect 5518 1703 5519 1714
rect 5604 1703 5605 1714
rect 6280 1703 6281 1714
rect 6470 1703 6471 1714
rect 6556 1703 6557 1714
rect 6829 1703 6830 1714
rect 7027 1703 7028 1714
rect 8913 1703 8914 1714
rect 9103 1703 9104 1714
rect 9189 1703 9190 1714
rect 9865 1703 9866 1714
rect 10055 1703 10056 1714
rect 10141 1703 10142 1714
rect 10414 1703 10415 1714
rect 10612 1703 10613 1714
rect 12498 1703 12499 1714
rect 12688 1703 12689 1714
rect 12774 1703 12775 1714
rect 13450 1703 13451 1714
rect 13640 1703 13641 1714
rect 13726 1703 13727 1714
rect 13999 1703 14000 1714
rect 14197 1703 14198 1714
rect 16083 1703 16084 1714
rect 16273 1703 16274 1714
rect 16359 1703 16360 1714
rect 17035 1703 17036 1714
rect 17225 1703 17226 1714
rect 17311 1703 17312 1714
rect 17584 1703 17585 1714
rect 17782 1703 17783 1714
rect 19668 1703 19669 1714
rect 19858 1703 19859 1714
rect 19944 1703 19945 1714
rect 20620 1703 20621 1714
rect 20810 1703 20811 1714
rect 20896 1703 20897 1714
rect 21169 1703 21170 1714
rect 21367 1703 21368 1714
rect 3133 1507 3134 1703
rect 3323 1507 3324 1703
rect 3409 1507 3410 1703
rect 5277 1671 5301 1677
rect 5305 1676 5329 1677
rect 5339 1507 5340 1703
rect 5529 1507 5530 1703
rect 5615 1507 5616 1703
rect 6291 1507 6292 1703
rect 6481 1507 6482 1703
rect 6567 1507 6568 1703
rect 6840 1507 6841 1703
rect 7038 1507 7039 1703
rect 8862 1671 8886 1677
rect 8890 1676 8914 1677
rect 8924 1507 8925 1703
rect 9114 1507 9115 1703
rect 9200 1507 9201 1703
rect 9876 1507 9877 1703
rect 10066 1507 10067 1703
rect 10152 1507 10153 1703
rect 10425 1507 10426 1703
rect 10623 1507 10624 1703
rect 12447 1671 12471 1677
rect 12475 1676 12499 1677
rect 12509 1507 12510 1703
rect 12699 1507 12700 1703
rect 12785 1507 12786 1703
rect 13461 1507 13462 1703
rect 13651 1507 13652 1703
rect 13737 1507 13738 1703
rect 14010 1507 14011 1703
rect 14208 1507 14209 1703
rect 16032 1671 16056 1677
rect 16060 1676 16084 1677
rect 16094 1507 16095 1703
rect 16284 1507 16285 1703
rect 16370 1507 16371 1703
rect 17046 1507 17047 1703
rect 17236 1507 17237 1703
rect 17322 1507 17323 1703
rect 17595 1507 17596 1703
rect 17793 1507 17794 1703
rect 19617 1671 19641 1677
rect 19645 1676 19669 1677
rect 19679 1507 19680 1703
rect 19869 1507 19870 1703
rect 19955 1507 19956 1703
rect 20631 1507 20632 1703
rect 20821 1507 20822 1703
rect 20907 1507 20908 1703
rect 21180 1507 21181 1703
rect 21378 1507 21379 1703
rect 3447 1403 3471 1437
rect 5653 1403 5677 1437
rect 6605 1403 6629 1437
rect 9238 1403 9262 1437
rect 10190 1403 10214 1437
rect 12823 1403 12847 1437
rect 13775 1403 13799 1437
rect 16408 1403 16432 1437
rect 17360 1403 17384 1437
rect 19993 1403 20017 1437
rect 20945 1403 20969 1437
rect 6605 1085 6629 1119
rect 10190 1085 10214 1119
rect 13775 1085 13799 1119
rect 17360 1085 17384 1119
rect 20945 1085 20969 1119
rect 3694 1057 3703 1066
rect 3741 1057 3750 1066
rect 4958 1057 4967 1066
rect 5005 1057 5014 1066
rect 5350 1057 5358 1066
rect 5397 1057 5406 1066
rect 5550 1057 5559 1066
rect 5597 1057 5606 1066
rect 7279 1057 7288 1066
rect 7326 1057 7335 1066
rect 8543 1057 8552 1066
rect 8590 1057 8599 1066
rect 8935 1057 8943 1066
rect 8982 1057 8991 1066
rect 9135 1057 9144 1066
rect 9182 1057 9191 1066
rect 10864 1057 10873 1066
rect 10911 1057 10920 1066
rect 12128 1057 12137 1066
rect 12175 1057 12184 1066
rect 12520 1057 12528 1066
rect 12567 1057 12576 1066
rect 12720 1057 12729 1066
rect 12767 1057 12776 1066
rect 14449 1057 14458 1066
rect 14496 1057 14505 1066
rect 15713 1057 15722 1066
rect 15760 1057 15769 1066
rect 16105 1057 16113 1066
rect 16152 1057 16161 1066
rect 16305 1057 16314 1066
rect 16352 1057 16361 1066
rect 18034 1057 18043 1066
rect 18081 1057 18090 1066
rect 19298 1057 19307 1066
rect 19345 1057 19354 1066
rect 19690 1057 19698 1066
rect 19737 1057 19746 1066
rect 19890 1057 19899 1066
rect 19937 1057 19946 1066
rect 3685 1048 3694 1057
rect 3750 1048 3759 1057
rect 4949 1048 4958 1057
rect 4664 1038 4670 1044
rect 4710 1038 4716 1044
rect 4972 1043 4984 1051
rect 4994 1043 5006 1051
rect 5014 1048 5023 1057
rect 5073 1051 5089 1052
rect 4968 1040 4970 1043
rect 5008 1040 5010 1043
rect 5067 1039 5078 1051
rect 5341 1048 5350 1057
rect 5406 1051 5415 1057
rect 5347 1045 5350 1047
rect 5354 1045 5360 1051
rect 5400 1048 5415 1051
rect 5541 1048 5550 1057
rect 5606 1050 5615 1057
rect 5400 1045 5406 1048
rect 4658 1032 4664 1038
rect 4716 1032 4722 1038
rect 4949 1031 4955 1037
rect 4960 1031 4968 1039
rect 4971 1037 5006 1039
rect 4971 1036 4972 1037
rect 4970 1031 4971 1035
rect 4972 1031 4973 1036
rect 5004 1031 5006 1037
rect 3692 1026 3694 1030
rect 3677 1023 3716 1026
rect 4718 1023 4757 1028
rect 4943 1025 4949 1031
rect 4969 1026 4970 1031
rect 4968 1024 4969 1026
rect 3674 1022 3677 1023
rect 3674 1015 3686 1022
rect 3690 1016 3692 1022
rect 3674 1013 3690 1015
rect 3696 1013 3708 1022
rect 3716 1020 3745 1023
rect 3745 1014 3749 1020
rect 4485 1018 4537 1020
rect 4757 1018 4771 1023
rect 4967 1020 4968 1023
rect 4457 1016 4537 1018
rect 4457 1015 4508 1016
rect 3749 1013 3750 1014
rect 4432 1013 4457 1015
rect 4479 1014 4485 1015
rect 4508 1014 4513 1015
rect 3670 1011 3674 1013
rect 3686 1010 3690 1013
rect 4398 1011 4428 1013
rect 4474 1012 4479 1014
rect 3662 998 3670 1010
rect 3669 988 3670 998
rect 3674 1007 3708 1010
rect 3674 1003 3676 1007
rect 3674 996 3675 1003
rect 3686 1001 3690 1007
rect 3705 1005 3708 1007
rect 3711 1004 3720 1010
rect 3673 994 3675 996
rect 3672 988 3678 994
rect 3683 988 3686 1001
rect 3666 982 3672 988
rect 3669 976 3670 982
rect 3673 962 3674 988
rect 3706 982 3708 1004
rect 3712 998 3720 1004
rect 3750 1001 3759 1010
rect 4281 1005 4295 1007
rect 4307 1005 4398 1011
rect 4470 1007 4474 1012
rect 4281 1004 4307 1005
rect 4281 1003 4295 1004
rect 4275 1002 4295 1003
rect 4316 1002 4321 1005
rect 4466 1002 4470 1007
rect 4513 1005 4530 1014
rect 4530 1004 4532 1005
rect 3718 988 3724 994
rect 3741 992 3750 1001
rect 4266 997 4290 1002
rect 4321 997 4327 1002
rect 4465 1001 4466 1002
rect 4537 1001 4554 1016
rect 4771 1015 4778 1018
rect 4966 1016 4967 1020
rect 4778 1014 4781 1015
rect 4781 1005 4803 1014
rect 4964 1012 4966 1016
rect 5004 1014 5008 1031
rect 5010 1027 5018 1039
rect 5276 1037 5288 1045
rect 5337 1041 5347 1045
rect 5348 1041 5354 1045
rect 5312 1037 5354 1041
rect 5406 1039 5412 1045
rect 5559 1044 5565 1050
rect 5605 1048 5615 1050
rect 7270 1048 7279 1057
rect 7335 1048 7344 1057
rect 8534 1048 8543 1057
rect 5568 1044 5580 1048
rect 5590 1044 5602 1048
rect 5605 1044 5611 1048
rect 5553 1038 5559 1044
rect 5611 1038 5617 1044
rect 8249 1038 8255 1044
rect 8295 1038 8301 1044
rect 8557 1043 8569 1051
rect 8579 1043 8591 1051
rect 8599 1048 8608 1057
rect 8658 1051 8674 1052
rect 8553 1040 8555 1043
rect 8593 1040 8595 1043
rect 8652 1039 8663 1051
rect 8926 1048 8935 1057
rect 8991 1051 9000 1057
rect 8932 1045 8935 1047
rect 8939 1045 8945 1051
rect 8985 1048 9000 1051
rect 9126 1048 9135 1057
rect 9191 1050 9200 1057
rect 8985 1045 8991 1048
rect 5057 1020 5067 1036
rect 5088 1034 5100 1037
rect 5282 1036 5288 1037
rect 5334 1036 5337 1037
rect 5082 1033 5102 1034
rect 5276 1033 5282 1036
rect 5318 1033 5348 1036
rect 5082 1031 5088 1033
rect 5102 1031 5132 1033
rect 5079 1025 5082 1031
rect 5076 1022 5082 1025
rect 5134 1024 5155 1031
rect 5182 1024 5188 1030
rect 4803 1004 4806 1005
rect 4663 1001 4664 1004
rect 4264 996 4266 997
rect 3724 982 3730 988
rect 3741 986 3745 992
rect 4253 989 4264 996
rect 4275 993 4290 997
rect 4327 996 4328 997
rect 3739 974 3740 979
rect 3897 976 3913 984
rect 4080 976 4096 989
rect 4163 979 4180 989
rect 4239 981 4253 989
rect 4233 979 4239 981
rect 4180 978 4233 979
rect 4264 977 4272 989
rect 4276 987 4281 989
rect 4328 987 4340 996
rect 3897 974 3954 976
rect 3735 957 3739 972
rect 3897 968 3942 974
rect 3954 968 3958 974
rect 3673 944 3680 957
rect 3734 953 3735 956
rect 3733 949 3734 952
rect 3736 944 3750 953
rect 3881 952 3897 968
rect 3958 961 3963 968
rect 3888 944 3897 952
rect 3666 936 3672 942
rect 3672 930 3678 936
rect 3680 934 3705 944
rect 3720 936 3736 944
rect 3718 934 3736 936
rect 3884 935 3888 944
rect 3891 940 3897 941
rect 3891 939 3933 940
rect 3937 939 3943 941
rect 3891 936 3902 939
rect 3891 935 3897 936
rect 3933 935 3943 939
rect 3884 934 3891 935
rect 3711 929 3714 934
rect 3718 930 3724 934
rect 3707 923 3710 928
rect 3881 925 3884 934
rect 3885 929 3891 934
rect 3943 929 3949 935
rect 3950 933 3962 941
rect 4023 934 4029 940
rect 4069 934 4075 940
rect 4080 934 4086 956
rect 4145 952 4151 958
rect 4191 952 4197 958
rect 4264 956 4272 967
rect 4276 958 4278 987
rect 4526 984 4528 1001
rect 4532 999 4554 1001
rect 4532 989 4540 999
rect 4658 992 4663 1001
rect 4806 996 4827 1004
rect 4961 1002 4964 1011
rect 5004 1007 5006 1014
rect 4995 1005 5006 1007
rect 5010 1010 5018 1017
rect 5010 1005 5023 1010
rect 5008 1004 5009 1005
rect 5014 1001 5023 1005
rect 5057 1002 5067 1018
rect 5076 1015 5079 1022
rect 5130 1018 5136 1024
rect 5188 1018 5194 1024
rect 5264 1021 5272 1033
rect 5276 1031 5310 1033
rect 5276 1030 5282 1031
rect 5276 1029 5279 1030
rect 5076 1014 5078 1015
rect 5076 1013 5080 1014
rect 5078 1001 5080 1013
rect 4960 996 4961 997
rect 4716 995 4749 996
rect 4827 995 4829 996
rect 4751 993 4757 995
rect 4658 986 4664 992
rect 4716 987 4722 992
rect 4757 991 4761 993
rect 4829 991 4839 995
rect 4959 991 4960 995
rect 5001 993 5014 1001
rect 5076 998 5080 1001
rect 5264 999 5272 1011
rect 5276 1002 5278 1029
rect 5556 1024 5559 1036
rect 5611 1032 5614 1036
rect 8243 1032 8249 1038
rect 8301 1032 8307 1038
rect 5564 1018 5568 1031
rect 5611 1021 5627 1032
rect 8534 1031 8540 1037
rect 8545 1031 8553 1039
rect 8556 1037 8591 1039
rect 8556 1036 8557 1037
rect 8555 1031 8556 1035
rect 8557 1031 8558 1036
rect 8589 1031 8591 1037
rect 7277 1026 7279 1030
rect 5627 1018 5643 1021
rect 5353 1007 5354 1008
rect 5354 1005 5355 1006
rect 5276 1001 5279 1002
rect 5322 1001 5350 1002
rect 5276 999 5288 1001
rect 5322 1000 5348 1001
rect 5006 992 5014 993
rect 5067 991 5071 996
rect 5076 991 5081 998
rect 5276 997 5277 999
rect 5322 998 5344 1000
rect 5350 999 5354 1001
rect 5277 996 5278 997
rect 5322 996 5337 998
rect 5278 995 5280 996
rect 5276 993 5282 995
rect 5322 994 5338 996
rect 5348 995 5354 999
rect 5357 997 5362 1003
rect 5406 1001 5415 1010
rect 5541 1001 5550 1010
rect 5550 1000 5556 1001
rect 4385 981 4401 984
rect 4403 981 4419 984
rect 4379 978 4399 981
rect 4520 979 4532 984
rect 4656 979 4657 983
rect 4664 980 4670 986
rect 4674 983 4742 987
rect 4761 986 4773 991
rect 4423 974 4424 978
rect 4381 972 4473 974
rect 4520 972 4540 979
rect 4655 974 4656 979
rect 4674 977 4700 983
rect 4710 980 4716 983
rect 4742 977 4755 983
rect 4773 978 4794 986
rect 4839 978 4873 991
rect 5005 988 5006 990
rect 4943 979 4949 985
rect 4959 983 4960 987
rect 5002 985 5005 986
rect 4654 972 4655 974
rect 4692 972 4700 977
rect 4285 963 4381 972
rect 4423 969 4424 972
rect 4382 963 4394 965
rect 4285 960 4382 963
rect 4276 957 4280 958
rect 4285 957 4381 960
rect 4276 956 4285 957
rect 4259 955 4283 956
rect 4287 955 4310 956
rect 4259 953 4278 955
rect 4327 954 4342 957
rect 4252 952 4259 953
rect 4272 952 4273 953
rect 4139 946 4145 952
rect 4197 946 4203 952
rect 4233 949 4252 952
rect 4320 951 4327 954
rect 4276 950 4287 951
rect 4318 950 4320 951
rect 4211 946 4233 949
rect 4203 945 4225 946
rect 4276 943 4288 950
rect 4339 944 4340 954
rect 4369 952 4379 957
rect 4378 944 4379 952
rect 4424 952 4435 968
rect 4424 951 4426 952
rect 4465 947 4466 968
rect 4473 965 4545 972
rect 4469 963 4545 965
rect 4473 956 4545 963
rect 4554 962 4555 968
rect 4548 956 4555 962
rect 4594 956 4600 962
rect 4649 956 4654 972
rect 4516 955 4557 956
rect 4542 950 4557 955
rect 4600 950 4606 956
rect 4396 942 4404 944
rect 4386 940 4396 942
rect 4384 939 4386 940
rect 3964 932 3966 933
rect 3937 927 3962 929
rect 3879 924 3881 925
rect 3702 914 3707 923
rect 3795 922 3825 924
rect 3875 922 3879 924
rect 3786 916 3795 922
rect 3825 916 3875 922
rect 3700 907 3702 914
rect 3668 895 3669 905
rect 3698 896 3700 907
rect 3771 906 3786 916
rect 3960 915 3962 927
rect 3966 917 3974 929
rect 4011 928 4023 934
rect 4075 928 4086 934
rect 4080 922 4086 928
rect 4197 926 4200 930
rect 4326 927 4384 939
rect 4426 938 4428 944
rect 4431 942 4477 944
rect 4477 940 4485 942
rect 4485 939 4488 940
rect 4396 930 4408 938
rect 4418 930 4430 938
rect 4321 926 4326 927
rect 3960 906 3963 915
rect 3999 910 4004 922
rect 4082 916 4089 922
rect 4089 914 4092 916
rect 4200 914 4214 926
rect 4307 923 4321 926
rect 4331 925 4339 927
rect 4428 926 4430 930
rect 4488 927 4535 939
rect 4548 935 4557 950
rect 4647 949 4649 956
rect 4665 952 4674 968
rect 4683 955 4692 972
rect 4755 968 4772 977
rect 4794 968 4833 978
rect 4646 946 4647 949
rect 4550 934 4552 935
rect 4600 933 4606 936
rect 4535 926 4540 927
rect 4548 926 4550 933
rect 4606 930 4613 933
rect 4623 930 4635 938
rect 4643 937 4645 942
rect 4665 937 4674 950
rect 4680 946 4683 955
rect 4725 954 4754 964
rect 4772 963 4833 968
rect 4772 957 4794 963
rect 4833 960 4843 963
rect 4718 945 4754 954
rect 4765 952 4774 954
rect 4677 937 4679 942
rect 4636 926 4643 937
rect 4665 934 4677 937
rect 4709 936 4718 945
rect 4725 944 4754 945
rect 4755 945 4774 952
rect 4794 950 4815 957
rect 4843 956 4853 960
rect 4873 956 4930 978
rect 4949 973 4955 979
rect 4960 977 4961 983
rect 5001 979 5007 985
rect 4961 972 4962 977
rect 4995 974 5001 979
rect 5002 974 5005 979
rect 4995 973 5002 974
rect 5001 972 5002 973
rect 4959 968 4962 972
rect 5010 971 5012 991
rect 5071 985 5077 991
rect 5082 988 5083 990
rect 5084 986 5087 987
rect 5087 985 5092 986
rect 5071 984 5127 985
rect 5276 984 5287 993
rect 5322 990 5334 994
rect 5348 993 5362 995
rect 5406 993 5412 999
rect 5550 998 5557 1000
rect 5559 998 5568 1018
rect 5643 1015 5656 1018
rect 6280 1015 6281 1026
rect 6470 1015 6471 1026
rect 6556 1015 6557 1026
rect 6829 1015 6830 1026
rect 7026 1015 7027 1026
rect 7262 1023 7301 1026
rect 8303 1023 8342 1028
rect 8528 1025 8534 1031
rect 8554 1026 8555 1031
rect 8553 1024 8554 1026
rect 7259 1022 7262 1023
rect 7259 1015 7271 1022
rect 7275 1016 7277 1022
rect 5656 1001 5720 1015
rect 5720 998 5730 1001
rect 5350 992 5360 993
rect 5397 992 5406 993
rect 5550 992 5568 998
rect 5611 992 5617 998
rect 5730 992 5775 998
rect 5870 994 5888 995
rect 5858 992 5870 994
rect 5322 986 5340 990
rect 5354 987 5360 992
rect 5400 987 5406 992
rect 5559 991 5565 992
rect 5559 989 5566 991
rect 5567 990 5568 992
rect 5597 991 5600 992
rect 5559 986 5565 989
rect 5567 987 5571 988
rect 5586 987 5597 991
rect 5602 986 5611 992
rect 5730 988 5858 992
rect 5071 983 5136 984
rect 5280 983 5288 984
rect 5088 981 5136 983
rect 5088 979 5100 981
rect 5282 978 5298 983
rect 5303 981 5304 984
rect 5130 972 5136 978
rect 5188 972 5194 978
rect 4959 967 4964 968
rect 5000 967 5001 971
rect 4950 958 4964 967
rect 4853 954 4858 956
rect 4930 955 4949 956
rect 4950 955 4962 958
rect 4858 951 4865 954
rect 4930 951 4962 955
rect 4964 951 4965 957
rect 4865 950 4867 951
rect 4755 944 4767 945
rect 4725 943 4732 944
rect 4774 943 4783 945
rect 4815 944 4853 950
rect 4868 949 4870 950
rect 4930 949 4950 951
rect 4953 949 4966 950
rect 4870 946 4879 949
rect 4943 948 4966 949
rect 4943 946 4950 948
rect 4953 945 4970 948
rect 4995 946 5000 967
rect 5012 951 5014 968
rect 5136 966 5142 972
rect 5145 967 5148 972
rect 5014 949 5019 950
rect 4953 944 4966 945
rect 4725 942 4730 943
rect 4725 941 4727 942
rect 4725 940 4771 941
rect 4772 940 4783 943
rect 4721 939 4726 940
rect 4733 939 4767 940
rect 4721 938 4767 939
rect 4721 937 4733 938
rect 4330 924 4331 925
rect 4298 921 4307 923
rect 4328 922 4330 924
rect 4286 920 4298 921
rect 4325 920 4328 922
rect 4256 916 4325 920
rect 4239 915 4256 916
rect 4227 914 4239 915
rect 4267 914 4286 916
rect 4384 914 4392 926
rect 4396 924 4430 926
rect 4092 913 4222 914
rect 4200 909 4214 913
rect 4256 911 4267 914
rect 4249 907 4255 911
rect 3767 900 3771 906
rect 3960 902 3962 906
rect 3697 891 3698 895
rect 3762 892 3767 899
rect 3945 898 3962 902
rect 3941 897 3962 898
rect 3937 896 3962 897
rect 3934 895 3962 896
rect 3966 895 3974 907
rect 4139 900 4145 906
rect 3949 891 3962 895
rect 3965 892 3966 894
rect 3696 888 3697 891
rect 3759 887 3762 891
rect 3936 889 3949 891
rect 3758 886 3759 887
rect 3885 886 3891 889
rect 3911 887 3949 889
rect 3911 886 3936 887
rect 3751 875 3758 885
rect 3850 875 3933 886
rect 3943 883 3949 887
rect 3950 883 3962 891
rect 3999 888 4004 900
rect 4145 894 4151 900
rect 4173 892 4186 900
rect 4216 892 4227 907
rect 4378 906 4383 913
rect 4241 900 4246 904
rect 4383 901 4387 906
rect 4387 899 4389 901
rect 4396 899 4398 924
rect 4173 889 4182 892
rect 4186 891 4188 892
rect 4228 889 4230 891
rect 4238 889 4247 898
rect 4389 892 4398 899
rect 4428 892 4430 924
rect 4434 914 4442 926
rect 4540 925 4550 926
rect 4540 923 4548 925
rect 4607 924 4635 926
rect 4546 922 4548 923
rect 4600 922 4601 924
rect 4633 922 4635 924
rect 4636 922 4647 926
rect 4545 921 4546 922
rect 4633 921 4647 922
rect 4466 916 4471 921
rect 4541 916 4545 921
rect 4599 917 4600 921
rect 4471 907 4480 916
rect 4535 907 4541 915
rect 4480 906 4535 907
rect 4542 904 4548 910
rect 4598 907 4599 916
rect 4633 915 4635 921
rect 4636 915 4647 921
rect 4670 925 4677 934
rect 4720 931 4733 937
rect 4764 936 4767 938
rect 4771 937 4783 940
rect 4853 937 4917 944
rect 4765 931 4767 936
rect 4778 931 4784 937
rect 4853 934 4949 937
rect 4953 934 4969 944
rect 4970 943 4980 945
rect 5012 944 5019 949
rect 5148 948 5155 967
rect 5182 966 5194 972
rect 5287 968 5298 978
rect 5322 980 5341 986
rect 5322 973 5359 980
rect 5483 976 5499 984
rect 5561 982 5564 986
rect 5560 976 5561 981
rect 5304 968 5307 972
rect 5188 945 5194 966
rect 5298 953 5310 968
rect 5326 965 5359 973
rect 5443 968 5446 976
rect 5484 975 5499 976
rect 5559 970 5560 975
rect 5602 969 5605 986
rect 5614 972 5715 977
rect 5715 969 5726 972
rect 5757 969 5858 988
rect 5888 980 5910 994
rect 5304 951 5307 953
rect 5310 951 5312 953
rect 5312 945 5325 951
rect 5341 948 5359 965
rect 5439 957 5443 968
rect 5434 955 5439 957
rect 5325 944 5327 945
rect 5397 944 5411 950
rect 5434 948 5446 955
rect 5433 947 5446 948
rect 5456 947 5468 955
rect 5499 952 5515 968
rect 5430 945 5439 947
rect 5007 943 5019 944
rect 4980 934 5044 943
rect 5327 942 5332 944
rect 5145 936 5227 942
rect 5128 934 5145 936
rect 4721 930 4733 931
rect 4670 924 4678 925
rect 4670 915 4677 924
rect 4678 922 4680 924
rect 4680 921 4682 922
rect 4681 918 4687 921
rect 4682 916 4687 918
rect 4633 911 4636 915
rect 4638 914 4647 915
rect 4638 912 4639 914
rect 4597 904 4598 906
rect 4600 904 4606 910
rect 4633 906 4635 911
rect 4639 907 4641 912
rect 4641 906 4642 907
rect 4632 904 4635 906
rect 4642 904 4643 906
rect 4548 898 4554 904
rect 4590 902 4593 904
rect 4594 902 4600 904
rect 4589 898 4600 902
rect 4631 901 4632 904
rect 4589 892 4596 898
rect 4630 897 4631 900
rect 4628 894 4630 895
rect 4633 894 4635 904
rect 4601 892 4635 894
rect 4639 899 4647 904
rect 4639 892 4653 899
rect 4628 891 4630 892
rect 4653 891 4654 892
rect 4654 890 4656 891
rect 3696 871 3697 875
rect 3749 871 3751 874
rect 3820 871 3850 875
rect 3748 870 3749 871
rect 3812 870 3820 871
rect 3810 869 3812 870
rect 3747 868 3748 869
rect 3808 868 3810 869
rect 3899 868 3901 875
rect 3934 868 3935 879
rect 3937 877 3943 883
rect 4017 882 4023 888
rect 4075 882 4081 888
rect 4011 876 4029 882
rect 4069 876 4075 882
rect 4182 880 4191 889
rect 4228 888 4238 889
rect 4626 888 4628 889
rect 4229 887 4238 888
rect 4229 880 4249 887
rect 4431 885 4432 888
rect 4392 882 4393 884
rect 4601 880 4613 888
rect 4623 882 4635 888
rect 4660 885 4670 915
rect 4687 912 4700 916
rect 4700 907 4712 912
rect 4715 906 4717 907
rect 4726 906 4733 930
rect 4778 928 4779 931
rect 4901 919 4949 934
rect 4969 932 5044 934
rect 5061 933 5112 934
rect 5114 933 5125 934
rect 5061 932 5122 933
rect 4969 930 5061 932
rect 4717 904 4722 906
rect 4726 904 4778 906
rect 4722 901 4778 904
rect 4726 899 4778 901
rect 4709 889 4718 898
rect 4726 896 4795 899
rect 4726 891 4783 896
rect 4795 892 4820 896
rect 4917 894 4925 919
rect 4949 916 4956 919
rect 4969 918 4985 930
rect 4987 918 5003 930
rect 5108 929 5123 932
rect 5104 927 5108 929
rect 5098 925 5104 927
rect 5114 926 5123 929
rect 5157 926 5164 936
rect 5094 924 5098 925
rect 5088 922 5094 924
rect 5117 920 5122 922
rect 4935 908 4937 916
rect 4956 914 4987 916
rect 4988 914 4990 918
rect 4956 909 4988 914
rect 4979 907 4996 909
rect 4937 900 4939 906
rect 4979 902 4988 907
rect 4996 906 5000 907
rect 4939 896 4940 899
rect 4959 898 4979 902
rect 4820 891 4826 892
rect 4720 889 4784 891
rect 4826 890 4832 891
rect 4916 890 4917 893
rect 4940 891 4941 896
rect 4954 891 4959 898
rect 5000 892 5057 906
rect 5057 891 5060 892
rect 4718 885 4784 889
rect 4832 887 4850 890
rect 4850 885 4862 887
rect 4915 885 4916 889
rect 4941 887 4942 891
rect 4656 884 4658 885
rect 4622 880 4635 882
rect 4192 875 4195 880
rect 4236 879 4249 880
rect 3734 864 3747 868
rect 3802 864 3808 868
rect 3728 862 3734 864
rect 3799 862 3802 864
rect 3724 856 3728 862
rect 3792 857 3799 862
rect 3791 856 3792 857
rect 3722 841 3724 855
rect 3788 849 3791 855
rect 3790 838 3799 842
rect 3837 838 3846 842
rect 3849 838 3865 854
rect 3867 838 3883 854
rect 3901 838 3905 867
rect 3932 847 3934 867
rect 3721 833 3722 838
rect 3788 833 3799 838
rect 3833 833 3849 838
rect 3781 832 3794 833
rect 3833 832 3855 833
rect 3720 825 3721 832
rect 3779 831 3788 832
rect 3719 819 3720 822
rect 3718 812 3719 816
rect 3718 804 3722 812
rect 3779 811 3781 831
rect 3782 826 3788 831
rect 3787 822 3788 826
rect 3820 824 3855 832
rect 3820 822 3849 824
rect 3894 822 3899 838
rect 3932 833 3933 838
rect 4040 833 4052 864
rect 4195 860 4202 875
rect 4234 873 4249 875
rect 4074 833 4086 838
rect 4097 837 4109 845
rect 4163 838 4179 854
rect 4202 842 4211 860
rect 4203 841 4211 842
rect 4215 845 4216 862
rect 4215 843 4219 845
rect 4247 844 4249 873
rect 4250 871 4252 874
rect 4253 871 4261 875
rect 4252 869 4261 871
rect 4253 863 4261 869
rect 4257 862 4258 863
rect 4258 859 4260 862
rect 4393 860 4397 879
rect 4430 866 4431 880
rect 4512 867 4518 873
rect 4558 867 4564 873
rect 4622 870 4626 880
rect 4655 870 4660 884
rect 4718 880 4732 885
rect 4726 871 4732 880
rect 4768 880 4778 885
rect 4768 870 4769 880
rect 4772 879 4778 880
rect 4862 879 4899 885
rect 4914 881 4915 885
rect 4900 874 4905 879
rect 4905 872 4907 874
rect 4911 871 4914 881
rect 4942 879 4944 885
rect 4951 881 4953 889
rect 5060 888 5074 891
rect 5120 890 5122 920
rect 5126 910 5134 922
rect 5164 914 5169 926
rect 5169 902 5174 914
rect 5194 910 5201 936
rect 5227 934 5231 936
rect 5308 935 5309 942
rect 5332 936 5344 942
rect 5231 933 5232 934
rect 5232 927 5235 933
rect 5235 925 5236 927
rect 5236 922 5238 924
rect 5238 919 5240 922
rect 5240 916 5241 919
rect 5091 888 5122 890
rect 5126 888 5134 900
rect 5174 899 5175 902
rect 5201 900 5203 910
rect 5241 906 5246 916
rect 5309 910 5313 935
rect 5344 934 5348 936
rect 5359 935 5360 942
rect 5346 933 5352 934
rect 5346 932 5354 933
rect 5360 932 5361 935
rect 5396 934 5411 944
rect 5429 943 5430 945
rect 5433 943 5439 945
rect 5472 943 5473 945
rect 5479 943 5485 948
rect 5422 942 5429 943
rect 5433 942 5468 943
rect 5472 942 5485 943
rect 5422 937 5433 942
rect 5434 941 5468 942
rect 5420 934 5426 937
rect 5427 936 5433 937
rect 5467 936 5468 941
rect 5485 936 5491 942
rect 5499 934 5515 950
rect 5553 944 5559 968
rect 5605 956 5606 968
rect 5610 965 5611 969
rect 5726 968 5745 969
rect 5753 968 5757 969
rect 5717 964 5753 968
rect 5803 965 5807 969
rect 5551 934 5553 943
rect 5416 932 5420 934
rect 5354 931 5395 932
rect 5360 918 5377 931
rect 5379 926 5395 931
rect 5413 930 5416 932
rect 5406 926 5413 930
rect 5379 918 5406 926
rect 5498 925 5499 931
rect 5550 927 5551 932
rect 5497 920 5499 925
rect 5549 924 5550 925
rect 5560 922 5568 934
rect 5572 922 5574 956
rect 5610 951 5611 964
rect 5717 960 5765 964
rect 5708 954 5717 960
rect 5605 945 5606 951
rect 5703 945 5708 954
rect 5746 949 5765 960
rect 5765 948 5767 949
rect 5807 948 5812 965
rect 5910 961 5913 980
rect 5913 954 5914 960
rect 5767 945 5771 948
rect 5812 945 5813 948
rect 5914 945 5916 954
rect 5611 936 5612 945
rect 5697 936 5703 944
rect 5612 928 5618 934
rect 5692 928 5704 936
rect 5714 928 5726 936
rect 5771 934 5786 945
rect 5813 934 5817 945
rect 5916 941 5917 944
rect 5914 934 5917 941
rect 5786 932 5787 934
rect 5787 928 5788 930
rect 5817 929 5819 934
rect 5613 922 5618 928
rect 5693 926 5697 928
rect 5730 926 5731 928
rect 5692 924 5693 925
rect 5732 924 5735 925
rect 5496 919 5499 920
rect 5246 902 5248 906
rect 5360 905 5361 918
rect 5388 916 5406 918
rect 5495 918 5499 919
rect 5495 916 5496 918
rect 5548 916 5549 919
rect 5568 916 5569 921
rect 5601 916 5606 922
rect 5613 916 5614 922
rect 5382 912 5388 916
rect 5491 909 5495 916
rect 5547 909 5548 916
rect 5569 912 5571 916
rect 5599 913 5601 916
rect 5594 911 5599 913
rect 5610 911 5614 916
rect 5680 912 5688 924
rect 5692 922 5726 924
rect 5692 921 5695 922
rect 5572 910 5610 911
rect 5361 902 5362 904
rect 5248 899 5250 902
rect 5203 894 5204 899
rect 5250 896 5251 899
rect 5251 892 5253 896
rect 5074 885 5085 888
rect 5088 887 5092 888
rect 5092 885 5101 887
rect 5085 884 5091 885
rect 4944 875 4945 879
rect 4945 872 4946 874
rect 4948 871 4951 881
rect 5101 879 5127 885
rect 5176 881 5178 889
rect 5110 876 5122 879
rect 5127 874 5149 879
rect 5178 874 5179 881
rect 5163 872 5168 874
rect 5168 871 5170 872
rect 5204 871 5208 890
rect 5253 888 5255 891
rect 5359 890 5362 896
rect 5368 891 5379 908
rect 5434 906 5440 909
rect 5546 908 5547 909
rect 5485 906 5491 908
rect 5594 906 5599 910
rect 5440 903 5446 906
rect 5475 903 5485 906
rect 5545 903 5546 906
rect 5592 903 5594 906
rect 5446 902 5475 903
rect 5590 899 5592 903
rect 5544 896 5545 899
rect 5427 890 5433 896
rect 5485 890 5491 896
rect 5543 892 5544 896
rect 5587 891 5590 898
rect 5255 886 5256 887
rect 5357 885 5359 889
rect 5365 886 5368 890
rect 5256 874 5263 885
rect 5263 871 5264 874
rect 5310 871 5313 885
rect 5347 881 5357 885
rect 5433 884 5439 890
rect 5443 887 5444 890
rect 5453 886 5460 890
rect 5444 883 5447 885
rect 5450 884 5452 885
rect 5479 884 5485 890
rect 5542 888 5543 891
rect 5680 890 5688 902
rect 5692 890 5694 921
rect 5725 920 5726 922
rect 5732 912 5738 924
rect 5788 913 5790 925
rect 5819 916 5835 928
rect 5905 925 5914 934
rect 5897 924 5905 925
rect 5885 922 5897 924
rect 5848 916 5885 922
rect 5819 913 5848 916
rect 5732 911 5735 912
rect 5735 899 5740 910
rect 5780 906 5835 913
rect 5773 905 5780 906
rect 5767 903 5773 905
rect 5754 899 5767 903
rect 5729 891 5754 899
rect 5726 890 5729 891
rect 5586 887 5587 890
rect 5735 888 5740 891
rect 5790 889 5792 906
rect 5585 885 5586 887
rect 5688 886 5691 888
rect 5740 886 5741 888
rect 5792 885 5793 888
rect 5444 882 5449 883
rect 5345 874 5363 881
rect 5339 871 5345 874
rect 4597 868 4598 869
rect 4621 867 4622 870
rect 4506 861 4512 867
rect 4564 861 4570 867
rect 4619 860 4621 867
rect 4260 854 4266 858
rect 4260 853 4275 854
rect 4246 843 4249 844
rect 4215 841 4249 843
rect 4253 850 4275 853
rect 4397 852 4398 858
rect 4431 854 4432 858
rect 4253 841 4261 850
rect 4266 840 4275 850
rect 3820 820 3840 822
rect 3848 820 3868 822
rect 3778 810 3781 811
rect 3779 804 3781 810
rect 3787 804 3803 820
rect 3840 819 3848 820
rect 3859 816 3894 817
rect 3893 812 3894 816
rect 3722 799 3741 804
rect 3752 799 3787 804
rect 3722 797 3752 799
rect 3771 788 3788 799
rect 3779 786 3788 788
rect 3781 780 3788 786
rect 3846 783 3855 786
rect 3859 785 3861 788
rect 3891 785 3893 788
rect 3904 786 3905 828
rect 3932 820 3937 833
rect 4032 831 4109 833
rect 3929 804 3945 820
rect 3932 789 3937 804
rect 3945 789 3961 803
rect 4004 795 4023 798
rect 3917 787 3942 789
rect 3945 788 3970 789
rect 3917 785 3919 787
rect 4032 786 4090 831
rect 4107 801 4109 831
rect 4113 821 4121 833
rect 4179 822 4195 838
rect 4249 837 4253 840
rect 4273 838 4275 840
rect 4297 838 4303 844
rect 4343 839 4349 844
rect 4339 838 4351 839
rect 4398 838 4401 850
rect 4433 841 4449 854
rect 4504 852 4512 858
rect 4502 850 4512 852
rect 4616 851 4619 860
rect 4565 848 4575 850
rect 4575 846 4581 848
rect 4614 847 4616 851
rect 4492 844 4506 846
rect 4581 844 4588 846
rect 4432 840 4449 841
rect 4432 838 4436 840
rect 4215 829 4227 837
rect 4237 829 4249 837
rect 4275 832 4355 838
rect 4215 828 4216 829
rect 4104 799 4109 801
rect 4110 812 4113 819
rect 4216 818 4218 828
rect 4275 822 4291 832
rect 4297 827 4349 832
rect 4143 812 4179 816
rect 4218 814 4220 818
rect 4110 805 4179 812
rect 4220 809 4221 812
rect 4221 805 4222 809
rect 3859 783 3893 785
rect 3840 782 3868 783
rect 3825 780 3868 782
rect 3781 777 3794 780
rect 3834 777 3840 780
rect 3846 777 3855 780
rect 3857 779 3868 780
rect 4023 780 4090 786
rect 4110 791 4171 805
rect 4179 791 4199 805
rect 4222 799 4223 803
rect 4223 795 4224 799
rect 4297 793 4317 827
rect 4357 815 4363 827
rect 4343 793 4351 795
rect 4357 793 4363 805
rect 4379 804 4387 820
rect 4402 814 4405 829
rect 4417 822 4436 838
rect 4470 833 4479 842
rect 4492 841 4512 844
rect 4588 843 4592 844
rect 4592 842 4597 843
rect 4613 842 4614 844
rect 4609 841 4620 842
rect 4645 841 4655 869
rect 4660 866 4661 868
rect 4661 856 4663 862
rect 4732 860 4737 870
rect 4908 868 4911 870
rect 4907 865 4911 868
rect 4908 860 4911 865
rect 4938 864 4948 870
rect 5170 869 5176 871
rect 5179 869 5185 870
rect 5176 868 5185 869
rect 5179 866 5185 868
rect 5179 864 5191 866
rect 4938 862 4949 864
rect 4663 854 4664 855
rect 4737 854 4738 860
rect 4907 858 4909 860
rect 4907 854 4908 858
rect 4663 852 4667 854
rect 4664 841 4667 852
rect 4729 849 4745 854
rect 4728 848 4742 849
rect 4747 848 4763 854
rect 4720 841 4728 848
rect 4742 842 4765 848
rect 4492 838 4506 841
rect 4612 839 4613 841
rect 4620 840 4655 841
rect 4666 840 4667 841
rect 4718 840 4720 841
rect 4645 839 4693 840
rect 4716 838 4718 840
rect 4732 839 4744 842
rect 4825 841 4841 854
rect 4843 841 4859 854
rect 4905 847 4907 853
rect 4909 852 4910 855
rect 4765 840 4766 841
rect 4818 840 4819 841
rect 4737 838 4744 839
rect 4486 834 4500 838
rect 4486 833 4497 834
rect 4461 824 4470 833
rect 4432 820 4436 822
rect 4417 814 4436 820
rect 4405 809 4406 812
rect 4406 799 4408 808
rect 4417 804 4433 814
rect 4492 812 4500 824
rect 4504 814 4506 838
rect 4609 832 4612 838
rect 4598 831 4612 832
rect 4598 822 4610 831
rect 4564 815 4570 821
rect 4605 818 4607 822
rect 4610 818 4616 822
rect 4604 815 4605 818
rect 4616 816 4618 818
rect 4558 814 4564 815
rect 4603 814 4604 815
rect 4504 812 4538 814
rect 4547 812 4606 814
rect 4618 813 4622 816
rect 4617 812 4623 813
rect 4436 808 4437 812
rect 4528 809 4538 812
rect 4542 810 4547 812
rect 4519 808 4528 809
rect 4531 808 4537 809
rect 4539 808 4542 810
rect 4558 809 4564 812
rect 4437 804 4438 808
rect 4504 805 4516 808
rect 4519 805 4538 808
rect 4504 804 4517 805
rect 4433 800 4438 804
rect 4495 800 4516 804
rect 4526 800 4538 805
rect 4594 800 4603 811
rect 4606 810 4614 812
rect 4617 810 4628 812
rect 4636 811 4645 838
rect 4667 822 4683 838
rect 4707 832 4715 838
rect 4614 809 4628 810
rect 4630 809 4636 810
rect 4614 808 4636 809
rect 4667 808 4683 820
rect 4736 811 4738 838
rect 4739 837 4744 838
rect 4741 836 4744 837
rect 4766 838 4767 840
rect 4817 838 4818 840
rect 4871 838 4874 841
rect 4903 839 4905 847
rect 4938 838 4948 862
rect 4949 855 4954 862
rect 4954 852 4956 855
rect 4956 848 4959 852
rect 5086 842 5092 844
rect 5086 838 5100 842
rect 5132 838 5138 844
rect 5139 838 5155 854
rect 5179 838 5185 864
rect 5191 863 5194 864
rect 5194 856 5196 862
rect 5196 853 5197 855
rect 5197 838 5202 852
rect 4742 834 4746 836
rect 4747 832 4748 834
rect 4740 828 4744 830
rect 4617 804 4683 808
rect 4626 800 4667 804
rect 4707 801 4708 804
rect 4433 797 4440 800
rect 4495 797 4515 800
rect 4433 794 4441 797
rect 4433 793 4443 794
rect 4224 792 4225 793
rect 4297 792 4349 793
rect 4355 792 4371 793
rect 4433 792 4445 793
rect 4110 784 4139 791
rect 4225 789 4231 792
rect 4231 784 4238 789
rect 4291 788 4371 792
rect 4409 790 4410 792
rect 4433 789 4454 792
rect 4433 788 4448 789
rect 4291 786 4355 788
rect 4443 786 4448 788
rect 4454 787 4459 789
rect 4459 786 4463 787
rect 4464 786 4495 797
rect 4527 793 4531 800
rect 4589 793 4594 799
rect 4526 790 4527 793
rect 4587 790 4589 793
rect 4238 783 4239 784
rect 4274 783 4275 785
rect 4023 777 4099 780
rect 4240 779 4246 783
rect 4271 779 4274 783
rect 4297 780 4303 786
rect 4339 781 4351 786
rect 4459 785 4470 786
rect 4461 783 4470 785
rect 4461 782 4473 783
rect 4343 780 4349 781
rect 4409 779 4410 781
rect 4246 777 4251 779
rect 4270 777 4271 779
rect 4408 777 4409 779
rect 4461 777 4470 782
rect 4476 779 4479 781
rect 4479 777 4498 779
rect 4526 777 4535 786
rect 4557 782 4563 788
rect 4584 786 4587 790
rect 4603 782 4609 788
rect 4621 786 4630 800
rect 4633 788 4649 800
rect 4651 796 4687 800
rect 4708 798 4709 801
rect 4735 800 4736 810
rect 4742 798 4744 828
rect 4748 818 4756 830
rect 4766 822 4779 838
rect 4809 836 4817 838
rect 4874 837 4875 838
rect 4809 823 4816 836
rect 4833 826 4845 832
rect 4830 825 4889 826
rect 4893 825 4903 838
rect 4830 823 4838 825
rect 4889 823 4903 825
rect 4910 824 4912 832
rect 4766 820 4768 822
rect 4829 821 4830 823
rect 4766 814 4779 820
rect 4710 797 4744 798
rect 4709 796 4744 797
rect 4748 796 4756 808
rect 4765 804 4779 814
rect 4821 816 4829 820
rect 4833 818 4840 820
rect 4821 808 4827 816
rect 4833 814 4834 818
rect 4893 816 4918 823
rect 4927 816 4938 837
rect 4959 822 4971 838
rect 5080 832 5086 838
rect 5096 832 5121 838
rect 5138 832 5144 838
rect 5155 832 5171 838
rect 5185 832 5186 838
rect 5202 832 5204 838
rect 5084 830 5086 832
rect 5088 830 5096 832
rect 5138 830 5171 832
rect 5204 830 5205 832
rect 5208 830 5220 870
rect 5264 869 5265 871
rect 5265 865 5267 868
rect 5267 863 5268 864
rect 5268 859 5270 862
rect 5294 838 5310 870
rect 5334 869 5339 871
rect 5347 870 5357 874
rect 5332 868 5334 869
rect 5328 866 5332 868
rect 5327 865 5328 866
rect 5326 863 5327 864
rect 5324 859 5326 862
rect 5340 859 5347 870
rect 5322 856 5324 859
rect 5320 854 5322 855
rect 5313 851 5322 854
rect 5313 839 5320 851
rect 5313 838 5314 839
rect 5294 830 5313 838
rect 5327 830 5340 859
rect 5357 846 5364 858
rect 5369 848 5370 880
rect 5436 876 5442 879
rect 5433 874 5436 876
rect 5424 869 5433 874
rect 5444 870 5447 882
rect 5481 870 5484 884
rect 5541 881 5542 885
rect 5540 874 5541 881
rect 5581 874 5585 885
rect 5691 884 5693 885
rect 5692 883 5694 884
rect 5692 879 5695 883
rect 5741 880 5742 882
rect 5692 878 5696 879
rect 5695 876 5696 878
rect 5742 876 5743 880
rect 5793 876 5794 879
rect 5819 878 5835 906
rect 5539 871 5540 874
rect 5580 872 5581 874
rect 5417 860 5418 863
rect 5447 860 5449 870
rect 5481 862 5495 870
rect 5579 869 5580 871
rect 5696 869 5699 874
rect 5538 868 5539 869
rect 5537 864 5538 867
rect 5577 864 5579 868
rect 5576 862 5577 864
rect 5699 863 5701 869
rect 5412 848 5417 860
rect 5369 847 5374 848
rect 5369 846 5403 847
rect 5410 846 5415 848
rect 5364 844 5365 846
rect 5409 844 5410 846
rect 5406 842 5408 843
rect 5369 834 5381 841
rect 5391 834 5403 841
rect 5449 830 5460 859
rect 5484 830 5495 862
rect 5634 861 5635 862
rect 5536 856 5537 859
rect 5574 856 5576 861
rect 5701 860 5702 863
rect 5535 855 5536 856
rect 5513 851 5529 854
rect 5533 851 5535 854
rect 5572 851 5574 855
rect 5615 854 5627 855
rect 5513 843 5533 851
rect 5569 843 5572 851
rect 5609 849 5627 854
rect 5637 849 5649 855
rect 5609 843 5700 849
rect 5702 848 5706 860
rect 5706 844 5707 847
rect 5723 843 5739 854
rect 5511 839 5514 843
rect 5567 839 5569 843
rect 5603 842 5608 843
rect 5603 840 5607 842
rect 5609 841 5649 843
rect 5596 839 5606 840
rect 5609 839 5615 841
rect 5590 838 5595 839
rect 5609 838 5610 839
rect 5497 830 5511 838
rect 5564 836 5567 838
rect 5586 837 5590 838
rect 5577 836 5583 837
rect 5564 834 5577 836
rect 5554 833 5558 834
rect 5548 832 5554 833
rect 5564 832 5567 834
rect 5535 830 5548 832
rect 5076 827 5084 830
rect 5088 828 5091 830
rect 5075 821 5085 827
rect 4764 802 4765 804
rect 4766 800 4768 804
rect 4893 801 4903 816
rect 4905 812 4913 816
rect 4905 804 4914 812
rect 4918 807 4950 816
rect 4959 807 4971 820
rect 5051 807 5075 821
rect 5076 818 5084 821
rect 4914 801 4915 803
rect 4651 788 4667 796
rect 4687 795 4692 796
rect 4692 793 4703 795
rect 4710 794 4717 796
rect 4717 793 4723 794
rect 4734 793 4735 796
rect 4703 792 4708 793
rect 4723 792 4743 793
rect 4746 792 4748 795
rect 4763 794 4764 796
rect 4723 786 4744 792
rect 4760 789 4763 793
rect 4745 788 4763 789
rect 4745 786 4760 788
rect 4816 786 4817 788
rect 4821 786 4827 798
rect 4875 789 4876 797
rect 4890 790 4893 800
rect 4915 797 4924 801
rect 4927 800 4938 807
rect 4950 804 4971 807
rect 4925 797 4927 800
rect 4950 797 4969 804
rect 5039 800 5051 807
rect 5037 799 5039 800
rect 4921 796 4969 797
rect 5030 796 5037 799
rect 5076 796 5084 808
rect 5088 796 5090 828
rect 5156 822 5385 830
rect 5156 821 5157 822
rect 5159 820 5385 822
rect 5157 814 5385 820
rect 5413 814 5535 830
rect 5560 822 5564 831
rect 5593 822 5609 838
rect 5558 818 5560 822
rect 5557 817 5558 818
rect 5557 816 5563 817
rect 5556 815 5563 816
rect 5157 812 5413 814
rect 5158 804 5171 812
rect 5188 807 5190 812
rect 5158 803 5159 804
rect 5159 801 5160 802
rect 5157 798 5159 801
rect 5189 800 5190 807
rect 5201 804 5213 812
rect 5213 803 5214 804
rect 5218 803 5220 808
rect 5237 803 5316 812
rect 5214 802 5316 803
rect 5217 799 5233 802
rect 5156 796 5157 797
rect 4921 793 4959 796
rect 4969 795 4971 796
rect 4834 787 4835 788
rect 4833 786 4839 787
rect 4615 782 4621 786
rect 4732 784 4744 786
rect 3668 755 3669 777
rect 3697 772 3698 777
rect 3788 774 3827 777
rect 3834 774 3846 777
rect 3698 759 3706 772
rect 3790 768 3827 774
rect 3837 768 3846 774
rect 3903 768 3904 777
rect 3698 755 3709 759
rect 3669 749 3670 755
rect 3706 753 3709 755
rect 3707 750 3712 753
rect 3681 747 3710 748
rect 3713 747 3714 749
rect 3663 713 3670 725
rect 3675 716 3676 747
rect 3704 745 3709 747
rect 3708 716 3709 745
rect 3710 738 3721 747
rect 3937 740 3941 777
rect 4032 768 4041 777
rect 4084 768 4090 777
rect 4246 776 4270 777
rect 4406 772 4408 777
rect 4470 772 4498 777
rect 4399 759 4406 772
rect 4470 768 4479 772
rect 4517 768 4526 777
rect 4551 776 4557 782
rect 4609 776 4621 782
rect 4733 776 4734 781
rect 4609 766 4613 773
rect 4765 772 4766 786
rect 4817 783 4818 786
rect 4828 784 4830 785
rect 4874 784 4875 788
rect 4889 787 4890 790
rect 4915 789 4959 793
rect 4971 792 4978 795
rect 5028 793 5030 796
rect 5127 795 5155 796
rect 4978 789 4982 792
rect 4915 788 4937 789
rect 4939 788 4955 789
rect 4982 788 4984 789
rect 5024 788 5028 793
rect 5139 792 5155 795
rect 5185 793 5189 799
rect 4896 787 4903 788
rect 4911 787 4925 788
rect 4984 787 4987 788
rect 4888 786 4896 787
rect 4883 785 4896 786
rect 4915 785 4925 787
rect 5080 786 5086 792
rect 5138 791 5155 792
rect 5182 791 5185 793
rect 5138 789 5194 791
rect 5215 789 5233 799
rect 5138 788 5155 789
rect 5182 788 5185 789
rect 5194 788 5233 789
rect 5235 788 5316 802
rect 5327 800 5340 812
rect 5403 804 5404 807
rect 5138 786 5144 788
rect 5181 786 5182 788
rect 4880 784 4889 785
rect 4818 780 4830 783
rect 4833 780 4834 781
rect 4842 780 4880 784
rect 4818 779 4877 780
rect 4833 774 4845 779
rect 4764 763 4766 772
rect 4883 763 4889 784
rect 4915 784 4929 785
rect 4389 756 4406 759
rect 4730 756 4733 763
rect 4389 755 4399 756
rect 4389 754 4396 755
rect 4729 754 4730 756
rect 4389 753 4393 754
rect 4378 749 4420 753
rect 4378 748 4405 749
rect 4420 748 4421 749
rect 4376 747 4378 748
rect 4421 747 4423 748
rect 4362 745 4376 747
rect 3894 738 3900 740
rect 3937 739 3946 740
rect 3714 735 3732 738
rect 3721 725 3732 735
rect 3894 734 3906 738
rect 3940 734 3946 739
rect 4329 738 4362 745
rect 4323 737 4328 738
rect 3888 728 3894 734
rect 3946 729 3952 734
rect 4300 733 4323 737
rect 4377 735 4385 747
rect 4389 746 4394 747
rect 4294 731 4300 733
rect 4288 729 4290 731
rect 3910 728 4041 729
rect 3894 726 3910 728
rect 3946 727 4249 728
rect 4276 727 4282 729
rect 4287 728 4288 729
rect 4041 726 4042 727
rect 4249 726 4282 727
rect 4285 726 4287 728
rect 3675 714 3679 716
rect 3706 714 3709 716
rect 3675 713 3709 714
rect 3714 713 3732 725
rect 3882 714 3890 726
rect 3894 724 3900 726
rect 3670 711 3671 713
rect 3671 708 3676 711
rect 3709 708 3714 711
rect 3675 707 3687 708
rect 3674 701 3687 707
rect 3697 701 3709 708
rect 3721 707 3732 713
rect 3732 706 3737 707
rect 3674 694 3676 701
rect 3732 694 3739 706
rect 3737 690 3739 694
rect 3882 692 3890 704
rect 3894 694 3896 724
rect 4043 719 4047 726
rect 4249 723 4284 726
rect 4322 723 4328 729
rect 4047 708 4054 719
rect 4270 717 4276 723
rect 4277 719 4284 723
rect 4328 719 4334 723
rect 4377 719 4385 725
rect 4389 719 4391 746
rect 4718 744 4724 750
rect 4726 744 4729 754
rect 4764 750 4765 763
rect 4870 757 4876 762
rect 4882 757 4883 762
rect 4915 758 4925 784
rect 4929 783 4933 784
rect 4988 783 4994 786
rect 5023 783 5024 786
rect 5086 784 5100 786
rect 5086 783 5092 784
rect 5124 783 5128 784
rect 4995 781 4997 782
rect 4997 780 5000 781
rect 5013 780 5023 783
rect 4942 775 4948 779
rect 4948 772 4953 775
rect 5000 772 5023 780
rect 4954 766 4978 772
rect 5013 769 5045 772
rect 5051 769 5124 783
rect 5132 780 5138 786
rect 5139 784 5140 785
rect 5180 784 5181 786
rect 5215 783 5218 788
rect 5224 787 5316 788
rect 5288 786 5316 787
rect 5265 785 5316 786
rect 5324 785 5327 799
rect 5402 797 5403 801
rect 5449 800 5460 814
rect 5484 804 5495 814
rect 5497 804 5513 814
rect 5550 807 5563 815
rect 5547 805 5563 807
rect 5593 805 5609 820
rect 5647 811 5649 841
rect 5653 831 5661 843
rect 5700 838 5740 843
rect 5743 842 5750 874
rect 5785 840 5793 852
rect 5797 842 5799 874
rect 5829 869 5831 874
rect 5829 868 5832 869
rect 5829 842 5831 868
rect 5832 862 5833 864
rect 5833 857 5834 862
rect 5834 852 5835 855
rect 5797 840 5831 842
rect 5835 840 5843 852
rect 5750 838 5751 840
rect 5740 837 5755 838
rect 5797 837 5798 838
rect 5749 836 5755 837
rect 5794 836 5796 837
rect 5631 809 5649 811
rect 5653 809 5661 821
rect 5710 805 5720 836
rect 5749 832 5764 836
rect 5752 808 5764 832
rect 5797 828 5809 836
rect 5819 828 5831 836
rect 5837 834 5851 838
rect 5838 828 5851 834
rect 5798 824 5799 828
rect 5839 822 5851 828
rect 5799 820 5800 822
rect 5751 807 5764 808
rect 5536 804 5649 805
rect 5513 803 5649 804
rect 5401 791 5402 796
rect 5400 788 5401 791
rect 5460 789 5463 799
rect 5495 794 5503 800
rect 5513 795 5529 803
rect 5531 797 5649 803
rect 5720 801 5724 805
rect 5750 804 5764 807
rect 5785 815 5800 820
rect 5839 820 5840 822
rect 5839 816 5851 820
rect 6291 819 6292 1015
rect 6481 819 6482 1015
rect 6567 819 6568 1015
rect 6840 819 6841 1015
rect 7037 819 7038 1015
rect 7259 1013 7275 1015
rect 7281 1013 7293 1022
rect 7301 1020 7330 1023
rect 7330 1014 7334 1020
rect 8070 1018 8122 1020
rect 8342 1018 8356 1023
rect 8552 1020 8553 1023
rect 8042 1016 8122 1018
rect 8042 1015 8093 1016
rect 7334 1013 7335 1014
rect 8017 1013 8042 1015
rect 8064 1014 8070 1015
rect 8093 1014 8098 1015
rect 7255 1011 7259 1013
rect 7271 1010 7275 1013
rect 7983 1011 8013 1013
rect 8059 1012 8064 1014
rect 7247 998 7255 1010
rect 7254 988 7255 998
rect 7259 1007 7293 1010
rect 7259 1003 7261 1007
rect 7259 996 7260 1003
rect 7271 1001 7275 1007
rect 7290 1005 7293 1007
rect 7296 1004 7305 1010
rect 7258 994 7260 996
rect 7257 988 7263 994
rect 7268 988 7271 1001
rect 7251 982 7257 988
rect 7254 976 7255 982
rect 7258 962 7259 988
rect 7291 982 7293 1004
rect 7297 998 7305 1004
rect 7335 1001 7344 1010
rect 7866 1005 7880 1007
rect 7892 1005 7983 1011
rect 8055 1007 8059 1012
rect 7866 1004 7892 1005
rect 7866 1003 7880 1004
rect 7860 1002 7880 1003
rect 7901 1002 7906 1005
rect 8051 1002 8055 1007
rect 8098 1005 8115 1014
rect 8115 1004 8117 1005
rect 7303 988 7309 994
rect 7326 992 7335 1001
rect 7851 997 7875 1002
rect 7906 997 7912 1002
rect 8050 1001 8051 1002
rect 8122 1001 8139 1016
rect 8356 1015 8363 1018
rect 8551 1016 8552 1020
rect 8363 1014 8366 1015
rect 8366 1005 8388 1014
rect 8549 1012 8551 1016
rect 8589 1014 8593 1031
rect 8595 1027 8603 1039
rect 8861 1037 8873 1045
rect 8922 1041 8932 1045
rect 8933 1041 8939 1045
rect 8897 1037 8939 1041
rect 8991 1039 8997 1045
rect 9144 1044 9150 1050
rect 9190 1048 9200 1050
rect 10855 1048 10864 1057
rect 10920 1048 10929 1057
rect 12119 1048 12128 1057
rect 9153 1044 9165 1048
rect 9175 1044 9187 1048
rect 9190 1044 9196 1048
rect 9138 1038 9144 1044
rect 9196 1038 9202 1044
rect 11834 1038 11840 1044
rect 11880 1038 11886 1044
rect 12142 1043 12154 1051
rect 12164 1043 12176 1051
rect 12184 1048 12193 1057
rect 12243 1051 12259 1052
rect 12138 1040 12140 1043
rect 12178 1040 12180 1043
rect 12237 1039 12248 1051
rect 12511 1048 12520 1057
rect 12576 1051 12585 1057
rect 12517 1045 12520 1047
rect 12524 1045 12530 1051
rect 12570 1048 12585 1051
rect 12711 1048 12720 1057
rect 12776 1050 12785 1057
rect 12570 1045 12576 1048
rect 8642 1020 8652 1036
rect 8673 1034 8685 1037
rect 8867 1036 8873 1037
rect 8919 1036 8922 1037
rect 8667 1033 8687 1034
rect 8861 1033 8867 1036
rect 8903 1033 8933 1036
rect 8667 1031 8673 1033
rect 8687 1031 8717 1033
rect 8664 1025 8667 1031
rect 8661 1022 8667 1025
rect 8719 1024 8740 1031
rect 8767 1024 8773 1030
rect 8388 1004 8391 1005
rect 8248 1001 8249 1004
rect 7849 996 7851 997
rect 7309 982 7315 988
rect 7326 986 7330 992
rect 7838 989 7849 996
rect 7860 993 7875 997
rect 7912 996 7913 997
rect 7324 974 7325 979
rect 7482 976 7498 984
rect 7665 976 7681 989
rect 7748 979 7765 989
rect 7824 981 7838 989
rect 7818 979 7824 981
rect 7765 978 7818 979
rect 7849 977 7857 989
rect 7861 987 7866 989
rect 7913 987 7925 996
rect 7482 974 7539 976
rect 7320 957 7324 972
rect 7482 968 7527 974
rect 7539 968 7543 974
rect 7258 944 7265 957
rect 7319 953 7320 956
rect 7318 949 7319 952
rect 7321 944 7335 953
rect 7466 952 7482 968
rect 7543 961 7548 968
rect 7473 944 7482 952
rect 7251 936 7257 942
rect 7257 930 7263 936
rect 7265 934 7290 944
rect 7305 936 7321 944
rect 7303 934 7321 936
rect 7469 935 7473 944
rect 7476 940 7482 941
rect 7476 939 7518 940
rect 7522 939 7528 941
rect 7476 936 7487 939
rect 7476 935 7482 936
rect 7518 935 7528 939
rect 7469 934 7476 935
rect 7296 929 7299 934
rect 7303 930 7309 934
rect 7292 923 7295 928
rect 7466 925 7469 934
rect 7470 929 7476 934
rect 7528 929 7534 935
rect 7535 933 7547 941
rect 7608 934 7614 940
rect 7654 934 7660 940
rect 7665 934 7671 956
rect 7730 952 7736 958
rect 7776 952 7782 958
rect 7849 956 7857 967
rect 7861 958 7863 987
rect 8111 984 8113 1001
rect 8117 999 8139 1001
rect 8117 989 8125 999
rect 8243 992 8248 1001
rect 8391 996 8412 1004
rect 8546 1002 8549 1011
rect 8589 1007 8591 1014
rect 8580 1005 8591 1007
rect 8595 1010 8603 1017
rect 8595 1005 8608 1010
rect 8593 1004 8594 1005
rect 8599 1001 8608 1005
rect 8642 1002 8652 1018
rect 8661 1015 8664 1022
rect 8715 1018 8721 1024
rect 8773 1018 8779 1024
rect 8849 1021 8857 1033
rect 8861 1031 8895 1033
rect 8861 1030 8867 1031
rect 8861 1029 8864 1030
rect 8661 1014 8663 1015
rect 8661 1013 8665 1014
rect 8663 1001 8665 1013
rect 8545 996 8546 997
rect 8301 995 8334 996
rect 8412 995 8414 996
rect 8336 993 8342 995
rect 8243 986 8249 992
rect 8301 987 8307 992
rect 8342 991 8346 993
rect 8414 991 8424 995
rect 8544 991 8545 995
rect 8586 993 8599 1001
rect 8661 998 8665 1001
rect 8849 999 8857 1011
rect 8861 1002 8863 1029
rect 9141 1024 9144 1036
rect 9196 1032 9199 1036
rect 11828 1032 11834 1038
rect 11886 1032 11892 1038
rect 9149 1018 9153 1031
rect 9196 1021 9212 1032
rect 12119 1031 12125 1037
rect 12130 1031 12138 1039
rect 12141 1037 12176 1039
rect 12141 1036 12142 1037
rect 12140 1031 12141 1035
rect 12142 1031 12143 1036
rect 12174 1031 12176 1037
rect 10862 1026 10864 1030
rect 9212 1018 9228 1021
rect 8938 1007 8939 1008
rect 8939 1005 8940 1006
rect 8861 1001 8864 1002
rect 8907 1001 8935 1002
rect 8861 999 8873 1001
rect 8907 1000 8933 1001
rect 8591 992 8599 993
rect 8652 991 8656 996
rect 8661 991 8666 998
rect 8861 997 8862 999
rect 8907 998 8929 1000
rect 8935 999 8939 1001
rect 8862 996 8863 997
rect 8907 996 8922 998
rect 8863 995 8865 996
rect 8861 993 8867 995
rect 8907 994 8923 996
rect 8933 995 8939 999
rect 8942 997 8947 1003
rect 8991 1001 9000 1010
rect 9126 1001 9135 1010
rect 9135 1000 9141 1001
rect 7970 981 7986 984
rect 7988 981 8004 984
rect 7964 978 7984 981
rect 8105 979 8117 984
rect 8241 979 8242 983
rect 8249 980 8255 986
rect 8259 983 8327 987
rect 8346 986 8358 991
rect 8008 974 8009 978
rect 7966 972 8058 974
rect 8105 972 8125 979
rect 8240 974 8241 979
rect 8259 977 8285 983
rect 8295 980 8301 983
rect 8327 977 8340 983
rect 8358 978 8379 986
rect 8424 978 8458 991
rect 8590 988 8591 990
rect 8528 979 8534 985
rect 8544 983 8545 987
rect 8587 985 8590 986
rect 8239 972 8240 974
rect 8277 972 8285 977
rect 7870 963 7966 972
rect 8008 969 8009 972
rect 7967 963 7979 965
rect 7870 960 7967 963
rect 7861 957 7865 958
rect 7870 957 7966 960
rect 7861 956 7870 957
rect 7844 955 7868 956
rect 7872 955 7895 956
rect 7844 953 7863 955
rect 7912 954 7927 957
rect 7837 952 7844 953
rect 7857 952 7858 953
rect 7724 946 7730 952
rect 7782 946 7788 952
rect 7818 949 7837 952
rect 7905 951 7912 954
rect 7861 950 7872 951
rect 7903 950 7905 951
rect 7796 946 7818 949
rect 7788 945 7810 946
rect 7861 943 7873 950
rect 7924 944 7925 954
rect 7954 952 7964 957
rect 7963 944 7964 952
rect 8009 952 8020 968
rect 8009 951 8011 952
rect 8050 947 8051 968
rect 8058 965 8130 972
rect 8054 963 8130 965
rect 8058 956 8130 963
rect 8139 962 8140 968
rect 8133 956 8140 962
rect 8179 956 8185 962
rect 8234 956 8239 972
rect 8101 955 8142 956
rect 8127 950 8142 955
rect 8185 950 8191 956
rect 7981 942 7989 944
rect 7971 940 7981 942
rect 7969 939 7971 940
rect 7549 932 7551 933
rect 7522 927 7547 929
rect 7464 924 7466 925
rect 7287 914 7292 923
rect 7380 922 7410 924
rect 7460 922 7464 924
rect 7371 916 7380 922
rect 7410 916 7460 922
rect 7285 907 7287 914
rect 7253 895 7254 905
rect 7283 896 7285 907
rect 7356 906 7371 916
rect 7545 915 7547 927
rect 7551 917 7559 929
rect 7596 928 7608 934
rect 7660 928 7671 934
rect 7665 922 7671 928
rect 7782 926 7785 930
rect 7911 927 7969 939
rect 8011 938 8013 944
rect 8016 942 8062 944
rect 8062 940 8070 942
rect 8070 939 8073 940
rect 7981 930 7993 938
rect 8003 930 8015 938
rect 7906 926 7911 927
rect 7545 906 7548 915
rect 7584 910 7589 922
rect 7667 916 7674 922
rect 7674 914 7677 916
rect 7785 914 7799 926
rect 7892 923 7906 926
rect 7916 925 7924 927
rect 8013 926 8015 930
rect 8073 927 8120 939
rect 8133 935 8142 950
rect 8232 949 8234 956
rect 8250 952 8259 968
rect 8268 955 8277 972
rect 8340 968 8357 977
rect 8379 968 8418 978
rect 8231 946 8232 949
rect 8135 934 8137 935
rect 8185 933 8191 936
rect 8120 926 8125 927
rect 8133 926 8135 933
rect 8191 930 8198 933
rect 8208 930 8220 938
rect 8228 937 8230 942
rect 8250 937 8259 950
rect 8265 946 8268 955
rect 8310 954 8339 964
rect 8357 963 8418 968
rect 8357 957 8379 963
rect 8418 960 8428 963
rect 8303 945 8339 954
rect 8350 952 8359 954
rect 8262 937 8264 942
rect 8221 926 8228 937
rect 8250 934 8262 937
rect 8294 936 8303 945
rect 8310 944 8339 945
rect 8340 945 8359 952
rect 8379 950 8400 957
rect 8428 956 8438 960
rect 8458 956 8515 978
rect 8534 973 8540 979
rect 8545 977 8546 983
rect 8586 979 8592 985
rect 8546 972 8547 977
rect 8580 974 8586 979
rect 8587 974 8590 979
rect 8580 973 8587 974
rect 8586 972 8587 973
rect 8544 968 8547 972
rect 8595 971 8597 991
rect 8656 985 8662 991
rect 8667 988 8668 990
rect 8669 986 8672 987
rect 8672 985 8677 986
rect 8656 984 8712 985
rect 8861 984 8872 993
rect 8907 990 8919 994
rect 8933 993 8947 995
rect 8991 993 8997 999
rect 9135 998 9142 1000
rect 9144 998 9153 1018
rect 9228 1015 9241 1018
rect 9865 1015 9866 1026
rect 10055 1015 10056 1026
rect 10141 1015 10142 1026
rect 10414 1015 10415 1026
rect 10611 1015 10612 1026
rect 10847 1023 10886 1026
rect 11888 1023 11927 1028
rect 12113 1025 12119 1031
rect 12139 1026 12140 1031
rect 12138 1024 12139 1026
rect 10844 1022 10847 1023
rect 10844 1015 10856 1022
rect 10860 1016 10862 1022
rect 9241 1001 9305 1015
rect 9305 998 9315 1001
rect 8935 992 8945 993
rect 8982 992 8991 993
rect 9135 992 9153 998
rect 9196 992 9202 998
rect 9315 992 9360 998
rect 9455 994 9473 995
rect 9443 992 9455 994
rect 8907 986 8925 990
rect 8939 987 8945 992
rect 8985 987 8991 992
rect 9144 991 9150 992
rect 9144 989 9151 991
rect 9152 990 9153 992
rect 9182 991 9185 992
rect 9144 986 9150 989
rect 9152 987 9156 988
rect 9171 987 9182 991
rect 9187 986 9196 992
rect 9315 988 9443 992
rect 8656 983 8721 984
rect 8865 983 8873 984
rect 8673 981 8721 983
rect 8673 979 8685 981
rect 8867 978 8883 983
rect 8888 981 8889 984
rect 8715 972 8721 978
rect 8773 972 8779 978
rect 8544 967 8549 968
rect 8585 967 8586 971
rect 8535 958 8549 967
rect 8438 954 8443 956
rect 8515 955 8534 956
rect 8535 955 8547 958
rect 8443 951 8450 954
rect 8515 951 8547 955
rect 8549 951 8550 957
rect 8450 950 8452 951
rect 8340 944 8352 945
rect 8310 943 8317 944
rect 8359 943 8368 945
rect 8400 944 8438 950
rect 8453 949 8455 950
rect 8515 949 8535 951
rect 8538 949 8551 950
rect 8455 946 8464 949
rect 8528 948 8551 949
rect 8528 946 8535 948
rect 8538 945 8555 948
rect 8580 946 8585 967
rect 8597 951 8599 968
rect 8721 966 8727 972
rect 8730 967 8733 972
rect 8599 949 8604 950
rect 8538 944 8551 945
rect 8310 942 8315 943
rect 8310 941 8312 942
rect 8310 940 8356 941
rect 8357 940 8368 943
rect 8306 939 8311 940
rect 8318 939 8352 940
rect 8306 938 8352 939
rect 8306 937 8318 938
rect 7915 924 7916 925
rect 7883 921 7892 923
rect 7913 922 7915 924
rect 7871 920 7883 921
rect 7910 920 7913 922
rect 7841 916 7910 920
rect 7824 915 7841 916
rect 7812 914 7824 915
rect 7852 914 7871 916
rect 7969 914 7977 926
rect 7981 924 8015 926
rect 7677 913 7807 914
rect 7785 909 7799 913
rect 7841 911 7852 914
rect 7834 907 7840 911
rect 7352 900 7356 906
rect 7545 902 7547 906
rect 7282 891 7283 895
rect 7347 892 7352 899
rect 7530 898 7547 902
rect 7526 897 7547 898
rect 7522 896 7547 897
rect 7519 895 7547 896
rect 7551 895 7559 907
rect 7724 900 7730 906
rect 7534 891 7547 895
rect 7550 892 7551 894
rect 7281 888 7282 891
rect 7344 887 7347 891
rect 7521 889 7534 891
rect 7343 886 7344 887
rect 7470 886 7476 889
rect 7496 887 7534 889
rect 7496 886 7521 887
rect 7336 875 7343 885
rect 7435 875 7518 886
rect 7528 883 7534 887
rect 7535 883 7547 891
rect 7584 888 7589 900
rect 7730 894 7736 900
rect 7758 892 7771 900
rect 7801 892 7812 907
rect 7963 906 7968 913
rect 7826 900 7831 904
rect 7968 901 7972 906
rect 7972 899 7974 901
rect 7981 899 7983 924
rect 7758 889 7767 892
rect 7771 891 7773 892
rect 7813 889 7815 891
rect 7823 889 7832 898
rect 7974 892 7983 899
rect 8013 892 8015 924
rect 8019 914 8027 926
rect 8125 925 8135 926
rect 8125 923 8133 925
rect 8192 924 8220 926
rect 8131 922 8133 923
rect 8185 922 8186 924
rect 8218 922 8220 924
rect 8221 922 8232 926
rect 8130 921 8131 922
rect 8218 921 8232 922
rect 8051 916 8056 921
rect 8126 916 8130 921
rect 8184 917 8185 921
rect 8056 907 8065 916
rect 8120 907 8126 915
rect 8065 906 8120 907
rect 8127 904 8133 910
rect 8183 907 8184 916
rect 8218 915 8220 921
rect 8221 915 8232 921
rect 8255 925 8262 934
rect 8305 931 8318 937
rect 8349 936 8352 938
rect 8356 937 8368 940
rect 8438 937 8502 944
rect 8350 931 8352 936
rect 8363 931 8369 937
rect 8438 934 8534 937
rect 8538 934 8554 944
rect 8555 943 8565 945
rect 8597 944 8604 949
rect 8733 948 8740 967
rect 8767 966 8779 972
rect 8872 968 8883 978
rect 8907 980 8926 986
rect 8907 973 8944 980
rect 9068 976 9084 984
rect 9146 982 9149 986
rect 9145 976 9146 981
rect 8889 968 8892 972
rect 8773 945 8779 966
rect 8883 953 8895 968
rect 8911 965 8944 973
rect 9028 968 9031 976
rect 9069 975 9084 976
rect 9144 970 9145 975
rect 9187 969 9190 986
rect 9199 972 9300 977
rect 9300 969 9311 972
rect 9342 969 9443 988
rect 9473 980 9495 994
rect 8889 951 8892 953
rect 8895 951 8897 953
rect 8897 945 8910 951
rect 8926 948 8944 965
rect 9024 957 9028 968
rect 9019 955 9024 957
rect 8910 944 8912 945
rect 8982 944 8996 950
rect 9019 948 9031 955
rect 9018 947 9031 948
rect 9041 947 9053 955
rect 9084 952 9100 968
rect 9015 945 9024 947
rect 8592 943 8604 944
rect 8565 934 8629 943
rect 8912 942 8917 944
rect 8730 936 8812 942
rect 8713 934 8730 936
rect 8306 930 8318 931
rect 8255 924 8263 925
rect 8255 915 8262 924
rect 8263 922 8265 924
rect 8265 921 8267 922
rect 8266 918 8272 921
rect 8267 916 8272 918
rect 8218 911 8221 915
rect 8223 914 8232 915
rect 8223 912 8224 914
rect 8182 904 8183 906
rect 8185 904 8191 910
rect 8218 906 8220 911
rect 8224 907 8226 912
rect 8226 906 8227 907
rect 8217 904 8220 906
rect 8227 904 8228 906
rect 8133 898 8139 904
rect 8175 902 8178 904
rect 8179 902 8185 904
rect 8174 898 8185 902
rect 8216 901 8217 904
rect 8174 892 8181 898
rect 8215 897 8216 900
rect 8213 894 8215 895
rect 8218 894 8220 904
rect 8186 892 8220 894
rect 8224 899 8232 904
rect 8224 892 8238 899
rect 8213 891 8215 892
rect 8238 891 8239 892
rect 8239 890 8241 891
rect 7281 871 7282 875
rect 7334 871 7336 874
rect 7405 871 7435 875
rect 7333 870 7334 871
rect 7397 870 7405 871
rect 7395 869 7397 870
rect 7332 868 7333 869
rect 7393 868 7395 869
rect 7484 868 7486 875
rect 7519 868 7520 879
rect 7522 877 7528 883
rect 7602 882 7608 888
rect 7660 882 7666 888
rect 7596 876 7614 882
rect 7654 876 7660 882
rect 7767 880 7776 889
rect 7813 888 7823 889
rect 8211 888 8213 889
rect 7814 887 7823 888
rect 7814 880 7834 887
rect 8016 885 8017 888
rect 7977 882 7978 884
rect 8186 880 8198 888
rect 8208 882 8220 888
rect 8245 885 8255 915
rect 8272 912 8285 916
rect 8285 907 8297 912
rect 8300 906 8302 907
rect 8311 906 8318 930
rect 8363 928 8364 931
rect 8486 919 8534 934
rect 8554 932 8629 934
rect 8646 933 8697 934
rect 8699 933 8710 934
rect 8646 932 8707 933
rect 8554 930 8646 932
rect 8302 904 8307 906
rect 8311 904 8363 906
rect 8307 901 8363 904
rect 8311 899 8363 901
rect 8294 889 8303 898
rect 8311 896 8380 899
rect 8311 891 8368 896
rect 8380 892 8405 896
rect 8502 894 8510 919
rect 8534 916 8541 919
rect 8554 918 8570 930
rect 8572 918 8588 930
rect 8693 929 8708 932
rect 8689 927 8693 929
rect 8683 925 8689 927
rect 8699 926 8708 929
rect 8742 926 8749 936
rect 8679 924 8683 925
rect 8673 922 8679 924
rect 8702 920 8707 922
rect 8520 908 8522 916
rect 8541 914 8572 916
rect 8573 914 8575 918
rect 8541 909 8573 914
rect 8564 907 8581 909
rect 8522 900 8524 906
rect 8564 902 8573 907
rect 8581 906 8585 907
rect 8524 896 8525 899
rect 8544 898 8564 902
rect 8405 891 8411 892
rect 8305 889 8369 891
rect 8411 890 8417 891
rect 8501 890 8502 893
rect 8525 891 8526 896
rect 8539 891 8544 898
rect 8585 892 8642 906
rect 8642 891 8645 892
rect 8303 885 8369 889
rect 8417 887 8435 890
rect 8435 885 8447 887
rect 8500 885 8501 889
rect 8526 887 8527 891
rect 8241 884 8243 885
rect 8207 880 8220 882
rect 7777 875 7780 880
rect 7821 879 7834 880
rect 7319 864 7332 868
rect 7387 864 7393 868
rect 7313 862 7319 864
rect 7384 862 7387 864
rect 7309 856 7313 862
rect 7377 857 7384 862
rect 7376 856 7377 857
rect 7307 841 7309 855
rect 7373 849 7376 855
rect 7375 838 7384 842
rect 7422 838 7431 842
rect 7434 838 7450 854
rect 7452 838 7468 854
rect 7486 838 7490 867
rect 7517 847 7519 867
rect 7306 833 7307 838
rect 7373 833 7384 838
rect 7418 833 7434 838
rect 7366 832 7379 833
rect 7418 832 7440 833
rect 7305 825 7306 832
rect 7364 831 7373 832
rect 7304 819 7305 822
rect 5785 804 5801 815
rect 5840 805 5851 816
rect 5841 804 5851 805
rect 7303 812 7304 816
rect 7303 804 7307 812
rect 7364 811 7366 831
rect 7367 826 7373 831
rect 7372 822 7373 826
rect 7405 824 7440 832
rect 7405 822 7434 824
rect 7479 822 7484 838
rect 7517 833 7518 838
rect 7625 833 7637 864
rect 7780 860 7787 875
rect 7819 873 7834 875
rect 7659 833 7671 838
rect 7682 837 7694 845
rect 7748 838 7764 854
rect 7787 842 7796 860
rect 7788 841 7796 842
rect 7800 845 7801 862
rect 7800 843 7804 845
rect 7832 844 7834 873
rect 7835 871 7837 874
rect 7838 871 7846 875
rect 7837 869 7846 871
rect 7838 863 7846 869
rect 7842 862 7843 863
rect 7843 859 7845 862
rect 7978 860 7982 879
rect 8015 866 8016 880
rect 8097 867 8103 873
rect 8143 867 8149 873
rect 8207 870 8211 880
rect 8240 870 8245 884
rect 8303 880 8317 885
rect 8311 871 8317 880
rect 8353 880 8363 885
rect 8353 870 8354 880
rect 8357 879 8363 880
rect 8447 879 8484 885
rect 8499 881 8500 885
rect 8485 874 8490 879
rect 8490 872 8492 874
rect 8496 871 8499 881
rect 8527 879 8529 885
rect 8536 881 8538 889
rect 8645 888 8659 891
rect 8705 890 8707 920
rect 8711 910 8719 922
rect 8749 914 8754 926
rect 8754 902 8759 914
rect 8779 910 8786 936
rect 8812 934 8816 936
rect 8893 935 8894 942
rect 8917 936 8929 942
rect 8816 933 8817 934
rect 8817 927 8820 933
rect 8820 925 8821 927
rect 8821 922 8823 924
rect 8823 919 8825 922
rect 8825 916 8826 919
rect 8676 888 8707 890
rect 8711 888 8719 900
rect 8759 899 8760 902
rect 8786 900 8788 910
rect 8826 906 8831 916
rect 8894 910 8898 935
rect 8929 934 8933 936
rect 8944 935 8945 942
rect 8931 933 8937 934
rect 8931 932 8939 933
rect 8945 932 8946 935
rect 8981 934 8996 944
rect 9014 943 9015 945
rect 9018 943 9024 945
rect 9057 943 9058 945
rect 9064 943 9070 948
rect 9007 942 9014 943
rect 9018 942 9053 943
rect 9057 942 9070 943
rect 9007 937 9018 942
rect 9019 941 9053 942
rect 9005 934 9011 937
rect 9012 936 9018 937
rect 9052 936 9053 941
rect 9070 936 9076 942
rect 9084 934 9100 950
rect 9138 944 9144 968
rect 9190 956 9191 968
rect 9195 965 9196 969
rect 9311 968 9330 969
rect 9338 968 9342 969
rect 9302 964 9338 968
rect 9388 965 9392 969
rect 9136 934 9138 943
rect 9001 932 9005 934
rect 8939 931 8980 932
rect 8945 918 8962 931
rect 8964 926 8980 931
rect 8998 930 9001 932
rect 8991 926 8998 930
rect 8964 918 8991 926
rect 9083 925 9084 931
rect 9135 927 9136 932
rect 9082 920 9084 925
rect 9134 924 9135 925
rect 9145 922 9153 934
rect 9157 922 9159 956
rect 9195 951 9196 964
rect 9302 960 9350 964
rect 9293 954 9302 960
rect 9190 945 9191 951
rect 9288 945 9293 954
rect 9331 949 9350 960
rect 9350 948 9352 949
rect 9392 948 9397 965
rect 9495 961 9498 980
rect 9498 954 9499 960
rect 9352 945 9356 948
rect 9397 945 9398 948
rect 9499 945 9501 954
rect 9196 936 9197 945
rect 9282 936 9288 944
rect 9197 928 9203 934
rect 9277 928 9289 936
rect 9299 928 9311 936
rect 9356 934 9371 945
rect 9398 934 9402 945
rect 9501 941 9502 944
rect 9499 934 9502 941
rect 9371 932 9372 934
rect 9372 928 9373 930
rect 9402 929 9404 934
rect 9198 922 9203 928
rect 9278 926 9282 928
rect 9315 926 9316 928
rect 9277 924 9278 925
rect 9317 924 9320 925
rect 9081 919 9084 920
rect 8831 902 8833 906
rect 8945 905 8946 918
rect 8973 916 8991 918
rect 9080 918 9084 919
rect 9080 916 9081 918
rect 9133 916 9134 919
rect 9153 916 9154 921
rect 9186 916 9191 922
rect 9198 916 9199 922
rect 8967 912 8973 916
rect 9076 909 9080 916
rect 9132 909 9133 916
rect 9154 912 9156 916
rect 9184 913 9186 916
rect 9179 911 9184 913
rect 9195 911 9199 916
rect 9265 912 9273 924
rect 9277 922 9311 924
rect 9277 921 9280 922
rect 9157 910 9195 911
rect 8946 902 8947 904
rect 8833 899 8835 902
rect 8788 894 8789 899
rect 8835 896 8836 899
rect 8836 892 8838 896
rect 8659 885 8670 888
rect 8673 887 8677 888
rect 8677 885 8686 887
rect 8670 884 8676 885
rect 8529 875 8530 879
rect 8530 872 8531 874
rect 8533 871 8536 881
rect 8686 879 8712 885
rect 8761 881 8763 889
rect 8695 876 8707 879
rect 8712 874 8734 879
rect 8763 874 8764 881
rect 8748 872 8753 874
rect 8753 871 8755 872
rect 8789 871 8793 890
rect 8838 888 8840 891
rect 8944 890 8947 896
rect 8953 891 8964 908
rect 9019 906 9025 909
rect 9131 908 9132 909
rect 9070 906 9076 908
rect 9179 906 9184 910
rect 9025 903 9031 906
rect 9060 903 9070 906
rect 9130 903 9131 906
rect 9177 903 9179 906
rect 9031 902 9060 903
rect 9175 899 9177 903
rect 9129 896 9130 899
rect 9012 890 9018 896
rect 9070 890 9076 896
rect 9128 892 9129 896
rect 9172 891 9175 898
rect 8840 886 8841 887
rect 8942 885 8944 889
rect 8950 886 8953 890
rect 8841 874 8848 885
rect 8848 871 8849 874
rect 8895 871 8898 885
rect 8932 881 8942 885
rect 9018 884 9024 890
rect 9028 887 9029 890
rect 9038 886 9045 890
rect 9029 883 9032 885
rect 9035 884 9037 885
rect 9064 884 9070 890
rect 9127 888 9128 891
rect 9265 890 9273 902
rect 9277 890 9279 921
rect 9310 920 9311 922
rect 9317 912 9323 924
rect 9373 913 9375 925
rect 9404 916 9420 928
rect 9490 925 9499 934
rect 9482 924 9490 925
rect 9470 922 9482 924
rect 9433 916 9470 922
rect 9404 913 9433 916
rect 9317 911 9320 912
rect 9320 899 9325 910
rect 9365 906 9420 913
rect 9358 905 9365 906
rect 9352 903 9358 905
rect 9339 899 9352 903
rect 9314 891 9339 899
rect 9311 890 9314 891
rect 9171 887 9172 890
rect 9320 888 9325 891
rect 9375 889 9377 906
rect 9170 885 9171 887
rect 9273 886 9276 888
rect 9325 886 9326 888
rect 9377 885 9378 888
rect 9029 882 9034 883
rect 8930 874 8948 881
rect 8924 871 8930 874
rect 8182 868 8183 869
rect 8206 867 8207 870
rect 8091 861 8097 867
rect 8149 861 8155 867
rect 8204 860 8206 867
rect 7845 854 7851 858
rect 7845 853 7860 854
rect 7831 843 7834 844
rect 7800 841 7834 843
rect 7838 850 7860 853
rect 7982 852 7983 858
rect 8016 854 8017 858
rect 7838 841 7846 850
rect 7851 840 7860 850
rect 7405 820 7425 822
rect 7433 820 7453 822
rect 7363 810 7366 811
rect 7364 804 7366 810
rect 7372 804 7388 820
rect 7425 819 7433 820
rect 7444 816 7479 817
rect 7478 812 7479 816
rect 5749 803 5750 804
rect 5748 801 5749 802
rect 5696 799 5739 801
rect 5657 797 5696 799
rect 5531 796 5657 797
rect 5531 795 5637 796
rect 5720 795 5739 799
rect 5513 794 5547 795
rect 5495 792 5529 794
rect 5474 789 5503 792
rect 5389 785 5400 788
rect 5449 787 5474 789
rect 5436 786 5449 787
rect 5432 785 5436 786
rect 5291 784 5294 785
rect 5312 784 5400 785
rect 5312 783 5389 784
rect 5405 783 5432 785
rect 5460 784 5463 787
rect 5134 779 5135 780
rect 5172 769 5180 783
rect 5214 778 5215 783
rect 5290 781 5291 783
rect 5313 782 5315 783
rect 5289 778 5290 781
rect 5315 780 5318 782
rect 5323 781 5324 783
rect 5381 782 5385 783
rect 5389 782 5405 783
rect 5370 779 5381 782
rect 5318 778 5321 779
rect 4870 756 4888 757
rect 4916 756 4922 758
rect 4864 750 4928 756
rect 4953 753 4983 766
rect 5013 763 5051 769
rect 5169 763 5172 769
rect 5013 759 5045 763
rect 5012 756 5013 758
rect 4953 750 4989 753
rect 5010 752 5012 756
rect 5014 755 5045 759
rect 5042 754 5044 755
rect 5045 754 5048 755
rect 5164 754 5169 763
rect 5041 752 5042 754
rect 5048 751 5053 754
rect 5163 752 5164 754
rect 4764 744 4770 750
rect 4870 745 4922 750
rect 4674 742 4718 744
rect 4523 741 4557 742
rect 4674 741 4680 742
rect 4486 740 4523 741
rect 4463 739 4486 740
rect 4460 737 4463 739
rect 4712 738 4718 742
rect 4770 738 4776 744
rect 4435 723 4460 737
rect 4551 730 4557 736
rect 4609 731 4615 736
rect 4864 733 4876 745
rect 4910 735 4915 745
rect 4640 731 4676 733
rect 4557 724 4563 730
rect 4581 729 4640 731
rect 4676 729 4682 731
rect 4579 726 4581 729
rect 4430 720 4435 723
rect 4328 717 4410 719
rect 4331 716 4410 717
rect 4427 716 4435 720
rect 4377 713 4385 716
rect 4389 715 4391 716
rect 4410 715 4439 716
rect 4389 713 4423 715
rect 4420 709 4423 713
rect 4427 713 4435 715
rect 4439 714 4467 715
rect 4427 711 4430 713
rect 4424 709 4427 711
rect 4467 710 4481 714
rect 4573 713 4579 726
rect 4603 724 4609 729
rect 4682 726 4693 729
rect 4870 726 4876 733
rect 4672 722 4674 723
rect 4693 722 4704 726
rect 4869 723 4876 726
rect 4704 721 4706 722
rect 4706 720 4710 721
rect 4054 707 4055 708
rect 4276 707 4277 708
rect 4389 701 4401 709
rect 4411 701 4423 709
rect 4481 705 4487 710
rect 4571 708 4573 713
rect 4570 707 4571 708
rect 4487 703 4498 705
rect 4115 697 4249 700
rect 4415 698 4419 701
rect 4498 699 4511 703
rect 4511 698 4516 699
rect 3991 695 4115 697
rect 4249 695 4255 697
rect 3894 692 3900 694
rect 3969 692 3991 695
rect 4255 692 4261 695
rect 4407 694 4415 698
rect 4516 694 4532 698
rect 4564 694 4570 706
rect 3676 688 3677 690
rect 3677 669 3687 688
rect 3739 674 3755 690
rect 3890 688 3892 691
rect 3946 689 3969 692
rect 4261 689 4267 692
rect 4399 690 4407 694
rect 4532 692 4548 694
rect 4664 693 4672 698
rect 4676 693 4678 720
rect 4864 711 4876 723
rect 4915 711 4917 726
rect 4953 723 4983 750
rect 5009 749 5010 751
rect 5053 750 5055 751
rect 4993 746 4995 747
rect 5007 745 5009 749
rect 4996 737 5010 745
rect 5038 744 5040 749
rect 5058 747 5061 749
rect 5061 746 5063 747
rect 5063 743 5067 746
rect 5087 743 5099 749
rect 5158 744 5161 749
rect 5193 744 5214 778
rect 5280 756 5289 778
rect 5318 776 5323 778
rect 5336 776 5370 779
rect 5463 778 5464 781
rect 5318 775 5336 776
rect 5318 756 5323 775
rect 5464 772 5468 778
rect 5464 756 5471 772
rect 5495 756 5503 789
rect 5513 788 5529 792
rect 5531 788 5547 794
rect 5609 788 5625 795
rect 5723 788 5739 795
rect 5726 787 5727 788
rect 5727 783 5728 785
rect 5729 772 5732 779
rect 5752 778 5764 804
rect 5801 797 5802 802
rect 5840 798 5841 800
rect 7307 799 7326 804
rect 7337 799 7372 804
rect 7307 797 7337 799
rect 5801 796 5803 797
rect 5839 796 5840 797
rect 5801 791 5809 796
rect 5836 791 5839 796
rect 5801 788 5817 791
rect 5819 788 5835 791
rect 7356 788 7373 799
rect 7364 786 7373 788
rect 7366 780 7373 786
rect 7431 783 7440 786
rect 7444 785 7446 788
rect 7476 785 7478 788
rect 7489 786 7490 828
rect 7517 820 7522 833
rect 7617 831 7694 833
rect 7514 804 7530 820
rect 7517 789 7522 804
rect 7530 789 7546 803
rect 7589 795 7608 798
rect 7502 787 7527 789
rect 7530 788 7555 789
rect 7502 785 7504 787
rect 7617 786 7675 831
rect 7692 801 7694 831
rect 7698 821 7706 833
rect 7764 822 7780 838
rect 7834 837 7838 840
rect 7858 838 7860 840
rect 7882 838 7888 844
rect 7928 839 7934 844
rect 7924 838 7936 839
rect 7983 838 7986 850
rect 8018 841 8034 854
rect 8089 852 8097 858
rect 8087 850 8097 852
rect 8201 851 8204 860
rect 8150 848 8160 850
rect 8160 846 8166 848
rect 8199 847 8201 851
rect 8077 844 8091 846
rect 8166 844 8173 846
rect 8017 840 8034 841
rect 8017 838 8021 840
rect 7800 829 7812 837
rect 7822 829 7834 837
rect 7860 832 7940 838
rect 7800 828 7801 829
rect 7689 799 7694 801
rect 7695 812 7698 819
rect 7801 818 7803 828
rect 7860 822 7876 832
rect 7882 827 7934 832
rect 7728 812 7764 816
rect 7803 814 7805 818
rect 7695 805 7764 812
rect 7805 809 7806 812
rect 7806 805 7807 809
rect 7444 783 7478 785
rect 7425 782 7453 783
rect 7410 780 7453 782
rect 5275 745 5280 756
rect 5315 744 5318 756
rect 5468 750 5471 756
rect 5468 744 5475 750
rect 5503 744 5505 756
rect 5533 751 5545 759
rect 5555 751 5567 759
rect 5732 755 5737 772
rect 5764 770 5768 778
rect 7366 777 7379 780
rect 7419 777 7425 780
rect 7431 777 7440 780
rect 7442 779 7453 780
rect 7608 780 7675 786
rect 7695 791 7756 805
rect 7764 791 7784 805
rect 7807 799 7808 803
rect 7808 795 7809 799
rect 7882 793 7902 827
rect 7942 815 7948 827
rect 7928 793 7936 795
rect 7942 793 7948 805
rect 7964 804 7972 820
rect 7987 814 7990 829
rect 8002 822 8021 838
rect 8055 833 8064 842
rect 8077 841 8097 844
rect 8173 843 8177 844
rect 8177 842 8182 843
rect 8198 842 8199 844
rect 8194 841 8205 842
rect 8230 841 8240 869
rect 8245 866 8246 868
rect 8246 856 8248 862
rect 8317 860 8322 870
rect 8493 868 8496 870
rect 8492 865 8496 868
rect 8493 860 8496 865
rect 8523 864 8533 870
rect 8755 869 8761 871
rect 8764 869 8770 870
rect 8761 868 8770 869
rect 8764 866 8770 868
rect 8764 864 8776 866
rect 8523 862 8534 864
rect 8248 854 8249 855
rect 8322 854 8323 860
rect 8492 858 8494 860
rect 8492 854 8493 858
rect 8248 852 8252 854
rect 8249 841 8252 852
rect 8314 849 8330 854
rect 8313 848 8327 849
rect 8332 848 8348 854
rect 8305 841 8313 848
rect 8327 842 8350 848
rect 8077 838 8091 841
rect 8197 839 8198 841
rect 8205 840 8240 841
rect 8251 840 8252 841
rect 8303 840 8305 841
rect 8230 839 8278 840
rect 8301 838 8303 840
rect 8317 839 8329 842
rect 8410 841 8426 854
rect 8428 841 8444 854
rect 8490 847 8492 853
rect 8494 852 8495 855
rect 8350 840 8351 841
rect 8403 840 8404 841
rect 8322 838 8329 839
rect 8071 834 8085 838
rect 8071 833 8082 834
rect 8046 824 8055 833
rect 8017 820 8021 822
rect 8002 814 8021 820
rect 7990 809 7991 812
rect 7991 799 7993 808
rect 8002 804 8018 814
rect 8077 812 8085 824
rect 8089 814 8091 838
rect 8194 832 8197 838
rect 8183 831 8197 832
rect 8183 822 8195 831
rect 8149 815 8155 821
rect 8190 818 8192 822
rect 8195 818 8201 822
rect 8189 815 8190 818
rect 8201 816 8203 818
rect 8143 814 8149 815
rect 8188 814 8189 815
rect 8089 812 8123 814
rect 8132 812 8191 814
rect 8203 813 8207 816
rect 8202 812 8208 813
rect 8021 808 8022 812
rect 8113 809 8123 812
rect 8127 810 8132 812
rect 8104 808 8113 809
rect 8116 808 8122 809
rect 8124 808 8127 810
rect 8143 809 8149 812
rect 8022 804 8023 808
rect 8089 805 8101 808
rect 8104 805 8123 808
rect 8089 804 8102 805
rect 8018 800 8023 804
rect 8080 800 8101 804
rect 8111 800 8123 805
rect 8179 800 8188 811
rect 8191 810 8199 812
rect 8202 810 8213 812
rect 8221 811 8230 838
rect 8252 822 8268 838
rect 8292 832 8300 838
rect 8199 809 8213 810
rect 8215 809 8221 810
rect 8199 808 8221 809
rect 8252 808 8268 820
rect 8321 811 8323 838
rect 8324 837 8329 838
rect 8326 836 8329 837
rect 8351 838 8352 840
rect 8402 838 8403 840
rect 8456 838 8459 841
rect 8488 839 8490 847
rect 8523 838 8533 862
rect 8534 855 8539 862
rect 8539 852 8541 855
rect 8541 848 8544 852
rect 8671 842 8677 844
rect 8671 838 8685 842
rect 8717 838 8723 844
rect 8724 838 8740 854
rect 8764 838 8770 864
rect 8776 863 8779 864
rect 8779 856 8781 862
rect 8781 853 8782 855
rect 8782 838 8787 852
rect 8327 834 8331 836
rect 8332 832 8333 834
rect 8325 828 8329 830
rect 8202 804 8268 808
rect 8211 800 8252 804
rect 8292 801 8293 804
rect 8018 797 8025 800
rect 8080 797 8100 800
rect 8018 794 8026 797
rect 8018 793 8028 794
rect 7809 792 7810 793
rect 7882 792 7934 793
rect 7940 792 7956 793
rect 8018 792 8030 793
rect 7695 784 7724 791
rect 7810 789 7816 792
rect 7816 784 7823 789
rect 7876 788 7956 792
rect 7994 790 7995 792
rect 8018 789 8039 792
rect 8018 788 8033 789
rect 7876 786 7940 788
rect 8028 786 8033 788
rect 8039 787 8044 789
rect 8044 786 8048 787
rect 8049 786 8080 797
rect 8112 793 8116 800
rect 8174 793 8179 799
rect 8111 790 8112 793
rect 8172 790 8174 793
rect 7823 783 7824 784
rect 7859 783 7860 785
rect 7608 777 7684 780
rect 7825 779 7831 783
rect 7856 779 7859 783
rect 7882 780 7888 786
rect 7924 781 7936 786
rect 8044 785 8055 786
rect 8046 783 8055 785
rect 8046 782 8058 783
rect 7928 780 7934 781
rect 7994 779 7995 781
rect 7831 777 7836 779
rect 7855 777 7856 779
rect 7993 777 7994 779
rect 8046 777 8055 782
rect 8061 779 8064 781
rect 8064 777 8083 779
rect 8111 777 8120 786
rect 8142 782 8148 788
rect 8169 786 8172 790
rect 8188 782 8194 788
rect 8206 786 8215 800
rect 8218 788 8234 800
rect 8236 796 8272 800
rect 8293 798 8294 801
rect 8320 800 8321 810
rect 8327 798 8329 828
rect 8333 818 8341 830
rect 8351 822 8364 838
rect 8394 836 8402 838
rect 8459 837 8460 838
rect 8394 823 8401 836
rect 8418 826 8430 832
rect 8415 825 8474 826
rect 8478 825 8488 838
rect 8415 823 8423 825
rect 8474 823 8488 825
rect 8495 824 8497 832
rect 8351 820 8353 822
rect 8414 821 8415 823
rect 8351 814 8364 820
rect 8295 797 8329 798
rect 8294 796 8329 797
rect 8333 796 8341 808
rect 8350 804 8364 814
rect 8406 816 8414 820
rect 8418 818 8425 820
rect 8406 808 8412 816
rect 8418 814 8419 818
rect 8478 816 8503 823
rect 8512 816 8523 837
rect 8544 822 8556 838
rect 8665 832 8671 838
rect 8681 832 8706 838
rect 8723 832 8729 838
rect 8740 832 8756 838
rect 8770 832 8771 838
rect 8787 832 8789 838
rect 8669 830 8671 832
rect 8673 830 8681 832
rect 8723 830 8756 832
rect 8789 830 8790 832
rect 8793 830 8805 870
rect 8849 869 8850 871
rect 8850 865 8852 868
rect 8852 863 8853 864
rect 8853 859 8855 862
rect 8879 838 8895 870
rect 8919 869 8924 871
rect 8932 870 8942 874
rect 8917 868 8919 869
rect 8913 866 8917 868
rect 8912 865 8913 866
rect 8911 863 8912 864
rect 8909 859 8911 862
rect 8925 859 8932 870
rect 8907 856 8909 859
rect 8905 854 8907 855
rect 8898 851 8907 854
rect 8898 839 8905 851
rect 8898 838 8899 839
rect 8879 830 8898 838
rect 8912 830 8925 859
rect 8942 846 8949 858
rect 8954 848 8955 880
rect 9021 876 9027 879
rect 9018 874 9021 876
rect 9009 869 9018 874
rect 9029 870 9032 882
rect 9066 870 9069 884
rect 9126 881 9127 885
rect 9125 874 9126 881
rect 9166 874 9170 885
rect 9276 884 9278 885
rect 9277 883 9279 884
rect 9277 879 9280 883
rect 9326 880 9327 882
rect 9277 878 9281 879
rect 9280 876 9281 878
rect 9327 876 9328 880
rect 9378 876 9379 879
rect 9404 878 9420 906
rect 9124 871 9125 874
rect 9165 872 9166 874
rect 9002 860 9003 863
rect 9032 860 9034 870
rect 9066 862 9080 870
rect 9164 869 9165 871
rect 9281 869 9284 874
rect 9123 868 9124 869
rect 9122 864 9123 867
rect 9162 864 9164 868
rect 9161 862 9162 864
rect 9284 863 9286 869
rect 8997 848 9002 860
rect 8954 847 8959 848
rect 8954 846 8988 847
rect 8995 846 9000 848
rect 8949 844 8950 846
rect 8994 844 8995 846
rect 8991 842 8993 843
rect 8954 834 8966 841
rect 8976 834 8988 841
rect 9034 830 9045 859
rect 9069 830 9080 862
rect 9219 861 9220 862
rect 9121 856 9122 859
rect 9159 856 9161 861
rect 9286 860 9287 863
rect 9120 855 9121 856
rect 9098 851 9114 854
rect 9118 851 9120 854
rect 9157 851 9159 855
rect 9200 854 9212 855
rect 9098 843 9118 851
rect 9154 843 9157 851
rect 9194 849 9212 854
rect 9222 849 9234 855
rect 9194 843 9285 849
rect 9287 848 9291 860
rect 9291 844 9292 847
rect 9308 843 9324 854
rect 9096 839 9099 843
rect 9152 839 9154 843
rect 9188 842 9193 843
rect 9188 840 9192 842
rect 9194 841 9234 843
rect 9181 839 9191 840
rect 9194 839 9200 841
rect 9175 838 9180 839
rect 9194 838 9195 839
rect 9082 830 9096 838
rect 9149 836 9152 838
rect 9171 837 9175 838
rect 9162 836 9168 837
rect 9149 834 9162 836
rect 9139 833 9143 834
rect 9133 832 9139 833
rect 9149 832 9152 834
rect 9120 830 9133 832
rect 8661 827 8669 830
rect 8673 828 8676 830
rect 8660 821 8670 827
rect 8349 802 8350 804
rect 8351 800 8353 804
rect 8478 801 8488 816
rect 8490 812 8498 816
rect 8490 804 8499 812
rect 8503 807 8535 816
rect 8544 807 8556 820
rect 8636 807 8660 821
rect 8661 818 8669 821
rect 8499 801 8500 803
rect 8236 788 8252 796
rect 8272 795 8277 796
rect 8277 793 8288 795
rect 8295 794 8302 796
rect 8302 793 8308 794
rect 8319 793 8320 796
rect 8288 792 8293 793
rect 8308 792 8328 793
rect 8331 792 8333 795
rect 8348 794 8349 796
rect 8308 786 8329 792
rect 8345 789 8348 793
rect 8330 788 8348 789
rect 8330 786 8345 788
rect 8401 786 8402 788
rect 8406 786 8412 798
rect 8460 789 8461 797
rect 8475 790 8478 800
rect 8500 797 8509 801
rect 8512 800 8523 807
rect 8535 804 8556 807
rect 8510 797 8512 800
rect 8535 797 8554 804
rect 8624 800 8636 807
rect 8622 799 8624 800
rect 8506 796 8554 797
rect 8615 796 8622 799
rect 8661 796 8669 808
rect 8673 796 8675 828
rect 8741 822 8970 830
rect 8741 821 8742 822
rect 8744 820 8970 822
rect 8742 814 8970 820
rect 8998 814 9120 830
rect 9145 822 9149 831
rect 9178 822 9194 838
rect 9143 818 9145 822
rect 9142 817 9143 818
rect 9142 816 9148 817
rect 9141 815 9148 816
rect 8742 812 8998 814
rect 8743 804 8756 812
rect 8773 807 8775 812
rect 8743 803 8744 804
rect 8744 801 8745 802
rect 8742 798 8744 801
rect 8774 800 8775 807
rect 8786 804 8798 812
rect 8798 803 8799 804
rect 8803 803 8805 808
rect 8822 803 8901 812
rect 8799 802 8901 803
rect 8802 799 8818 802
rect 8741 796 8742 797
rect 8506 793 8544 796
rect 8554 795 8556 796
rect 8419 787 8420 788
rect 8418 786 8424 787
rect 8200 782 8206 786
rect 8317 784 8329 786
rect 5515 747 5521 750
rect 5569 749 5571 750
rect 5524 747 5528 749
rect 5515 746 5524 747
rect 5514 744 5522 746
rect 5533 745 5569 747
rect 5571 745 5579 747
rect 5036 738 5038 743
rect 5067 741 5099 743
rect 5095 740 5100 741
rect 5102 737 5105 739
rect 5155 738 5158 744
rect 5190 739 5193 744
rect 5273 740 5275 744
rect 5290 740 5302 742
rect 5003 734 5004 737
rect 5010 734 5014 737
rect 5002 732 5003 734
rect 5014 732 5018 734
rect 5034 732 5036 737
rect 5064 736 5065 737
rect 5094 734 5104 737
rect 5105 734 5111 737
rect 5117 734 5123 737
rect 5099 732 5104 734
rect 4999 725 5002 731
rect 5018 729 5022 732
rect 5032 729 5034 731
rect 4998 722 4999 724
rect 4994 711 4998 721
rect 5022 712 5050 729
rect 5063 726 5064 731
rect 5104 727 5108 732
rect 5110 731 5123 734
rect 5148 732 5152 734
rect 5146 731 5148 732
rect 5163 731 5169 737
rect 5253 734 5259 740
rect 5271 734 5272 736
rect 5290 734 5305 740
rect 5314 738 5315 742
rect 5463 738 5469 744
rect 5521 738 5527 744
rect 5533 743 5535 745
rect 5313 734 5314 737
rect 5186 732 5187 734
rect 5247 732 5311 734
rect 5108 726 5110 727
rect 5111 726 5117 731
rect 4865 710 4869 711
rect 4870 710 4922 711
rect 4864 706 4928 710
rect 4860 704 4928 706
rect 4991 704 4994 711
rect 4718 698 4724 699
rect 4732 698 4770 699
rect 4712 695 4724 698
rect 4728 695 4776 698
rect 4712 693 4718 695
rect 4728 693 4766 695
rect 4770 693 4776 695
rect 4860 694 4864 704
rect 4870 699 4888 704
rect 4870 698 4876 699
rect 4916 698 4922 704
rect 4989 699 4991 704
rect 4917 696 4918 698
rect 4987 695 4989 698
rect 5023 695 5031 712
rect 5051 709 5054 711
rect 5059 709 5063 726
rect 5110 717 5120 726
rect 5169 725 5175 731
rect 5182 725 5186 732
rect 5247 730 5305 732
rect 5306 730 5311 732
rect 5312 730 5313 732
rect 5247 728 5303 730
rect 5180 722 5181 724
rect 5120 709 5122 717
rect 5174 711 5180 721
rect 5054 708 5056 709
rect 5053 707 5057 708
rect 5053 703 5059 707
rect 5065 705 5066 707
rect 5065 703 5082 705
rect 5057 695 5059 703
rect 5062 699 5064 700
rect 5065 696 5089 699
rect 5122 698 5124 706
rect 5169 702 5174 711
rect 4984 694 4987 695
rect 4548 691 4557 692
rect 4563 691 4564 693
rect 4664 692 4776 693
rect 4664 691 4758 692
rect 4267 688 4270 689
rect 4274 688 4275 690
rect 4395 688 4399 690
rect 4557 689 4579 691
rect 4664 689 4754 691
rect 3888 682 3894 688
rect 3946 682 3952 688
rect 4270 686 4276 688
rect 3893 680 3906 682
rect 3893 676 3900 680
rect 3940 676 3946 682
rect 4274 677 4276 686
rect 4376 681 4395 688
rect 4376 679 4446 681
rect 3687 658 3697 669
rect 3689 656 3703 658
rect 3739 656 3755 672
rect 3893 669 3894 676
rect 4270 671 4276 677
rect 4328 678 4395 679
rect 4328 676 4392 678
rect 4446 676 4455 679
rect 4328 671 4334 676
rect 4273 669 4282 671
rect 3893 658 3903 668
rect 4273 658 4275 669
rect 4276 665 4282 669
rect 4322 665 4328 671
rect 4365 669 4376 676
rect 4455 675 4459 676
rect 4459 672 4461 675
rect 4563 671 4567 688
rect 4579 686 4614 689
rect 4664 686 4748 689
rect 4764 686 4770 692
rect 4859 690 4860 693
rect 4980 692 4984 694
rect 4978 691 4980 692
rect 4974 689 4978 691
rect 4970 688 4974 689
rect 5020 688 5023 695
rect 5056 690 5057 694
rect 5065 691 5077 696
rect 5089 693 5103 696
rect 5123 695 5124 698
rect 5253 696 5268 728
rect 5300 726 5303 728
rect 5306 726 5314 730
rect 5300 724 5302 726
rect 5301 700 5302 724
rect 5303 718 5314 726
rect 5303 714 5307 718
rect 5303 710 5306 714
rect 5309 712 5311 718
rect 5565 715 5567 745
rect 5569 742 5579 745
rect 5739 743 5741 749
rect 5749 743 5755 749
rect 5768 746 5791 770
rect 7253 755 7254 777
rect 7282 772 7283 777
rect 7373 774 7412 777
rect 7419 774 7431 777
rect 7283 759 7291 772
rect 7375 768 7412 774
rect 7422 768 7431 774
rect 7488 768 7489 777
rect 7283 755 7294 759
rect 7254 749 7255 755
rect 7291 753 7294 755
rect 7292 750 7297 753
rect 5795 743 5801 749
rect 7266 747 7295 748
rect 7298 747 7299 749
rect 5743 742 5749 743
rect 5571 738 5579 742
rect 5571 735 5589 738
rect 5579 731 5589 735
rect 5741 731 5749 742
rect 5754 738 5755 742
rect 5787 739 5793 742
rect 5752 731 5754 738
rect 5788 737 5793 739
rect 5801 737 5807 743
rect 5539 714 5567 715
rect 5534 713 5567 714
rect 5571 713 5579 725
rect 5589 721 5595 731
rect 5741 721 5752 731
rect 5733 720 5752 721
rect 5733 712 5742 720
rect 5308 710 5309 711
rect 5306 707 5309 710
rect 5568 709 5571 711
rect 5542 708 5545 709
rect 5305 702 5309 707
rect 5530 706 5540 708
rect 5521 704 5530 706
rect 5300 696 5302 699
rect 5306 696 5309 702
rect 5555 701 5567 709
rect 5746 707 5752 720
rect 5789 717 5793 737
rect 5745 706 5746 707
rect 5122 693 5123 694
rect 5103 692 5169 693
rect 5109 691 5169 692
rect 5115 690 5169 691
rect 4614 684 4633 686
rect 4672 684 4736 686
rect 4633 683 4641 684
rect 4641 681 4662 683
rect 4672 681 4731 684
rect 4662 679 4731 681
rect 4855 679 4859 688
rect 4918 686 4920 688
rect 4943 686 4970 688
rect 5019 686 5020 688
rect 4918 684 4950 686
rect 4908 683 4950 684
rect 4881 681 4950 683
rect 4863 679 4950 681
rect 5016 679 5019 684
rect 4672 678 4731 679
rect 4675 677 4710 678
rect 4836 677 4950 679
rect 4675 676 4707 677
rect 4709 676 4710 677
rect 4676 674 4688 676
rect 4690 675 4703 676
rect 4704 675 4709 676
rect 4814 675 4836 677
rect 4842 676 4950 677
rect 4855 675 4859 676
rect 4690 671 4717 675
rect 4766 671 4814 675
rect 5013 673 5016 679
rect 5053 672 5056 688
rect 5117 687 5169 690
rect 5253 688 5305 696
rect 5309 692 5310 694
rect 5463 693 5469 698
rect 5521 693 5527 698
rect 5742 697 5745 706
rect 5793 697 5795 717
rect 6556 703 6578 722
rect 7248 713 7255 725
rect 7260 716 7261 747
rect 7289 745 7294 747
rect 7293 716 7294 745
rect 7295 738 7306 747
rect 7522 740 7526 777
rect 7617 768 7626 777
rect 7669 768 7675 777
rect 7831 776 7855 777
rect 7991 772 7993 777
rect 8055 772 8083 777
rect 7984 759 7991 772
rect 8055 768 8064 772
rect 8102 768 8111 777
rect 8136 776 8142 782
rect 8194 776 8206 782
rect 8318 776 8319 781
rect 8194 766 8198 773
rect 8350 772 8351 786
rect 8402 783 8403 786
rect 8413 784 8415 785
rect 8459 784 8460 788
rect 8474 787 8475 790
rect 8500 789 8544 793
rect 8556 792 8563 795
rect 8613 793 8615 796
rect 8712 795 8740 796
rect 8563 789 8567 792
rect 8500 788 8522 789
rect 8524 788 8540 789
rect 8567 788 8569 789
rect 8609 788 8613 793
rect 8724 792 8740 795
rect 8770 793 8774 799
rect 8481 787 8488 788
rect 8496 787 8510 788
rect 8569 787 8572 788
rect 8473 786 8481 787
rect 8468 785 8481 786
rect 8500 785 8510 787
rect 8665 786 8671 792
rect 8723 791 8740 792
rect 8767 791 8770 793
rect 8723 789 8779 791
rect 8800 789 8818 799
rect 8723 788 8740 789
rect 8767 788 8770 789
rect 8779 788 8818 789
rect 8820 788 8901 802
rect 8912 800 8925 812
rect 8988 804 8989 807
rect 8723 786 8729 788
rect 8766 786 8767 788
rect 8465 784 8474 785
rect 8403 780 8415 783
rect 8418 780 8419 781
rect 8427 780 8465 784
rect 8403 779 8462 780
rect 8418 774 8430 779
rect 8349 763 8351 772
rect 8468 763 8474 784
rect 8500 784 8514 785
rect 7974 756 7991 759
rect 8315 756 8318 763
rect 7974 755 7984 756
rect 7974 754 7981 755
rect 8314 754 8315 756
rect 7974 753 7978 754
rect 7963 749 8005 753
rect 7963 748 7990 749
rect 8005 748 8006 749
rect 7961 747 7963 748
rect 8006 747 8008 748
rect 7947 745 7961 747
rect 7479 738 7485 740
rect 7522 739 7531 740
rect 7299 735 7317 738
rect 7306 725 7317 735
rect 7479 734 7491 738
rect 7525 734 7531 739
rect 7914 738 7947 745
rect 7908 737 7913 738
rect 7473 728 7479 734
rect 7531 729 7537 734
rect 7885 733 7908 737
rect 7962 735 7970 747
rect 7974 746 7979 747
rect 7879 731 7885 733
rect 7873 729 7875 731
rect 7495 728 7626 729
rect 7479 726 7495 728
rect 7531 727 7834 728
rect 7861 727 7867 729
rect 7872 728 7873 729
rect 7626 726 7627 727
rect 7834 726 7867 727
rect 7870 726 7872 728
rect 7260 714 7264 716
rect 7291 714 7294 716
rect 7260 713 7294 714
rect 7299 713 7317 725
rect 7467 714 7475 726
rect 7479 724 7485 726
rect 7255 711 7256 713
rect 7256 708 7261 711
rect 7294 708 7299 711
rect 7260 707 7272 708
rect 6527 697 6550 698
rect 6555 697 6578 703
rect 7259 701 7272 707
rect 7282 701 7294 708
rect 7306 707 7317 713
rect 7317 706 7322 707
rect 5742 694 5749 697
rect 5463 692 5527 693
rect 5116 685 5169 687
rect 5111 679 5175 685
rect 5247 682 5312 688
rect 5469 686 5475 692
rect 5515 686 5521 692
rect 5533 690 5534 694
rect 5741 690 5742 694
rect 5743 693 5749 694
rect 5801 693 5807 697
rect 7259 694 7261 701
rect 7317 694 7324 706
rect 5743 691 5807 693
rect 5740 688 5741 690
rect 5116 673 5123 679
rect 5163 673 5169 679
rect 5253 676 5259 682
rect 5299 676 5305 682
rect 4690 670 4728 671
rect 4755 670 4798 671
rect 4357 662 4365 669
rect 4463 667 4464 669
rect 4353 659 4357 662
rect 4464 660 4479 667
rect 4567 662 4569 669
rect 4690 664 4798 670
rect 5116 669 5121 673
rect 5256 672 5258 676
rect 5249 670 5258 672
rect 4692 662 4702 664
rect 4855 662 4856 669
rect 4569 660 4570 662
rect 4351 658 4353 659
rect 3903 656 3905 658
rect 4053 656 4055 657
rect 4273 656 4274 658
rect 4349 656 4351 658
rect 3705 640 3721 656
rect 3723 640 3739 656
rect 3906 653 3908 656
rect 4046 653 4052 656
rect 4275 653 4278 656
rect 4345 653 4349 656
rect 3908 651 3910 653
rect 4045 652 4046 653
rect 4343 652 4345 653
rect 4479 652 4591 660
rect 4683 658 4692 662
rect 4920 659 4923 669
rect 5052 666 5053 669
rect 4679 656 4683 658
rect 4856 656 4857 658
rect 4921 657 4923 659
rect 4919 656 4923 657
rect 4674 653 4679 656
rect 4857 653 4860 656
rect 4918 653 4919 656
rect 4953 654 4983 663
rect 4987 654 5000 660
rect 5052 659 5054 666
rect 5115 665 5123 669
rect 5113 658 5123 665
rect 5054 656 5055 658
rect 5112 656 5123 658
rect 5249 660 5256 670
rect 5311 669 5312 682
rect 5534 675 5535 688
rect 5527 669 5535 675
rect 5736 674 5740 686
rect 5749 685 5755 691
rect 5795 685 5801 691
rect 7322 690 7324 694
rect 7467 692 7475 704
rect 7479 694 7481 724
rect 7628 719 7632 726
rect 7834 723 7869 726
rect 7907 723 7913 729
rect 7632 708 7639 719
rect 7855 717 7861 723
rect 7862 719 7869 723
rect 7913 719 7919 723
rect 7962 719 7970 725
rect 7974 719 7976 746
rect 8303 744 8309 750
rect 8311 744 8314 754
rect 8349 750 8350 763
rect 8455 757 8461 762
rect 8467 757 8468 762
rect 8500 758 8510 784
rect 8514 783 8518 784
rect 8573 783 8579 786
rect 8608 783 8609 786
rect 8671 784 8685 786
rect 8671 783 8677 784
rect 8709 783 8713 784
rect 8580 781 8582 782
rect 8582 780 8585 781
rect 8598 780 8608 783
rect 8527 775 8533 779
rect 8533 772 8538 775
rect 8585 772 8608 780
rect 8539 766 8563 772
rect 8598 769 8630 772
rect 8636 769 8709 783
rect 8717 780 8723 786
rect 8724 784 8725 785
rect 8765 784 8766 786
rect 8800 783 8803 788
rect 8809 787 8901 788
rect 8873 786 8901 787
rect 8850 785 8901 786
rect 8909 785 8912 799
rect 8987 797 8988 801
rect 9034 800 9045 814
rect 9069 804 9080 814
rect 9082 804 9098 814
rect 9135 807 9148 815
rect 9132 805 9148 807
rect 9178 805 9194 820
rect 9232 811 9234 841
rect 9238 831 9246 843
rect 9285 838 9325 843
rect 9328 842 9335 874
rect 9370 840 9378 852
rect 9382 842 9384 874
rect 9414 869 9416 874
rect 9414 868 9417 869
rect 9414 842 9416 868
rect 9417 862 9418 864
rect 9418 857 9419 862
rect 9419 852 9420 855
rect 9382 840 9416 842
rect 9420 840 9428 852
rect 9335 838 9336 840
rect 9325 837 9340 838
rect 9382 837 9383 838
rect 9334 836 9340 837
rect 9379 836 9381 837
rect 9216 809 9234 811
rect 9238 809 9246 821
rect 9295 805 9305 836
rect 9334 832 9349 836
rect 9337 808 9349 832
rect 9382 828 9394 836
rect 9404 828 9416 836
rect 9422 834 9436 838
rect 9423 828 9436 834
rect 9383 824 9384 828
rect 9424 822 9436 828
rect 9384 820 9385 822
rect 9336 807 9349 808
rect 9121 804 9234 805
rect 9098 803 9234 804
rect 8986 791 8987 796
rect 8985 788 8986 791
rect 9045 789 9048 799
rect 9080 794 9088 800
rect 9098 795 9114 803
rect 9116 797 9234 803
rect 9305 801 9309 805
rect 9335 804 9349 807
rect 9370 815 9385 820
rect 9424 820 9425 822
rect 9424 816 9436 820
rect 9876 819 9877 1015
rect 10066 819 10067 1015
rect 10152 819 10153 1015
rect 10425 819 10426 1015
rect 10622 819 10623 1015
rect 10844 1013 10860 1015
rect 10866 1013 10878 1022
rect 10886 1020 10915 1023
rect 10915 1014 10919 1020
rect 11655 1018 11707 1020
rect 11927 1018 11941 1023
rect 12137 1020 12138 1023
rect 11627 1016 11707 1018
rect 11627 1015 11678 1016
rect 10919 1013 10920 1014
rect 11602 1013 11627 1015
rect 11649 1014 11655 1015
rect 11678 1014 11683 1015
rect 10840 1011 10844 1013
rect 10856 1010 10860 1013
rect 11568 1011 11598 1013
rect 11644 1012 11649 1014
rect 10832 998 10840 1010
rect 10839 988 10840 998
rect 10844 1007 10878 1010
rect 10844 1003 10846 1007
rect 10844 996 10845 1003
rect 10856 1001 10860 1007
rect 10875 1005 10878 1007
rect 10881 1004 10890 1010
rect 10843 994 10845 996
rect 10842 988 10848 994
rect 10853 988 10856 1001
rect 10836 982 10842 988
rect 10839 976 10840 982
rect 10843 962 10844 988
rect 10876 982 10878 1004
rect 10882 998 10890 1004
rect 10920 1001 10929 1010
rect 11451 1005 11465 1007
rect 11477 1005 11568 1011
rect 11640 1007 11644 1012
rect 11451 1004 11477 1005
rect 11451 1003 11465 1004
rect 11445 1002 11465 1003
rect 11486 1002 11491 1005
rect 11636 1002 11640 1007
rect 11683 1005 11700 1014
rect 11700 1004 11702 1005
rect 10888 988 10894 994
rect 10911 992 10920 1001
rect 11436 997 11460 1002
rect 11491 997 11497 1002
rect 11635 1001 11636 1002
rect 11707 1001 11724 1016
rect 11941 1015 11948 1018
rect 12136 1016 12137 1020
rect 11948 1014 11951 1015
rect 11951 1005 11973 1014
rect 12134 1012 12136 1016
rect 12174 1014 12178 1031
rect 12180 1027 12188 1039
rect 12446 1037 12458 1045
rect 12507 1041 12517 1045
rect 12518 1041 12524 1045
rect 12482 1037 12524 1041
rect 12576 1039 12582 1045
rect 12729 1044 12735 1050
rect 12775 1048 12785 1050
rect 14440 1048 14449 1057
rect 14505 1048 14514 1057
rect 15704 1048 15713 1057
rect 12738 1044 12750 1048
rect 12760 1044 12772 1048
rect 12775 1044 12781 1048
rect 12723 1038 12729 1044
rect 12781 1038 12787 1044
rect 15419 1038 15425 1044
rect 15465 1038 15471 1044
rect 15727 1043 15739 1051
rect 15749 1043 15761 1051
rect 15769 1048 15778 1057
rect 15828 1051 15844 1052
rect 15723 1040 15725 1043
rect 15763 1040 15765 1043
rect 15822 1039 15833 1051
rect 16096 1048 16105 1057
rect 16161 1051 16170 1057
rect 16102 1045 16105 1047
rect 16109 1045 16115 1051
rect 16155 1048 16170 1051
rect 16296 1048 16305 1057
rect 16361 1050 16370 1057
rect 16155 1045 16161 1048
rect 12227 1020 12237 1036
rect 12258 1034 12270 1037
rect 12452 1036 12458 1037
rect 12504 1036 12507 1037
rect 12252 1033 12272 1034
rect 12446 1033 12452 1036
rect 12488 1033 12518 1036
rect 12252 1031 12258 1033
rect 12272 1031 12302 1033
rect 12249 1025 12252 1031
rect 12246 1022 12252 1025
rect 12304 1024 12325 1031
rect 12352 1024 12358 1030
rect 11973 1004 11976 1005
rect 11833 1001 11834 1004
rect 11434 996 11436 997
rect 10894 982 10900 988
rect 10911 986 10915 992
rect 11423 989 11434 996
rect 11445 993 11460 997
rect 11497 996 11498 997
rect 10909 974 10910 979
rect 11067 976 11083 984
rect 11250 976 11266 989
rect 11333 979 11350 989
rect 11409 981 11423 989
rect 11403 979 11409 981
rect 11350 978 11403 979
rect 11434 977 11442 989
rect 11446 987 11451 989
rect 11498 987 11510 996
rect 11067 974 11124 976
rect 10905 957 10909 972
rect 11067 968 11112 974
rect 11124 968 11128 974
rect 10843 944 10850 957
rect 10904 953 10905 956
rect 10903 949 10904 952
rect 10906 944 10920 953
rect 11051 952 11067 968
rect 11128 961 11133 968
rect 11058 944 11067 952
rect 10836 936 10842 942
rect 10842 930 10848 936
rect 10850 934 10875 944
rect 10890 936 10906 944
rect 10888 934 10906 936
rect 11054 935 11058 944
rect 11061 940 11067 941
rect 11061 939 11103 940
rect 11107 939 11113 941
rect 11061 936 11072 939
rect 11061 935 11067 936
rect 11103 935 11113 939
rect 11054 934 11061 935
rect 10881 929 10884 934
rect 10888 930 10894 934
rect 10877 923 10880 928
rect 11051 925 11054 934
rect 11055 929 11061 934
rect 11113 929 11119 935
rect 11120 933 11132 941
rect 11193 934 11199 940
rect 11239 934 11245 940
rect 11250 934 11256 956
rect 11315 952 11321 958
rect 11361 952 11367 958
rect 11434 956 11442 967
rect 11446 958 11448 987
rect 11696 984 11698 1001
rect 11702 999 11724 1001
rect 11702 989 11710 999
rect 11828 992 11833 1001
rect 11976 996 11997 1004
rect 12131 1002 12134 1011
rect 12174 1007 12176 1014
rect 12165 1005 12176 1007
rect 12180 1010 12188 1017
rect 12180 1005 12193 1010
rect 12178 1004 12179 1005
rect 12184 1001 12193 1005
rect 12227 1002 12237 1018
rect 12246 1015 12249 1022
rect 12300 1018 12306 1024
rect 12358 1018 12364 1024
rect 12434 1021 12442 1033
rect 12446 1031 12480 1033
rect 12446 1030 12452 1031
rect 12446 1029 12449 1030
rect 12246 1014 12248 1015
rect 12246 1013 12250 1014
rect 12248 1001 12250 1013
rect 12130 996 12131 997
rect 11886 995 11919 996
rect 11997 995 11999 996
rect 11921 993 11927 995
rect 11828 986 11834 992
rect 11886 987 11892 992
rect 11927 991 11931 993
rect 11999 991 12009 995
rect 12129 991 12130 995
rect 12171 993 12184 1001
rect 12246 998 12250 1001
rect 12434 999 12442 1011
rect 12446 1002 12448 1029
rect 12726 1024 12729 1036
rect 12781 1032 12784 1036
rect 15413 1032 15419 1038
rect 15471 1032 15477 1038
rect 12734 1018 12738 1031
rect 12781 1021 12797 1032
rect 15704 1031 15710 1037
rect 15715 1031 15723 1039
rect 15726 1037 15761 1039
rect 15726 1036 15727 1037
rect 15725 1031 15726 1035
rect 15727 1031 15728 1036
rect 15759 1031 15761 1037
rect 14447 1026 14449 1030
rect 12797 1018 12813 1021
rect 12523 1007 12524 1008
rect 12524 1005 12525 1006
rect 12446 1001 12449 1002
rect 12492 1001 12520 1002
rect 12446 999 12458 1001
rect 12492 1000 12518 1001
rect 12176 992 12184 993
rect 12237 991 12241 996
rect 12246 991 12251 998
rect 12446 997 12447 999
rect 12492 998 12514 1000
rect 12520 999 12524 1001
rect 12447 996 12448 997
rect 12492 996 12507 998
rect 12448 995 12450 996
rect 12446 993 12452 995
rect 12492 994 12508 996
rect 12518 995 12524 999
rect 12527 997 12532 1003
rect 12576 1001 12585 1010
rect 12711 1001 12720 1010
rect 12720 1000 12726 1001
rect 11555 981 11571 984
rect 11573 981 11589 984
rect 11549 978 11569 981
rect 11690 979 11702 984
rect 11826 979 11827 983
rect 11834 980 11840 986
rect 11844 983 11912 987
rect 11931 986 11943 991
rect 11593 974 11594 978
rect 11551 972 11643 974
rect 11690 972 11710 979
rect 11825 974 11826 979
rect 11844 977 11870 983
rect 11880 980 11886 983
rect 11912 977 11925 983
rect 11943 978 11964 986
rect 12009 978 12043 991
rect 12175 988 12176 990
rect 12113 979 12119 985
rect 12129 983 12130 987
rect 12172 985 12175 986
rect 11824 972 11825 974
rect 11862 972 11870 977
rect 11455 963 11551 972
rect 11593 969 11594 972
rect 11552 963 11564 965
rect 11455 960 11552 963
rect 11446 957 11450 958
rect 11455 957 11551 960
rect 11446 956 11455 957
rect 11429 955 11453 956
rect 11457 955 11480 956
rect 11429 953 11448 955
rect 11497 954 11512 957
rect 11422 952 11429 953
rect 11442 952 11443 953
rect 11309 946 11315 952
rect 11367 946 11373 952
rect 11403 949 11422 952
rect 11490 951 11497 954
rect 11446 950 11457 951
rect 11488 950 11490 951
rect 11381 946 11403 949
rect 11373 945 11395 946
rect 11446 943 11458 950
rect 11509 944 11510 954
rect 11539 952 11549 957
rect 11548 944 11549 952
rect 11594 952 11605 968
rect 11594 951 11596 952
rect 11635 947 11636 968
rect 11643 965 11715 972
rect 11639 963 11715 965
rect 11643 956 11715 963
rect 11724 962 11725 968
rect 11718 956 11725 962
rect 11764 956 11770 962
rect 11819 956 11824 972
rect 11686 955 11727 956
rect 11712 950 11727 955
rect 11770 950 11776 956
rect 11566 942 11574 944
rect 11556 940 11566 942
rect 11554 939 11556 940
rect 11134 932 11136 933
rect 11107 927 11132 929
rect 11049 924 11051 925
rect 10872 914 10877 923
rect 10965 922 10995 924
rect 11045 922 11049 924
rect 10956 916 10965 922
rect 10995 916 11045 922
rect 10870 907 10872 914
rect 10838 895 10839 905
rect 10868 896 10870 907
rect 10941 906 10956 916
rect 11130 915 11132 927
rect 11136 917 11144 929
rect 11181 928 11193 934
rect 11245 928 11256 934
rect 11250 922 11256 928
rect 11367 926 11370 930
rect 11496 927 11554 939
rect 11596 938 11598 944
rect 11601 942 11647 944
rect 11647 940 11655 942
rect 11655 939 11658 940
rect 11566 930 11578 938
rect 11588 930 11600 938
rect 11491 926 11496 927
rect 11130 906 11133 915
rect 11169 910 11174 922
rect 11252 916 11259 922
rect 11259 914 11262 916
rect 11370 914 11384 926
rect 11477 923 11491 926
rect 11501 925 11509 927
rect 11598 926 11600 930
rect 11658 927 11705 939
rect 11718 935 11727 950
rect 11817 949 11819 956
rect 11835 952 11844 968
rect 11853 955 11862 972
rect 11925 968 11942 977
rect 11964 968 12003 978
rect 11816 946 11817 949
rect 11720 934 11722 935
rect 11770 933 11776 936
rect 11705 926 11710 927
rect 11718 926 11720 933
rect 11776 930 11783 933
rect 11793 930 11805 938
rect 11813 937 11815 942
rect 11835 937 11844 950
rect 11850 946 11853 955
rect 11895 954 11924 964
rect 11942 963 12003 968
rect 11942 957 11964 963
rect 12003 960 12013 963
rect 11888 945 11924 954
rect 11935 952 11944 954
rect 11847 937 11849 942
rect 11806 926 11813 937
rect 11835 934 11847 937
rect 11879 936 11888 945
rect 11895 944 11924 945
rect 11925 945 11944 952
rect 11964 950 11985 957
rect 12013 956 12023 960
rect 12043 956 12100 978
rect 12119 973 12125 979
rect 12130 977 12131 983
rect 12171 979 12177 985
rect 12131 972 12132 977
rect 12165 974 12171 979
rect 12172 974 12175 979
rect 12165 973 12172 974
rect 12171 972 12172 973
rect 12129 968 12132 972
rect 12180 971 12182 991
rect 12241 985 12247 991
rect 12252 988 12253 990
rect 12254 986 12257 987
rect 12257 985 12262 986
rect 12241 984 12297 985
rect 12446 984 12457 993
rect 12492 990 12504 994
rect 12518 993 12532 995
rect 12576 993 12582 999
rect 12720 998 12727 1000
rect 12729 998 12738 1018
rect 12813 1015 12826 1018
rect 13450 1015 13451 1026
rect 13640 1015 13641 1026
rect 13726 1015 13727 1026
rect 13999 1015 14000 1026
rect 14196 1015 14197 1026
rect 14432 1023 14471 1026
rect 15473 1023 15512 1028
rect 15698 1025 15704 1031
rect 15724 1026 15725 1031
rect 15723 1024 15724 1026
rect 14429 1022 14432 1023
rect 14429 1015 14441 1022
rect 14445 1016 14447 1022
rect 12826 1001 12890 1015
rect 12890 998 12900 1001
rect 12520 992 12530 993
rect 12567 992 12576 993
rect 12720 992 12738 998
rect 12781 992 12787 998
rect 12900 992 12945 998
rect 13040 994 13058 995
rect 13028 992 13040 994
rect 12492 986 12510 990
rect 12524 987 12530 992
rect 12570 987 12576 992
rect 12729 991 12735 992
rect 12729 989 12736 991
rect 12737 990 12738 992
rect 12767 991 12770 992
rect 12729 986 12735 989
rect 12737 987 12741 988
rect 12756 987 12767 991
rect 12772 986 12781 992
rect 12900 988 13028 992
rect 12241 983 12306 984
rect 12450 983 12458 984
rect 12258 981 12306 983
rect 12258 979 12270 981
rect 12452 978 12468 983
rect 12473 981 12474 984
rect 12300 972 12306 978
rect 12358 972 12364 978
rect 12129 967 12134 968
rect 12170 967 12171 971
rect 12120 958 12134 967
rect 12023 954 12028 956
rect 12100 955 12119 956
rect 12120 955 12132 958
rect 12028 951 12035 954
rect 12100 951 12132 955
rect 12134 951 12135 957
rect 12035 950 12037 951
rect 11925 944 11937 945
rect 11895 943 11902 944
rect 11944 943 11953 945
rect 11985 944 12023 950
rect 12038 949 12040 950
rect 12100 949 12120 951
rect 12123 949 12136 950
rect 12040 946 12049 949
rect 12113 948 12136 949
rect 12113 946 12120 948
rect 12123 945 12140 948
rect 12165 946 12170 967
rect 12182 951 12184 968
rect 12306 966 12312 972
rect 12315 967 12318 972
rect 12184 949 12189 950
rect 12123 944 12136 945
rect 11895 942 11900 943
rect 11895 941 11897 942
rect 11895 940 11941 941
rect 11942 940 11953 943
rect 11891 939 11896 940
rect 11903 939 11937 940
rect 11891 938 11937 939
rect 11891 937 11903 938
rect 11500 924 11501 925
rect 11468 921 11477 923
rect 11498 922 11500 924
rect 11456 920 11468 921
rect 11495 920 11498 922
rect 11426 916 11495 920
rect 11409 915 11426 916
rect 11397 914 11409 915
rect 11437 914 11456 916
rect 11554 914 11562 926
rect 11566 924 11600 926
rect 11262 913 11392 914
rect 11370 909 11384 913
rect 11426 911 11437 914
rect 11419 907 11425 911
rect 10937 900 10941 906
rect 11130 902 11132 906
rect 10867 891 10868 895
rect 10932 892 10937 899
rect 11115 898 11132 902
rect 11111 897 11132 898
rect 11107 896 11132 897
rect 11104 895 11132 896
rect 11136 895 11144 907
rect 11309 900 11315 906
rect 11119 891 11132 895
rect 11135 892 11136 894
rect 10866 888 10867 891
rect 10929 887 10932 891
rect 11106 889 11119 891
rect 10928 886 10929 887
rect 11055 886 11061 889
rect 11081 887 11119 889
rect 11081 886 11106 887
rect 10921 875 10928 885
rect 11020 875 11103 886
rect 11113 883 11119 887
rect 11120 883 11132 891
rect 11169 888 11174 900
rect 11315 894 11321 900
rect 11343 892 11356 900
rect 11386 892 11397 907
rect 11548 906 11553 913
rect 11411 900 11416 904
rect 11553 901 11557 906
rect 11557 899 11559 901
rect 11566 899 11568 924
rect 11343 889 11352 892
rect 11356 891 11358 892
rect 11398 889 11400 891
rect 11408 889 11417 898
rect 11559 892 11568 899
rect 11598 892 11600 924
rect 11604 914 11612 926
rect 11710 925 11720 926
rect 11710 923 11718 925
rect 11777 924 11805 926
rect 11716 922 11718 923
rect 11770 922 11771 924
rect 11803 922 11805 924
rect 11806 922 11817 926
rect 11715 921 11716 922
rect 11803 921 11817 922
rect 11636 916 11641 921
rect 11711 916 11715 921
rect 11769 917 11770 921
rect 11641 907 11650 916
rect 11705 907 11711 915
rect 11650 906 11705 907
rect 11712 904 11718 910
rect 11768 907 11769 916
rect 11803 915 11805 921
rect 11806 915 11817 921
rect 11840 925 11847 934
rect 11890 931 11903 937
rect 11934 936 11937 938
rect 11941 937 11953 940
rect 12023 937 12087 944
rect 11935 931 11937 936
rect 11948 931 11954 937
rect 12023 934 12119 937
rect 12123 934 12139 944
rect 12140 943 12150 945
rect 12182 944 12189 949
rect 12318 948 12325 967
rect 12352 966 12364 972
rect 12457 968 12468 978
rect 12492 980 12511 986
rect 12492 973 12529 980
rect 12653 976 12669 984
rect 12731 982 12734 986
rect 12730 976 12731 981
rect 12474 968 12477 972
rect 12358 945 12364 966
rect 12468 953 12480 968
rect 12496 965 12529 973
rect 12613 968 12616 976
rect 12654 975 12669 976
rect 12729 970 12730 975
rect 12772 969 12775 986
rect 12784 972 12885 977
rect 12885 969 12896 972
rect 12927 969 13028 988
rect 13058 980 13080 994
rect 12474 951 12477 953
rect 12480 951 12482 953
rect 12482 945 12495 951
rect 12511 948 12529 965
rect 12609 957 12613 968
rect 12604 955 12609 957
rect 12495 944 12497 945
rect 12567 944 12581 950
rect 12604 948 12616 955
rect 12603 947 12616 948
rect 12626 947 12638 955
rect 12669 952 12685 968
rect 12600 945 12609 947
rect 12177 943 12189 944
rect 12150 934 12214 943
rect 12497 942 12502 944
rect 12315 936 12397 942
rect 12298 934 12315 936
rect 11891 930 11903 931
rect 11840 924 11848 925
rect 11840 915 11847 924
rect 11848 922 11850 924
rect 11850 921 11852 922
rect 11851 918 11857 921
rect 11852 916 11857 918
rect 11803 911 11806 915
rect 11808 914 11817 915
rect 11808 912 11809 914
rect 11767 904 11768 906
rect 11770 904 11776 910
rect 11803 906 11805 911
rect 11809 907 11811 912
rect 11811 906 11812 907
rect 11802 904 11805 906
rect 11812 904 11813 906
rect 11718 898 11724 904
rect 11760 902 11763 904
rect 11764 902 11770 904
rect 11759 898 11770 902
rect 11801 901 11802 904
rect 11759 892 11766 898
rect 11800 897 11801 900
rect 11798 894 11800 895
rect 11803 894 11805 904
rect 11771 892 11805 894
rect 11809 899 11817 904
rect 11809 892 11823 899
rect 11798 891 11800 892
rect 11823 891 11824 892
rect 11824 890 11826 891
rect 10866 871 10867 875
rect 10919 871 10921 874
rect 10990 871 11020 875
rect 10918 870 10919 871
rect 10982 870 10990 871
rect 10980 869 10982 870
rect 10917 868 10918 869
rect 10978 868 10980 869
rect 11069 868 11071 875
rect 11104 868 11105 879
rect 11107 877 11113 883
rect 11187 882 11193 888
rect 11245 882 11251 888
rect 11181 876 11199 882
rect 11239 876 11245 882
rect 11352 880 11361 889
rect 11398 888 11408 889
rect 11796 888 11798 889
rect 11399 887 11408 888
rect 11399 880 11419 887
rect 11601 885 11602 888
rect 11562 882 11563 884
rect 11771 880 11783 888
rect 11793 882 11805 888
rect 11830 885 11840 915
rect 11857 912 11870 916
rect 11870 907 11882 912
rect 11885 906 11887 907
rect 11896 906 11903 930
rect 11948 928 11949 931
rect 12071 919 12119 934
rect 12139 932 12214 934
rect 12231 933 12282 934
rect 12284 933 12295 934
rect 12231 932 12292 933
rect 12139 930 12231 932
rect 11887 904 11892 906
rect 11896 904 11948 906
rect 11892 901 11948 904
rect 11896 899 11948 901
rect 11879 889 11888 898
rect 11896 896 11965 899
rect 11896 891 11953 896
rect 11965 892 11990 896
rect 12087 894 12095 919
rect 12119 916 12126 919
rect 12139 918 12155 930
rect 12157 918 12173 930
rect 12278 929 12293 932
rect 12274 927 12278 929
rect 12268 925 12274 927
rect 12284 926 12293 929
rect 12327 926 12334 936
rect 12264 924 12268 925
rect 12258 922 12264 924
rect 12287 920 12292 922
rect 12105 908 12107 916
rect 12126 914 12157 916
rect 12158 914 12160 918
rect 12126 909 12158 914
rect 12149 907 12166 909
rect 12107 900 12109 906
rect 12149 902 12158 907
rect 12166 906 12170 907
rect 12109 896 12110 899
rect 12129 898 12149 902
rect 11990 891 11996 892
rect 11890 889 11954 891
rect 11996 890 12002 891
rect 12086 890 12087 893
rect 12110 891 12111 896
rect 12124 891 12129 898
rect 12170 892 12227 906
rect 12227 891 12230 892
rect 11888 885 11954 889
rect 12002 887 12020 890
rect 12020 885 12032 887
rect 12085 885 12086 889
rect 12111 887 12112 891
rect 11826 884 11828 885
rect 11792 880 11805 882
rect 11362 875 11365 880
rect 11406 879 11419 880
rect 10904 864 10917 868
rect 10972 864 10978 868
rect 10898 862 10904 864
rect 10969 862 10972 864
rect 10894 856 10898 862
rect 10962 857 10969 862
rect 10961 856 10962 857
rect 10892 841 10894 855
rect 10958 849 10961 855
rect 10960 838 10969 842
rect 11007 838 11016 842
rect 11019 838 11035 854
rect 11037 838 11053 854
rect 11071 838 11075 867
rect 11102 847 11104 867
rect 10891 833 10892 838
rect 10958 833 10969 838
rect 11003 833 11019 838
rect 10951 832 10964 833
rect 11003 832 11025 833
rect 10890 825 10891 832
rect 10949 831 10958 832
rect 10889 819 10890 822
rect 9370 804 9386 815
rect 9425 805 9436 816
rect 9426 804 9436 805
rect 10888 812 10889 816
rect 10888 804 10892 812
rect 10949 811 10951 831
rect 10952 826 10958 831
rect 10957 822 10958 826
rect 10990 824 11025 832
rect 10990 822 11019 824
rect 11064 822 11069 838
rect 11102 833 11103 838
rect 11210 833 11222 864
rect 11365 860 11372 875
rect 11404 873 11419 875
rect 11244 833 11256 838
rect 11267 837 11279 845
rect 11333 838 11349 854
rect 11372 842 11381 860
rect 11373 841 11381 842
rect 11385 845 11386 862
rect 11385 843 11389 845
rect 11417 844 11419 873
rect 11420 871 11422 874
rect 11423 871 11431 875
rect 11422 869 11431 871
rect 11423 863 11431 869
rect 11427 862 11428 863
rect 11428 859 11430 862
rect 11563 860 11567 879
rect 11600 866 11601 880
rect 11682 867 11688 873
rect 11728 867 11734 873
rect 11792 870 11796 880
rect 11825 870 11830 884
rect 11888 880 11902 885
rect 11896 871 11902 880
rect 11938 880 11948 885
rect 11938 870 11939 880
rect 11942 879 11948 880
rect 12032 879 12069 885
rect 12084 881 12085 885
rect 12070 874 12075 879
rect 12075 872 12077 874
rect 12081 871 12084 881
rect 12112 879 12114 885
rect 12121 881 12123 889
rect 12230 888 12244 891
rect 12290 890 12292 920
rect 12296 910 12304 922
rect 12334 914 12339 926
rect 12339 902 12344 914
rect 12364 910 12371 936
rect 12397 934 12401 936
rect 12478 935 12479 942
rect 12502 936 12514 942
rect 12401 933 12402 934
rect 12402 927 12405 933
rect 12405 925 12406 927
rect 12406 922 12408 924
rect 12408 919 12410 922
rect 12410 916 12411 919
rect 12261 888 12292 890
rect 12296 888 12304 900
rect 12344 899 12345 902
rect 12371 900 12373 910
rect 12411 906 12416 916
rect 12479 910 12483 935
rect 12514 934 12518 936
rect 12529 935 12530 942
rect 12516 933 12522 934
rect 12516 932 12524 933
rect 12530 932 12531 935
rect 12566 934 12581 944
rect 12599 943 12600 945
rect 12603 943 12609 945
rect 12642 943 12643 945
rect 12649 943 12655 948
rect 12592 942 12599 943
rect 12603 942 12638 943
rect 12642 942 12655 943
rect 12592 937 12603 942
rect 12604 941 12638 942
rect 12590 934 12596 937
rect 12597 936 12603 937
rect 12637 936 12638 941
rect 12655 936 12661 942
rect 12669 934 12685 950
rect 12723 944 12729 968
rect 12775 956 12776 968
rect 12780 965 12781 969
rect 12896 968 12915 969
rect 12923 968 12927 969
rect 12887 964 12923 968
rect 12973 965 12977 969
rect 12721 934 12723 943
rect 12586 932 12590 934
rect 12524 931 12565 932
rect 12530 918 12547 931
rect 12549 926 12565 931
rect 12583 930 12586 932
rect 12576 926 12583 930
rect 12549 918 12576 926
rect 12668 925 12669 931
rect 12720 927 12721 932
rect 12667 920 12669 925
rect 12719 924 12720 925
rect 12730 922 12738 934
rect 12742 922 12744 956
rect 12780 951 12781 964
rect 12887 960 12935 964
rect 12878 954 12887 960
rect 12775 945 12776 951
rect 12873 945 12878 954
rect 12916 949 12935 960
rect 12935 948 12937 949
rect 12977 948 12982 965
rect 13080 961 13083 980
rect 13083 954 13084 960
rect 12937 945 12941 948
rect 12982 945 12983 948
rect 13084 945 13086 954
rect 12781 936 12782 945
rect 12867 936 12873 944
rect 12782 928 12788 934
rect 12862 928 12874 936
rect 12884 928 12896 936
rect 12941 934 12956 945
rect 12983 934 12987 945
rect 13086 941 13087 944
rect 13084 934 13087 941
rect 12956 932 12957 934
rect 12957 928 12958 930
rect 12987 929 12989 934
rect 12783 922 12788 928
rect 12863 926 12867 928
rect 12900 926 12901 928
rect 12862 924 12863 925
rect 12902 924 12905 925
rect 12666 919 12669 920
rect 12416 902 12418 906
rect 12530 905 12531 918
rect 12558 916 12576 918
rect 12665 918 12669 919
rect 12665 916 12666 918
rect 12718 916 12719 919
rect 12738 916 12739 921
rect 12771 916 12776 922
rect 12783 916 12784 922
rect 12552 912 12558 916
rect 12661 909 12665 916
rect 12717 909 12718 916
rect 12739 912 12741 916
rect 12769 913 12771 916
rect 12764 911 12769 913
rect 12780 911 12784 916
rect 12850 912 12858 924
rect 12862 922 12896 924
rect 12862 921 12865 922
rect 12742 910 12780 911
rect 12531 902 12532 904
rect 12418 899 12420 902
rect 12373 894 12374 899
rect 12420 896 12421 899
rect 12421 892 12423 896
rect 12244 885 12255 888
rect 12258 887 12262 888
rect 12262 885 12271 887
rect 12255 884 12261 885
rect 12114 875 12115 879
rect 12115 872 12116 874
rect 12118 871 12121 881
rect 12271 879 12297 885
rect 12346 881 12348 889
rect 12280 876 12292 879
rect 12297 874 12319 879
rect 12348 874 12349 881
rect 12333 872 12338 874
rect 12338 871 12340 872
rect 12374 871 12378 890
rect 12423 888 12425 891
rect 12529 890 12532 896
rect 12538 891 12549 908
rect 12604 906 12610 909
rect 12716 908 12717 909
rect 12655 906 12661 908
rect 12764 906 12769 910
rect 12610 903 12616 906
rect 12645 903 12655 906
rect 12715 903 12716 906
rect 12762 903 12764 906
rect 12616 902 12645 903
rect 12760 899 12762 903
rect 12714 896 12715 899
rect 12597 890 12603 896
rect 12655 890 12661 896
rect 12713 892 12714 896
rect 12757 891 12760 898
rect 12425 886 12426 887
rect 12527 885 12529 889
rect 12535 886 12538 890
rect 12426 874 12433 885
rect 12433 871 12434 874
rect 12480 871 12483 885
rect 12517 881 12527 885
rect 12603 884 12609 890
rect 12613 887 12614 890
rect 12623 886 12630 890
rect 12614 883 12617 885
rect 12620 884 12622 885
rect 12649 884 12655 890
rect 12712 888 12713 891
rect 12850 890 12858 902
rect 12862 890 12864 921
rect 12895 920 12896 922
rect 12902 912 12908 924
rect 12958 913 12960 925
rect 12989 916 13005 928
rect 13075 925 13084 934
rect 13067 924 13075 925
rect 13055 922 13067 924
rect 13018 916 13055 922
rect 12989 913 13018 916
rect 12902 911 12905 912
rect 12905 899 12910 910
rect 12950 906 13005 913
rect 12943 905 12950 906
rect 12937 903 12943 905
rect 12924 899 12937 903
rect 12899 891 12924 899
rect 12896 890 12899 891
rect 12756 887 12757 890
rect 12905 888 12910 891
rect 12960 889 12962 906
rect 12755 885 12756 887
rect 12858 886 12861 888
rect 12910 886 12911 888
rect 12962 885 12963 888
rect 12614 882 12619 883
rect 12515 874 12533 881
rect 12509 871 12515 874
rect 11767 868 11768 869
rect 11791 867 11792 870
rect 11676 861 11682 867
rect 11734 861 11740 867
rect 11789 860 11791 867
rect 11430 854 11436 858
rect 11430 853 11445 854
rect 11416 843 11419 844
rect 11385 841 11419 843
rect 11423 850 11445 853
rect 11567 852 11568 858
rect 11601 854 11602 858
rect 11423 841 11431 850
rect 11436 840 11445 850
rect 10990 820 11010 822
rect 11018 820 11038 822
rect 10948 810 10951 811
rect 10949 804 10951 810
rect 10957 804 10973 820
rect 11010 819 11018 820
rect 11029 816 11064 817
rect 11063 812 11064 816
rect 9334 803 9335 804
rect 9333 801 9334 802
rect 9281 799 9324 801
rect 9242 797 9281 799
rect 9116 796 9242 797
rect 9116 795 9222 796
rect 9305 795 9324 799
rect 9098 794 9132 795
rect 9080 792 9114 794
rect 9059 789 9088 792
rect 8974 785 8985 788
rect 9034 787 9059 789
rect 9021 786 9034 787
rect 9017 785 9021 786
rect 8876 784 8879 785
rect 8897 784 8985 785
rect 8897 783 8974 784
rect 8990 783 9017 785
rect 9045 784 9048 787
rect 8719 779 8720 780
rect 8757 769 8765 783
rect 8799 778 8800 783
rect 8875 781 8876 783
rect 8898 782 8900 783
rect 8874 778 8875 781
rect 8900 780 8903 782
rect 8908 781 8909 783
rect 8966 782 8970 783
rect 8974 782 8990 783
rect 8955 779 8966 782
rect 8903 778 8906 779
rect 8455 756 8473 757
rect 8501 756 8507 758
rect 8449 750 8513 756
rect 8538 753 8568 766
rect 8598 763 8636 769
rect 8754 763 8757 769
rect 8598 759 8630 763
rect 8597 756 8598 758
rect 8538 750 8574 753
rect 8595 752 8597 756
rect 8599 755 8630 759
rect 8627 754 8629 755
rect 8630 754 8633 755
rect 8749 754 8754 763
rect 8626 752 8627 754
rect 8633 751 8638 754
rect 8748 752 8749 754
rect 8349 744 8355 750
rect 8455 745 8507 750
rect 8259 742 8303 744
rect 8108 741 8142 742
rect 8259 741 8265 742
rect 8071 740 8108 741
rect 8048 739 8071 740
rect 8045 737 8048 739
rect 8297 738 8303 742
rect 8355 738 8361 744
rect 8020 723 8045 737
rect 8136 730 8142 736
rect 8194 731 8200 736
rect 8449 733 8461 745
rect 8495 735 8500 745
rect 8225 731 8261 733
rect 8142 724 8148 730
rect 8166 729 8225 731
rect 8261 729 8267 731
rect 8164 726 8166 729
rect 8015 720 8020 723
rect 7913 717 7995 719
rect 7916 716 7995 717
rect 8012 716 8020 720
rect 7962 713 7970 716
rect 7974 715 7976 716
rect 7995 715 8024 716
rect 7974 713 8008 715
rect 8005 709 8008 713
rect 8012 713 8020 715
rect 8024 714 8052 715
rect 8012 711 8015 713
rect 8009 709 8012 711
rect 8052 710 8066 714
rect 8158 713 8164 726
rect 8188 724 8194 729
rect 8267 726 8278 729
rect 8455 726 8461 733
rect 8257 722 8259 723
rect 8278 722 8289 726
rect 8454 723 8461 726
rect 8289 721 8291 722
rect 8291 720 8295 721
rect 7639 707 7640 708
rect 7861 707 7862 708
rect 7974 701 7986 709
rect 7996 701 8008 709
rect 8066 705 8072 710
rect 8156 708 8158 713
rect 8155 707 8156 708
rect 8072 703 8083 705
rect 7700 697 7834 700
rect 8000 698 8004 701
rect 8083 699 8096 703
rect 8096 698 8101 699
rect 7576 695 7700 697
rect 7834 695 7840 697
rect 7479 692 7485 694
rect 7554 692 7576 695
rect 7840 692 7846 695
rect 7992 694 8000 698
rect 8101 694 8117 698
rect 8149 694 8155 706
rect 7261 688 7262 690
rect 5795 674 5797 685
rect 5249 656 5255 660
rect 5311 656 5315 669
rect 5527 660 5536 669
rect 5527 658 5537 660
rect 5527 656 5538 658
rect 5595 656 5611 672
rect 5733 665 5742 674
rect 5798 669 5807 674
rect 7262 669 7272 688
rect 7324 674 7340 690
rect 7475 688 7477 691
rect 7531 689 7554 692
rect 7846 689 7852 692
rect 7984 690 7992 694
rect 8117 692 8133 694
rect 8249 693 8257 698
rect 8261 693 8263 720
rect 8449 711 8461 723
rect 8500 711 8502 726
rect 8538 723 8568 750
rect 8594 749 8595 751
rect 8638 750 8640 751
rect 8578 746 8580 747
rect 8592 745 8594 749
rect 8581 737 8595 745
rect 8623 744 8625 749
rect 8643 747 8646 749
rect 8646 746 8648 747
rect 8648 743 8652 746
rect 8672 743 8684 749
rect 8743 744 8746 749
rect 8778 744 8799 778
rect 8865 756 8874 778
rect 8903 776 8908 778
rect 8921 776 8955 779
rect 9048 778 9049 781
rect 8903 775 8921 776
rect 8903 756 8908 775
rect 9049 772 9053 778
rect 9049 756 9056 772
rect 9080 756 9088 789
rect 9098 788 9114 792
rect 9116 788 9132 794
rect 9194 788 9210 795
rect 9308 788 9324 795
rect 9311 787 9312 788
rect 9312 783 9313 785
rect 9314 772 9317 779
rect 9337 778 9349 804
rect 9386 797 9387 802
rect 9425 798 9426 800
rect 10892 799 10911 804
rect 10922 799 10957 804
rect 10892 797 10922 799
rect 9386 796 9388 797
rect 9424 796 9425 797
rect 9386 791 9394 796
rect 9421 791 9424 796
rect 9386 788 9402 791
rect 9404 788 9420 791
rect 10941 788 10958 799
rect 10949 786 10958 788
rect 10951 780 10958 786
rect 11016 783 11025 786
rect 11029 785 11031 788
rect 11061 785 11063 788
rect 11074 786 11075 828
rect 11102 820 11107 833
rect 11202 831 11279 833
rect 11099 804 11115 820
rect 11102 789 11107 804
rect 11115 789 11131 803
rect 11174 795 11193 798
rect 11087 787 11112 789
rect 11115 788 11140 789
rect 11087 785 11089 787
rect 11202 786 11260 831
rect 11277 801 11279 831
rect 11283 821 11291 833
rect 11349 822 11365 838
rect 11419 837 11423 840
rect 11443 838 11445 840
rect 11467 838 11473 844
rect 11513 839 11519 844
rect 11509 838 11521 839
rect 11568 838 11571 850
rect 11603 841 11619 854
rect 11674 852 11682 858
rect 11672 850 11682 852
rect 11786 851 11789 860
rect 11735 848 11745 850
rect 11745 846 11751 848
rect 11784 847 11786 851
rect 11662 844 11676 846
rect 11751 844 11758 846
rect 11602 840 11619 841
rect 11602 838 11606 840
rect 11385 829 11397 837
rect 11407 829 11419 837
rect 11445 832 11525 838
rect 11385 828 11386 829
rect 11274 799 11279 801
rect 11280 812 11283 819
rect 11386 818 11388 828
rect 11445 822 11461 832
rect 11467 827 11519 832
rect 11313 812 11349 816
rect 11388 814 11390 818
rect 11280 805 11349 812
rect 11390 809 11391 812
rect 11391 805 11392 809
rect 11029 783 11063 785
rect 11010 782 11038 783
rect 10995 780 11038 782
rect 8860 745 8865 756
rect 8900 744 8903 756
rect 9053 750 9056 756
rect 9053 744 9060 750
rect 9088 744 9090 756
rect 9118 751 9130 759
rect 9140 751 9152 759
rect 9317 755 9322 772
rect 9349 770 9353 778
rect 10951 777 10964 780
rect 11004 777 11010 780
rect 11016 777 11025 780
rect 11027 779 11038 780
rect 11193 780 11260 786
rect 11280 791 11341 805
rect 11349 791 11369 805
rect 11392 799 11393 803
rect 11393 795 11394 799
rect 11467 793 11487 827
rect 11527 815 11533 827
rect 11513 793 11521 795
rect 11527 793 11533 805
rect 11549 804 11557 820
rect 11572 814 11575 829
rect 11587 822 11606 838
rect 11640 833 11649 842
rect 11662 841 11682 844
rect 11758 843 11762 844
rect 11762 842 11767 843
rect 11783 842 11784 844
rect 11779 841 11790 842
rect 11815 841 11825 869
rect 11830 866 11831 868
rect 11831 856 11833 862
rect 11902 860 11907 870
rect 12078 868 12081 870
rect 12077 865 12081 868
rect 12078 860 12081 865
rect 12108 864 12118 870
rect 12340 869 12346 871
rect 12349 869 12355 870
rect 12346 868 12355 869
rect 12349 866 12355 868
rect 12349 864 12361 866
rect 12108 862 12119 864
rect 11833 854 11834 855
rect 11907 854 11908 860
rect 12077 858 12079 860
rect 12077 854 12078 858
rect 11833 852 11837 854
rect 11834 841 11837 852
rect 11899 849 11915 854
rect 11898 848 11912 849
rect 11917 848 11933 854
rect 11890 841 11898 848
rect 11912 842 11935 848
rect 11662 838 11676 841
rect 11782 839 11783 841
rect 11790 840 11825 841
rect 11836 840 11837 841
rect 11888 840 11890 841
rect 11815 839 11863 840
rect 11886 838 11888 840
rect 11902 839 11914 842
rect 11995 841 12011 854
rect 12013 841 12029 854
rect 12075 847 12077 853
rect 12079 852 12080 855
rect 11935 840 11936 841
rect 11988 840 11989 841
rect 11907 838 11914 839
rect 11656 834 11670 838
rect 11656 833 11667 834
rect 11631 824 11640 833
rect 11602 820 11606 822
rect 11587 814 11606 820
rect 11575 809 11576 812
rect 11576 799 11578 808
rect 11587 804 11603 814
rect 11662 812 11670 824
rect 11674 814 11676 838
rect 11779 832 11782 838
rect 11768 831 11782 832
rect 11768 822 11780 831
rect 11734 815 11740 821
rect 11775 818 11777 822
rect 11780 818 11786 822
rect 11774 815 11775 818
rect 11786 816 11788 818
rect 11728 814 11734 815
rect 11773 814 11774 815
rect 11674 812 11708 814
rect 11717 812 11776 814
rect 11788 813 11792 816
rect 11787 812 11793 813
rect 11606 808 11607 812
rect 11698 809 11708 812
rect 11712 810 11717 812
rect 11689 808 11698 809
rect 11701 808 11707 809
rect 11709 808 11712 810
rect 11728 809 11734 812
rect 11607 804 11608 808
rect 11674 805 11686 808
rect 11689 805 11708 808
rect 11674 804 11687 805
rect 11603 800 11608 804
rect 11665 800 11686 804
rect 11696 800 11708 805
rect 11764 800 11773 811
rect 11776 810 11784 812
rect 11787 810 11798 812
rect 11806 811 11815 838
rect 11837 822 11853 838
rect 11877 832 11885 838
rect 11784 809 11798 810
rect 11800 809 11806 810
rect 11784 808 11806 809
rect 11837 808 11853 820
rect 11906 811 11908 838
rect 11909 837 11914 838
rect 11911 836 11914 837
rect 11936 838 11937 840
rect 11987 838 11988 840
rect 12041 838 12044 841
rect 12073 839 12075 847
rect 12108 838 12118 862
rect 12119 855 12124 862
rect 12124 852 12126 855
rect 12126 848 12129 852
rect 12256 842 12262 844
rect 12256 838 12270 842
rect 12302 838 12308 844
rect 12309 838 12325 854
rect 12349 838 12355 864
rect 12361 863 12364 864
rect 12364 856 12366 862
rect 12366 853 12367 855
rect 12367 838 12372 852
rect 11912 834 11916 836
rect 11917 832 11918 834
rect 11910 828 11914 830
rect 11787 804 11853 808
rect 11796 800 11837 804
rect 11877 801 11878 804
rect 11603 797 11610 800
rect 11665 797 11685 800
rect 11603 794 11611 797
rect 11603 793 11613 794
rect 11394 792 11395 793
rect 11467 792 11519 793
rect 11525 792 11541 793
rect 11603 792 11615 793
rect 11280 784 11309 791
rect 11395 789 11401 792
rect 11401 784 11408 789
rect 11461 788 11541 792
rect 11579 790 11580 792
rect 11603 789 11624 792
rect 11603 788 11618 789
rect 11461 786 11525 788
rect 11613 786 11618 788
rect 11624 787 11629 789
rect 11629 786 11633 787
rect 11634 786 11665 797
rect 11697 793 11701 800
rect 11759 793 11764 799
rect 11696 790 11697 793
rect 11757 790 11759 793
rect 11408 783 11409 784
rect 11444 783 11445 785
rect 11193 777 11269 780
rect 11410 779 11416 783
rect 11441 779 11444 783
rect 11467 780 11473 786
rect 11509 781 11521 786
rect 11629 785 11640 786
rect 11631 783 11640 785
rect 11631 782 11643 783
rect 11513 780 11519 781
rect 11579 779 11580 781
rect 11416 777 11421 779
rect 11440 777 11441 779
rect 11578 777 11579 779
rect 11631 777 11640 782
rect 11646 779 11649 781
rect 11649 777 11668 779
rect 11696 777 11705 786
rect 11727 782 11733 788
rect 11754 786 11757 790
rect 11773 782 11779 788
rect 11791 786 11800 800
rect 11803 788 11819 800
rect 11821 796 11857 800
rect 11878 798 11879 801
rect 11905 800 11906 810
rect 11912 798 11914 828
rect 11918 818 11926 830
rect 11936 822 11949 838
rect 11979 836 11987 838
rect 12044 837 12045 838
rect 11979 823 11986 836
rect 12003 826 12015 832
rect 12000 825 12059 826
rect 12063 825 12073 838
rect 12000 823 12008 825
rect 12059 823 12073 825
rect 12080 824 12082 832
rect 11936 820 11938 822
rect 11999 821 12000 823
rect 11936 814 11949 820
rect 11880 797 11914 798
rect 11879 796 11914 797
rect 11918 796 11926 808
rect 11935 804 11949 814
rect 11991 816 11999 820
rect 12003 818 12010 820
rect 11991 808 11997 816
rect 12003 814 12004 818
rect 12063 816 12088 823
rect 12097 816 12108 837
rect 12129 822 12141 838
rect 12250 832 12256 838
rect 12266 832 12291 838
rect 12308 832 12314 838
rect 12325 832 12341 838
rect 12355 832 12356 838
rect 12372 832 12374 838
rect 12254 830 12256 832
rect 12258 830 12266 832
rect 12308 830 12341 832
rect 12374 830 12375 832
rect 12378 830 12390 870
rect 12434 869 12435 871
rect 12435 865 12437 868
rect 12437 863 12438 864
rect 12438 859 12440 862
rect 12464 838 12480 870
rect 12504 869 12509 871
rect 12517 870 12527 874
rect 12502 868 12504 869
rect 12498 866 12502 868
rect 12497 865 12498 866
rect 12496 863 12497 864
rect 12494 859 12496 862
rect 12510 859 12517 870
rect 12492 856 12494 859
rect 12490 854 12492 855
rect 12483 851 12492 854
rect 12483 839 12490 851
rect 12483 838 12484 839
rect 12464 830 12483 838
rect 12497 830 12510 859
rect 12527 846 12534 858
rect 12539 848 12540 880
rect 12606 876 12612 879
rect 12603 874 12606 876
rect 12594 869 12603 874
rect 12614 870 12617 882
rect 12651 870 12654 884
rect 12711 881 12712 885
rect 12710 874 12711 881
rect 12751 874 12755 885
rect 12861 884 12863 885
rect 12862 883 12864 884
rect 12862 879 12865 883
rect 12911 880 12912 882
rect 12862 878 12866 879
rect 12865 876 12866 878
rect 12912 876 12913 880
rect 12963 876 12964 879
rect 12989 878 13005 906
rect 12709 871 12710 874
rect 12750 872 12751 874
rect 12587 860 12588 863
rect 12617 860 12619 870
rect 12651 862 12665 870
rect 12749 869 12750 871
rect 12866 869 12869 874
rect 12708 868 12709 869
rect 12707 864 12708 867
rect 12747 864 12749 868
rect 12746 862 12747 864
rect 12869 863 12871 869
rect 12582 848 12587 860
rect 12539 847 12544 848
rect 12539 846 12573 847
rect 12580 846 12585 848
rect 12534 844 12535 846
rect 12579 844 12580 846
rect 12576 842 12578 843
rect 12539 834 12551 841
rect 12561 834 12573 841
rect 12619 830 12630 859
rect 12654 830 12665 862
rect 12804 861 12805 862
rect 12706 856 12707 859
rect 12744 856 12746 861
rect 12871 860 12872 863
rect 12705 855 12706 856
rect 12683 851 12699 854
rect 12703 851 12705 854
rect 12742 851 12744 855
rect 12785 854 12797 855
rect 12683 843 12703 851
rect 12739 843 12742 851
rect 12779 849 12797 854
rect 12807 849 12819 855
rect 12779 843 12870 849
rect 12872 848 12876 860
rect 12876 844 12877 847
rect 12893 843 12909 854
rect 12681 839 12684 843
rect 12737 839 12739 843
rect 12773 842 12778 843
rect 12773 840 12777 842
rect 12779 841 12819 843
rect 12766 839 12776 840
rect 12779 839 12785 841
rect 12760 838 12765 839
rect 12779 838 12780 839
rect 12667 830 12681 838
rect 12734 836 12737 838
rect 12756 837 12760 838
rect 12747 836 12753 837
rect 12734 834 12747 836
rect 12724 833 12728 834
rect 12718 832 12724 833
rect 12734 832 12737 834
rect 12705 830 12718 832
rect 12246 827 12254 830
rect 12258 828 12261 830
rect 12245 821 12255 827
rect 11934 802 11935 804
rect 11936 800 11938 804
rect 12063 801 12073 816
rect 12075 812 12083 816
rect 12075 804 12084 812
rect 12088 807 12120 816
rect 12129 807 12141 820
rect 12221 807 12245 821
rect 12246 818 12254 821
rect 12084 801 12085 803
rect 11821 788 11837 796
rect 11857 795 11862 796
rect 11862 793 11873 795
rect 11880 794 11887 796
rect 11887 793 11893 794
rect 11904 793 11905 796
rect 11873 792 11878 793
rect 11893 792 11913 793
rect 11916 792 11918 795
rect 11933 794 11934 796
rect 11893 786 11914 792
rect 11930 789 11933 793
rect 11915 788 11933 789
rect 11915 786 11930 788
rect 11986 786 11987 788
rect 11991 786 11997 798
rect 12045 789 12046 797
rect 12060 790 12063 800
rect 12085 797 12094 801
rect 12097 800 12108 807
rect 12120 804 12141 807
rect 12095 797 12097 800
rect 12120 797 12139 804
rect 12209 800 12221 807
rect 12207 799 12209 800
rect 12091 796 12139 797
rect 12200 796 12207 799
rect 12246 796 12254 808
rect 12258 796 12260 828
rect 12326 822 12555 830
rect 12326 821 12327 822
rect 12329 820 12555 822
rect 12327 814 12555 820
rect 12583 814 12705 830
rect 12730 822 12734 831
rect 12763 822 12779 838
rect 12728 818 12730 822
rect 12727 817 12728 818
rect 12727 816 12733 817
rect 12726 815 12733 816
rect 12327 812 12583 814
rect 12328 804 12341 812
rect 12358 807 12360 812
rect 12328 803 12329 804
rect 12329 801 12330 802
rect 12327 798 12329 801
rect 12359 800 12360 807
rect 12371 804 12383 812
rect 12383 803 12384 804
rect 12388 803 12390 808
rect 12407 803 12486 812
rect 12384 802 12486 803
rect 12387 799 12403 802
rect 12326 796 12327 797
rect 12091 793 12129 796
rect 12139 795 12141 796
rect 12004 787 12005 788
rect 12003 786 12009 787
rect 11785 782 11791 786
rect 11902 784 11914 786
rect 9100 747 9106 750
rect 9154 749 9156 750
rect 9109 747 9113 749
rect 9100 746 9109 747
rect 9099 744 9107 746
rect 9118 745 9154 747
rect 9156 745 9164 747
rect 8621 738 8623 743
rect 8652 741 8684 743
rect 8680 740 8685 741
rect 8687 737 8690 739
rect 8740 738 8743 744
rect 8775 739 8778 744
rect 8858 740 8860 744
rect 8875 740 8887 742
rect 8588 734 8589 737
rect 8595 734 8599 737
rect 8587 732 8588 734
rect 8599 732 8603 734
rect 8619 732 8621 737
rect 8649 736 8650 737
rect 8679 734 8689 737
rect 8690 734 8696 737
rect 8702 734 8708 737
rect 8684 732 8689 734
rect 8584 725 8587 731
rect 8603 729 8607 732
rect 8617 729 8619 731
rect 8583 722 8584 724
rect 8579 711 8583 721
rect 8607 712 8635 729
rect 8648 726 8649 731
rect 8689 727 8693 732
rect 8695 731 8708 734
rect 8733 732 8737 734
rect 8731 731 8733 732
rect 8748 731 8754 737
rect 8838 734 8844 740
rect 8856 734 8857 736
rect 8875 734 8890 740
rect 8899 738 8900 742
rect 9048 738 9054 744
rect 9106 738 9112 744
rect 9118 743 9120 745
rect 8898 734 8899 737
rect 8771 732 8772 734
rect 8832 732 8896 734
rect 8693 726 8695 727
rect 8696 726 8702 731
rect 8450 710 8454 711
rect 8455 710 8507 711
rect 8449 706 8513 710
rect 8445 704 8513 706
rect 8576 704 8579 711
rect 8303 698 8309 699
rect 8317 698 8355 699
rect 8297 695 8309 698
rect 8313 695 8361 698
rect 8297 693 8303 695
rect 8313 693 8351 695
rect 8355 693 8361 695
rect 8445 694 8449 704
rect 8455 699 8473 704
rect 8455 698 8461 699
rect 8501 698 8507 704
rect 8574 699 8576 704
rect 8502 696 8503 698
rect 8572 695 8574 698
rect 8608 695 8616 712
rect 8636 709 8639 711
rect 8644 709 8648 726
rect 8695 717 8705 726
rect 8754 725 8760 731
rect 8767 725 8771 732
rect 8832 730 8890 732
rect 8891 730 8896 732
rect 8897 730 8898 732
rect 8832 728 8888 730
rect 8765 722 8766 724
rect 8705 709 8707 717
rect 8759 711 8765 721
rect 8639 708 8641 709
rect 8638 707 8642 708
rect 8638 703 8644 707
rect 8650 705 8651 707
rect 8650 703 8667 705
rect 8642 695 8644 703
rect 8647 699 8649 700
rect 8650 696 8674 699
rect 8707 698 8709 706
rect 8754 702 8759 711
rect 8569 694 8572 695
rect 8133 691 8142 692
rect 8148 691 8149 693
rect 8249 692 8361 693
rect 8249 691 8343 692
rect 7852 688 7855 689
rect 7859 688 7860 690
rect 7980 688 7984 690
rect 8142 689 8164 691
rect 8249 689 8339 691
rect 7473 682 7479 688
rect 7531 682 7537 688
rect 7855 686 7861 688
rect 7478 680 7491 682
rect 7478 676 7485 680
rect 7525 676 7531 682
rect 7859 677 7861 686
rect 7961 681 7980 688
rect 7961 679 8031 681
rect 5797 667 5807 669
rect 5798 665 5807 667
rect 5735 656 5736 658
rect 5742 656 5751 665
rect 5789 656 5803 665
rect 7272 658 7282 669
rect 7274 656 7288 658
rect 7324 656 7340 672
rect 7478 669 7479 676
rect 7855 671 7861 677
rect 7913 678 7980 679
rect 7913 676 7977 678
rect 8031 676 8040 679
rect 7913 671 7919 676
rect 7858 669 7867 671
rect 7478 658 7488 668
rect 7858 658 7860 669
rect 7861 665 7867 669
rect 7907 665 7913 671
rect 7950 669 7961 676
rect 8040 675 8044 676
rect 8044 672 8046 675
rect 8148 671 8152 688
rect 8164 686 8199 689
rect 8249 686 8333 689
rect 8349 686 8355 692
rect 8444 690 8445 693
rect 8565 692 8569 694
rect 8563 691 8565 692
rect 8559 689 8563 691
rect 8555 688 8559 689
rect 8605 688 8608 695
rect 8641 690 8642 694
rect 8650 691 8662 696
rect 8674 693 8688 696
rect 8708 695 8709 698
rect 8838 696 8853 728
rect 8885 726 8888 728
rect 8891 726 8899 730
rect 8885 724 8887 726
rect 8886 700 8887 724
rect 8888 718 8899 726
rect 8888 714 8892 718
rect 8888 710 8891 714
rect 8894 712 8896 718
rect 9150 715 9152 745
rect 9154 742 9164 745
rect 9324 743 9326 749
rect 9334 743 9340 749
rect 9353 746 9376 770
rect 10838 755 10839 777
rect 10867 772 10868 777
rect 10958 774 10997 777
rect 11004 774 11016 777
rect 10868 759 10876 772
rect 10960 768 10997 774
rect 11007 768 11016 774
rect 11073 768 11074 777
rect 10868 755 10879 759
rect 10839 749 10840 755
rect 10876 753 10879 755
rect 10877 750 10882 753
rect 9380 743 9386 749
rect 10851 747 10880 748
rect 10883 747 10884 749
rect 9328 742 9334 743
rect 9156 738 9164 742
rect 9156 735 9174 738
rect 9164 731 9174 735
rect 9326 731 9334 742
rect 9339 738 9340 742
rect 9372 739 9378 742
rect 9337 731 9339 738
rect 9373 737 9378 739
rect 9386 737 9392 743
rect 9124 714 9152 715
rect 9119 713 9152 714
rect 9156 713 9164 725
rect 9174 721 9180 731
rect 9326 721 9337 731
rect 9318 720 9337 721
rect 9318 712 9327 720
rect 8893 710 8894 711
rect 8891 707 8894 710
rect 9153 709 9156 711
rect 9127 708 9130 709
rect 8890 702 8894 707
rect 9115 706 9125 708
rect 9106 704 9115 706
rect 8885 696 8887 699
rect 8891 696 8894 702
rect 9140 701 9152 709
rect 9331 707 9337 720
rect 9374 717 9378 737
rect 9330 706 9331 707
rect 8707 693 8708 694
rect 8688 692 8754 693
rect 8694 691 8754 692
rect 8700 690 8754 691
rect 8199 684 8218 686
rect 8257 684 8321 686
rect 8218 683 8226 684
rect 8226 681 8247 683
rect 8257 681 8316 684
rect 8247 679 8316 681
rect 8440 679 8444 688
rect 8503 686 8505 688
rect 8528 686 8555 688
rect 8604 686 8605 688
rect 8503 684 8535 686
rect 8493 683 8535 684
rect 8466 681 8535 683
rect 8448 679 8535 681
rect 8601 679 8604 684
rect 8257 678 8316 679
rect 8260 677 8295 678
rect 8421 677 8535 679
rect 8260 676 8292 677
rect 8294 676 8295 677
rect 8261 674 8273 676
rect 8275 675 8288 676
rect 8289 675 8294 676
rect 8399 675 8421 677
rect 8427 676 8535 677
rect 8440 675 8444 676
rect 8275 671 8302 675
rect 8351 671 8399 675
rect 8598 673 8601 679
rect 8638 672 8641 688
rect 8702 687 8754 690
rect 8838 688 8890 696
rect 8894 692 8895 694
rect 9048 693 9054 698
rect 9106 693 9112 698
rect 9327 697 9330 706
rect 9378 697 9380 717
rect 10141 703 10163 722
rect 10833 713 10840 725
rect 10845 716 10846 747
rect 10874 745 10879 747
rect 10878 716 10879 745
rect 10880 738 10891 747
rect 11107 740 11111 777
rect 11202 768 11211 777
rect 11254 768 11260 777
rect 11416 776 11440 777
rect 11576 772 11578 777
rect 11640 772 11668 777
rect 11569 759 11576 772
rect 11640 768 11649 772
rect 11687 768 11696 777
rect 11721 776 11727 782
rect 11779 776 11791 782
rect 11903 776 11904 781
rect 11779 766 11783 773
rect 11935 772 11936 786
rect 11987 783 11988 786
rect 11998 784 12000 785
rect 12044 784 12045 788
rect 12059 787 12060 790
rect 12085 789 12129 793
rect 12141 792 12148 795
rect 12198 793 12200 796
rect 12297 795 12325 796
rect 12148 789 12152 792
rect 12085 788 12107 789
rect 12109 788 12125 789
rect 12152 788 12154 789
rect 12194 788 12198 793
rect 12309 792 12325 795
rect 12355 793 12359 799
rect 12066 787 12073 788
rect 12081 787 12095 788
rect 12154 787 12157 788
rect 12058 786 12066 787
rect 12053 785 12066 786
rect 12085 785 12095 787
rect 12250 786 12256 792
rect 12308 791 12325 792
rect 12352 791 12355 793
rect 12308 789 12364 791
rect 12385 789 12403 799
rect 12308 788 12325 789
rect 12352 788 12355 789
rect 12364 788 12403 789
rect 12405 788 12486 802
rect 12497 800 12510 812
rect 12573 804 12574 807
rect 12308 786 12314 788
rect 12351 786 12352 788
rect 12050 784 12059 785
rect 11988 780 12000 783
rect 12003 780 12004 781
rect 12012 780 12050 784
rect 11988 779 12047 780
rect 12003 774 12015 779
rect 11934 763 11936 772
rect 12053 763 12059 784
rect 12085 784 12099 785
rect 11559 756 11576 759
rect 11900 756 11903 763
rect 11559 755 11569 756
rect 11559 754 11566 755
rect 11899 754 11900 756
rect 11559 753 11563 754
rect 11548 749 11590 753
rect 11548 748 11575 749
rect 11590 748 11591 749
rect 11546 747 11548 748
rect 11591 747 11593 748
rect 11532 745 11546 747
rect 11064 738 11070 740
rect 11107 739 11116 740
rect 10884 735 10902 738
rect 10891 725 10902 735
rect 11064 734 11076 738
rect 11110 734 11116 739
rect 11499 738 11532 745
rect 11493 737 11498 738
rect 11058 728 11064 734
rect 11116 729 11122 734
rect 11470 733 11493 737
rect 11547 735 11555 747
rect 11559 746 11564 747
rect 11464 731 11470 733
rect 11458 729 11460 731
rect 11080 728 11211 729
rect 11064 726 11080 728
rect 11116 727 11419 728
rect 11446 727 11452 729
rect 11457 728 11458 729
rect 11211 726 11212 727
rect 11419 726 11452 727
rect 11455 726 11457 728
rect 10845 714 10849 716
rect 10876 714 10879 716
rect 10845 713 10879 714
rect 10884 713 10902 725
rect 11052 714 11060 726
rect 11064 724 11070 726
rect 10840 711 10841 713
rect 10841 708 10846 711
rect 10879 708 10884 711
rect 10845 707 10857 708
rect 10112 697 10135 698
rect 10140 697 10163 703
rect 10844 701 10857 707
rect 10867 701 10879 708
rect 10891 707 10902 713
rect 10902 706 10907 707
rect 9327 694 9334 697
rect 9048 692 9112 693
rect 8701 685 8754 687
rect 8696 679 8760 685
rect 8832 682 8897 688
rect 9054 686 9060 692
rect 9100 686 9106 692
rect 9118 690 9119 694
rect 9326 690 9327 694
rect 9328 693 9334 694
rect 9386 693 9392 697
rect 10844 694 10846 701
rect 10902 694 10909 706
rect 9328 691 9392 693
rect 9325 688 9326 690
rect 8701 673 8708 679
rect 8748 673 8754 679
rect 8838 676 8844 682
rect 8884 676 8890 682
rect 8275 670 8313 671
rect 8340 670 8383 671
rect 7942 662 7950 669
rect 8048 667 8049 669
rect 7938 659 7942 662
rect 8049 660 8064 667
rect 8152 662 8154 669
rect 8275 664 8383 670
rect 8701 669 8706 673
rect 8841 672 8843 676
rect 8834 670 8843 672
rect 8277 662 8287 664
rect 8440 662 8441 669
rect 8154 660 8155 662
rect 7936 658 7938 659
rect 7488 656 7490 658
rect 7638 656 7640 657
rect 7858 656 7859 658
rect 7934 656 7936 658
rect 4669 652 4670 653
rect 4917 652 4918 653
rect 4950 652 4987 654
rect 5055 653 5056 656
rect 5111 653 5112 655
rect 5254 654 5255 656
rect 4043 651 4045 652
rect 3910 649 3986 651
rect 4038 649 4043 651
rect 4278 649 4282 652
rect 4341 650 4343 652
rect 4331 649 4341 650
rect 3993 648 4037 649
rect 4289 640 4305 649
rect 4306 648 4307 649
rect 4571 647 4573 651
rect 4591 647 4703 652
rect 4585 644 4703 647
rect 4801 644 4950 652
rect 4585 640 4601 644
rect 4703 641 4714 644
rect 4754 641 4801 644
rect 4714 640 4754 641
rect 4891 640 4907 644
rect 4953 636 4983 652
rect 5091 640 5107 653
rect 5254 644 5264 654
rect 5527 652 5540 656
rect 5562 652 5595 656
rect 5795 652 5798 656
rect 5542 651 5561 652
rect 5310 645 5311 651
rect 5265 640 5281 644
rect 5283 640 5299 644
rect 5579 640 5595 652
rect 5736 645 5746 652
rect 5790 646 5795 652
rect 5784 645 5790 646
rect 5746 644 5787 645
rect 5771 640 5787 644
rect 7290 640 7306 656
rect 7308 640 7324 656
rect 7491 653 7493 656
rect 7631 653 7637 656
rect 7860 653 7863 656
rect 7930 653 7934 656
rect 7493 651 7495 653
rect 7630 652 7631 653
rect 7928 652 7930 653
rect 8064 652 8176 660
rect 8268 658 8277 662
rect 8505 659 8508 669
rect 8637 666 8638 669
rect 8264 656 8268 658
rect 8441 656 8442 658
rect 8506 657 8508 659
rect 8504 656 8508 657
rect 8259 653 8264 656
rect 8442 653 8445 656
rect 8503 653 8504 656
rect 8538 654 8568 663
rect 8572 654 8585 660
rect 8637 659 8639 666
rect 8700 665 8708 669
rect 8698 658 8708 665
rect 8639 656 8640 658
rect 8697 656 8708 658
rect 8834 660 8841 670
rect 8896 669 8897 682
rect 9119 675 9120 688
rect 9112 669 9120 675
rect 9321 674 9325 686
rect 9334 685 9340 691
rect 9380 685 9386 691
rect 10907 690 10909 694
rect 11052 692 11060 704
rect 11064 694 11066 724
rect 11213 719 11217 726
rect 11419 723 11454 726
rect 11492 723 11498 729
rect 11217 708 11224 719
rect 11440 717 11446 723
rect 11447 719 11454 723
rect 11498 719 11504 723
rect 11547 719 11555 725
rect 11559 719 11561 746
rect 11888 744 11894 750
rect 11896 744 11899 754
rect 11934 750 11935 763
rect 12040 757 12046 762
rect 12052 757 12053 762
rect 12085 758 12095 784
rect 12099 783 12103 784
rect 12158 783 12164 786
rect 12193 783 12194 786
rect 12256 784 12270 786
rect 12256 783 12262 784
rect 12294 783 12298 784
rect 12165 781 12167 782
rect 12167 780 12170 781
rect 12183 780 12193 783
rect 12112 775 12118 779
rect 12118 772 12123 775
rect 12170 772 12193 780
rect 12124 766 12148 772
rect 12183 769 12215 772
rect 12221 769 12294 783
rect 12302 780 12308 786
rect 12309 784 12310 785
rect 12350 784 12351 786
rect 12385 783 12388 788
rect 12394 787 12486 788
rect 12458 786 12486 787
rect 12435 785 12486 786
rect 12494 785 12497 799
rect 12572 797 12573 801
rect 12619 800 12630 814
rect 12654 804 12665 814
rect 12667 804 12683 814
rect 12720 807 12733 815
rect 12717 805 12733 807
rect 12763 805 12779 820
rect 12817 811 12819 841
rect 12823 831 12831 843
rect 12870 838 12910 843
rect 12913 842 12920 874
rect 12955 840 12963 852
rect 12967 842 12969 874
rect 12999 869 13001 874
rect 12999 868 13002 869
rect 12999 842 13001 868
rect 13002 862 13003 864
rect 13003 857 13004 862
rect 13004 852 13005 855
rect 12967 840 13001 842
rect 13005 840 13013 852
rect 12920 838 12921 840
rect 12910 837 12925 838
rect 12967 837 12968 838
rect 12919 836 12925 837
rect 12964 836 12966 837
rect 12801 809 12819 811
rect 12823 809 12831 821
rect 12880 805 12890 836
rect 12919 832 12934 836
rect 12922 808 12934 832
rect 12967 828 12979 836
rect 12989 828 13001 836
rect 13007 834 13021 838
rect 13008 828 13021 834
rect 12968 824 12969 828
rect 13009 822 13021 828
rect 12969 820 12970 822
rect 12921 807 12934 808
rect 12706 804 12819 805
rect 12683 803 12819 804
rect 12571 791 12572 796
rect 12570 788 12571 791
rect 12630 789 12633 799
rect 12665 794 12673 800
rect 12683 795 12699 803
rect 12701 797 12819 803
rect 12890 801 12894 805
rect 12920 804 12934 807
rect 12955 815 12970 820
rect 13009 820 13010 822
rect 13009 816 13021 820
rect 13461 819 13462 1015
rect 13651 819 13652 1015
rect 13737 819 13738 1015
rect 14010 819 14011 1015
rect 14207 819 14208 1015
rect 14429 1013 14445 1015
rect 14451 1013 14463 1022
rect 14471 1020 14500 1023
rect 14500 1014 14504 1020
rect 15240 1018 15292 1020
rect 15512 1018 15526 1023
rect 15722 1020 15723 1023
rect 15212 1016 15292 1018
rect 15212 1015 15263 1016
rect 14504 1013 14505 1014
rect 15187 1013 15212 1015
rect 15234 1014 15240 1015
rect 15263 1014 15268 1015
rect 14425 1011 14429 1013
rect 14441 1010 14445 1013
rect 15153 1011 15183 1013
rect 15229 1012 15234 1014
rect 14417 998 14425 1010
rect 14424 988 14425 998
rect 14429 1007 14463 1010
rect 14429 1003 14431 1007
rect 14429 996 14430 1003
rect 14441 1001 14445 1007
rect 14460 1005 14463 1007
rect 14466 1004 14475 1010
rect 14428 994 14430 996
rect 14427 988 14433 994
rect 14438 988 14441 1001
rect 14421 982 14427 988
rect 14424 976 14425 982
rect 14428 962 14429 988
rect 14461 982 14463 1004
rect 14467 998 14475 1004
rect 14505 1001 14514 1010
rect 15036 1005 15050 1007
rect 15062 1005 15153 1011
rect 15225 1007 15229 1012
rect 15036 1004 15062 1005
rect 15036 1003 15050 1004
rect 15030 1002 15050 1003
rect 15071 1002 15076 1005
rect 15221 1002 15225 1007
rect 15268 1005 15285 1014
rect 15285 1004 15287 1005
rect 14473 988 14479 994
rect 14496 992 14505 1001
rect 15021 997 15045 1002
rect 15076 997 15082 1002
rect 15220 1001 15221 1002
rect 15292 1001 15309 1016
rect 15526 1015 15533 1018
rect 15721 1016 15722 1020
rect 15533 1014 15536 1015
rect 15536 1005 15558 1014
rect 15719 1012 15721 1016
rect 15759 1014 15763 1031
rect 15765 1027 15773 1039
rect 16031 1037 16043 1045
rect 16092 1041 16102 1045
rect 16103 1041 16109 1045
rect 16067 1037 16109 1041
rect 16161 1039 16167 1045
rect 16314 1044 16320 1050
rect 16360 1048 16370 1050
rect 18025 1048 18034 1057
rect 18090 1048 18099 1057
rect 19289 1048 19298 1057
rect 16323 1044 16335 1048
rect 16345 1044 16357 1048
rect 16360 1044 16366 1048
rect 16308 1038 16314 1044
rect 16366 1038 16372 1044
rect 19004 1038 19010 1044
rect 19050 1038 19056 1044
rect 19312 1043 19324 1051
rect 19334 1043 19346 1051
rect 19354 1048 19363 1057
rect 19413 1051 19429 1052
rect 19308 1040 19310 1043
rect 19348 1040 19350 1043
rect 19407 1039 19418 1051
rect 19681 1048 19690 1057
rect 19746 1051 19755 1057
rect 19687 1045 19690 1047
rect 19694 1045 19700 1051
rect 19740 1048 19755 1051
rect 19881 1048 19890 1057
rect 19946 1050 19955 1057
rect 19740 1045 19746 1048
rect 15812 1020 15822 1036
rect 15843 1034 15855 1037
rect 16037 1036 16043 1037
rect 16089 1036 16092 1037
rect 15837 1033 15857 1034
rect 16031 1033 16037 1036
rect 16073 1033 16103 1036
rect 15837 1031 15843 1033
rect 15857 1031 15887 1033
rect 15834 1025 15837 1031
rect 15831 1022 15837 1025
rect 15889 1024 15910 1031
rect 15937 1024 15943 1030
rect 15558 1004 15561 1005
rect 15418 1001 15419 1004
rect 14479 982 14485 988
rect 14496 986 14500 992
rect 15008 989 15021 997
rect 15030 993 15045 997
rect 14494 974 14495 979
rect 14652 976 14668 984
rect 14835 976 14851 989
rect 14918 979 14935 989
rect 14994 981 15008 989
rect 14988 979 14994 981
rect 14935 978 14988 979
rect 15019 977 15027 989
rect 15031 987 15036 989
rect 15082 987 15095 997
rect 14652 974 14709 976
rect 14490 957 14494 972
rect 14652 968 14697 974
rect 14709 968 14713 974
rect 14428 944 14435 957
rect 14489 953 14490 956
rect 14488 949 14489 952
rect 14491 944 14505 953
rect 14636 952 14652 968
rect 14713 961 14718 968
rect 14643 944 14652 952
rect 14421 936 14427 942
rect 14427 930 14433 936
rect 14435 934 14460 944
rect 14475 936 14491 944
rect 14473 934 14491 936
rect 14639 935 14643 944
rect 14646 940 14652 941
rect 14646 939 14688 940
rect 14692 939 14698 941
rect 14646 936 14657 939
rect 14646 935 14652 936
rect 14688 935 14698 939
rect 14639 934 14646 935
rect 14466 929 14469 934
rect 14473 930 14479 934
rect 14462 923 14465 928
rect 14636 925 14639 934
rect 14640 929 14646 934
rect 14698 929 14704 935
rect 14705 933 14717 941
rect 14778 934 14784 940
rect 14824 934 14830 940
rect 14835 934 14841 956
rect 14900 952 14906 958
rect 14946 952 14952 958
rect 15019 956 15027 967
rect 15031 958 15033 987
rect 15281 984 15283 1001
rect 15287 999 15309 1001
rect 15287 989 15295 999
rect 15413 992 15418 1001
rect 15561 996 15582 1004
rect 15716 1002 15719 1011
rect 15759 1007 15761 1014
rect 15750 1005 15761 1007
rect 15765 1010 15773 1017
rect 15765 1005 15778 1010
rect 15763 1004 15764 1005
rect 15769 1001 15778 1005
rect 15812 1002 15822 1018
rect 15831 1015 15834 1022
rect 15885 1018 15891 1024
rect 15943 1018 15949 1024
rect 16019 1021 16027 1033
rect 16031 1031 16065 1033
rect 16031 1030 16037 1031
rect 16031 1029 16034 1030
rect 15831 1014 15833 1015
rect 15831 1013 15835 1014
rect 15833 1001 15835 1013
rect 15471 995 15504 996
rect 15582 995 15584 996
rect 15506 993 15512 995
rect 15413 986 15419 992
rect 15471 987 15477 992
rect 15512 991 15516 993
rect 15584 991 15594 995
rect 15714 991 15716 997
rect 15756 993 15769 1001
rect 15831 998 15835 1001
rect 16019 999 16027 1011
rect 16031 1002 16033 1029
rect 16311 1024 16314 1036
rect 16366 1032 16369 1036
rect 18998 1032 19004 1038
rect 19056 1032 19062 1038
rect 16319 1018 16323 1031
rect 16366 1021 16382 1032
rect 19289 1031 19295 1037
rect 19300 1031 19308 1039
rect 19311 1037 19346 1039
rect 19311 1036 19312 1037
rect 19310 1031 19311 1035
rect 19312 1031 19313 1036
rect 19344 1031 19346 1037
rect 18032 1026 18034 1030
rect 16382 1018 16398 1021
rect 16108 1007 16109 1008
rect 16109 1005 16110 1006
rect 16031 1001 16034 1002
rect 16077 1001 16105 1002
rect 16031 999 16043 1001
rect 16077 1000 16103 1001
rect 15761 992 15769 993
rect 15822 991 15826 996
rect 15831 991 15836 998
rect 16031 997 16032 999
rect 16077 998 16099 1000
rect 16105 999 16109 1001
rect 16032 995 16035 997
rect 16077 996 16092 998
rect 16031 993 16037 995
rect 16077 994 16093 996
rect 16103 995 16109 999
rect 16112 997 16117 1003
rect 16161 1001 16170 1010
rect 16296 1001 16305 1010
rect 16305 1000 16311 1001
rect 15140 981 15156 984
rect 15158 981 15174 984
rect 15134 978 15154 981
rect 15275 979 15287 984
rect 15411 979 15412 983
rect 15419 980 15425 986
rect 15429 983 15497 987
rect 15516 986 15528 991
rect 15178 974 15179 978
rect 15136 972 15228 974
rect 15275 972 15295 979
rect 15410 974 15411 979
rect 15429 977 15455 983
rect 15465 980 15471 983
rect 15497 977 15510 983
rect 15528 978 15549 986
rect 15594 978 15628 991
rect 15760 988 15761 990
rect 15698 979 15704 985
rect 15714 983 15715 987
rect 15757 985 15760 986
rect 15409 972 15410 974
rect 15447 972 15455 977
rect 15040 963 15136 972
rect 15178 969 15179 972
rect 15137 963 15149 965
rect 15040 960 15137 963
rect 15031 957 15035 958
rect 15040 957 15136 960
rect 15031 956 15040 957
rect 15014 955 15038 956
rect 15042 955 15065 956
rect 15014 953 15033 955
rect 15082 954 15097 957
rect 15007 952 15014 953
rect 15027 952 15028 953
rect 14894 946 14900 952
rect 14952 946 14958 952
rect 14988 949 15007 952
rect 15075 951 15082 954
rect 15031 950 15042 951
rect 15073 950 15075 951
rect 14966 946 14988 949
rect 14958 945 14980 946
rect 15031 943 15043 950
rect 15094 939 15095 954
rect 15124 952 15134 957
rect 15133 939 15134 952
rect 15179 952 15190 968
rect 15151 942 15159 944
rect 15141 940 15151 942
rect 15139 939 15141 940
rect 14719 932 14721 933
rect 14692 927 14717 929
rect 14634 924 14636 925
rect 14457 914 14462 923
rect 14550 922 14580 924
rect 14630 922 14634 924
rect 14541 916 14550 922
rect 14580 916 14630 922
rect 14455 907 14457 914
rect 14423 895 14424 905
rect 14453 896 14455 907
rect 14526 906 14541 916
rect 14715 915 14717 927
rect 14721 917 14729 929
rect 14766 928 14778 934
rect 14830 928 14841 934
rect 14835 922 14841 928
rect 14952 926 14955 930
rect 15081 927 15139 939
rect 15179 938 15183 952
rect 15220 947 15221 968
rect 15228 965 15300 972
rect 15224 963 15300 965
rect 15228 956 15300 963
rect 15309 962 15310 968
rect 15303 956 15310 962
rect 15349 956 15355 962
rect 15404 956 15409 972
rect 15271 955 15312 956
rect 15297 950 15312 955
rect 15355 950 15361 956
rect 15186 942 15232 944
rect 15232 940 15240 942
rect 15240 939 15243 940
rect 15151 930 15163 938
rect 15173 930 15185 938
rect 15076 926 15081 927
rect 14715 906 14718 915
rect 14754 910 14759 922
rect 14837 916 14844 922
rect 14844 914 14847 916
rect 14955 914 14969 926
rect 15062 923 15076 926
rect 15085 924 15094 927
rect 15183 926 15185 930
rect 15243 927 15290 939
rect 15303 935 15312 950
rect 15402 949 15404 956
rect 15420 952 15429 968
rect 15438 955 15447 972
rect 15510 968 15527 977
rect 15549 968 15588 978
rect 15401 946 15402 949
rect 15305 934 15310 935
rect 15355 933 15361 936
rect 15290 926 15295 927
rect 15303 926 15305 933
rect 15361 930 15368 933
rect 15378 930 15390 938
rect 15398 937 15400 942
rect 15420 937 15429 950
rect 15435 946 15438 955
rect 15480 954 15509 964
rect 15527 963 15588 968
rect 15527 957 15549 963
rect 15588 960 15598 963
rect 15473 945 15509 954
rect 15520 952 15529 954
rect 15432 937 15434 942
rect 15391 926 15398 937
rect 15420 934 15432 937
rect 15464 936 15473 945
rect 15480 944 15509 945
rect 15510 945 15529 952
rect 15549 950 15570 957
rect 15598 956 15608 960
rect 15628 956 15685 978
rect 15704 973 15710 979
rect 15715 977 15716 983
rect 15756 979 15762 985
rect 15716 972 15717 977
rect 15750 974 15756 979
rect 15757 974 15760 979
rect 15750 973 15757 974
rect 15756 972 15757 973
rect 15714 968 15717 972
rect 15765 971 15767 991
rect 15826 985 15832 991
rect 15837 988 15838 990
rect 15839 986 15842 987
rect 15842 985 15847 986
rect 15826 984 15882 985
rect 16031 984 16042 993
rect 16077 990 16089 994
rect 16103 993 16117 995
rect 16161 993 16167 999
rect 16305 998 16312 1000
rect 16314 998 16323 1018
rect 16398 1015 16411 1018
rect 17035 1015 17036 1026
rect 17225 1015 17226 1026
rect 17311 1015 17312 1026
rect 17584 1015 17585 1026
rect 17781 1015 17782 1026
rect 18017 1023 18056 1026
rect 19058 1023 19097 1028
rect 19283 1025 19289 1031
rect 19309 1026 19310 1031
rect 19308 1024 19309 1026
rect 18014 1022 18017 1023
rect 18014 1015 18026 1022
rect 18030 1016 18032 1022
rect 16411 1001 16475 1015
rect 16475 998 16485 1001
rect 16105 992 16115 993
rect 16152 992 16161 993
rect 16305 992 16323 998
rect 16366 992 16372 998
rect 16485 992 16530 998
rect 16625 994 16643 995
rect 16613 992 16625 994
rect 16077 986 16095 990
rect 16109 987 16115 992
rect 16155 987 16161 992
rect 16314 991 16320 992
rect 16314 989 16321 991
rect 16322 990 16323 992
rect 16352 991 16355 992
rect 16314 986 16320 989
rect 16322 987 16326 988
rect 16341 987 16352 991
rect 16357 986 16366 992
rect 16485 988 16613 992
rect 15826 983 15891 984
rect 16035 983 16043 984
rect 15843 981 15891 983
rect 15843 979 15855 981
rect 16037 978 16053 983
rect 16058 981 16059 984
rect 15885 972 15891 978
rect 15943 972 15949 978
rect 15714 967 15719 968
rect 15755 967 15756 971
rect 15705 958 15719 967
rect 15608 954 15613 956
rect 15685 955 15704 956
rect 15705 955 15717 958
rect 15613 951 15620 954
rect 15685 951 15717 955
rect 15719 951 15720 957
rect 15620 950 15622 951
rect 15510 944 15522 945
rect 15480 943 15487 944
rect 15529 943 15538 945
rect 15480 942 15485 943
rect 15480 941 15482 942
rect 15480 940 15526 941
rect 15527 940 15538 943
rect 15476 939 15481 940
rect 15488 939 15522 940
rect 15476 938 15522 939
rect 15476 937 15488 938
rect 15425 926 15432 934
rect 15475 931 15488 937
rect 15519 936 15522 938
rect 15526 937 15538 940
rect 15570 937 15672 950
rect 15685 949 15705 951
rect 15708 949 15724 950
rect 15698 948 15724 949
rect 15698 946 15705 948
rect 15708 945 15725 948
rect 15750 946 15755 967
rect 15767 951 15769 968
rect 15891 966 15897 972
rect 15900 967 15903 972
rect 15769 949 15774 950
rect 15520 931 15522 936
rect 15533 931 15539 937
rect 15570 934 15704 937
rect 15708 934 15724 945
rect 15725 943 15735 945
rect 15762 943 15774 949
rect 15903 948 15910 967
rect 15937 966 15949 972
rect 16042 968 16053 978
rect 16077 980 16096 986
rect 16077 973 16114 980
rect 16238 976 16254 984
rect 16316 982 16319 986
rect 16315 976 16316 981
rect 16059 968 16062 972
rect 15943 945 15949 966
rect 16053 953 16065 968
rect 16081 965 16114 973
rect 16198 968 16201 976
rect 16239 975 16254 976
rect 16314 970 16315 975
rect 16357 969 16360 986
rect 16369 972 16470 977
rect 16470 969 16481 972
rect 16512 969 16613 988
rect 16643 980 16665 994
rect 16059 951 16062 953
rect 16065 951 16067 953
rect 15735 934 15799 943
rect 16067 942 16087 951
rect 16096 948 16114 965
rect 16194 957 16198 968
rect 16189 955 16194 957
rect 16151 950 16152 953
rect 15900 936 15982 942
rect 15883 934 15900 936
rect 15476 930 15488 931
rect 15053 921 15062 923
rect 15041 920 15053 921
rect 15080 920 15085 924
rect 14994 915 15080 920
rect 14982 914 14994 915
rect 15022 914 15041 915
rect 15139 914 15147 926
rect 15151 924 15185 926
rect 14847 913 14977 914
rect 14955 909 14969 913
rect 15011 911 15022 914
rect 15004 907 15010 911
rect 14522 900 14526 906
rect 14715 902 14717 906
rect 14452 891 14453 895
rect 14517 892 14522 899
rect 14700 898 14717 902
rect 14696 897 14717 898
rect 14692 896 14717 897
rect 14689 895 14717 896
rect 14721 895 14729 907
rect 14894 900 14900 906
rect 14704 891 14717 895
rect 14720 892 14721 894
rect 14451 888 14452 891
rect 14514 887 14517 891
rect 14691 889 14704 891
rect 14513 886 14514 887
rect 14640 886 14646 889
rect 14666 887 14704 889
rect 14666 886 14691 887
rect 14506 875 14513 885
rect 14605 875 14688 886
rect 14698 883 14704 887
rect 14705 883 14717 891
rect 14754 888 14759 900
rect 14900 894 14906 900
rect 14928 892 14941 900
rect 14971 892 14982 907
rect 14996 900 15001 904
rect 15133 901 15142 913
rect 15151 901 15153 924
rect 14928 889 14937 892
rect 14941 891 14943 892
rect 14983 889 14985 891
rect 14993 889 15002 898
rect 15142 892 15153 901
rect 15183 892 15185 924
rect 15189 914 15197 926
rect 15295 924 15305 926
rect 15362 924 15390 926
rect 15391 924 15402 926
rect 15295 923 15303 924
rect 15300 921 15303 923
rect 15355 921 15356 924
rect 15388 921 15402 924
rect 15221 907 15235 921
rect 15290 910 15300 921
rect 15354 917 15355 921
rect 15290 907 15303 910
rect 15353 907 15354 916
rect 15388 915 15390 921
rect 15391 915 15402 921
rect 15425 924 15433 926
rect 15425 915 15432 924
rect 15433 921 15437 924
rect 15436 918 15442 921
rect 15437 916 15442 918
rect 15388 911 15391 915
rect 15393 914 15402 915
rect 15393 912 15394 914
rect 15235 906 15290 907
rect 15297 904 15303 907
rect 15352 904 15353 906
rect 15355 904 15361 910
rect 15388 906 15390 911
rect 15394 907 15396 912
rect 15396 906 15397 907
rect 15387 904 15390 906
rect 15397 904 15398 906
rect 15303 898 15309 904
rect 15345 902 15348 904
rect 15349 902 15355 904
rect 15344 898 15355 902
rect 15386 901 15387 904
rect 15344 892 15351 898
rect 15385 897 15386 900
rect 15383 894 15385 895
rect 15388 894 15390 904
rect 15356 892 15390 894
rect 15394 901 15402 904
rect 15394 892 15408 901
rect 15383 891 15385 892
rect 15408 890 15411 892
rect 14451 871 14452 875
rect 14504 871 14506 874
rect 14575 871 14605 875
rect 14503 870 14504 871
rect 14567 870 14575 871
rect 14565 869 14567 870
rect 14502 868 14503 869
rect 14563 868 14565 869
rect 14654 868 14656 875
rect 14689 868 14690 879
rect 14692 877 14698 883
rect 14772 882 14778 888
rect 14830 882 14836 888
rect 14766 876 14784 882
rect 14824 876 14830 882
rect 14937 880 14946 889
rect 14983 888 14993 889
rect 15381 888 15383 889
rect 14984 887 14993 888
rect 14984 880 15004 887
rect 15186 885 15187 888
rect 15147 882 15148 884
rect 15356 880 15368 888
rect 15378 882 15390 888
rect 15411 884 15413 890
rect 15415 885 15425 915
rect 15442 912 15455 916
rect 15455 907 15467 912
rect 15470 906 15472 907
rect 15481 906 15488 930
rect 15533 928 15534 931
rect 15656 919 15704 934
rect 15724 932 15799 934
rect 15816 933 15867 934
rect 15869 933 15880 934
rect 15816 932 15877 933
rect 15724 930 15816 932
rect 15472 904 15477 906
rect 15481 904 15533 906
rect 15477 901 15533 904
rect 15481 899 15533 901
rect 15464 889 15473 898
rect 15481 896 15550 899
rect 15481 891 15538 896
rect 15550 892 15575 896
rect 15672 894 15680 919
rect 15704 916 15711 919
rect 15724 918 15740 930
rect 15742 918 15758 930
rect 15863 929 15878 932
rect 15859 927 15863 929
rect 15843 922 15859 927
rect 15869 926 15878 929
rect 15912 926 15919 936
rect 15872 920 15877 922
rect 15690 900 15694 916
rect 15711 914 15742 916
rect 15743 914 15745 918
rect 15711 909 15743 914
rect 15734 907 15751 909
rect 15734 902 15743 907
rect 15751 906 15755 907
rect 15694 896 15695 899
rect 15714 898 15734 902
rect 15475 889 15539 891
rect 15575 890 15587 892
rect 15671 890 15672 893
rect 15473 885 15539 889
rect 15377 880 15390 882
rect 14947 875 14950 880
rect 14991 879 15004 880
rect 14489 864 14502 868
rect 14557 864 14563 868
rect 14483 862 14489 864
rect 14554 862 14557 864
rect 14479 856 14483 862
rect 14547 857 14554 862
rect 14546 856 14547 857
rect 14477 841 14479 855
rect 14543 849 14546 855
rect 14545 838 14554 842
rect 14592 838 14601 842
rect 14604 838 14620 854
rect 14622 838 14638 854
rect 14656 838 14660 867
rect 14687 847 14689 867
rect 14476 833 14477 838
rect 14543 833 14554 838
rect 14588 833 14604 838
rect 14536 832 14549 833
rect 14588 832 14610 833
rect 14475 825 14476 832
rect 14534 831 14543 832
rect 14474 819 14475 822
rect 12955 804 12971 815
rect 13010 805 13021 816
rect 13011 804 13021 805
rect 14473 812 14474 816
rect 14473 804 14477 812
rect 14534 811 14536 831
rect 14537 826 14543 831
rect 14542 822 14543 826
rect 14575 824 14610 832
rect 14575 822 14604 824
rect 14649 822 14654 838
rect 14687 833 14688 838
rect 14795 833 14807 864
rect 14950 860 14957 875
rect 14989 873 15004 875
rect 14829 833 14841 838
rect 14852 837 14864 845
rect 14918 838 14934 854
rect 14957 842 14966 860
rect 14958 841 14966 842
rect 14970 845 14971 862
rect 14970 843 14974 845
rect 15002 844 15004 873
rect 15005 869 15016 875
rect 15008 863 15016 869
rect 15012 859 15015 863
rect 15148 860 15152 879
rect 15185 866 15186 880
rect 15267 867 15273 873
rect 15313 867 15319 873
rect 15377 870 15381 880
rect 15410 870 15415 884
rect 15473 880 15487 885
rect 15481 871 15487 880
rect 15523 880 15533 885
rect 15523 870 15524 880
rect 15527 879 15533 880
rect 15587 879 15654 890
rect 15670 885 15671 889
rect 15669 881 15670 885
rect 15655 875 15659 879
rect 15659 872 15662 875
rect 15666 871 15669 881
rect 15695 879 15699 896
rect 15709 891 15714 898
rect 15755 892 15812 906
rect 15812 891 15815 892
rect 15706 881 15708 889
rect 15815 888 15829 891
rect 15875 890 15877 920
rect 15881 910 15889 922
rect 15919 914 15924 926
rect 15924 902 15929 914
rect 15949 910 15956 936
rect 15982 934 15986 936
rect 16063 935 16064 942
rect 16087 936 16099 942
rect 15986 933 15987 934
rect 15987 927 15990 933
rect 15990 922 15993 927
rect 15993 919 15995 922
rect 15995 916 15996 919
rect 15846 888 15877 890
rect 15881 888 15889 900
rect 15929 899 15930 902
rect 15956 900 15958 910
rect 15996 902 16003 916
rect 16064 910 16068 935
rect 16099 934 16103 936
rect 16114 935 16115 942
rect 16101 933 16107 934
rect 16101 932 16109 933
rect 16115 932 16116 935
rect 16151 934 16166 950
rect 16189 948 16201 955
rect 16188 947 16201 948
rect 16211 947 16223 955
rect 16254 952 16270 968
rect 16185 945 16194 947
rect 16184 943 16185 945
rect 16188 943 16194 945
rect 16227 943 16228 945
rect 16234 943 16240 948
rect 16177 942 16184 943
rect 16188 942 16223 943
rect 16227 942 16240 943
rect 16177 937 16188 942
rect 16189 941 16223 942
rect 16175 934 16181 937
rect 16182 936 16188 937
rect 16222 936 16223 941
rect 16240 936 16246 942
rect 16254 934 16270 950
rect 16306 934 16314 968
rect 16360 956 16361 968
rect 16365 965 16366 969
rect 16481 968 16500 969
rect 16508 968 16512 969
rect 16472 964 16508 968
rect 16558 965 16562 969
rect 16171 932 16175 934
rect 16109 931 16150 932
rect 16115 918 16132 931
rect 16134 926 16150 931
rect 16168 930 16171 932
rect 16161 926 16168 930
rect 16253 927 16254 931
rect 16305 927 16306 932
rect 16134 918 16161 926
rect 16252 920 16254 927
rect 16304 922 16305 927
rect 16315 922 16323 934
rect 16327 922 16329 956
rect 16365 951 16366 964
rect 16472 960 16520 964
rect 16463 954 16472 960
rect 16360 945 16361 951
rect 16366 936 16367 945
rect 16452 936 16463 954
rect 16501 949 16520 960
rect 16520 948 16522 949
rect 16562 948 16567 965
rect 16665 961 16668 980
rect 16668 954 16669 960
rect 16522 945 16526 948
rect 16567 945 16568 948
rect 16447 934 16463 936
rect 16367 928 16373 934
rect 16368 922 16373 928
rect 16447 928 16459 934
rect 16469 928 16481 936
rect 16526 934 16541 945
rect 16568 934 16572 945
rect 16669 934 16672 954
rect 16541 932 16542 934
rect 16542 928 16543 930
rect 16572 929 16574 934
rect 16447 924 16452 928
rect 16485 926 16486 928
rect 16487 924 16490 925
rect 16251 919 16254 920
rect 16115 905 16116 918
rect 16143 916 16161 918
rect 16250 918 16254 919
rect 16250 916 16251 918
rect 16303 916 16304 919
rect 16323 916 16324 921
rect 16137 912 16143 916
rect 16246 909 16250 916
rect 16302 909 16303 916
rect 16324 912 16326 916
rect 16354 913 16361 922
rect 16368 916 16369 922
rect 16347 911 16354 913
rect 16365 911 16369 916
rect 16435 912 16443 924
rect 16447 922 16481 924
rect 16447 921 16450 922
rect 16327 910 16365 911
rect 16116 902 16117 904
rect 16003 899 16005 902
rect 15958 894 15959 899
rect 16005 896 16006 899
rect 15829 885 15840 888
rect 15843 885 15882 888
rect 15840 884 15882 885
rect 15699 872 15701 879
rect 15701 870 15702 872
rect 15703 871 15706 881
rect 15843 879 15882 884
rect 15931 881 15933 889
rect 15865 876 15877 879
rect 15882 874 15904 879
rect 15933 874 15934 881
rect 15918 872 15923 874
rect 15352 868 15353 869
rect 15376 867 15377 870
rect 15261 861 15267 867
rect 15319 861 15325 867
rect 15374 860 15376 867
rect 15015 854 15021 858
rect 15015 853 15030 854
rect 15001 843 15004 844
rect 14970 841 15004 843
rect 15008 850 15030 853
rect 15152 852 15153 858
rect 15186 854 15187 858
rect 15008 841 15016 850
rect 15021 840 15030 850
rect 14575 820 14595 822
rect 14603 820 14623 822
rect 14533 810 14536 811
rect 14534 804 14536 810
rect 14542 804 14558 820
rect 14595 819 14603 820
rect 14614 816 14649 817
rect 14648 812 14649 816
rect 12919 803 12920 804
rect 12918 801 12919 802
rect 12866 799 12909 801
rect 12827 797 12866 799
rect 12701 796 12827 797
rect 12701 795 12807 796
rect 12890 795 12909 799
rect 12683 794 12717 795
rect 12665 792 12699 794
rect 12644 789 12673 792
rect 12559 785 12570 788
rect 12619 787 12644 789
rect 12606 786 12619 787
rect 12602 785 12606 786
rect 12461 784 12464 785
rect 12482 784 12570 785
rect 12482 783 12559 784
rect 12575 783 12602 785
rect 12630 784 12633 787
rect 12304 779 12305 780
rect 12342 769 12350 783
rect 12384 778 12385 783
rect 12460 781 12461 783
rect 12483 782 12485 783
rect 12459 778 12460 781
rect 12485 780 12488 782
rect 12493 781 12494 783
rect 12551 782 12555 783
rect 12559 782 12575 783
rect 12540 779 12551 782
rect 12488 778 12491 779
rect 12040 756 12058 757
rect 12086 756 12092 758
rect 12034 750 12098 756
rect 12123 753 12153 766
rect 12183 763 12221 769
rect 12339 763 12342 769
rect 12183 759 12215 763
rect 12182 756 12183 758
rect 12123 750 12159 753
rect 12180 752 12182 756
rect 12184 755 12215 759
rect 12212 754 12214 755
rect 12215 754 12218 755
rect 12334 754 12339 763
rect 12211 752 12212 754
rect 12218 751 12223 754
rect 12333 752 12334 754
rect 11934 744 11940 750
rect 12040 745 12092 750
rect 11844 742 11888 744
rect 11693 741 11727 742
rect 11844 741 11850 742
rect 11656 740 11693 741
rect 11633 739 11656 740
rect 11630 737 11633 739
rect 11882 738 11888 742
rect 11940 738 11946 744
rect 11605 723 11630 737
rect 11721 730 11727 736
rect 11779 731 11785 736
rect 12034 733 12046 745
rect 12080 735 12085 745
rect 11810 731 11846 733
rect 11727 724 11733 730
rect 11751 729 11810 731
rect 11846 729 11852 731
rect 11749 726 11751 729
rect 11600 720 11605 723
rect 11498 717 11580 719
rect 11501 716 11580 717
rect 11597 716 11605 720
rect 11547 713 11555 716
rect 11559 715 11561 716
rect 11580 715 11609 716
rect 11559 713 11593 715
rect 11590 709 11593 713
rect 11597 713 11605 715
rect 11609 714 11637 715
rect 11597 711 11600 713
rect 11594 709 11597 711
rect 11637 710 11651 714
rect 11743 713 11749 726
rect 11773 724 11779 729
rect 11852 726 11863 729
rect 12040 726 12046 733
rect 11842 722 11844 723
rect 11863 722 11874 726
rect 12039 723 12046 726
rect 11874 721 11876 722
rect 11876 720 11880 721
rect 11224 707 11225 708
rect 11446 707 11447 708
rect 11559 701 11571 709
rect 11581 701 11593 709
rect 11651 705 11657 710
rect 11741 708 11743 713
rect 11740 707 11741 708
rect 11657 703 11668 705
rect 11285 697 11419 700
rect 11585 698 11589 701
rect 11668 699 11681 703
rect 11681 698 11686 699
rect 11161 695 11285 697
rect 11419 695 11425 697
rect 11064 692 11070 694
rect 11139 692 11161 695
rect 11425 692 11431 695
rect 11577 694 11585 698
rect 11686 694 11702 698
rect 11734 694 11740 706
rect 10846 688 10847 690
rect 9380 674 9382 685
rect 8834 656 8840 660
rect 8896 656 8900 669
rect 9112 660 9121 669
rect 9112 658 9122 660
rect 9112 656 9123 658
rect 9180 656 9196 672
rect 9318 665 9327 674
rect 9383 669 9392 674
rect 10847 669 10857 688
rect 10909 674 10925 690
rect 11060 688 11062 691
rect 11116 689 11139 692
rect 11431 689 11437 692
rect 11569 690 11577 694
rect 11702 692 11718 694
rect 11834 693 11842 698
rect 11846 693 11848 720
rect 12034 711 12046 723
rect 12085 711 12087 726
rect 12123 723 12153 750
rect 12179 749 12180 751
rect 12223 750 12225 751
rect 12163 746 12165 747
rect 12177 745 12179 749
rect 12166 737 12180 745
rect 12208 744 12210 749
rect 12228 747 12231 749
rect 12231 746 12233 747
rect 12233 743 12237 746
rect 12257 743 12269 749
rect 12328 744 12331 749
rect 12363 744 12384 778
rect 12450 756 12459 778
rect 12488 776 12493 778
rect 12506 776 12540 779
rect 12633 778 12634 781
rect 12488 775 12506 776
rect 12488 756 12493 775
rect 12634 772 12638 778
rect 12634 756 12641 772
rect 12665 756 12673 789
rect 12683 788 12699 792
rect 12701 788 12717 794
rect 12779 788 12795 795
rect 12893 788 12909 795
rect 12896 787 12897 788
rect 12897 783 12898 785
rect 12899 772 12902 779
rect 12922 778 12934 804
rect 12971 797 12972 802
rect 13010 798 13011 800
rect 14477 799 14496 804
rect 14507 799 14542 804
rect 14477 797 14507 799
rect 12971 796 12973 797
rect 13009 796 13010 797
rect 12971 791 12979 796
rect 13006 791 13009 796
rect 12971 788 12987 791
rect 12989 788 13005 791
rect 14526 788 14543 799
rect 14534 786 14543 788
rect 14536 780 14543 786
rect 14601 783 14610 786
rect 14614 785 14616 788
rect 14646 785 14648 788
rect 14659 786 14660 828
rect 14687 820 14692 833
rect 14787 831 14864 833
rect 14684 804 14700 820
rect 14687 789 14692 804
rect 14700 789 14716 803
rect 14759 795 14778 798
rect 14672 787 14697 789
rect 14700 788 14725 789
rect 14672 785 14674 787
rect 14787 786 14845 831
rect 14862 801 14864 831
rect 14868 821 14876 833
rect 14934 822 14950 838
rect 15004 837 15008 840
rect 15028 838 15030 840
rect 15052 838 15058 844
rect 15098 839 15104 844
rect 15094 838 15106 839
rect 15153 838 15156 850
rect 15188 841 15204 854
rect 15259 852 15267 858
rect 15257 850 15267 852
rect 15371 851 15374 860
rect 15320 848 15330 850
rect 15330 846 15336 848
rect 15369 847 15371 851
rect 15247 844 15261 846
rect 15336 844 15343 846
rect 15187 840 15204 841
rect 15187 838 15191 840
rect 14970 829 14982 837
rect 14992 829 15004 837
rect 15030 832 15110 838
rect 14970 828 14971 829
rect 14859 799 14864 801
rect 14865 812 14868 819
rect 14971 818 14973 828
rect 15030 822 15046 832
rect 15052 827 15104 832
rect 14898 812 14934 816
rect 14973 814 14975 818
rect 14865 805 14934 812
rect 14975 809 14976 812
rect 14976 805 14977 809
rect 14614 783 14648 785
rect 14595 782 14623 783
rect 14580 780 14623 782
rect 12445 745 12450 756
rect 12485 744 12488 756
rect 12638 750 12641 756
rect 12638 744 12645 750
rect 12673 744 12675 756
rect 12703 751 12715 759
rect 12725 751 12737 759
rect 12902 755 12907 772
rect 12934 770 12938 778
rect 14536 777 14549 780
rect 14589 777 14595 780
rect 14601 777 14610 780
rect 14612 779 14623 780
rect 14778 780 14845 786
rect 14865 791 14926 805
rect 14934 791 14954 805
rect 14977 799 14978 803
rect 14978 795 14979 799
rect 15052 793 15072 827
rect 15112 815 15118 827
rect 15098 793 15106 795
rect 15112 793 15118 805
rect 15134 804 15142 820
rect 15157 814 15160 829
rect 15172 822 15191 838
rect 15225 833 15234 842
rect 15247 841 15267 844
rect 15343 843 15347 844
rect 15347 842 15352 843
rect 15368 842 15369 844
rect 15364 841 15375 842
rect 15400 841 15410 869
rect 15415 866 15416 869
rect 15416 854 15419 865
rect 15487 860 15492 870
rect 15663 869 15666 870
rect 15662 865 15666 869
rect 15663 860 15666 865
rect 15693 866 15703 870
rect 15923 866 15940 872
rect 15959 871 15963 890
rect 16006 888 16010 896
rect 16114 890 16117 896
rect 16123 891 16134 908
rect 16189 903 16201 909
rect 16301 908 16302 909
rect 16230 903 16246 908
rect 16300 903 16301 908
rect 16347 903 16354 910
rect 16201 902 16230 903
rect 16299 896 16300 899
rect 16182 890 16188 896
rect 16240 890 16246 896
rect 16010 874 16018 888
rect 16112 885 16114 889
rect 16120 886 16123 890
rect 15492 854 15493 860
rect 15662 854 15665 860
rect 15416 852 15422 854
rect 15419 841 15422 852
rect 15484 849 15500 854
rect 15483 848 15497 849
rect 15502 848 15518 854
rect 15475 841 15483 848
rect 15497 842 15520 848
rect 15247 838 15261 841
rect 15367 839 15368 841
rect 15375 840 15410 841
rect 15421 840 15422 841
rect 15473 840 15475 841
rect 15400 839 15448 840
rect 15471 838 15473 840
rect 15487 839 15499 842
rect 15580 841 15596 854
rect 15598 841 15614 854
rect 15660 847 15662 853
rect 15663 852 15665 854
rect 15693 852 15711 866
rect 15934 863 15949 866
rect 15520 840 15521 841
rect 15573 840 15574 841
rect 15492 838 15499 839
rect 15241 834 15255 838
rect 15241 833 15252 834
rect 15216 824 15225 833
rect 15187 820 15191 822
rect 15172 814 15191 820
rect 15160 809 15161 812
rect 15161 799 15163 808
rect 15172 804 15188 814
rect 15247 812 15255 824
rect 15259 814 15261 838
rect 15364 832 15367 838
rect 15319 815 15325 821
rect 15353 818 15371 832
rect 15359 815 15360 818
rect 15313 814 15319 815
rect 15358 814 15359 815
rect 15259 812 15293 814
rect 15302 812 15361 814
rect 15371 813 15377 818
rect 15372 812 15378 813
rect 15191 808 15192 812
rect 15283 809 15293 812
rect 15297 810 15302 812
rect 15274 808 15283 809
rect 15286 808 15292 809
rect 15294 808 15297 810
rect 15313 809 15319 812
rect 15192 804 15193 808
rect 15259 805 15271 808
rect 15274 805 15293 808
rect 15259 804 15272 805
rect 15188 794 15196 804
rect 15219 800 15271 804
rect 15281 800 15293 805
rect 15349 800 15358 811
rect 15361 810 15369 812
rect 15372 810 15383 812
rect 15391 811 15400 838
rect 15422 822 15438 838
rect 15462 832 15470 838
rect 15369 809 15383 810
rect 15385 809 15391 810
rect 15369 808 15391 809
rect 15422 808 15438 820
rect 15491 811 15493 838
rect 15494 837 15499 838
rect 15496 836 15499 837
rect 15521 838 15522 840
rect 15572 838 15573 840
rect 15497 834 15501 836
rect 15502 832 15503 834
rect 15521 832 15534 838
rect 15495 828 15499 830
rect 15372 804 15438 808
rect 15381 800 15422 804
rect 15462 801 15463 804
rect 15188 793 15198 794
rect 14979 792 14980 793
rect 15052 792 15104 793
rect 15110 792 15126 793
rect 15188 792 15200 793
rect 14865 784 14894 791
rect 14980 789 14986 792
rect 14986 784 14993 789
rect 15046 788 15126 792
rect 15164 790 15165 792
rect 15188 789 15209 792
rect 15188 788 15203 789
rect 15046 786 15110 788
rect 15198 786 15203 788
rect 15209 787 15214 789
rect 15214 786 15218 787
rect 15219 786 15270 800
rect 15282 793 15286 800
rect 15344 793 15349 799
rect 15281 790 15282 793
rect 15342 790 15344 793
rect 14993 783 14994 784
rect 15029 783 15030 785
rect 14778 777 14854 780
rect 14995 779 15001 783
rect 15026 779 15029 783
rect 15052 780 15058 786
rect 15094 781 15106 786
rect 15214 785 15225 786
rect 15216 783 15225 785
rect 15216 782 15228 783
rect 15098 780 15104 781
rect 15164 779 15165 781
rect 15001 777 15006 779
rect 15025 777 15026 779
rect 15163 777 15164 779
rect 15216 777 15225 782
rect 15231 779 15234 781
rect 15234 777 15253 779
rect 15281 777 15290 786
rect 15312 782 15318 788
rect 15339 786 15342 790
rect 15358 782 15364 788
rect 15376 786 15385 800
rect 15388 788 15404 800
rect 15406 796 15442 800
rect 15463 798 15465 801
rect 15490 800 15491 810
rect 15497 798 15499 828
rect 15503 818 15511 830
rect 15520 822 15534 832
rect 15564 836 15572 838
rect 15626 837 15630 841
rect 15658 839 15660 847
rect 15693 838 15703 852
rect 15711 848 15714 852
rect 15841 842 15847 844
rect 15841 838 15855 842
rect 15887 838 15893 844
rect 15894 838 15910 854
rect 15934 838 15940 863
rect 15949 853 15952 863
rect 15952 838 15957 852
rect 15564 822 15571 836
rect 15588 826 15600 832
rect 15585 825 15644 826
rect 15648 825 15658 838
rect 15585 823 15593 825
rect 15644 823 15658 825
rect 15665 823 15668 838
rect 15520 820 15523 822
rect 15584 821 15585 823
rect 15463 796 15499 798
rect 15503 796 15511 808
rect 15520 804 15534 820
rect 15576 816 15584 820
rect 15588 818 15595 820
rect 15576 808 15582 816
rect 15588 814 15589 818
rect 15648 816 15673 823
rect 15682 816 15693 837
rect 15714 822 15726 838
rect 15835 832 15841 838
rect 15839 830 15841 832
rect 15843 830 15876 838
rect 15893 832 15899 838
rect 15910 832 15926 838
rect 15940 832 15941 838
rect 15893 830 15926 832
rect 15957 830 15960 838
rect 15963 830 15975 870
rect 16018 863 16023 874
rect 16065 871 16068 885
rect 16102 881 16112 885
rect 16188 884 16194 890
rect 16198 887 16199 890
rect 16208 886 16215 890
rect 16199 883 16202 885
rect 16205 884 16207 885
rect 16234 884 16240 890
rect 16297 888 16299 896
rect 16199 882 16204 883
rect 16100 874 16118 881
rect 16083 870 16100 874
rect 16102 870 16112 874
rect 16023 859 16025 863
rect 16049 838 16065 870
rect 16083 866 16102 870
rect 16081 863 16083 866
rect 16079 859 16081 863
rect 16095 859 16102 866
rect 16077 856 16079 859
rect 16075 854 16077 856
rect 16068 851 16077 854
rect 16068 839 16075 851
rect 16068 838 16069 839
rect 16025 830 16026 838
rect 16049 830 16068 838
rect 16082 830 16095 859
rect 16112 846 16119 858
rect 16124 848 16125 880
rect 16191 876 16197 879
rect 16188 874 16191 876
rect 16179 869 16188 874
rect 16199 870 16202 882
rect 16236 870 16239 884
rect 16296 881 16297 888
rect 16295 874 16296 881
rect 16172 860 16173 863
rect 16202 860 16204 870
rect 16236 862 16250 870
rect 16292 863 16295 874
rect 16167 848 16172 860
rect 16124 847 16129 848
rect 16124 846 16158 847
rect 16165 846 16170 848
rect 16119 844 16120 846
rect 16164 844 16165 846
rect 16161 842 16163 843
rect 16124 834 16136 841
rect 16146 834 16158 841
rect 16204 830 16215 859
rect 16239 830 16250 862
rect 16291 856 16292 859
rect 16329 856 16347 903
rect 16435 890 16443 902
rect 16447 890 16449 921
rect 16480 920 16481 922
rect 16487 912 16493 924
rect 16543 913 16545 925
rect 16574 924 16590 928
rect 16660 925 16669 934
rect 16652 924 16660 925
rect 16574 913 16652 924
rect 16487 911 16490 912
rect 16490 903 16495 910
rect 16528 905 16590 913
rect 16522 903 16528 905
rect 16481 890 16522 903
rect 16490 888 16495 890
rect 16545 889 16547 905
rect 16443 886 16446 888
rect 16495 886 16496 888
rect 16547 885 16548 888
rect 16446 884 16448 885
rect 16447 883 16449 884
rect 16447 879 16450 883
rect 16496 880 16497 882
rect 16447 878 16451 879
rect 16450 876 16451 878
rect 16497 876 16498 880
rect 16548 876 16549 879
rect 16574 878 16590 905
rect 16451 869 16454 874
rect 16454 863 16456 869
rect 16389 861 16390 862
rect 16456 860 16457 863
rect 16268 851 16284 854
rect 16288 851 16291 856
rect 16327 851 16329 856
rect 16370 854 16382 855
rect 16268 843 16288 851
rect 16324 843 16327 851
rect 16364 849 16382 854
rect 16392 849 16404 855
rect 16364 843 16455 849
rect 16457 848 16461 860
rect 16461 844 16462 847
rect 16478 843 16494 854
rect 16266 839 16269 843
rect 16322 839 16324 843
rect 16358 842 16363 843
rect 16358 840 16362 842
rect 16364 841 16404 843
rect 16351 839 16361 840
rect 16364 839 16370 841
rect 16345 838 16350 839
rect 16364 838 16365 839
rect 16252 830 16266 838
rect 16319 836 16322 838
rect 16341 837 16345 838
rect 16332 836 16338 837
rect 16319 834 16332 836
rect 16309 833 16313 834
rect 16303 832 16309 833
rect 16290 830 16303 832
rect 16319 831 16322 834
rect 15831 827 15839 830
rect 15843 828 15846 830
rect 15830 821 15840 827
rect 15519 802 15520 804
rect 15521 800 15523 804
rect 15648 801 15658 816
rect 15660 812 15668 816
rect 15660 804 15669 812
rect 15673 807 15705 816
rect 15714 807 15726 820
rect 15806 807 15830 821
rect 15831 818 15839 821
rect 15669 801 15670 803
rect 15682 801 15693 807
rect 15705 804 15726 807
rect 15406 788 15422 796
rect 15442 795 15447 796
rect 15447 793 15458 795
rect 15465 794 15472 796
rect 15472 793 15478 794
rect 15489 793 15490 796
rect 15458 792 15463 793
rect 15478 792 15498 793
rect 15501 792 15503 795
rect 15518 794 15519 796
rect 15478 786 15499 792
rect 15515 789 15518 793
rect 15500 788 15518 789
rect 15500 786 15515 788
rect 15571 786 15572 788
rect 15576 786 15582 798
rect 15630 789 15631 801
rect 15645 790 15648 800
rect 15670 797 15698 801
rect 15705 797 15724 804
rect 15794 800 15806 807
rect 15792 799 15794 800
rect 15670 796 15724 797
rect 15785 796 15792 799
rect 15831 796 15839 808
rect 15843 796 15845 828
rect 15911 822 16140 830
rect 15911 820 15913 822
rect 15914 820 16140 822
rect 15911 814 16140 820
rect 16168 814 16290 830
rect 16313 818 16319 831
rect 16348 822 16364 838
rect 16311 815 16318 818
rect 15911 812 16168 814
rect 15913 804 15926 812
rect 15943 807 15945 812
rect 15913 803 15914 804
rect 15914 801 15915 802
rect 15911 796 15914 801
rect 15944 800 15945 807
rect 15956 804 15968 812
rect 15968 803 15969 804
rect 15973 803 15975 808
rect 15992 803 16071 812
rect 15969 802 16071 803
rect 15972 799 15988 802
rect 15589 787 15590 788
rect 15588 786 15594 787
rect 15370 782 15376 786
rect 15487 784 15499 786
rect 12685 747 12691 750
rect 12739 749 12741 750
rect 12694 747 12698 749
rect 12685 746 12694 747
rect 12684 744 12692 746
rect 12703 745 12739 747
rect 12741 745 12749 747
rect 12206 738 12208 743
rect 12237 741 12269 743
rect 12265 740 12270 741
rect 12272 737 12275 739
rect 12325 738 12328 744
rect 12360 739 12363 744
rect 12443 740 12445 744
rect 12460 740 12472 742
rect 12173 734 12174 737
rect 12180 734 12184 737
rect 12172 732 12173 734
rect 12184 732 12188 734
rect 12204 732 12206 737
rect 12234 736 12235 737
rect 12264 734 12274 737
rect 12275 734 12281 737
rect 12287 734 12293 737
rect 12269 732 12274 734
rect 12169 725 12172 731
rect 12188 729 12192 732
rect 12202 729 12204 731
rect 12168 722 12169 724
rect 12164 711 12168 721
rect 12192 712 12220 729
rect 12233 726 12234 731
rect 12274 727 12278 732
rect 12280 731 12293 734
rect 12318 732 12322 734
rect 12316 731 12318 732
rect 12333 731 12339 737
rect 12423 734 12429 740
rect 12441 734 12442 736
rect 12460 734 12475 740
rect 12484 738 12485 742
rect 12633 738 12639 744
rect 12691 738 12697 744
rect 12703 743 12705 745
rect 12483 734 12484 737
rect 12356 732 12357 734
rect 12417 732 12481 734
rect 12278 726 12280 727
rect 12281 726 12287 731
rect 12035 710 12039 711
rect 12040 710 12092 711
rect 12034 706 12098 710
rect 12030 704 12098 706
rect 12161 704 12164 711
rect 11888 698 11894 699
rect 11902 698 11940 699
rect 11882 695 11894 698
rect 11898 695 11946 698
rect 11882 693 11888 695
rect 11898 693 11936 695
rect 11940 693 11946 695
rect 12030 694 12034 704
rect 12040 699 12058 704
rect 12040 698 12046 699
rect 12086 698 12092 704
rect 12159 699 12161 704
rect 12087 696 12088 698
rect 12157 695 12159 698
rect 12193 695 12201 712
rect 12221 709 12224 711
rect 12229 709 12233 726
rect 12280 717 12290 726
rect 12339 725 12345 731
rect 12352 725 12356 732
rect 12417 730 12475 732
rect 12476 730 12481 732
rect 12482 730 12483 732
rect 12417 728 12473 730
rect 12350 722 12351 724
rect 12290 709 12292 717
rect 12344 711 12350 721
rect 12224 708 12226 709
rect 12223 707 12227 708
rect 12223 703 12229 707
rect 12235 705 12236 707
rect 12235 703 12252 705
rect 12227 695 12229 703
rect 12232 699 12234 700
rect 12235 696 12259 699
rect 12292 698 12294 706
rect 12339 702 12344 711
rect 12154 694 12157 695
rect 11718 691 11727 692
rect 11733 691 11734 693
rect 11834 692 11946 693
rect 11834 691 11928 692
rect 11437 688 11440 689
rect 11444 688 11445 690
rect 11565 688 11569 690
rect 11727 689 11749 691
rect 11834 689 11924 691
rect 11058 682 11064 688
rect 11116 682 11122 688
rect 11440 686 11446 688
rect 11063 680 11076 682
rect 11063 676 11070 680
rect 11110 676 11116 682
rect 11444 677 11446 686
rect 11546 681 11565 688
rect 11546 679 11616 681
rect 9382 667 9392 669
rect 9383 665 9392 667
rect 9320 656 9321 658
rect 9327 656 9336 665
rect 9374 656 9388 665
rect 10857 658 10867 669
rect 10859 656 10873 658
rect 10909 656 10925 672
rect 11063 669 11064 676
rect 11440 671 11446 677
rect 11498 678 11565 679
rect 11498 676 11562 678
rect 11616 676 11625 679
rect 11498 671 11504 676
rect 11443 669 11452 671
rect 11063 658 11073 668
rect 11443 658 11445 669
rect 11446 665 11452 669
rect 11492 665 11498 671
rect 11535 669 11546 676
rect 11625 675 11629 676
rect 11629 672 11631 675
rect 11733 671 11737 688
rect 11749 686 11784 689
rect 11834 686 11918 689
rect 11934 686 11940 692
rect 12029 690 12030 693
rect 12150 692 12154 694
rect 12148 691 12150 692
rect 12144 689 12148 691
rect 12140 688 12144 689
rect 12190 688 12193 695
rect 12226 690 12227 694
rect 12235 691 12247 696
rect 12259 693 12273 696
rect 12293 695 12294 698
rect 12423 696 12438 728
rect 12470 726 12473 728
rect 12476 726 12484 730
rect 12470 724 12472 726
rect 12471 700 12472 724
rect 12473 718 12484 726
rect 12473 714 12477 718
rect 12473 710 12476 714
rect 12479 712 12481 718
rect 12735 715 12737 745
rect 12739 742 12749 745
rect 12909 743 12911 749
rect 12919 743 12925 749
rect 12938 746 12961 770
rect 14423 755 14424 777
rect 14452 772 14453 777
rect 14543 774 14582 777
rect 14589 774 14601 777
rect 14453 759 14461 772
rect 14545 768 14582 774
rect 14592 768 14601 774
rect 14658 768 14659 777
rect 14453 755 14464 759
rect 14424 749 14425 755
rect 14461 753 14464 755
rect 14462 750 14467 753
rect 12965 743 12971 749
rect 14436 747 14465 748
rect 14468 747 14469 749
rect 12913 742 12919 743
rect 12741 738 12749 742
rect 12741 735 12759 738
rect 12749 731 12759 735
rect 12911 731 12919 742
rect 12924 738 12925 742
rect 12957 739 12963 742
rect 12922 731 12924 738
rect 12958 737 12963 739
rect 12971 737 12977 743
rect 12709 714 12737 715
rect 12704 713 12737 714
rect 12741 713 12749 725
rect 12759 721 12765 731
rect 12911 721 12922 731
rect 12903 720 12922 721
rect 12903 712 12912 720
rect 12478 710 12479 711
rect 12476 707 12479 710
rect 12738 709 12741 711
rect 12712 708 12715 709
rect 12475 702 12479 707
rect 12700 706 12710 708
rect 12691 704 12700 706
rect 12470 696 12472 699
rect 12476 696 12479 702
rect 12725 701 12737 709
rect 12916 707 12922 720
rect 12959 717 12963 737
rect 12915 706 12916 707
rect 12292 693 12293 694
rect 12273 692 12339 693
rect 12279 691 12339 692
rect 12285 690 12339 691
rect 11784 684 11803 686
rect 11842 684 11906 686
rect 11803 683 11811 684
rect 11811 681 11832 683
rect 11842 681 11901 684
rect 11832 679 11901 681
rect 12025 679 12029 688
rect 12088 686 12090 688
rect 12113 686 12140 688
rect 12189 686 12190 688
rect 12088 684 12120 686
rect 12078 683 12120 684
rect 12051 681 12120 683
rect 12033 679 12120 681
rect 12186 679 12189 684
rect 11842 678 11901 679
rect 11845 677 11880 678
rect 12006 677 12120 679
rect 11845 676 11877 677
rect 11879 676 11880 677
rect 11846 674 11858 676
rect 11860 675 11873 676
rect 11874 675 11879 676
rect 11984 675 12006 677
rect 12012 676 12120 677
rect 12025 675 12029 676
rect 11860 671 11887 675
rect 11936 671 11984 675
rect 12183 673 12186 679
rect 12223 672 12226 688
rect 12287 687 12339 690
rect 12423 688 12475 696
rect 12479 692 12480 694
rect 12633 693 12639 698
rect 12691 693 12697 698
rect 12912 697 12915 706
rect 12963 697 12965 717
rect 13726 703 13748 722
rect 14418 713 14425 725
rect 14430 716 14431 747
rect 14459 745 14464 747
rect 14463 716 14464 745
rect 14465 738 14476 747
rect 14692 740 14696 777
rect 14787 768 14796 777
rect 14839 768 14845 777
rect 15001 776 15025 777
rect 15161 772 15163 777
rect 15225 772 15253 777
rect 15154 759 15161 772
rect 15225 768 15234 772
rect 15272 768 15281 777
rect 15306 776 15312 782
rect 15364 776 15376 782
rect 15488 776 15489 781
rect 15364 766 15368 773
rect 15520 772 15521 786
rect 15572 783 15573 786
rect 15583 784 15585 785
rect 15629 784 15630 788
rect 15644 787 15645 790
rect 15670 789 15714 796
rect 15724 795 15726 796
rect 15726 792 15733 795
rect 15783 793 15785 796
rect 15882 795 15910 796
rect 15733 789 15737 792
rect 15670 788 15692 789
rect 15694 788 15710 789
rect 15737 788 15739 789
rect 15779 788 15783 793
rect 15894 792 15910 795
rect 15940 793 15944 799
rect 15651 787 15658 788
rect 15666 787 15680 788
rect 15739 787 15742 788
rect 15643 786 15651 787
rect 15638 785 15651 786
rect 15670 785 15680 787
rect 15835 786 15841 792
rect 15893 791 15910 792
rect 15937 791 15940 793
rect 15893 789 15949 791
rect 15970 789 15988 799
rect 15893 788 15910 789
rect 15937 788 15940 789
rect 15949 788 15988 789
rect 15990 788 16071 802
rect 16082 800 16095 812
rect 16158 804 16159 807
rect 15893 786 15899 788
rect 15936 786 15937 788
rect 15635 784 15644 785
rect 15573 780 15585 783
rect 15588 780 15589 781
rect 15597 780 15635 784
rect 15573 779 15632 780
rect 15588 774 15600 779
rect 15519 763 15521 772
rect 15638 763 15644 784
rect 15670 784 15684 785
rect 15144 756 15161 759
rect 15485 756 15488 763
rect 15144 755 15154 756
rect 15144 754 15151 755
rect 15484 754 15485 756
rect 15144 753 15148 754
rect 15133 749 15175 753
rect 15133 748 15160 749
rect 15131 747 15133 748
rect 15175 747 15178 749
rect 15117 745 15131 747
rect 14649 738 14655 740
rect 14692 739 14701 740
rect 14469 735 14487 738
rect 14476 725 14487 735
rect 14649 734 14661 738
rect 14695 734 14701 739
rect 15084 738 15117 745
rect 15078 737 15083 738
rect 14643 728 14649 734
rect 14701 729 14707 734
rect 15055 733 15078 737
rect 15132 735 15140 747
rect 15144 746 15149 747
rect 15049 731 15055 733
rect 15043 729 15045 731
rect 14665 728 14796 729
rect 14649 726 14665 728
rect 14701 727 15004 728
rect 15031 727 15037 729
rect 15042 728 15043 729
rect 14796 726 14797 727
rect 15004 726 15037 727
rect 15040 726 15042 728
rect 14430 714 14434 716
rect 14461 714 14464 716
rect 14430 713 14464 714
rect 14469 713 14487 725
rect 14637 714 14645 726
rect 14649 724 14655 726
rect 14425 711 14426 713
rect 14426 708 14431 711
rect 14464 708 14469 711
rect 14430 707 14442 708
rect 13697 697 13720 698
rect 13725 697 13748 703
rect 14429 701 14442 707
rect 14452 701 14464 708
rect 14476 707 14487 713
rect 12912 694 12919 697
rect 12633 692 12697 693
rect 12286 685 12339 687
rect 12281 679 12345 685
rect 12417 682 12482 688
rect 12639 686 12645 692
rect 12685 686 12691 692
rect 12703 690 12704 694
rect 12911 690 12912 694
rect 12913 693 12919 694
rect 12971 693 12977 697
rect 14429 694 14431 701
rect 12913 691 12977 693
rect 12910 688 12911 690
rect 12286 673 12293 679
rect 12333 673 12339 679
rect 12423 676 12429 682
rect 12469 676 12475 682
rect 11860 670 11898 671
rect 11925 670 11968 671
rect 11527 662 11535 669
rect 11633 667 11634 669
rect 11523 659 11527 662
rect 11634 660 11649 667
rect 11737 662 11739 669
rect 11860 664 11968 670
rect 12286 669 12291 673
rect 12426 672 12428 676
rect 12419 670 12428 672
rect 11862 662 11872 664
rect 12025 662 12026 669
rect 11739 660 11740 662
rect 11521 658 11523 659
rect 11073 656 11075 658
rect 11223 656 11225 657
rect 11443 656 11444 658
rect 11519 656 11521 658
rect 8254 652 8255 653
rect 8502 652 8503 653
rect 8535 652 8572 654
rect 8640 653 8641 656
rect 8696 653 8697 655
rect 8839 654 8840 656
rect 7628 651 7630 652
rect 7495 649 7571 651
rect 7623 649 7628 651
rect 7863 649 7867 652
rect 7926 650 7928 652
rect 7916 649 7926 650
rect 7578 648 7622 649
rect 7874 640 7890 649
rect 7891 648 7892 649
rect 8156 647 8158 651
rect 8176 647 8288 652
rect 8170 644 8288 647
rect 8386 644 8535 652
rect 8170 640 8186 644
rect 8288 641 8299 644
rect 8339 641 8386 644
rect 8299 640 8339 641
rect 8476 640 8492 644
rect 5284 639 5285 640
rect 8538 636 8568 652
rect 8676 640 8692 653
rect 8839 644 8849 654
rect 9112 652 9125 656
rect 9147 652 9180 656
rect 9380 652 9383 656
rect 9127 651 9146 652
rect 8895 645 8896 651
rect 8850 640 8866 644
rect 8868 640 8884 644
rect 9164 640 9180 652
rect 9321 645 9331 652
rect 9375 646 9380 652
rect 9369 645 9375 646
rect 9331 644 9372 645
rect 9356 640 9372 644
rect 10875 640 10891 656
rect 10893 640 10909 656
rect 11076 653 11078 656
rect 11216 653 11222 656
rect 11445 653 11448 656
rect 11515 653 11519 656
rect 11078 651 11080 653
rect 11215 652 11216 653
rect 11513 652 11515 653
rect 11649 652 11761 660
rect 11853 658 11862 662
rect 12090 659 12093 669
rect 12222 666 12223 669
rect 11849 656 11853 658
rect 12026 656 12027 658
rect 12091 657 12093 659
rect 12089 656 12093 657
rect 11844 653 11849 656
rect 12027 653 12030 656
rect 12088 653 12089 656
rect 12123 654 12153 663
rect 12157 654 12170 660
rect 12222 659 12224 666
rect 12285 665 12293 669
rect 12283 658 12293 665
rect 12224 656 12225 658
rect 12282 656 12293 658
rect 12419 660 12426 670
rect 12481 669 12482 682
rect 12704 675 12705 688
rect 12697 669 12705 675
rect 12906 674 12910 686
rect 12919 685 12925 691
rect 12965 685 12971 691
rect 14487 690 14494 707
rect 14637 692 14645 704
rect 14649 694 14651 724
rect 14798 719 14802 726
rect 15004 723 15039 726
rect 15077 723 15083 729
rect 14802 708 14809 719
rect 15025 717 15031 723
rect 15032 719 15039 723
rect 15083 719 15089 723
rect 15132 719 15140 725
rect 15144 719 15146 746
rect 15473 744 15479 750
rect 15481 744 15484 754
rect 15519 750 15520 763
rect 15625 757 15631 762
rect 15637 757 15638 762
rect 15670 758 15680 784
rect 15684 783 15688 784
rect 15743 783 15749 786
rect 15778 783 15779 786
rect 15841 784 15855 786
rect 15841 783 15847 784
rect 15879 783 15883 784
rect 15750 781 15752 782
rect 15752 780 15755 781
rect 15768 780 15778 783
rect 15697 775 15703 779
rect 15703 772 15708 775
rect 15755 772 15778 780
rect 15709 766 15733 772
rect 15768 769 15800 772
rect 15806 769 15879 783
rect 15887 780 15893 786
rect 15894 784 15895 785
rect 15935 784 15936 786
rect 15970 783 15973 788
rect 15979 787 16071 788
rect 16043 786 16071 787
rect 16020 785 16071 786
rect 16079 785 16082 799
rect 16157 797 16158 801
rect 16204 800 16215 814
rect 16239 804 16250 814
rect 16252 804 16268 814
rect 16305 807 16318 815
rect 16302 805 16318 807
rect 16348 805 16364 820
rect 16402 811 16404 841
rect 16408 831 16416 843
rect 16455 838 16495 843
rect 16498 842 16505 874
rect 16540 840 16548 852
rect 16552 842 16554 874
rect 16584 857 16589 874
rect 16584 842 16586 857
rect 16589 852 16590 856
rect 16552 840 16586 842
rect 16590 840 16598 852
rect 16505 838 16506 840
rect 16592 838 16594 840
rect 16495 837 16510 838
rect 16552 837 16553 838
rect 16504 836 16510 837
rect 16549 836 16551 837
rect 16386 809 16404 811
rect 16408 809 16416 821
rect 16465 805 16475 836
rect 16504 832 16519 836
rect 16507 808 16519 832
rect 16552 828 16564 836
rect 16574 828 16586 836
rect 16592 828 16606 838
rect 16553 820 16555 828
rect 16506 807 16519 808
rect 16291 804 16404 805
rect 16268 803 16404 804
rect 16156 791 16157 796
rect 16155 788 16156 791
rect 16215 789 16218 799
rect 16250 794 16258 800
rect 16268 795 16284 803
rect 16286 799 16404 803
rect 16475 801 16479 805
rect 16505 804 16519 807
rect 16540 815 16555 820
rect 16594 822 16606 828
rect 16594 820 16596 822
rect 16540 804 16556 815
rect 16594 805 16606 820
rect 17046 819 17047 1015
rect 17236 819 17237 1015
rect 17322 819 17323 1015
rect 17595 819 17596 1015
rect 17792 819 17793 1015
rect 18014 1013 18030 1015
rect 18036 1013 18048 1022
rect 18056 1020 18085 1023
rect 18085 1014 18089 1020
rect 18825 1018 18877 1020
rect 19097 1018 19111 1023
rect 19307 1020 19308 1023
rect 18797 1016 18877 1018
rect 18797 1015 18848 1016
rect 18089 1013 18090 1014
rect 18772 1013 18797 1015
rect 18819 1014 18825 1015
rect 18848 1014 18853 1015
rect 18010 1011 18014 1013
rect 18026 1010 18030 1013
rect 18738 1011 18768 1013
rect 18814 1012 18819 1014
rect 18002 998 18010 1010
rect 18009 988 18010 998
rect 18014 1007 18048 1010
rect 18014 1003 18016 1007
rect 18014 996 18015 1003
rect 18026 1001 18030 1007
rect 18045 1005 18048 1007
rect 18051 1004 18060 1010
rect 18013 994 18015 996
rect 18012 988 18018 994
rect 18023 988 18026 1001
rect 18006 982 18012 988
rect 18013 986 18014 988
rect 18013 976 18015 986
rect 18046 982 18048 1004
rect 18052 998 18060 1004
rect 18090 1001 18099 1010
rect 18621 1005 18635 1007
rect 18647 1005 18738 1011
rect 18810 1007 18814 1012
rect 18621 1004 18647 1005
rect 18621 1003 18635 1004
rect 18615 1002 18635 1003
rect 18656 1002 18661 1005
rect 18806 1002 18810 1007
rect 18853 1005 18870 1014
rect 18870 1004 18872 1005
rect 18058 988 18064 994
rect 18081 992 18090 1001
rect 18606 997 18630 1002
rect 18661 997 18667 1002
rect 18805 1001 18806 1002
rect 18877 1001 18894 1016
rect 19111 1015 19118 1018
rect 19306 1016 19307 1020
rect 19118 1014 19121 1015
rect 19121 1005 19143 1014
rect 19304 1012 19306 1016
rect 19344 1014 19348 1031
rect 19350 1027 19358 1039
rect 19616 1037 19628 1045
rect 19677 1041 19687 1045
rect 19688 1041 19694 1045
rect 19652 1037 19694 1041
rect 19746 1039 19752 1045
rect 19899 1044 19905 1050
rect 19945 1048 19955 1050
rect 19908 1044 19920 1048
rect 19930 1044 19942 1048
rect 19945 1044 19951 1048
rect 19893 1038 19899 1044
rect 19951 1038 19957 1044
rect 19397 1020 19407 1036
rect 19428 1034 19440 1037
rect 19622 1036 19628 1037
rect 19674 1036 19677 1037
rect 19422 1033 19442 1034
rect 19616 1033 19622 1036
rect 19658 1033 19688 1036
rect 19422 1031 19428 1033
rect 19442 1031 19472 1033
rect 19419 1025 19422 1031
rect 19416 1022 19422 1025
rect 19474 1024 19495 1031
rect 19522 1024 19528 1030
rect 19143 1004 19146 1005
rect 19003 1001 19004 1004
rect 18064 982 18070 988
rect 18081 986 18085 992
rect 18593 989 18606 997
rect 18615 993 18630 997
rect 18013 962 18014 976
rect 18079 974 18080 979
rect 18237 976 18253 984
rect 18420 976 18436 989
rect 18503 979 18520 989
rect 18579 981 18593 989
rect 18573 979 18579 981
rect 18520 978 18573 979
rect 18604 977 18612 989
rect 18616 987 18621 989
rect 18667 987 18680 997
rect 18237 974 18294 976
rect 18075 957 18079 972
rect 18237 968 18282 974
rect 18294 968 18298 974
rect 18013 944 18020 957
rect 18074 953 18075 956
rect 18073 949 18074 952
rect 18076 944 18090 953
rect 18221 952 18237 968
rect 18298 961 18303 968
rect 18228 944 18237 952
rect 18006 936 18012 942
rect 18012 930 18018 936
rect 18020 934 18045 944
rect 18060 936 18076 944
rect 18058 934 18076 936
rect 18224 935 18228 944
rect 18231 940 18237 941
rect 18231 939 18273 940
rect 18277 939 18283 941
rect 18231 936 18242 939
rect 18231 935 18237 936
rect 18273 935 18283 939
rect 18224 934 18231 935
rect 18051 929 18054 934
rect 18058 930 18064 934
rect 18047 923 18050 928
rect 18221 925 18224 934
rect 18225 929 18231 934
rect 18283 929 18289 935
rect 18290 933 18302 941
rect 18363 934 18369 940
rect 18409 934 18415 940
rect 18420 934 18426 956
rect 18485 952 18491 958
rect 18531 952 18537 958
rect 18604 956 18612 967
rect 18616 958 18618 987
rect 18866 984 18868 1001
rect 18872 999 18894 1001
rect 18872 989 18880 999
rect 18998 992 19003 1001
rect 19146 996 19167 1004
rect 19301 1002 19304 1011
rect 19344 1007 19346 1014
rect 19335 1005 19346 1007
rect 19350 1010 19358 1017
rect 19350 1005 19363 1010
rect 19348 1004 19349 1005
rect 19354 1001 19363 1005
rect 19397 1002 19407 1018
rect 19416 1015 19419 1022
rect 19470 1018 19476 1024
rect 19528 1018 19534 1024
rect 19604 1021 19612 1033
rect 19616 1031 19650 1033
rect 19616 1030 19622 1031
rect 19616 1029 19619 1030
rect 19416 1014 19418 1015
rect 19416 1013 19420 1014
rect 19418 1001 19420 1013
rect 19056 995 19089 996
rect 19167 995 19169 996
rect 19091 993 19097 995
rect 18998 986 19004 992
rect 19056 987 19062 992
rect 19097 991 19101 993
rect 19169 991 19179 995
rect 19299 991 19301 997
rect 19341 993 19354 1001
rect 19416 998 19420 1001
rect 19604 999 19612 1011
rect 19616 1002 19618 1029
rect 19896 1024 19899 1036
rect 19951 1032 19954 1036
rect 19904 1018 19908 1031
rect 19951 1021 19967 1032
rect 19967 1018 19983 1021
rect 19693 1007 19694 1008
rect 19694 1005 19695 1006
rect 19616 1001 19619 1002
rect 19662 1001 19690 1002
rect 19616 999 19628 1001
rect 19662 1000 19688 1001
rect 19346 992 19354 993
rect 19407 991 19411 996
rect 19416 991 19421 998
rect 19616 997 19617 999
rect 19662 998 19684 1000
rect 19690 999 19694 1001
rect 19617 995 19620 997
rect 19662 996 19677 998
rect 19616 993 19622 995
rect 19662 994 19678 996
rect 19688 995 19694 999
rect 19697 997 19702 1003
rect 19746 1001 19755 1010
rect 19881 1001 19890 1010
rect 19890 1000 19896 1001
rect 18725 981 18741 984
rect 18743 981 18759 984
rect 18719 978 18739 981
rect 18860 979 18872 984
rect 18996 979 18997 983
rect 19004 980 19010 986
rect 19014 983 19082 987
rect 19101 986 19113 991
rect 18763 974 18764 978
rect 18721 972 18813 974
rect 18860 972 18880 979
rect 18995 974 18996 979
rect 19014 977 19040 983
rect 19050 980 19056 983
rect 19082 977 19095 983
rect 19113 978 19134 986
rect 19179 978 19213 991
rect 19345 988 19346 990
rect 19283 979 19289 985
rect 19299 983 19300 987
rect 19342 985 19345 986
rect 18994 972 18995 974
rect 19032 972 19040 977
rect 18625 963 18721 972
rect 18763 969 18764 972
rect 18722 963 18734 965
rect 18625 960 18722 963
rect 18616 957 18620 958
rect 18625 957 18721 960
rect 18616 956 18625 957
rect 18599 955 18623 956
rect 18627 955 18650 956
rect 18599 953 18618 955
rect 18667 954 18682 957
rect 18592 952 18599 953
rect 18612 952 18613 953
rect 18479 946 18485 952
rect 18537 946 18543 952
rect 18573 949 18592 952
rect 18660 951 18667 954
rect 18616 950 18627 951
rect 18658 950 18660 951
rect 18551 946 18573 949
rect 18543 945 18565 946
rect 18616 943 18628 950
rect 18679 939 18680 954
rect 18709 952 18719 957
rect 18718 939 18719 952
rect 18764 952 18775 968
rect 18736 942 18744 944
rect 18726 940 18736 942
rect 18724 939 18726 940
rect 18304 932 18306 933
rect 18277 927 18302 929
rect 18219 924 18221 925
rect 18042 914 18047 923
rect 18135 922 18165 924
rect 18215 922 18219 924
rect 18126 916 18135 922
rect 18165 916 18215 922
rect 18040 907 18042 914
rect 18008 895 18009 905
rect 18038 896 18040 907
rect 18111 906 18126 916
rect 18300 915 18302 927
rect 18306 917 18314 929
rect 18351 928 18363 934
rect 18415 928 18426 934
rect 18420 922 18426 928
rect 18537 926 18540 930
rect 18666 927 18724 939
rect 18764 938 18768 952
rect 18805 947 18806 968
rect 18813 965 18885 972
rect 18809 963 18885 965
rect 18813 956 18885 963
rect 18894 962 18895 968
rect 18888 956 18895 962
rect 18934 956 18940 962
rect 18989 956 18994 972
rect 18856 955 18897 956
rect 18882 950 18897 955
rect 18940 950 18946 956
rect 18771 942 18817 944
rect 18817 940 18825 942
rect 18825 939 18828 940
rect 18736 930 18748 938
rect 18758 930 18770 938
rect 18661 926 18666 927
rect 18300 906 18303 915
rect 18339 910 18344 922
rect 18422 916 18429 922
rect 18429 914 18432 916
rect 18540 914 18554 926
rect 18647 923 18661 926
rect 18670 924 18679 927
rect 18768 926 18770 930
rect 18828 927 18875 939
rect 18888 935 18897 950
rect 18987 949 18989 956
rect 19005 952 19014 968
rect 19023 955 19032 972
rect 19095 968 19112 977
rect 19134 968 19173 978
rect 18986 946 18987 949
rect 18890 934 18895 935
rect 18940 933 18946 936
rect 18875 926 18880 927
rect 18888 926 18890 933
rect 18946 930 18953 933
rect 18963 930 18975 938
rect 18983 937 18985 942
rect 19005 937 19014 950
rect 19020 946 19023 955
rect 19065 954 19094 964
rect 19112 963 19173 968
rect 19112 957 19134 963
rect 19173 960 19183 963
rect 19058 945 19094 954
rect 19105 952 19114 954
rect 19017 937 19019 942
rect 18976 926 18983 937
rect 19005 934 19017 937
rect 19049 936 19058 945
rect 19065 944 19094 945
rect 19095 945 19114 952
rect 19134 950 19155 957
rect 19183 956 19193 960
rect 19213 956 19270 978
rect 19289 973 19295 979
rect 19300 977 19301 983
rect 19341 979 19347 985
rect 19301 972 19302 977
rect 19335 974 19341 979
rect 19342 974 19345 979
rect 19335 973 19342 974
rect 19341 972 19342 973
rect 19299 968 19302 972
rect 19350 971 19352 991
rect 19411 985 19417 991
rect 19422 988 19423 990
rect 19424 986 19427 987
rect 19427 985 19432 986
rect 19411 984 19467 985
rect 19616 984 19627 993
rect 19662 990 19674 994
rect 19688 993 19702 995
rect 19746 993 19752 999
rect 19890 998 19897 1000
rect 19899 998 19908 1018
rect 19983 1015 19996 1018
rect 20620 1015 20621 1026
rect 20810 1015 20811 1026
rect 20896 1015 20897 1026
rect 21169 1015 21170 1026
rect 21366 1015 21367 1026
rect 19996 1001 20060 1015
rect 20060 998 20070 1001
rect 19690 992 19700 993
rect 19737 992 19746 993
rect 19890 992 19908 998
rect 19951 992 19957 998
rect 20070 992 20115 998
rect 20210 994 20228 995
rect 20198 992 20210 994
rect 19662 986 19680 990
rect 19694 987 19700 992
rect 19740 987 19746 992
rect 19899 991 19905 992
rect 19899 989 19906 991
rect 19907 990 19908 992
rect 19937 991 19940 992
rect 19899 986 19905 989
rect 19907 987 19911 988
rect 19926 987 19937 991
rect 19942 986 19951 992
rect 20070 988 20198 992
rect 19411 983 19476 984
rect 19620 983 19628 984
rect 19428 981 19476 983
rect 19428 979 19440 981
rect 19622 978 19638 983
rect 19643 981 19644 984
rect 19470 972 19476 978
rect 19528 972 19534 978
rect 19299 967 19304 968
rect 19340 967 19341 971
rect 19290 958 19304 967
rect 19193 954 19198 956
rect 19270 955 19289 956
rect 19290 955 19302 958
rect 19198 951 19205 954
rect 19270 951 19302 955
rect 19304 951 19305 957
rect 19205 950 19207 951
rect 19095 944 19107 945
rect 19065 943 19072 944
rect 19114 943 19123 945
rect 19065 942 19070 943
rect 19065 941 19067 942
rect 19065 940 19111 941
rect 19112 940 19123 943
rect 19061 939 19066 940
rect 19073 939 19107 940
rect 19061 938 19107 939
rect 19061 937 19073 938
rect 19010 926 19017 934
rect 19060 931 19073 937
rect 19104 936 19107 938
rect 19111 937 19123 940
rect 19155 937 19257 950
rect 19270 949 19290 951
rect 19293 949 19309 950
rect 19283 948 19309 949
rect 19283 946 19290 948
rect 19293 945 19310 948
rect 19335 946 19340 967
rect 19352 951 19354 968
rect 19476 966 19482 972
rect 19485 967 19488 972
rect 19354 949 19359 950
rect 19105 931 19107 936
rect 19118 931 19124 937
rect 19155 934 19289 937
rect 19293 934 19309 945
rect 19310 943 19320 945
rect 19347 943 19359 949
rect 19488 948 19495 967
rect 19522 966 19534 972
rect 19627 968 19638 978
rect 19662 980 19681 986
rect 19662 973 19699 980
rect 19823 976 19839 984
rect 19901 982 19904 986
rect 19900 976 19901 981
rect 19644 968 19647 972
rect 19528 945 19534 966
rect 19638 953 19650 968
rect 19666 965 19699 973
rect 19783 968 19786 976
rect 19824 975 19839 976
rect 19899 970 19900 975
rect 19942 969 19945 986
rect 19954 972 20055 977
rect 20055 969 20066 972
rect 20097 969 20198 988
rect 20228 980 20250 994
rect 19644 951 19647 953
rect 19650 951 19652 953
rect 19320 934 19384 943
rect 19652 942 19672 951
rect 19681 948 19699 965
rect 19779 957 19783 968
rect 19774 955 19779 957
rect 19736 950 19737 953
rect 19485 936 19567 942
rect 19468 934 19485 936
rect 19061 930 19073 931
rect 18638 921 18647 923
rect 18626 920 18638 921
rect 18665 920 18670 924
rect 18579 915 18665 920
rect 18567 914 18579 915
rect 18607 914 18626 915
rect 18724 914 18732 926
rect 18736 924 18770 926
rect 18432 913 18562 914
rect 18540 909 18554 913
rect 18596 911 18607 914
rect 18589 907 18595 911
rect 18107 900 18111 906
rect 18300 902 18302 906
rect 18037 891 18038 895
rect 18102 892 18107 899
rect 18285 898 18302 902
rect 18281 897 18302 898
rect 18277 896 18302 897
rect 18274 895 18302 896
rect 18306 895 18314 907
rect 18479 900 18485 906
rect 18289 891 18302 895
rect 18305 892 18306 894
rect 18036 888 18037 891
rect 18099 887 18102 891
rect 18276 889 18289 891
rect 18098 886 18099 887
rect 18225 886 18231 889
rect 18251 887 18289 889
rect 18251 886 18276 887
rect 18091 875 18098 885
rect 18190 875 18273 886
rect 18283 883 18289 887
rect 18290 883 18302 891
rect 18339 888 18344 900
rect 18485 894 18491 900
rect 18513 892 18526 900
rect 18556 892 18567 907
rect 18581 900 18586 904
rect 18718 901 18727 913
rect 18736 901 18738 924
rect 18513 889 18522 892
rect 18526 891 18528 892
rect 18568 889 18570 891
rect 18578 889 18587 898
rect 18727 892 18738 901
rect 18768 892 18770 924
rect 18774 914 18782 926
rect 18880 924 18890 926
rect 18947 924 18975 926
rect 18976 924 18987 926
rect 18880 923 18888 924
rect 18885 921 18888 923
rect 18940 921 18941 924
rect 18973 921 18987 924
rect 18806 907 18820 921
rect 18875 910 18885 921
rect 18939 917 18940 921
rect 18875 907 18888 910
rect 18938 907 18939 916
rect 18973 915 18975 921
rect 18976 915 18987 921
rect 19010 924 19018 926
rect 19010 915 19017 924
rect 19018 921 19022 924
rect 19021 918 19027 921
rect 19022 916 19027 918
rect 18973 911 18976 915
rect 18978 914 18987 915
rect 18978 912 18979 914
rect 18820 906 18875 907
rect 18882 904 18888 907
rect 18937 904 18938 906
rect 18940 904 18946 910
rect 18973 906 18975 911
rect 18979 907 18981 912
rect 18981 906 18982 907
rect 18972 904 18975 906
rect 18982 904 18983 906
rect 18888 898 18894 904
rect 18930 902 18933 904
rect 18934 902 18940 904
rect 18929 898 18940 902
rect 18971 901 18972 904
rect 18929 892 18936 898
rect 18970 897 18971 900
rect 18968 894 18970 895
rect 18973 894 18975 904
rect 18941 892 18975 894
rect 18979 901 18987 904
rect 18979 892 18993 901
rect 18968 891 18970 892
rect 18993 890 18996 892
rect 18036 871 18037 875
rect 18089 871 18091 874
rect 18160 871 18190 875
rect 18088 870 18089 871
rect 18152 870 18160 871
rect 18150 869 18152 870
rect 18087 868 18088 869
rect 18148 868 18150 869
rect 18239 868 18241 875
rect 18274 868 18275 879
rect 18277 877 18283 883
rect 18357 882 18363 888
rect 18415 882 18421 888
rect 18351 876 18369 882
rect 18409 876 18415 882
rect 18522 880 18531 889
rect 18568 888 18578 889
rect 18966 888 18968 889
rect 18569 887 18578 888
rect 18569 880 18589 887
rect 18771 885 18772 888
rect 18732 882 18733 884
rect 18941 880 18953 888
rect 18963 882 18975 888
rect 18996 884 18998 890
rect 19000 885 19010 915
rect 19027 912 19040 916
rect 19040 907 19052 912
rect 19055 906 19057 907
rect 19066 906 19073 930
rect 19118 928 19119 931
rect 19241 919 19289 934
rect 19309 932 19384 934
rect 19401 933 19452 934
rect 19454 933 19465 934
rect 19401 932 19462 933
rect 19309 930 19401 932
rect 19057 904 19062 906
rect 19066 904 19118 906
rect 19062 901 19118 904
rect 19066 899 19118 901
rect 19049 889 19058 898
rect 19066 896 19135 899
rect 19066 891 19123 896
rect 19135 892 19160 896
rect 19257 894 19265 919
rect 19289 916 19296 919
rect 19309 918 19325 930
rect 19327 918 19343 930
rect 19448 929 19463 932
rect 19444 927 19448 929
rect 19428 922 19444 927
rect 19454 926 19463 929
rect 19497 926 19504 936
rect 19457 920 19462 922
rect 19275 900 19279 916
rect 19296 914 19327 916
rect 19328 914 19330 918
rect 19296 909 19328 914
rect 19319 907 19336 909
rect 19319 902 19328 907
rect 19336 906 19340 907
rect 19279 896 19280 899
rect 19299 898 19319 902
rect 19060 889 19124 891
rect 19160 890 19172 892
rect 19256 890 19257 893
rect 19058 885 19124 889
rect 18962 880 18975 882
rect 18532 875 18535 880
rect 18576 879 18589 880
rect 18074 864 18087 868
rect 18142 864 18148 868
rect 18068 862 18074 864
rect 18139 862 18142 864
rect 18064 856 18068 862
rect 18132 857 18139 862
rect 18131 856 18132 857
rect 18062 841 18064 855
rect 18128 849 18131 855
rect 18130 838 18139 842
rect 18177 838 18186 842
rect 18189 838 18205 854
rect 18207 838 18223 854
rect 18241 838 18245 867
rect 18272 847 18274 867
rect 18061 833 18062 838
rect 18128 833 18139 838
rect 18173 833 18189 838
rect 18121 832 18134 833
rect 18173 832 18195 833
rect 18060 825 18061 832
rect 18119 831 18128 832
rect 18059 819 18060 822
rect 16596 804 16606 805
rect 18058 812 18059 816
rect 18058 804 18062 812
rect 18119 811 18121 831
rect 18122 826 18128 831
rect 18127 822 18128 826
rect 18160 824 18195 832
rect 18160 822 18189 824
rect 18234 822 18239 838
rect 18272 833 18273 838
rect 18380 833 18392 864
rect 18535 860 18542 875
rect 18574 873 18589 875
rect 18414 833 18426 838
rect 18437 837 18449 845
rect 18503 838 18519 854
rect 18542 842 18551 860
rect 18543 841 18551 842
rect 18555 845 18556 862
rect 18555 843 18559 845
rect 18587 844 18589 873
rect 18590 869 18601 875
rect 18593 863 18601 869
rect 18597 859 18600 863
rect 18733 860 18737 879
rect 18770 866 18771 880
rect 18852 867 18858 873
rect 18898 867 18904 873
rect 18962 870 18966 880
rect 18995 870 19000 884
rect 19058 880 19072 885
rect 19066 871 19072 880
rect 19108 880 19118 885
rect 19108 870 19109 880
rect 19112 879 19118 880
rect 19172 879 19239 890
rect 19255 885 19256 889
rect 19254 881 19255 885
rect 19240 875 19244 879
rect 19244 872 19247 875
rect 19251 871 19254 881
rect 19280 879 19284 896
rect 19294 891 19299 898
rect 19340 892 19397 906
rect 19397 891 19400 892
rect 19291 881 19293 889
rect 19400 888 19414 891
rect 19460 890 19462 920
rect 19466 910 19474 922
rect 19504 914 19509 926
rect 19509 902 19514 914
rect 19534 910 19541 936
rect 19567 934 19571 936
rect 19648 935 19649 942
rect 19672 936 19684 942
rect 19571 933 19572 934
rect 19572 927 19575 933
rect 19575 922 19578 927
rect 19578 919 19580 922
rect 19580 916 19581 919
rect 19431 888 19462 890
rect 19466 888 19474 900
rect 19514 899 19515 902
rect 19541 900 19543 910
rect 19581 902 19588 916
rect 19649 910 19653 935
rect 19684 934 19688 936
rect 19699 935 19700 942
rect 19686 933 19692 934
rect 19686 932 19694 933
rect 19700 932 19701 935
rect 19736 934 19751 950
rect 19774 948 19786 955
rect 19773 947 19786 948
rect 19796 947 19808 955
rect 19839 952 19855 968
rect 19770 945 19779 947
rect 19769 943 19770 945
rect 19773 943 19779 945
rect 19812 943 19813 945
rect 19819 943 19825 948
rect 19762 942 19769 943
rect 19773 942 19808 943
rect 19812 942 19825 943
rect 19762 937 19773 942
rect 19774 941 19808 942
rect 19760 934 19766 937
rect 19767 936 19773 937
rect 19807 936 19808 941
rect 19825 936 19831 942
rect 19839 934 19855 950
rect 19891 934 19899 968
rect 19945 956 19946 968
rect 19950 965 19951 969
rect 20066 968 20085 969
rect 20093 968 20097 969
rect 20057 964 20093 968
rect 20143 965 20147 969
rect 19756 932 19760 934
rect 19694 931 19735 932
rect 19700 918 19717 931
rect 19719 926 19735 931
rect 19753 930 19756 932
rect 19746 926 19753 930
rect 19838 927 19839 931
rect 19890 927 19891 932
rect 19719 918 19746 926
rect 19837 920 19839 927
rect 19889 922 19890 927
rect 19900 922 19908 934
rect 19912 922 19914 956
rect 19950 951 19951 964
rect 20057 960 20105 964
rect 20048 954 20057 960
rect 19945 945 19946 951
rect 19951 936 19952 945
rect 20037 936 20048 954
rect 20086 949 20105 960
rect 20105 948 20107 949
rect 20147 948 20152 965
rect 20250 961 20253 980
rect 20253 954 20254 960
rect 20107 945 20111 948
rect 20152 945 20153 948
rect 20032 934 20048 936
rect 19952 928 19958 934
rect 19953 922 19958 928
rect 20032 928 20044 934
rect 20054 928 20066 936
rect 20111 934 20126 945
rect 20153 934 20157 945
rect 20254 934 20257 954
rect 20126 932 20127 934
rect 20127 928 20128 930
rect 20157 929 20159 934
rect 20032 924 20037 928
rect 20070 926 20071 928
rect 20072 924 20075 925
rect 19836 919 19839 920
rect 19700 905 19701 918
rect 19728 916 19746 918
rect 19835 918 19839 919
rect 19835 916 19836 918
rect 19888 916 19889 919
rect 19908 916 19909 921
rect 19722 912 19728 916
rect 19831 909 19835 916
rect 19887 909 19888 916
rect 19909 912 19911 916
rect 19939 913 19946 922
rect 19953 916 19954 922
rect 19932 911 19939 913
rect 19950 911 19954 916
rect 20020 912 20028 924
rect 20032 922 20066 924
rect 20032 921 20035 922
rect 19912 910 19950 911
rect 19701 902 19702 904
rect 19588 899 19590 902
rect 19543 894 19544 899
rect 19590 896 19591 899
rect 19414 885 19425 888
rect 19428 885 19467 888
rect 19425 884 19467 885
rect 19284 872 19286 879
rect 19286 870 19287 872
rect 19288 871 19291 881
rect 19428 879 19467 884
rect 19516 881 19518 889
rect 19450 876 19462 879
rect 19467 874 19489 879
rect 19518 874 19519 881
rect 19503 872 19508 874
rect 18937 868 18938 869
rect 18961 867 18962 870
rect 18846 861 18852 867
rect 18904 861 18910 867
rect 18959 860 18961 867
rect 18600 854 18606 858
rect 18600 853 18615 854
rect 18586 843 18589 844
rect 18555 841 18589 843
rect 18593 850 18615 853
rect 18737 852 18738 858
rect 18771 854 18772 858
rect 18593 841 18601 850
rect 18606 840 18615 850
rect 18160 820 18180 822
rect 18188 820 18208 822
rect 18118 810 18121 811
rect 18119 804 18121 810
rect 18127 804 18143 820
rect 18180 819 18188 820
rect 18199 816 18234 817
rect 18233 812 18234 816
rect 16504 803 16505 804
rect 16503 801 16504 802
rect 16451 799 16494 801
rect 16286 796 16451 799
rect 16286 795 16392 796
rect 16475 795 16494 799
rect 16268 794 16302 795
rect 16250 792 16284 794
rect 16229 789 16258 792
rect 16144 785 16155 788
rect 16204 787 16229 789
rect 16191 786 16204 787
rect 16187 785 16191 786
rect 16046 784 16049 785
rect 16067 784 16155 785
rect 16067 783 16144 784
rect 16160 783 16187 785
rect 16215 784 16218 787
rect 15889 779 15890 780
rect 15927 769 15935 783
rect 15969 778 15970 783
rect 16045 781 16046 783
rect 16068 782 16070 783
rect 16044 778 16045 781
rect 16070 780 16073 782
rect 16078 781 16079 783
rect 16136 782 16160 783
rect 16125 779 16136 782
rect 16073 778 16076 779
rect 15625 756 15643 757
rect 15671 756 15677 758
rect 15619 750 15683 756
rect 15708 753 15738 766
rect 15768 763 15806 769
rect 15924 763 15927 769
rect 15768 759 15800 763
rect 15767 756 15768 758
rect 15708 750 15744 753
rect 15765 752 15767 756
rect 15769 755 15800 759
rect 15797 754 15799 755
rect 15800 754 15803 755
rect 15919 754 15924 763
rect 15796 752 15797 754
rect 15803 751 15808 754
rect 15918 752 15919 754
rect 15519 744 15525 750
rect 15625 745 15677 750
rect 15429 742 15473 744
rect 15278 741 15312 742
rect 15429 741 15435 742
rect 15241 740 15278 741
rect 15218 739 15241 740
rect 15215 737 15218 739
rect 15467 738 15473 742
rect 15525 738 15531 744
rect 15190 723 15215 737
rect 15306 730 15312 736
rect 15364 731 15370 736
rect 15619 733 15631 745
rect 15665 735 15670 745
rect 15395 731 15431 733
rect 15312 724 15318 730
rect 15336 729 15395 731
rect 15431 729 15437 731
rect 15334 726 15336 729
rect 15185 720 15190 723
rect 15083 717 15165 719
rect 15086 716 15165 717
rect 15182 716 15190 720
rect 15132 713 15140 716
rect 15144 715 15146 716
rect 15165 715 15194 716
rect 15144 713 15178 715
rect 15175 709 15178 713
rect 15182 713 15190 715
rect 15194 714 15222 715
rect 15182 711 15185 713
rect 15179 709 15182 711
rect 15222 710 15236 714
rect 15328 713 15334 726
rect 15358 724 15364 729
rect 15437 726 15448 729
rect 15625 726 15631 733
rect 15427 722 15429 723
rect 15448 722 15459 726
rect 15624 723 15631 726
rect 15459 721 15461 722
rect 15461 720 15465 721
rect 14809 707 14810 708
rect 15031 707 15032 708
rect 15144 701 15156 709
rect 15166 701 15178 709
rect 15236 705 15242 710
rect 15326 708 15328 713
rect 15325 707 15326 708
rect 15242 703 15253 705
rect 14870 697 15004 700
rect 15170 698 15174 701
rect 15253 699 15266 703
rect 15266 698 15271 699
rect 14746 695 14870 697
rect 15004 695 15010 697
rect 14649 692 14655 694
rect 14724 692 14746 695
rect 15010 692 15016 695
rect 14431 688 14432 690
rect 14645 688 14647 691
rect 14648 688 14649 690
rect 14701 689 14724 692
rect 15016 689 15022 692
rect 15154 690 15170 698
rect 15271 694 15287 698
rect 15287 692 15303 694
rect 15303 691 15312 692
rect 15318 691 15325 706
rect 15419 693 15427 698
rect 15431 693 15433 720
rect 15619 711 15631 723
rect 15670 711 15672 726
rect 15708 723 15738 750
rect 15764 749 15765 751
rect 15808 750 15810 751
rect 15748 746 15750 747
rect 15762 745 15764 749
rect 15751 737 15765 745
rect 15793 744 15795 749
rect 15813 747 15816 749
rect 15816 746 15818 747
rect 15818 743 15822 746
rect 15842 743 15854 749
rect 15913 744 15916 749
rect 15948 744 15969 778
rect 16035 756 16044 778
rect 16073 776 16078 778
rect 16079 776 16125 779
rect 16218 778 16219 781
rect 16073 775 16125 776
rect 16073 756 16078 775
rect 16219 772 16223 778
rect 16219 756 16226 772
rect 16250 756 16258 789
rect 16268 788 16284 792
rect 16286 788 16302 794
rect 16364 788 16380 795
rect 16478 788 16494 795
rect 16481 787 16482 788
rect 16482 783 16483 785
rect 16484 772 16487 779
rect 16507 778 16519 804
rect 16556 799 16557 802
rect 16556 796 16558 799
rect 16594 796 16596 800
rect 18062 799 18081 804
rect 18092 799 18127 804
rect 18062 797 18092 799
rect 16556 791 16564 796
rect 16591 791 16594 796
rect 16556 788 16572 791
rect 16574 788 16590 791
rect 18111 788 18128 799
rect 18119 786 18128 788
rect 18121 780 18128 786
rect 18186 783 18195 786
rect 18199 785 18201 788
rect 18231 785 18233 788
rect 18244 786 18245 828
rect 18272 820 18277 833
rect 18372 831 18449 833
rect 18269 804 18285 820
rect 18272 789 18277 804
rect 18285 789 18301 803
rect 18344 795 18363 798
rect 18257 787 18282 789
rect 18285 788 18310 789
rect 18257 785 18259 787
rect 18372 786 18430 831
rect 18447 801 18449 831
rect 18453 821 18461 833
rect 18519 822 18535 838
rect 18589 837 18593 840
rect 18613 838 18615 840
rect 18637 838 18643 844
rect 18683 839 18689 844
rect 18679 838 18691 839
rect 18738 838 18741 850
rect 18773 841 18789 854
rect 18844 852 18852 858
rect 18842 850 18852 852
rect 18956 851 18959 860
rect 18905 848 18915 850
rect 18915 846 18921 848
rect 18954 847 18956 851
rect 18832 844 18846 846
rect 18921 844 18928 846
rect 18772 840 18789 841
rect 18772 838 18776 840
rect 18555 829 18567 837
rect 18577 829 18589 837
rect 18615 832 18695 838
rect 18555 828 18556 829
rect 18444 799 18449 801
rect 18450 812 18453 819
rect 18556 818 18558 828
rect 18615 822 18631 832
rect 18637 827 18689 832
rect 18483 812 18519 816
rect 18558 814 18560 818
rect 18450 805 18519 812
rect 18560 809 18561 812
rect 18561 805 18562 809
rect 18199 783 18233 785
rect 18180 782 18208 783
rect 18165 780 18208 782
rect 16030 745 16035 756
rect 16070 744 16073 756
rect 16223 750 16226 756
rect 16223 744 16230 750
rect 16258 744 16260 756
rect 16288 751 16300 759
rect 16310 751 16322 759
rect 16487 755 16492 772
rect 16519 770 16523 778
rect 18121 777 18134 780
rect 18174 777 18180 780
rect 18186 777 18195 780
rect 18197 779 18208 780
rect 18363 780 18430 786
rect 18450 791 18511 805
rect 18519 791 18539 805
rect 18562 799 18563 803
rect 18563 795 18564 799
rect 18637 793 18657 827
rect 18697 815 18703 827
rect 18683 793 18691 795
rect 18697 793 18703 805
rect 18719 804 18727 820
rect 18742 814 18745 829
rect 18757 822 18776 838
rect 18810 833 18819 842
rect 18832 841 18852 844
rect 18928 843 18932 844
rect 18932 842 18937 843
rect 18953 842 18954 844
rect 18949 841 18960 842
rect 18985 841 18995 869
rect 19000 866 19001 869
rect 19001 854 19004 865
rect 19072 860 19077 870
rect 19248 869 19251 870
rect 19247 865 19251 869
rect 19248 860 19251 865
rect 19278 866 19288 870
rect 19508 866 19525 872
rect 19544 871 19548 890
rect 19591 888 19595 896
rect 19699 890 19702 896
rect 19708 891 19719 908
rect 19774 903 19786 909
rect 19886 908 19887 909
rect 19815 903 19831 908
rect 19885 903 19886 908
rect 19932 903 19939 910
rect 19786 902 19815 903
rect 19884 896 19885 899
rect 19767 890 19773 896
rect 19825 890 19831 896
rect 19595 874 19603 888
rect 19697 885 19699 889
rect 19705 886 19708 890
rect 19077 854 19078 860
rect 19247 854 19250 860
rect 19001 852 19007 854
rect 19004 841 19007 852
rect 19069 849 19085 854
rect 19068 848 19082 849
rect 19087 848 19103 854
rect 19060 841 19068 848
rect 19082 842 19105 848
rect 18832 838 18846 841
rect 18952 839 18953 841
rect 18960 840 18995 841
rect 19006 840 19007 841
rect 19058 840 19060 841
rect 18985 839 19033 840
rect 19056 838 19058 840
rect 19072 839 19084 842
rect 19165 841 19181 854
rect 19183 841 19199 854
rect 19245 847 19247 853
rect 19248 852 19250 854
rect 19278 852 19296 866
rect 19519 863 19534 866
rect 19105 840 19106 841
rect 19158 840 19159 841
rect 19077 838 19084 839
rect 18826 834 18840 838
rect 18826 833 18837 834
rect 18801 824 18810 833
rect 18772 820 18776 822
rect 18757 814 18776 820
rect 18745 809 18746 812
rect 18746 799 18748 808
rect 18757 804 18773 814
rect 18832 812 18840 824
rect 18844 814 18846 838
rect 18949 832 18952 838
rect 18904 815 18910 821
rect 18938 818 18956 832
rect 18944 815 18945 818
rect 18898 814 18904 815
rect 18943 814 18944 815
rect 18844 812 18878 814
rect 18887 812 18946 814
rect 18956 813 18962 818
rect 18957 812 18963 813
rect 18776 808 18777 812
rect 18868 809 18878 812
rect 18882 810 18887 812
rect 18859 808 18868 809
rect 18871 808 18877 809
rect 18879 808 18882 810
rect 18898 809 18904 812
rect 18777 804 18778 808
rect 18844 805 18856 808
rect 18859 805 18878 808
rect 18844 804 18857 805
rect 18773 794 18781 804
rect 18804 800 18856 804
rect 18866 800 18878 805
rect 18934 800 18943 811
rect 18946 810 18954 812
rect 18957 810 18968 812
rect 18976 811 18985 838
rect 19007 822 19023 838
rect 19047 832 19055 838
rect 18954 809 18968 810
rect 18970 809 18976 810
rect 18954 808 18976 809
rect 19007 808 19023 820
rect 19076 811 19078 838
rect 19079 837 19084 838
rect 19081 836 19084 837
rect 19106 838 19107 840
rect 19157 838 19158 840
rect 19082 834 19086 836
rect 19087 832 19088 834
rect 19106 832 19119 838
rect 19080 828 19084 830
rect 18957 804 19023 808
rect 18966 800 19007 804
rect 19047 801 19048 804
rect 18773 793 18783 794
rect 18564 792 18565 793
rect 18637 792 18689 793
rect 18695 792 18711 793
rect 18773 792 18785 793
rect 18450 784 18479 791
rect 18565 789 18571 792
rect 18571 784 18578 789
rect 18631 788 18711 792
rect 18749 790 18750 792
rect 18773 789 18794 792
rect 18773 788 18788 789
rect 18631 786 18695 788
rect 18783 786 18788 788
rect 18794 787 18799 789
rect 18799 786 18803 787
rect 18804 786 18855 800
rect 18867 793 18871 800
rect 18929 793 18934 799
rect 18866 790 18867 793
rect 18927 790 18929 793
rect 18578 783 18579 784
rect 18614 783 18615 785
rect 18363 777 18439 780
rect 18580 779 18586 783
rect 18611 779 18614 783
rect 18637 780 18643 786
rect 18679 781 18691 786
rect 18799 785 18810 786
rect 18801 783 18810 785
rect 18801 782 18813 783
rect 18683 780 18689 781
rect 18749 779 18750 781
rect 18586 777 18591 779
rect 18610 777 18611 779
rect 18748 777 18749 779
rect 18801 777 18810 782
rect 18816 779 18819 781
rect 18819 777 18838 779
rect 18866 777 18875 786
rect 18897 782 18903 788
rect 18924 786 18927 790
rect 18943 782 18949 788
rect 18961 786 18970 800
rect 18973 788 18989 800
rect 18991 796 19027 800
rect 19048 798 19050 801
rect 19075 800 19076 810
rect 19082 798 19084 828
rect 19088 818 19096 830
rect 19105 822 19119 832
rect 19149 836 19157 838
rect 19211 837 19215 841
rect 19243 839 19245 847
rect 19278 838 19288 852
rect 19296 848 19299 852
rect 19426 842 19432 844
rect 19426 838 19440 842
rect 19472 838 19478 844
rect 19479 838 19495 854
rect 19519 838 19525 863
rect 19534 853 19537 863
rect 19537 838 19542 852
rect 19149 822 19156 836
rect 19173 826 19185 832
rect 19170 825 19229 826
rect 19233 825 19243 838
rect 19170 823 19178 825
rect 19229 823 19243 825
rect 19250 823 19253 838
rect 19105 820 19108 822
rect 19169 821 19170 823
rect 19048 796 19084 798
rect 19088 796 19096 808
rect 19105 804 19119 820
rect 19161 816 19169 820
rect 19173 818 19180 820
rect 19161 808 19167 816
rect 19173 814 19174 818
rect 19233 816 19258 823
rect 19267 816 19278 837
rect 19299 822 19311 838
rect 19420 832 19426 838
rect 19424 830 19426 832
rect 19428 830 19461 838
rect 19478 832 19484 838
rect 19495 832 19511 838
rect 19525 832 19526 838
rect 19478 830 19511 832
rect 19542 830 19545 838
rect 19548 830 19560 870
rect 19603 863 19608 874
rect 19650 871 19653 885
rect 19687 881 19697 885
rect 19773 884 19779 890
rect 19783 887 19784 890
rect 19793 886 19800 890
rect 19784 883 19787 885
rect 19790 884 19792 885
rect 19819 884 19825 890
rect 19882 888 19884 896
rect 19784 882 19789 883
rect 19685 874 19703 881
rect 19668 870 19685 874
rect 19687 870 19697 874
rect 19608 859 19610 863
rect 19634 838 19650 870
rect 19668 866 19687 870
rect 19666 863 19668 866
rect 19664 859 19666 863
rect 19680 859 19687 866
rect 19662 856 19664 859
rect 19660 854 19662 856
rect 19653 851 19662 854
rect 19653 839 19660 851
rect 19653 838 19654 839
rect 19610 830 19611 838
rect 19634 830 19653 838
rect 19667 830 19680 859
rect 19697 846 19704 858
rect 19709 848 19710 880
rect 19776 876 19782 879
rect 19773 874 19776 876
rect 19764 869 19773 874
rect 19784 870 19787 882
rect 19821 870 19824 884
rect 19881 881 19882 888
rect 19880 874 19881 881
rect 19757 860 19758 863
rect 19787 860 19789 870
rect 19821 862 19835 870
rect 19877 863 19880 874
rect 19752 848 19757 860
rect 19709 847 19714 848
rect 19709 846 19743 847
rect 19750 846 19755 848
rect 19704 844 19705 846
rect 19749 844 19750 846
rect 19746 842 19748 843
rect 19709 834 19721 841
rect 19731 834 19743 841
rect 19789 830 19800 859
rect 19824 830 19835 862
rect 19876 856 19877 859
rect 19914 856 19932 903
rect 20020 890 20028 902
rect 20032 890 20034 921
rect 20065 920 20066 922
rect 20072 912 20078 924
rect 20128 913 20130 925
rect 20159 924 20175 928
rect 20245 925 20254 934
rect 20237 924 20245 925
rect 20159 913 20237 924
rect 20072 911 20075 912
rect 20075 903 20080 910
rect 20113 905 20175 913
rect 20107 903 20113 905
rect 20066 890 20107 903
rect 20075 888 20080 890
rect 20130 889 20132 905
rect 20028 886 20031 888
rect 20080 886 20081 888
rect 20132 885 20133 888
rect 20031 884 20033 885
rect 20032 883 20034 884
rect 20032 879 20035 883
rect 20081 880 20082 882
rect 20032 878 20036 879
rect 20035 876 20036 878
rect 20082 876 20083 880
rect 20133 876 20134 879
rect 20159 878 20175 905
rect 20036 869 20039 874
rect 20039 863 20041 869
rect 19974 861 19975 862
rect 20041 860 20042 863
rect 19853 851 19869 854
rect 19873 851 19876 856
rect 19912 851 19914 856
rect 19955 854 19967 855
rect 19853 843 19873 851
rect 19909 843 19912 851
rect 19949 849 19967 854
rect 19977 849 19989 855
rect 19949 843 20040 849
rect 20042 848 20046 860
rect 20046 844 20047 847
rect 20063 843 20079 854
rect 19851 839 19854 843
rect 19907 839 19909 843
rect 19943 842 19948 843
rect 19943 840 19947 842
rect 19949 841 19989 843
rect 19936 839 19946 840
rect 19949 839 19955 841
rect 19930 838 19935 839
rect 19949 838 19950 839
rect 19837 830 19851 838
rect 19904 836 19907 838
rect 19926 837 19930 838
rect 19917 836 19923 837
rect 19904 834 19917 836
rect 19894 833 19898 834
rect 19888 832 19894 833
rect 19875 830 19888 832
rect 19904 831 19907 834
rect 19416 827 19424 830
rect 19428 828 19431 830
rect 19415 821 19425 827
rect 19104 802 19105 804
rect 19106 800 19108 804
rect 19233 801 19243 816
rect 19245 812 19253 816
rect 19245 804 19254 812
rect 19258 807 19290 816
rect 19299 807 19311 820
rect 19391 807 19415 821
rect 19416 818 19424 821
rect 19254 801 19255 803
rect 19267 801 19278 807
rect 19290 804 19311 807
rect 18991 788 19007 796
rect 19027 795 19032 796
rect 19032 793 19043 795
rect 19050 794 19057 796
rect 19057 793 19063 794
rect 19074 793 19075 796
rect 19043 792 19048 793
rect 19063 792 19083 793
rect 19086 792 19088 795
rect 19103 794 19104 796
rect 19063 786 19084 792
rect 19100 789 19103 793
rect 19085 788 19103 789
rect 19085 786 19100 788
rect 19156 786 19157 788
rect 19161 786 19167 798
rect 19215 789 19216 801
rect 19230 790 19233 800
rect 19255 797 19283 801
rect 19290 797 19309 804
rect 19379 800 19391 807
rect 19377 799 19379 800
rect 19255 796 19309 797
rect 19370 796 19377 799
rect 19416 796 19424 808
rect 19428 796 19430 828
rect 19496 822 19725 830
rect 19496 820 19498 822
rect 19499 820 19725 822
rect 19496 814 19725 820
rect 19753 814 19875 830
rect 19898 818 19904 831
rect 19933 822 19949 838
rect 19896 815 19903 818
rect 19496 812 19753 814
rect 19498 804 19511 812
rect 19528 807 19530 812
rect 19498 803 19499 804
rect 19499 801 19500 802
rect 19496 796 19499 801
rect 19529 800 19530 807
rect 19541 804 19553 812
rect 19553 803 19554 804
rect 19558 803 19560 808
rect 19577 803 19656 812
rect 19554 802 19656 803
rect 19557 799 19573 802
rect 19174 787 19175 788
rect 19173 786 19179 787
rect 18955 782 18961 786
rect 19072 784 19084 786
rect 16270 747 16276 750
rect 16324 749 16326 750
rect 16279 747 16283 749
rect 16270 746 16279 747
rect 16269 744 16277 746
rect 16288 745 16324 747
rect 16326 745 16334 747
rect 15791 738 15793 743
rect 15822 741 15854 743
rect 15850 740 15855 741
rect 15857 737 15860 739
rect 15910 738 15913 744
rect 15945 739 15948 744
rect 16028 740 16030 744
rect 16045 740 16057 742
rect 15758 734 15759 737
rect 15765 734 15769 737
rect 15757 732 15758 734
rect 15769 732 15773 734
rect 15789 732 15791 737
rect 15819 736 15820 737
rect 15849 734 15859 737
rect 15860 734 15866 737
rect 15872 734 15878 737
rect 15854 732 15859 734
rect 15754 725 15757 731
rect 15773 729 15777 732
rect 15787 729 15789 731
rect 15753 722 15754 724
rect 15749 711 15753 721
rect 15777 712 15805 729
rect 15818 726 15819 731
rect 15859 727 15863 732
rect 15865 731 15878 734
rect 15903 732 15907 734
rect 15901 731 15903 732
rect 15918 731 15924 737
rect 16008 734 16014 740
rect 16026 734 16027 736
rect 16045 734 16060 740
rect 16069 738 16070 742
rect 16218 738 16224 744
rect 16276 738 16282 744
rect 16288 743 16290 745
rect 16068 734 16069 737
rect 15941 732 15942 734
rect 16002 732 16066 734
rect 15863 726 15865 727
rect 15866 726 15872 731
rect 15620 710 15624 711
rect 15625 710 15677 711
rect 15619 706 15683 710
rect 15614 704 15683 706
rect 15746 704 15749 711
rect 15473 698 15479 699
rect 15487 698 15525 699
rect 15467 695 15479 698
rect 15483 695 15531 698
rect 15467 693 15473 695
rect 15483 693 15521 695
rect 15525 693 15531 695
rect 15419 692 15531 693
rect 15419 691 15513 692
rect 15022 688 15025 689
rect 15029 688 15031 690
rect 12965 674 12967 685
rect 12419 656 12425 660
rect 12481 656 12485 669
rect 12697 660 12706 669
rect 12697 658 12707 660
rect 12697 656 12708 658
rect 12765 656 12781 672
rect 12903 665 12912 674
rect 12968 669 12977 674
rect 14432 669 14442 688
rect 14643 682 14649 688
rect 14701 682 14707 688
rect 15025 686 15031 688
rect 14648 680 14661 682
rect 14648 676 14655 680
rect 14695 676 14701 682
rect 15029 677 15031 686
rect 15131 681 15154 690
rect 15312 689 15334 691
rect 15419 689 15509 691
rect 15131 679 15201 681
rect 12967 667 12977 669
rect 12968 665 12977 667
rect 12905 656 12906 658
rect 12912 656 12921 665
rect 12959 656 12973 665
rect 14442 658 14452 669
rect 14444 656 14458 658
rect 14494 656 14510 672
rect 14648 668 14649 676
rect 15025 671 15031 677
rect 15083 678 15154 679
rect 15083 676 15147 678
rect 15201 676 15210 679
rect 15083 671 15089 676
rect 14648 656 14660 668
rect 15028 665 15037 671
rect 15077 665 15083 671
rect 15028 662 15031 665
rect 15112 662 15131 676
rect 15210 675 15214 676
rect 15214 672 15216 675
rect 15218 667 15219 669
rect 15028 658 15030 662
rect 15108 659 15112 662
rect 15219 660 15234 667
rect 15318 662 15324 689
rect 15334 686 15369 689
rect 15419 686 15503 689
rect 15519 686 15525 692
rect 15614 690 15619 704
rect 15625 699 15643 704
rect 15625 698 15631 699
rect 15671 698 15677 704
rect 15744 699 15746 704
rect 15672 696 15673 698
rect 15742 695 15744 698
rect 15778 695 15786 712
rect 15806 709 15809 711
rect 15814 709 15818 726
rect 15865 717 15875 726
rect 15924 725 15930 731
rect 15937 725 15941 732
rect 16002 730 16060 732
rect 16061 730 16066 732
rect 16067 730 16068 732
rect 16002 728 16058 730
rect 15935 722 15936 724
rect 15875 709 15877 717
rect 15929 711 15935 721
rect 15809 708 15811 709
rect 15808 707 15812 708
rect 15808 703 15814 707
rect 15820 705 15821 707
rect 15820 703 15837 705
rect 15739 694 15742 695
rect 15735 692 15739 694
rect 15733 691 15735 692
rect 15369 684 15388 686
rect 15427 684 15491 686
rect 15388 683 15396 684
rect 15396 681 15417 683
rect 15427 681 15486 684
rect 15417 679 15486 681
rect 15610 679 15614 689
rect 15673 686 15675 690
rect 15729 689 15733 691
rect 15725 688 15729 689
rect 15775 688 15778 695
rect 15811 690 15814 703
rect 15817 699 15819 700
rect 15820 696 15844 699
rect 15820 691 15832 696
rect 15844 693 15858 696
rect 15877 693 15879 706
rect 15924 702 15929 711
rect 16008 696 16023 728
rect 16055 726 16058 728
rect 16061 726 16069 730
rect 16055 724 16057 726
rect 16056 700 16057 724
rect 16058 718 16069 726
rect 16058 714 16062 718
rect 16058 710 16061 714
rect 16064 712 16066 718
rect 16320 715 16322 745
rect 16324 742 16334 745
rect 16494 743 16496 749
rect 16504 743 16510 749
rect 16523 746 16546 770
rect 18008 755 18009 777
rect 18037 772 18038 777
rect 18128 774 18167 777
rect 18174 774 18186 777
rect 18038 759 18046 772
rect 18130 768 18167 774
rect 18177 768 18186 774
rect 18243 768 18244 777
rect 18038 755 18049 759
rect 18009 749 18010 755
rect 18046 753 18049 755
rect 18047 750 18052 753
rect 16550 743 16556 749
rect 18021 747 18050 748
rect 18053 747 18054 749
rect 16498 742 16504 743
rect 16326 738 16334 742
rect 16326 735 16344 738
rect 16334 731 16344 735
rect 16496 731 16504 742
rect 16509 738 16510 742
rect 16542 739 16548 742
rect 16507 731 16509 738
rect 16543 737 16548 739
rect 16556 737 16562 743
rect 16294 714 16322 715
rect 16289 713 16322 714
rect 16326 713 16334 725
rect 16344 721 16350 731
rect 16496 721 16507 731
rect 16488 720 16507 721
rect 16488 712 16497 720
rect 16063 710 16064 711
rect 16061 707 16065 710
rect 16323 709 16326 711
rect 16297 708 16300 709
rect 16060 702 16065 707
rect 16285 706 16295 708
rect 16276 704 16285 706
rect 16055 696 16057 699
rect 15858 692 15924 693
rect 15864 691 15924 692
rect 15698 686 15725 688
rect 15774 686 15775 688
rect 15673 684 15705 686
rect 15663 683 15705 684
rect 15636 681 15705 683
rect 15618 679 15705 681
rect 15771 679 15774 684
rect 15427 678 15486 679
rect 15430 677 15465 678
rect 15591 677 15705 679
rect 15430 676 15462 677
rect 15464 676 15465 677
rect 15431 674 15443 676
rect 15445 675 15464 676
rect 15569 675 15591 677
rect 15597 676 15705 677
rect 15610 675 15614 676
rect 15445 671 15472 675
rect 15521 671 15569 675
rect 15445 670 15483 671
rect 15510 670 15553 671
rect 15445 664 15553 670
rect 15447 662 15457 664
rect 15610 662 15611 675
rect 15675 672 15677 675
rect 15768 673 15771 679
rect 15324 660 15325 662
rect 15106 658 15108 659
rect 14808 656 14810 657
rect 15028 656 15029 658
rect 15104 656 15106 658
rect 11839 652 11840 653
rect 12087 652 12088 653
rect 12120 652 12157 654
rect 12225 653 12226 656
rect 12281 653 12282 655
rect 12424 654 12425 656
rect 11213 651 11215 652
rect 11080 649 11156 651
rect 11208 649 11213 651
rect 11448 649 11452 652
rect 11511 650 11513 652
rect 11501 649 11511 650
rect 11163 648 11207 649
rect 11459 640 11475 649
rect 11476 648 11477 649
rect 11741 647 11743 651
rect 11761 647 11873 652
rect 11755 644 11873 647
rect 11971 644 12120 652
rect 11755 640 11771 644
rect 11873 641 11884 644
rect 11924 641 11971 644
rect 11884 640 11924 641
rect 12061 640 12077 644
rect 8869 639 8870 640
rect 12123 636 12153 652
rect 12261 640 12277 653
rect 12424 644 12434 654
rect 12697 652 12710 656
rect 12732 652 12765 656
rect 12965 652 12968 656
rect 12712 651 12731 652
rect 12480 645 12481 651
rect 12435 640 12451 644
rect 12453 640 12469 644
rect 12749 640 12765 652
rect 12906 645 12916 652
rect 12960 646 12965 652
rect 12954 645 12960 646
rect 12916 644 12957 645
rect 12941 640 12957 644
rect 14460 640 14476 656
rect 14478 640 14494 656
rect 14661 653 14663 656
rect 14801 653 14807 656
rect 15030 653 15033 656
rect 15100 653 15104 656
rect 14663 651 14665 653
rect 14800 652 14801 653
rect 15098 652 15100 653
rect 15234 652 15346 660
rect 15438 658 15447 662
rect 15675 659 15678 672
rect 15807 666 15811 689
rect 15870 685 15924 691
rect 16008 688 16060 696
rect 16061 692 16065 702
rect 16218 693 16224 698
rect 16276 693 16282 698
rect 16218 692 16282 693
rect 16065 688 16067 690
rect 15866 679 15930 685
rect 16002 682 16067 688
rect 16224 686 16230 692
rect 16270 686 16276 692
rect 16288 690 16289 706
rect 16310 701 16322 709
rect 16501 707 16507 720
rect 16544 717 16548 737
rect 16500 706 16501 707
rect 16496 697 16500 706
rect 16548 697 16550 717
rect 17311 703 17333 722
rect 18003 713 18010 725
rect 18015 716 18016 747
rect 18044 745 18049 747
rect 18048 716 18049 745
rect 18050 738 18061 747
rect 18277 740 18281 777
rect 18372 768 18381 777
rect 18424 768 18430 777
rect 18586 776 18610 777
rect 18746 772 18748 777
rect 18810 772 18838 777
rect 18739 759 18746 772
rect 18810 768 18819 772
rect 18857 768 18866 777
rect 18891 776 18897 782
rect 18949 776 18961 782
rect 19073 776 19074 781
rect 18949 766 18953 773
rect 19105 772 19106 786
rect 19157 783 19158 786
rect 19168 784 19170 785
rect 19214 784 19215 788
rect 19229 787 19230 790
rect 19255 789 19299 796
rect 19309 795 19311 796
rect 19311 792 19318 795
rect 19368 793 19370 796
rect 19467 795 19495 796
rect 19318 789 19322 792
rect 19255 788 19277 789
rect 19279 788 19295 789
rect 19322 788 19324 789
rect 19364 788 19368 793
rect 19479 792 19495 795
rect 19525 793 19529 799
rect 19236 787 19243 788
rect 19251 787 19265 788
rect 19324 787 19327 788
rect 19228 786 19236 787
rect 19223 785 19236 786
rect 19255 785 19265 787
rect 19420 786 19426 792
rect 19478 791 19495 792
rect 19522 791 19525 793
rect 19478 789 19534 791
rect 19555 789 19573 799
rect 19478 788 19495 789
rect 19522 788 19525 789
rect 19534 788 19573 789
rect 19575 788 19656 802
rect 19667 800 19680 812
rect 19743 804 19744 807
rect 19478 786 19484 788
rect 19521 786 19522 788
rect 19220 784 19229 785
rect 19158 780 19170 783
rect 19173 780 19174 781
rect 19182 780 19220 784
rect 19158 779 19217 780
rect 19173 774 19185 779
rect 19104 763 19106 772
rect 19223 763 19229 784
rect 19255 784 19269 785
rect 18729 756 18746 759
rect 19070 756 19073 763
rect 18729 755 18739 756
rect 18729 754 18736 755
rect 19069 754 19070 756
rect 18729 753 18733 754
rect 18718 749 18760 753
rect 18718 748 18745 749
rect 18716 747 18718 748
rect 18760 747 18763 749
rect 18702 745 18716 747
rect 18234 738 18240 740
rect 18277 739 18286 740
rect 18054 735 18072 738
rect 18061 725 18072 735
rect 18234 734 18246 738
rect 18280 734 18286 739
rect 18669 738 18702 745
rect 18663 737 18668 738
rect 18228 728 18234 734
rect 18286 729 18292 734
rect 18640 733 18663 737
rect 18717 735 18725 747
rect 18729 746 18734 747
rect 18634 731 18640 733
rect 18628 729 18630 731
rect 18250 728 18381 729
rect 18234 726 18250 728
rect 18286 727 18589 728
rect 18616 727 18622 729
rect 18627 728 18628 729
rect 18381 726 18382 727
rect 18589 726 18622 727
rect 18625 726 18627 728
rect 18015 714 18019 716
rect 18046 714 18049 716
rect 18015 713 18049 714
rect 18054 713 18072 725
rect 18222 714 18230 726
rect 18234 724 18240 726
rect 18010 711 18011 713
rect 18011 708 18016 711
rect 18049 708 18054 711
rect 18015 707 18027 708
rect 17282 697 17305 698
rect 17310 697 17333 703
rect 18014 701 18027 707
rect 18037 701 18049 708
rect 18061 707 18072 713
rect 16496 693 16504 697
rect 16556 693 16562 697
rect 18014 694 18016 701
rect 16496 691 16562 693
rect 16496 690 16500 691
rect 16289 686 16291 690
rect 15870 673 15878 679
rect 15918 673 15924 679
rect 16008 676 16014 682
rect 16054 676 16060 682
rect 15870 666 15877 673
rect 16010 672 16013 676
rect 15434 656 15438 658
rect 15611 656 15612 658
rect 15676 657 15678 659
rect 15674 656 15678 657
rect 15429 653 15434 656
rect 15612 653 15615 656
rect 15673 653 15674 656
rect 15708 654 15738 663
rect 15742 654 15755 660
rect 15807 659 15809 666
rect 15870 665 15878 666
rect 15424 652 15425 653
rect 15672 652 15673 653
rect 15705 652 15742 654
rect 15809 653 15811 659
rect 15867 656 15878 665
rect 16004 660 16013 672
rect 16066 672 16067 682
rect 16004 656 16010 660
rect 16066 656 16070 672
rect 16282 660 16291 686
rect 16490 674 16496 690
rect 16504 685 16510 691
rect 16550 685 16556 691
rect 18072 690 18079 707
rect 18222 692 18230 704
rect 18234 694 18236 724
rect 18383 719 18387 726
rect 18589 723 18624 726
rect 18662 723 18668 729
rect 18387 708 18394 719
rect 18610 717 18616 723
rect 18617 719 18624 723
rect 18668 719 18674 723
rect 18717 719 18725 725
rect 18729 719 18731 746
rect 19058 744 19064 750
rect 19066 744 19069 754
rect 19104 750 19105 763
rect 19210 757 19216 762
rect 19222 757 19223 762
rect 19255 758 19265 784
rect 19269 783 19273 784
rect 19328 783 19334 786
rect 19363 783 19364 786
rect 19426 784 19440 786
rect 19426 783 19432 784
rect 19464 783 19468 784
rect 19335 781 19337 782
rect 19337 780 19340 781
rect 19353 780 19363 783
rect 19282 775 19288 779
rect 19288 772 19293 775
rect 19340 772 19363 780
rect 19294 766 19318 772
rect 19353 769 19385 772
rect 19391 769 19464 783
rect 19472 780 19478 786
rect 19479 784 19480 785
rect 19520 784 19521 786
rect 19555 783 19558 788
rect 19564 787 19656 788
rect 19628 786 19656 787
rect 19605 785 19656 786
rect 19664 785 19667 799
rect 19742 797 19743 801
rect 19789 800 19800 814
rect 19824 804 19835 814
rect 19837 804 19853 814
rect 19890 807 19903 815
rect 19887 805 19903 807
rect 19933 805 19949 820
rect 19987 811 19989 841
rect 19993 831 20001 843
rect 20040 838 20080 843
rect 20083 842 20090 874
rect 20125 840 20133 852
rect 20137 842 20139 874
rect 20169 857 20174 874
rect 20169 842 20171 857
rect 20174 852 20175 856
rect 20137 840 20171 842
rect 20175 840 20183 852
rect 20090 838 20091 840
rect 20177 838 20179 840
rect 20080 837 20095 838
rect 20137 837 20138 838
rect 20089 836 20095 837
rect 20134 836 20136 837
rect 19971 809 19989 811
rect 19993 809 20001 821
rect 20050 805 20060 836
rect 20089 832 20104 836
rect 20092 808 20104 832
rect 20137 828 20149 836
rect 20159 828 20171 836
rect 20177 828 20191 838
rect 20138 820 20140 828
rect 20091 807 20104 808
rect 19876 804 19989 805
rect 19853 803 19989 804
rect 19741 791 19742 796
rect 19740 788 19741 791
rect 19800 789 19803 799
rect 19835 794 19843 800
rect 19853 795 19869 803
rect 19871 799 19989 803
rect 20060 801 20064 805
rect 20090 804 20104 807
rect 20125 815 20140 820
rect 20179 822 20191 828
rect 20179 820 20181 822
rect 20125 804 20141 815
rect 20179 805 20191 820
rect 20631 819 20632 1015
rect 20821 819 20822 1015
rect 20907 819 20908 1015
rect 21180 819 21181 1015
rect 21377 819 21378 1015
rect 20181 804 20191 805
rect 20089 803 20090 804
rect 20088 801 20089 802
rect 20036 799 20079 801
rect 19871 796 20036 799
rect 19871 795 19977 796
rect 20060 795 20079 799
rect 19853 794 19887 795
rect 19835 792 19869 794
rect 19814 789 19843 792
rect 19729 785 19740 788
rect 19789 787 19814 789
rect 19776 786 19789 787
rect 19772 785 19776 786
rect 19631 784 19634 785
rect 19652 784 19740 785
rect 19652 783 19729 784
rect 19745 783 19772 785
rect 19800 784 19803 787
rect 19474 779 19475 780
rect 19512 769 19520 783
rect 19554 778 19555 783
rect 19630 781 19631 783
rect 19653 782 19655 783
rect 19629 778 19630 781
rect 19655 780 19658 782
rect 19663 781 19664 783
rect 19721 782 19745 783
rect 19710 779 19721 782
rect 19658 778 19661 779
rect 19210 756 19228 757
rect 19256 756 19262 758
rect 19204 750 19268 756
rect 19293 753 19323 766
rect 19353 763 19391 769
rect 19509 763 19512 769
rect 19353 759 19385 763
rect 19352 756 19353 758
rect 19293 750 19329 753
rect 19350 752 19352 756
rect 19354 755 19385 759
rect 19382 754 19384 755
rect 19385 754 19388 755
rect 19504 754 19509 763
rect 19381 752 19382 754
rect 19388 751 19393 754
rect 19503 752 19504 754
rect 19104 744 19110 750
rect 19210 745 19262 750
rect 19014 742 19058 744
rect 18863 741 18897 742
rect 19014 741 19020 742
rect 18826 740 18863 741
rect 18803 739 18826 740
rect 18800 737 18803 739
rect 19052 738 19058 742
rect 19110 738 19116 744
rect 18775 723 18800 737
rect 18891 730 18897 736
rect 18949 731 18955 736
rect 19204 733 19216 745
rect 19250 735 19255 745
rect 18980 731 19016 733
rect 18897 724 18903 730
rect 18921 729 18980 731
rect 19016 729 19022 731
rect 18919 726 18921 729
rect 18770 720 18775 723
rect 18668 717 18750 719
rect 18671 716 18750 717
rect 18767 716 18775 720
rect 18717 713 18725 716
rect 18729 715 18731 716
rect 18750 715 18779 716
rect 18729 713 18763 715
rect 18760 709 18763 713
rect 18767 713 18775 715
rect 18779 714 18807 715
rect 18767 711 18770 713
rect 18764 709 18767 711
rect 18807 710 18821 714
rect 18913 713 18919 726
rect 18943 724 18949 729
rect 19022 726 19033 729
rect 19210 726 19216 733
rect 19012 722 19014 723
rect 19033 722 19044 726
rect 19209 723 19216 726
rect 19044 721 19046 722
rect 19046 720 19050 721
rect 18394 707 18395 708
rect 18616 707 18617 708
rect 18729 701 18741 709
rect 18751 701 18763 709
rect 18821 705 18827 710
rect 18911 708 18913 713
rect 18910 707 18911 708
rect 18827 703 18838 705
rect 18455 697 18589 700
rect 18755 698 18759 701
rect 18838 699 18851 703
rect 18851 698 18856 699
rect 18331 695 18455 697
rect 18589 695 18595 697
rect 18234 692 18240 694
rect 18309 692 18331 695
rect 18595 692 18601 695
rect 18016 688 18017 690
rect 18230 688 18232 691
rect 18233 688 18234 690
rect 18286 689 18309 692
rect 18601 689 18607 692
rect 18739 690 18755 698
rect 18856 694 18872 698
rect 18872 692 18888 694
rect 18888 691 18897 692
rect 18903 691 18910 706
rect 19004 693 19012 698
rect 19016 693 19018 720
rect 19204 711 19216 723
rect 19255 711 19257 726
rect 19293 723 19323 750
rect 19349 749 19350 751
rect 19393 750 19395 751
rect 19333 746 19335 747
rect 19347 745 19349 749
rect 19336 737 19350 745
rect 19378 744 19380 749
rect 19398 747 19401 749
rect 19401 746 19403 747
rect 19403 743 19407 746
rect 19427 743 19439 749
rect 19498 744 19501 749
rect 19533 744 19554 778
rect 19620 756 19629 778
rect 19658 776 19663 778
rect 19664 776 19710 779
rect 19803 778 19804 781
rect 19658 775 19710 776
rect 19658 756 19663 775
rect 19804 772 19808 778
rect 19804 756 19811 772
rect 19835 756 19843 789
rect 19853 788 19869 792
rect 19871 788 19887 794
rect 19949 788 19965 795
rect 20063 788 20079 795
rect 20066 787 20067 788
rect 20067 783 20068 785
rect 20069 772 20072 779
rect 20092 778 20104 804
rect 20141 799 20142 802
rect 20141 796 20143 799
rect 20179 796 20181 800
rect 20141 791 20149 796
rect 20176 791 20179 796
rect 20141 788 20157 791
rect 20160 788 20175 791
rect 19615 745 19620 756
rect 19655 744 19658 756
rect 19808 750 19811 756
rect 19808 744 19815 750
rect 19843 744 19845 756
rect 19873 751 19885 759
rect 19895 751 19907 759
rect 20072 755 20077 772
rect 20104 770 20108 778
rect 19855 747 19861 750
rect 19909 749 19911 750
rect 19864 747 19868 749
rect 19855 746 19864 747
rect 19854 744 19862 746
rect 19873 745 19909 747
rect 19911 745 19919 747
rect 19376 738 19378 743
rect 19407 741 19439 743
rect 19435 740 19440 741
rect 19442 737 19445 739
rect 19495 738 19498 744
rect 19530 739 19533 744
rect 19613 740 19615 744
rect 19630 740 19642 742
rect 19343 734 19344 737
rect 19350 734 19354 737
rect 19342 732 19343 734
rect 19354 732 19358 734
rect 19374 732 19376 737
rect 19404 736 19405 737
rect 19434 734 19444 737
rect 19445 734 19451 737
rect 19457 734 19463 737
rect 19439 732 19444 734
rect 19339 725 19342 731
rect 19358 729 19362 732
rect 19372 729 19374 731
rect 19338 722 19339 724
rect 19334 711 19338 721
rect 19362 712 19390 729
rect 19403 726 19404 731
rect 19444 727 19448 732
rect 19450 731 19463 734
rect 19488 732 19492 734
rect 19486 731 19488 732
rect 19503 731 19509 737
rect 19593 734 19599 740
rect 19611 734 19612 736
rect 19630 734 19645 740
rect 19654 738 19655 742
rect 19803 738 19809 744
rect 19861 738 19867 744
rect 19873 743 19875 745
rect 19653 734 19654 737
rect 19526 732 19527 734
rect 19587 732 19651 734
rect 19448 726 19450 727
rect 19451 726 19457 731
rect 19205 710 19209 711
rect 19210 710 19262 711
rect 19204 706 19268 710
rect 19199 704 19268 706
rect 19331 704 19334 711
rect 19058 698 19064 699
rect 19072 698 19110 699
rect 19052 695 19064 698
rect 19068 695 19116 698
rect 19052 693 19058 695
rect 19068 693 19106 695
rect 19110 693 19116 695
rect 19004 692 19116 693
rect 19004 691 19098 692
rect 18607 688 18610 689
rect 18614 688 18616 690
rect 16550 674 16553 685
rect 15866 653 15867 655
rect 16009 654 16010 656
rect 14798 651 14800 652
rect 14665 649 14741 651
rect 14793 649 14798 651
rect 15033 649 15037 652
rect 15096 650 15098 652
rect 15086 649 15096 650
rect 14748 648 14792 649
rect 15044 640 15060 649
rect 15061 648 15062 649
rect 15326 647 15328 651
rect 15346 647 15458 652
rect 15340 644 15458 647
rect 15556 644 15705 652
rect 15340 640 15356 644
rect 15458 641 15469 644
rect 15509 641 15556 644
rect 15469 640 15509 641
rect 15646 640 15662 644
rect 12454 639 12455 640
rect 15708 636 15738 652
rect 15846 640 15862 653
rect 16009 644 16019 654
rect 16282 652 16295 660
rect 16350 656 16366 672
rect 16488 665 16497 674
rect 16550 667 16562 674
rect 18017 669 18027 688
rect 18228 682 18234 688
rect 18286 682 18292 688
rect 18610 686 18616 688
rect 18233 680 18246 682
rect 18233 676 18240 680
rect 18280 676 18286 682
rect 18614 677 18616 686
rect 18716 681 18739 690
rect 18897 689 18919 691
rect 19004 689 19094 691
rect 18716 679 18786 681
rect 16553 665 16562 667
rect 16490 656 16491 665
rect 16497 656 16506 665
rect 16544 656 16558 665
rect 18027 658 18037 669
rect 18029 656 18043 658
rect 18079 656 18095 672
rect 18233 668 18234 676
rect 18610 671 18616 677
rect 18668 678 18739 679
rect 18668 676 18732 678
rect 18786 676 18795 679
rect 18668 671 18674 676
rect 18233 656 18245 668
rect 18613 665 18622 671
rect 18662 665 18668 671
rect 18613 662 18616 665
rect 18697 662 18716 676
rect 18795 675 18799 676
rect 18799 672 18801 675
rect 18803 667 18804 669
rect 18613 658 18615 662
rect 18693 659 18697 662
rect 18804 660 18819 667
rect 18903 662 18909 689
rect 18919 686 18954 689
rect 19004 686 19088 689
rect 19104 686 19110 692
rect 19199 690 19204 704
rect 19210 699 19228 704
rect 19210 698 19216 699
rect 19256 698 19262 704
rect 19329 699 19331 704
rect 19257 696 19258 698
rect 19327 695 19329 698
rect 19363 695 19371 712
rect 19391 709 19394 711
rect 19399 709 19403 726
rect 19450 717 19460 726
rect 19509 725 19515 731
rect 19522 725 19526 732
rect 19587 730 19645 732
rect 19646 730 19651 732
rect 19652 730 19653 732
rect 19587 728 19643 730
rect 19520 722 19521 724
rect 19460 709 19462 717
rect 19514 711 19520 721
rect 19394 708 19396 709
rect 19393 707 19397 708
rect 19393 703 19399 707
rect 19405 705 19406 707
rect 19405 703 19422 705
rect 19324 694 19327 695
rect 19320 692 19324 694
rect 19318 691 19320 692
rect 18954 684 18973 686
rect 19012 684 19076 686
rect 18973 683 18981 684
rect 18981 681 19002 683
rect 19012 681 19071 684
rect 19002 679 19071 681
rect 19195 679 19199 689
rect 19258 686 19260 690
rect 19314 689 19318 691
rect 19310 688 19314 689
rect 19360 688 19363 695
rect 19396 690 19399 703
rect 19402 699 19404 700
rect 19405 696 19429 699
rect 19405 691 19417 696
rect 19429 693 19443 696
rect 19462 693 19464 706
rect 19509 702 19514 711
rect 19593 696 19608 728
rect 19640 726 19643 728
rect 19646 726 19654 730
rect 19640 724 19642 726
rect 19641 700 19642 724
rect 19643 718 19654 726
rect 19643 714 19647 718
rect 19643 710 19646 714
rect 19649 712 19651 718
rect 19905 715 19907 745
rect 19909 742 19919 745
rect 20079 743 20081 749
rect 20089 743 20095 749
rect 20108 746 20131 770
rect 20135 743 20141 749
rect 20083 742 20089 743
rect 19911 738 19919 742
rect 19911 735 19929 738
rect 19919 731 19929 735
rect 20081 731 20089 742
rect 20094 738 20095 742
rect 20127 739 20133 742
rect 20092 731 20094 738
rect 20128 737 20133 739
rect 20141 737 20147 743
rect 19879 714 19907 715
rect 19874 713 19907 714
rect 19911 713 19919 725
rect 19929 721 19935 731
rect 20081 721 20092 731
rect 20073 720 20092 721
rect 20073 712 20082 720
rect 19648 710 19649 711
rect 19646 707 19650 710
rect 19908 709 19911 711
rect 19882 708 19885 709
rect 19645 702 19650 707
rect 19870 706 19880 708
rect 19861 704 19870 706
rect 19640 696 19642 699
rect 19443 692 19509 693
rect 19449 691 19509 692
rect 19283 686 19310 688
rect 19359 686 19360 688
rect 19258 684 19290 686
rect 19248 683 19290 684
rect 19221 681 19290 683
rect 19203 679 19290 681
rect 19356 679 19359 684
rect 19012 678 19071 679
rect 19015 677 19050 678
rect 19176 677 19290 679
rect 19015 676 19047 677
rect 19049 676 19050 677
rect 19016 674 19028 676
rect 19030 675 19049 676
rect 19154 675 19176 677
rect 19182 676 19290 677
rect 19195 675 19199 676
rect 19030 671 19057 675
rect 19106 671 19154 675
rect 19030 670 19068 671
rect 19095 670 19138 671
rect 19030 664 19138 670
rect 19032 662 19042 664
rect 19195 662 19196 675
rect 19260 672 19262 675
rect 19353 673 19356 679
rect 18909 660 18910 662
rect 18691 658 18693 659
rect 18393 656 18395 657
rect 18613 656 18614 658
rect 18689 656 18691 658
rect 16317 652 16350 656
rect 16550 652 16553 656
rect 16297 651 16316 652
rect 16065 645 16066 651
rect 16020 640 16036 644
rect 16038 640 16054 644
rect 16334 640 16350 652
rect 16491 645 16501 652
rect 16545 646 16550 652
rect 16539 645 16545 646
rect 16501 644 16542 645
rect 16526 640 16542 644
rect 18045 640 18061 656
rect 18063 640 18079 656
rect 18246 653 18248 656
rect 18386 653 18392 656
rect 18615 653 18618 656
rect 18685 653 18689 656
rect 18248 651 18250 653
rect 18385 652 18386 653
rect 18683 652 18685 653
rect 18819 652 18931 660
rect 19023 658 19032 662
rect 19260 659 19263 672
rect 19392 666 19396 689
rect 19455 685 19509 691
rect 19593 688 19645 696
rect 19646 692 19650 702
rect 19803 693 19809 698
rect 19861 693 19867 698
rect 19803 692 19867 693
rect 19650 688 19652 690
rect 19451 679 19515 685
rect 19587 682 19652 688
rect 19809 686 19815 692
rect 19855 686 19861 692
rect 19873 690 19874 706
rect 19895 701 19907 709
rect 20086 707 20092 720
rect 20129 717 20133 737
rect 20085 706 20086 707
rect 20081 697 20085 706
rect 20133 697 20135 717
rect 20896 703 20918 722
rect 20867 697 20890 698
rect 20895 697 20918 703
rect 20081 693 20089 697
rect 20141 693 20147 697
rect 20081 691 20147 693
rect 20081 690 20085 691
rect 19874 686 19876 690
rect 19455 673 19463 679
rect 19503 673 19509 679
rect 19593 676 19599 682
rect 19639 676 19645 682
rect 19455 666 19462 673
rect 19595 672 19598 676
rect 19019 656 19023 658
rect 19196 656 19197 658
rect 19261 657 19263 659
rect 19259 656 19263 657
rect 19014 653 19019 656
rect 19197 653 19200 656
rect 19258 653 19259 656
rect 19293 654 19323 663
rect 19327 654 19340 660
rect 19392 659 19394 666
rect 19455 665 19463 666
rect 19009 652 19010 653
rect 19257 652 19258 653
rect 19290 652 19327 654
rect 19394 653 19396 659
rect 19452 656 19463 665
rect 19589 660 19598 672
rect 19651 672 19652 682
rect 19589 656 19595 660
rect 19651 656 19655 672
rect 19867 660 19876 686
rect 20075 674 20081 690
rect 20089 685 20095 691
rect 20135 685 20141 691
rect 20135 674 20138 685
rect 19451 653 19452 655
rect 19594 654 19595 656
rect 18383 651 18385 652
rect 18250 649 18326 651
rect 18378 649 18383 651
rect 18618 649 18622 652
rect 18681 650 18683 652
rect 18671 649 18681 650
rect 18333 648 18377 649
rect 18629 640 18645 649
rect 18646 648 18647 649
rect 18911 647 18913 651
rect 18931 647 19043 652
rect 18925 644 19043 647
rect 19141 644 19290 652
rect 18925 640 18941 644
rect 19043 641 19054 644
rect 19094 641 19141 644
rect 19054 640 19094 641
rect 19231 640 19247 644
rect 16039 639 16040 640
rect 19293 636 19323 652
rect 19431 640 19447 653
rect 19594 644 19604 654
rect 19867 652 19880 660
rect 19935 656 19951 672
rect 20073 665 20082 674
rect 20135 667 20147 674
rect 20138 665 20147 667
rect 20075 656 20076 665
rect 20082 656 20091 665
rect 20129 656 20143 665
rect 19902 652 19935 656
rect 20135 652 20138 656
rect 19882 651 19901 652
rect 19650 645 19651 651
rect 19605 640 19621 644
rect 19623 640 19639 644
rect 19919 640 19935 652
rect 20076 645 20086 652
rect 20130 646 20135 652
rect 20124 645 20130 646
rect 20086 644 20127 645
rect 20111 640 20127 644
rect 19624 639 19625 640
rect 6500 623 6527 629
rect 6528 623 6555 624
rect 10085 623 10112 629
rect 10113 623 10140 624
rect 13670 623 13697 629
rect 13698 623 13725 624
rect 17255 623 17282 629
rect 17283 623 17310 624
rect 20840 623 20867 629
rect 20868 623 20895 624
rect 7071 481 7072 487
rect 10656 481 10657 487
rect 14241 481 14242 487
rect 17826 481 17827 487
rect 21411 481 21412 487
rect 7037 441 7072 475
rect 7083 463 7084 475
rect 7083 441 7084 453
rect 10622 441 10657 475
rect 10668 463 10669 475
rect 10668 441 10669 453
rect 14207 441 14242 475
rect 14253 463 14254 475
rect 14253 441 14254 453
rect 17792 441 17827 475
rect 17838 463 17839 475
rect 17838 441 17839 453
rect 21377 441 21412 475
rect 21423 463 21424 475
rect 21423 441 21424 453
rect 6280 429 6281 440
rect 6470 429 6471 440
rect 6556 429 6557 440
rect 6829 429 6830 440
rect 7026 429 7027 440
rect 7060 429 7072 435
rect 9865 429 9866 440
rect 10055 429 10056 440
rect 10141 429 10142 440
rect 10414 429 10415 440
rect 10611 429 10612 440
rect 10645 429 10657 435
rect 13450 429 13451 440
rect 13640 429 13641 440
rect 13726 429 13727 440
rect 13999 429 14000 440
rect 14196 429 14197 440
rect 14230 429 14242 435
rect 17035 429 17036 440
rect 17225 429 17226 440
rect 17311 429 17312 440
rect 17584 429 17585 440
rect 17781 429 17782 440
rect 17815 429 17827 435
rect 20620 429 20621 440
rect 20810 429 20811 440
rect 20896 429 20897 440
rect 21169 429 21170 440
rect 21366 429 21367 440
rect 21400 429 21412 435
rect 6291 389 6292 429
rect 6481 389 6482 429
rect 6567 389 6568 429
rect 6840 389 6841 429
rect 7037 389 7038 429
rect 9876 389 9877 429
rect 10066 389 10067 429
rect 10152 389 10153 429
rect 10425 389 10426 429
rect 10622 389 10623 429
rect 13461 389 13462 429
rect 13651 389 13652 429
rect 13737 389 13738 429
rect 14010 389 14011 429
rect 14207 389 14208 429
rect 17046 389 17047 429
rect 17236 389 17237 429
rect 17322 389 17323 429
rect 17595 389 17596 429
rect 17792 389 17793 429
rect 20631 389 20632 429
rect 20821 389 20822 429
rect 20907 389 20908 429
rect 21180 389 21181 429
rect 21377 389 21378 429
<< nwell >>
rect 3002 1436 6166 1778
rect 8841 1676 8875 1710
rect 12426 1676 12460 1710
rect 16011 1676 16045 1710
rect 19596 1676 19630 1710
rect 3002 1116 21487 1436
rect 3002 1078 6166 1116
rect 3002 850 4489 1078
<< ndiff >>
rect 7038 441 7072 475
rect 10623 441 10657 475
rect 14208 441 14242 475
rect 17793 441 17827 475
rect 21378 441 21412 475
<< pdiff >>
rect 5256 1676 5290 1710
rect 8841 1676 8875 1710
rect 12426 1676 12460 1710
rect 16011 1676 16045 1710
rect 19596 1676 19630 1710
<< locali >>
rect 0 2202 21488 2522
rect 3410 1436 3444 1506
rect 3 1116 21487 1436
rect 4012 487 4041 548
rect 3 0 21487 320
<< metal1 >>
rect 0 2202 21488 2522
rect 21409 2012 21413 2041
rect 21372 2006 21442 2012
rect 3306 1892 3312 1950
rect 3370 1892 3376 1950
rect 21372 1948 21378 2006
rect 21436 1948 21442 2006
rect 21372 1942 21442 1948
rect 7037 1883 7107 1889
rect 5640 1872 5710 1878
rect 5640 1814 5646 1872
rect 5704 1814 5710 1872
rect 7037 1825 7043 1883
rect 7101 1825 7107 1883
rect 10621 1883 10692 1890
rect 7037 1819 7107 1825
rect 9231 1874 9301 1880
rect 5640 1808 5710 1814
rect 9231 1816 9237 1874
rect 9295 1816 9301 1874
rect 10621 1825 10628 1883
rect 10686 1825 10692 1883
rect 14198 1883 14268 1889
rect 10621 1819 10692 1825
rect 12817 1874 12887 1880
rect 9231 1810 9301 1816
rect 12817 1816 12823 1874
rect 12881 1816 12887 1874
rect 14198 1825 14204 1883
rect 14262 1825 14268 1883
rect 17783 1883 17853 1889
rect 14198 1819 14268 1825
rect 16391 1874 16461 1880
rect 12817 1810 12887 1816
rect 16391 1816 16397 1874
rect 16455 1816 16461 1874
rect 17783 1825 17789 1883
rect 17847 1825 17853 1883
rect 17783 1819 17853 1825
rect 20032 1874 20102 1880
rect 16391 1810 16461 1816
rect 20032 1816 20038 1874
rect 20096 1816 20102 1874
rect 20032 1810 20102 1816
rect 3231 1744 3237 1802
rect 3295 1744 3301 1802
rect 3038 1670 3096 1716
rect 5256 1676 5290 1710
rect 8841 1676 8875 1710
rect 12426 1676 12460 1710
rect 16011 1676 16045 1710
rect 19596 1676 19630 1710
rect 3 1116 21487 1436
rect 4012 487 4041 548
rect 7038 441 7072 475
rect 10623 441 10657 475
rect 14208 441 14242 475
rect 17793 441 17827 475
rect 21378 441 21412 475
rect 3 0 21487 320
<< via1 >>
rect 3312 1892 3370 1950
rect 21378 1948 21436 2006
rect 5646 1814 5704 1872
rect 7043 1825 7101 1883
rect 9237 1816 9295 1874
rect 10628 1825 10686 1883
rect 12823 1816 12881 1874
rect 14204 1825 14262 1883
rect 16397 1816 16455 1874
rect 17789 1825 17847 1883
rect 20038 1816 20096 1874
rect 3237 1744 3295 1802
<< metal2 >>
rect 3248 2167 21412 2201
rect 3248 1808 3282 2167
rect 21378 2012 21412 2167
rect 21372 2006 21442 2012
rect 3312 1950 3370 1956
rect 21372 1948 21378 2006
rect 21436 1948 21442 2006
rect 21372 1942 21442 1948
rect 3370 1898 3539 1932
rect 3312 1886 3370 1892
rect 3505 1858 3539 1898
rect 7037 1883 7107 1889
rect 5650 1878 5684 1879
rect 5640 1872 5710 1878
rect 5640 1858 5646 1872
rect 3505 1824 5646 1858
rect 5640 1814 5646 1824
rect 5704 1814 5710 1872
rect 7037 1825 7043 1883
rect 7101 1865 7107 1883
rect 10622 1883 10692 1889
rect 9231 1874 9301 1880
rect 9231 1865 9237 1874
rect 7101 1825 9237 1865
rect 7037 1819 7107 1825
rect 5640 1808 5710 1814
rect 9231 1816 9237 1825
rect 9295 1816 9301 1874
rect 10622 1825 10628 1883
rect 10686 1865 10692 1883
rect 14198 1883 14268 1889
rect 12817 1874 12887 1880
rect 12817 1865 12823 1874
rect 10686 1825 12823 1865
rect 10622 1819 10692 1825
rect 9231 1810 9301 1816
rect 12817 1816 12823 1825
rect 12881 1816 12887 1874
rect 14198 1825 14204 1883
rect 14262 1865 14268 1883
rect 17783 1883 17853 1889
rect 16391 1874 16461 1880
rect 16391 1865 16397 1874
rect 14262 1825 16397 1865
rect 14198 1819 14268 1825
rect 12817 1810 12887 1816
rect 16391 1816 16397 1825
rect 16455 1816 16461 1874
rect 17783 1825 17789 1883
rect 17847 1865 17853 1883
rect 20032 1874 20102 1880
rect 20032 1865 20038 1874
rect 17847 1825 20038 1865
rect 17783 1819 17853 1825
rect 16391 1810 16461 1816
rect 20032 1816 20038 1825
rect 20096 1816 20102 1874
rect 20032 1810 20102 1816
rect 3237 1802 3295 1808
rect 3237 1738 3295 1744
use sky130_osu_sc_12T_hs__mux2_1  sky130_osu_sc_12T_hs__mux2_1_0
timestamp 1698882961
transform 1 0 3013 0 -1 2263
box -8 0 552 902
use sky130_osu_single_mpr2at_8_b0r1  sky130_osu_single_mpr2at_8_b0r1_0
timestamp 1708006426
transform 1 0 17901 0 1 0
box 0 0 3587 2522
use sky130_osu_single_mpr2at_8_b0r1  sky130_osu_single_mpr2at_8_b0r1_1
timestamp 1708006426
transform 1 0 3561 0 1 0
box 0 0 3587 2522
use sky130_osu_single_mpr2at_8_b0r1  sky130_osu_single_mpr2at_8_b0r1_2
timestamp 1708006426
transform 1 0 7146 0 1 0
box 0 0 3587 2522
use sky130_osu_single_mpr2at_8_b0r1  sky130_osu_single_mpr2at_8_b0r1_3
timestamp 1708006426
transform 1 0 10731 0 1 0
box 0 0 3587 2522
use sky130_osu_single_mpr2at_8_b0r1  sky130_osu_single_mpr2at_8_b0r1_4
timestamp 1708006426
transform 1 0 14316 0 1 0
box 0 0 3587 2522
<< labels >>
flabel metal1 s 3038 1670 3096 1716 0 FreeSans 100 0 0 0 start
port 13 nsew signal input
flabel metal1 s 5256 1676 5290 1710 0 FreeSans 100 0 0 0 s1
port 1 nsew signal input
flabel metal1 s 8841 1676 8875 1710 0 FreeSans 100 0 0 0 s2
port 2 nsew signal input
flabel metal1 s 12426 1676 12460 1710 0 FreeSans 100 0 0 0 s3
port 3 nsew signal input
flabel metal1 s 16011 1676 16045 1710 0 FreeSans 100 0 0 0 s4
port 4 nsew signal input
flabel metal1 s 19596 1676 19630 1710 0 FreeSans 100 0 0 0 s5
port 5 nsew signal input
flabel metal1 s 7038 441 7072 475 0 FreeSans 100 0 0 0 X1_Y1
port 6 nsew signal output
flabel metal1 s 10623 441 10657 475 0 FreeSans 100 0 0 0 X2_Y1
port 7 nsew signal output
flabel metal1 s 14208 441 14242 475 0 FreeSans 100 0 0 0 X3_Y1
port 8 nsew signal output
flabel metal1 s 17793 441 17827 475 0 FreeSans 100 0 0 0 X4_Y1
port 9 nsew signal output
flabel metal1 s 21378 441 21412 475 0 FreeSans 100 0 0 0 X5_Y1
port 10 nsew signal output
flabel metal1 s 0 2202 21488 2522 0 FreeSans 100 0 0 0 vssd1
port 14 nsew ground bidirectional
flabel metal1 s 3 1116 21487 1436 0 FreeSans 100 0 0 0 vccd1
port 15 nsew power bidirectional
flabel metal1 s 3 0 21487 320 0 FreeSans 100 0 0 0 vssd1
port 14 nsew ground bidirectional
<< end >>
