magic
tech sky130A
magscale 1 2
timestamp 1713287902
<< nwell >>
rect -9 485 179 897
<< locali >>
rect 0 827 176 888
rect 0 0 176 61
<< metal1 >>
rect 0 827 176 888
rect 0 0 176 61
<< labels >>
rlabel metal1 111 859 111 859 1 vccd1
rlabel metal1 112 28 112 28 1 vssd1
<< end >>
