* NGSPICE file created from user_project_wrapper.ext - technology: sky130A

.subckt sky130_ef_sc_hd__decap_12 VGND VPWR  
X0 VPWR VGND VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1 VGND VPWR VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
.ends

.subckt sky130_fd_sc_hd__decap_4 VGND VPWR  
X0 VPWR VGND VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1 VGND VPWR VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
.ends

.subckt sky130_fd_sc_hd__buf_12   VGND VPWR A X
X0 VGND a_109_47# X sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15 M=12
X1 X a_109_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15 M=12
X2 VPWR A a_109_47# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15 M=4
X3 VGND A a_109_47# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15 M=4
.ends

.subckt sky130_fd_sc_hd__decap_3 VPWR VGND  
X0 VPWR VGND VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1 VGND VPWR VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
.ends

.subckt sky130_fd_sc_hd__decap_6 VPWR VGND  
X0 VPWR VGND VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X1 VGND VPWR VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1    
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2    
.ends

.subckt sky130_fd_sc_hd__decap_8 VPWR VGND  
X0 VPWR VGND VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X1 VGND VPWR VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
.ends

.subckt sky130_fd_sc_hd__a21oi_2   VGND VPWR A2 A1 Y B1
X0 VGND A2 a_285_47# sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.06825 ps=0.86 w=0.65 l=0.15
X1 VGND B1 Y sky130_fd_pr__nfet_01v8 ad=0.26 pd=2.1 as=0.08775 ps=0.92 w=0.65 l=0.15 M=2
X2 Y A1 a_114_47# sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X3 a_114_47# A2 VGND sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.18525 ps=1.87 w=0.65 l=0.15
X4 a_27_297# B1 Y sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.135 ps=1.27 w=1 l=0.15 M=2
X5 a_27_297# A1 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15 M=2
X6 VPWR A2 a_27_297# sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.15 M=2
X7 a_285_47# A1 Y sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.091 ps=0.93 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor2_1   VGND VPWR A B Y
X0 VPWR A a_109_297# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1 VGND A Y sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_109_297# B Y sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3 Y B VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__mux2_1 VGND VPWR   X A1 S A0
X0 VPWR a_505_21# a_535_374# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1 a_505_21# S VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_218_374# S VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X3 VGND a_505_21# a_439_47# sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_76_199# A0 a_218_374# sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X5 a_505_21# S VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X6 a_439_47# A0 a_76_199# sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X7 a_535_374# A1 a_76_199# sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X8 a_76_199# A1 a_218_47# sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X9 a_218_47# S VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X10 VPWR a_76_199# X sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X11 VGND a_76_199# X sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__mux4_1   VGND VPWR A1 A0 S0 A3 A2 S1 X
X0 a_277_47# a_247_21# a_27_413# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 VGND S0 a_247_21# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 a_834_97# a_247_21# a_750_97# sky130_fd_pr__nfet_01v8 ad=0.10795 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 VGND A3 a_668_97# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1079 ps=1.36 w=0.42 l=0.15
X4 a_1290_413# S1 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 a_834_97# A2 VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 a_750_97# S0 a_757_363# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1079 ps=1.36 w=0.42 l=0.15
X7 a_27_47# S0 a_277_47# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.085225 ps=0.925 w=0.42 l=0.15
X8 X a_1478_413# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X9 VPWR A1 a_27_413# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X10 VPWR S0 a_247_21# sky130_fd_pr__pfet_01v8_hvt ad=0.1079 pd=1.36 as=0.1083 ps=1.36 w=0.42 l=0.15
X11 X a_1478_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X12 a_193_47# A0 VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X13 a_750_97# a_1290_413# a_1478_413# sky130_fd_pr__pfet_01v8_hvt ad=0.2688 pd=2.12 as=0.092075 ps=0.99 w=0.42 l=0.15
X14 a_1478_413# S1 a_277_47# sky130_fd_pr__pfet_01v8_hvt ad=0.092075 pd=0.99 as=0.1092 ps=1.36 w=0.42 l=0.15
X15 a_1290_413# S1 VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X16 a_277_47# a_247_21# a_193_47# sky130_fd_pr__nfet_01v8 ad=0.085225 pd=0.925 as=0.0567 ps=0.69 w=0.42 l=0.15
X17 a_750_97# S0 a_668_97# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X18 a_923_363# a_247_21# a_750_97# sky130_fd_pr__pfet_01v8_hvt ad=0.090125 pd=0.995 as=0.0567 ps=0.69 w=0.42 l=0.15
X19 a_757_363# A2 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X20 VPWR A3 a_923_363# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.090125 ps=0.995 w=0.42 l=0.15
X21 a_277_47# a_1290_413# a_1478_413# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.151025 ps=1.285 w=0.42 l=0.15
X22 a_193_413# A0 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X23 a_193_413# S0 a_277_47# sky130_fd_pr__pfet_01v8_hvt ad=0.1079 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X24 VGND A1 a_27_47# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X25 a_1478_413# S1 a_750_97# sky130_fd_pr__nfet_01v8 ad=0.151025 pd=1.285 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a41o_1 VGND VPWR A3 A4 A2 X B1 A1  
X0 a_465_47# A2 a_381_47# sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 VGND A4 a_561_47# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X2 VPWR A3 a_297_297# sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X3 a_297_297# A2 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X4 a_297_297# A4 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X5 VPWR A1 a_297_297# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_381_47# A1 a_79_21# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.183625 ps=1.215 w=0.65 l=0.15
X7 a_297_297# B1 a_79_21# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8 VPWR a_79_21# X sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X9 a_79_21# B1 VGND sky130_fd_pr__nfet_01v8 ad=0.183625 pd=1.215 as=0.160875 ps=1.145 w=0.65 l=0.15
X10 VGND a_79_21# X sky130_fd_pr__nfet_01v8 ad=0.160875 pd=1.145 as=0.169 ps=1.82 w=0.65 l=0.15
X11 a_561_47# A3 a_465_47# sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or3b_1 VGND VPWR   B C_N A X
X0 a_109_93# C_N VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 a_215_53# B VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 VGND a_109_93# a_215_53# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 VGND A a_215_53# sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 VPWR A a_369_297# sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.06825 ps=0.745 w=0.42 l=0.15
X5 a_369_297# B a_297_297# sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 X a_215_53# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.14825 ps=1.34 w=1 l=0.15
X7 a_297_297# a_109_93# a_215_53# sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X8 a_109_93# C_N VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 X a_215_53# VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.10025 ps=0.985 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_1 VGND VPWR X A  
X0 VPWR a_75_212# X sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1 a_75_212# A VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 a_75_212# A VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X3 VGND a_75_212# X sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1  
.ends

.subckt sky130_fd_sc_hd__buf_1 VGND VPWR X A  
X0 VPWR A a_27_47# sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1 X a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 X a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X3 VGND A a_27_47# sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand3b_1   VGND VPWR Y B C A_N
X0 Y a_53_93# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.1925 ps=1.385 w=1 l=0.15
X1 a_232_47# C VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X2 VPWR B Y sky130_fd_pr__pfet_01v8_hvt ad=0.1925 pd=1.385 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR A_N a_53_93# sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X4 VGND A_N a_53_93# sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 a_316_47# B a_232_47# sky130_fd_pr__nfet_01v8 ad=0.125125 pd=1.035 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 Y a_53_93# a_316_47# sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.125125 ps=1.035 w=0.65 l=0.15
X7 Y C VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand2_1   VGND VPWR A Y B
X0 VPWR A Y sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A a_113_47# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_113_47# B VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 Y B VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_2 VGND VPWR A X  
X0 VPWR A a_27_47# sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X1 VPWR a_27_47# X sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15 M=2
X2 VGND A a_27_47# sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X3 X a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15 M=2
.ends

.subckt sky130_fd_sc_hd__a2111oi_1  VPWR VGND  D1 C1 B1 A1 Y A2
X0 a_316_297# C1 a_217_297# sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.1725 ps=1.345 w=1 l=0.15
X1 Y D1 VGND sky130_fd_pr__nfet_01v8 ad=0.125125 pd=1.035 as=0.481 ps=2.78 w=0.65 l=0.15
X2 VGND C1 Y sky130_fd_pr__nfet_01v8 ad=0.12025 pd=1.02 as=0.125125 ps=1.035 w=0.65 l=0.15
X3 a_420_297# B1 a_316_297# sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=1.58 as=0.185 ps=1.37 w=1 l=0.15
X4 VPWR A1 a_420_297# sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.29 ps=1.58 w=1 l=0.15
X5 VGND A2 a_568_47# sky130_fd_pr__nfet_01v8 ad=0.19175 pd=1.89 as=0.0845 ps=0.91 w=0.65 l=0.15
X6 Y B1 VGND sky130_fd_pr__nfet_01v8 ad=0.19175 pd=1.24 as=0.12025 ps=1.02 w=0.65 l=0.15
X7 a_420_297# A2 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.1375 ps=1.275 w=1 l=0.15
X8 a_217_297# D1 Y sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.755 ps=3.51 w=1 l=0.15
X9 a_568_47# A1 Y sky130_fd_pr__nfet_01v8 ad=0.0845 pd=0.91 as=0.19175 ps=1.24 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor3b_1   VGND VPWR C_N B Y A
X0 VGND a_91_199# Y sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.221 ps=1.98 w=0.65 l=0.15
X1 Y B VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 VPWR A a_245_297# sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X3 a_91_199# C_N VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X4 VGND A Y sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 a_245_297# B a_161_297# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_91_199# C_N VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X7 a_161_297# a_91_199# Y sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.32 ps=2.64 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_2 VPWR VGND X A  
X0 VPWR a_27_47# X sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15 M=2
X1 VPWR A a_27_47# sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X2 X a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15 M=2
X3 VGND A a_27_47# sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__and3b_1 A_N B X C VGND VPWR  
X0 a_109_93# A_N VGND sky130_fd_pr__nfet_01v8 ad=0.10785 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 X a_209_311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X2 a_109_93# A_N VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1087 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 a_296_53# a_109_93# a_209_311# sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.107825 ps=1.36 w=0.42 l=0.15
X4 VPWR C a_209_311# sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.074375 ps=0.815 w=0.42 l=0.15
X5 a_368_53# B a_296_53# sky130_fd_pr__nfet_01v8 ad=0.05355 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 X a_209_311# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.122275 ps=1.08 w=0.65 l=0.15
X7 a_209_311# B VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.074375 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 VPWR a_109_93# a_209_311# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1085 ps=1.36 w=0.42 l=0.15
X9 VGND C a_368_53# sky130_fd_pr__nfet_01v8 ad=0.122275 pd=1.08 as=0.05355 ps=0.675 w=0.42 l=0.15
.ends

.subckt mux16x1_project data_in[0] data_in[10] data_in[11] data_in[12] data_in[13]
+ data_in[14] data_in[15] data_in[1] data_in[2] data_in[3] data_in[4] data_in[5] data_in[6]
+ data_in[7] data_in[8] data_in[9] select[0] select[1] select[2] select[3] y vssd1
+ vccd1
XFILLER_0_3_39 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_18_29 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_0_29 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_10_41 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_29_39 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_21_51 vssd1 vccd1   sky130_fd_sc_hd__decap_4
XFILLER_0_26_29 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_10_53 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_19_51 vssd1 vccd1   sky130_fd_sc_hd__decap_4
XFILLER_0_1_51 vssd1 vccd1   sky130_fd_sc_hd__decap_4
XFILLER_0_6_29 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_13_9 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_16_41 vssd1 vccd1   sky130_ef_sc_hd__decap_12
Xoutput21   vssd1 vccd1 _26_/Y y sky130_fd_sc_hd__buf_12
XFILLER_0_13_53 vccd1 vssd1   sky130_fd_sc_hd__decap_3
XFILLER_0_9_18 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_10_10 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_10_65 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_24_41 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_16_53 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_27_30 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_4_41 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_13_21 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_24_53 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_10_22 vccd1 vssd1   sky130_fd_sc_hd__decap_6
XFILLER_0_10_77 vssd1 vccd1   sky130_fd_sc_hd__decap_4
XFILLER_0_7_30 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_13_33 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_27_42 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_4_53 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_24_65 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_27_6 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_7_42 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_0_9 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_13_45 vccd1 vssd1   sky130_fd_sc_hd__decap_8
XFILLER_0_24_77 vssd1 vccd1   sky130_fd_sc_hd__decap_4
XFILLER_0_4_65 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_18_3 vccd1 vssd1   sky130_fd_sc_hd__decap_8
XPHY_0 vccd1 vssd1   sky130_fd_sc_hd__decap_3
XFILLER_0_9_6 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_13_57 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_4_77 vssd1 vccd1   sky130_fd_sc_hd__decap_4
X_26_   vssd1 vccd1 _21_/X _25_/A _26_/Y _25_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_21_57 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XPHY_1 vccd1 vssd1   sky130_fd_sc_hd__decap_3
XFILLER_0_13_69 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_19_57 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_1_57 vssd1 vccd1   sky130_ef_sc_hd__decap_12
X_25_   vssd1 vccd1 _25_/A _25_/B _25_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_21_69 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XPHY_2 vccd1 vssd1   sky130_fd_sc_hd__decap_3
XFILLER_0_27_57 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_1_69 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_19_69 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_21_15 vssd1 vccd1   sky130_ef_sc_hd__decap_12
X_24_ vssd1 vccd1   _25_/B _22_/X _24_/S _23_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_16_15 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_27_69 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XPHY_3 vccd1 vssd1   sky130_fd_sc_hd__decap_3
XFILLER_0_7_57 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_16_3 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_19_15 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_1_15 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_21_27 vssd1 vccd1   sky130_ef_sc_hd__decap_12
X_23_   vssd1 vccd1 _23_/A1 _23_/A0 _20_/B _23_/A3 _23_/A2 _23_/S1 _23_/X
+ sky130_fd_sc_hd__mux4_1
XPHY_4 vccd1 vssd1   sky130_fd_sc_hd__decap_3
XFILLER_0_7_69 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_30_6 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_1_27 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_10_29 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_19_27 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_21_39 vssd1 vccd1   sky130_ef_sc_hd__decap_12
X_22_   vssd1 vccd1 _22_/A1 _22_/A0 _20_/B _22_/A3 _22_/A2 _23_/S1 _22_/X
+ sky130_fd_sc_hd__mux4_1
XPHY_5 vccd1 vssd1   sky130_fd_sc_hd__decap_3
XFILLER_0_21_3 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_19_39 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_1_39 vssd1 vccd1   sky130_ef_sc_hd__decap_12
X_21_ vssd1 vccd1 _19_/Y _20_/X _18_/Y _21_/X _16_/Y _23_/S1   sky130_fd_sc_hd__a41o_1
XFILLER_0_16_29 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XPHY_6 vccd1 vssd1   sky130_fd_sc_hd__decap_3
XFILLER_0_14_3 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_24_29 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_24_18 vccd1 vssd1   sky130_fd_sc_hd__decap_8
XFILLER_0_3_3 vssd1 vccd1   sky130_ef_sc_hd__decap_12
X_20_ vssd1 vccd1   _20_/B input4/X _24_/S _20_/X sky130_fd_sc_hd__or3b_1
Xinput1 vssd1 vccd1 _23_/A0 data_in[0]   sky130_fd_sc_hd__clkbuf_1
XPHY_7 vccd1 vssd1   sky130_fd_sc_hd__decap_3
XFILLER_0_27_18 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_4_18 vccd1 vssd1   sky130_fd_sc_hd__decap_8
XFILLER_0_4_29 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_14_41 vssd1 vccd1   sky130_ef_sc_hd__decap_12
Xinput2 vssd1 vccd1 _14_/C data_in[10]   sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_20 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XPHY_8 vccd1 vssd1   sky130_fd_sc_hd__decap_3
XFILLER_0_7_18 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_22_41 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_14_53 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_30_41 vssd1 vccd1   sky130_ef_sc_hd__decap_12
Xinput3 vssd1 vccd1 _13_/A1 data_in[11]   sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_32 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_22_53 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_2_41 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XPHY_9 vccd1 vssd1   sky130_fd_sc_hd__decap_3
XFILLER_0_17_53 vccd1 vssd1   sky130_fd_sc_hd__decap_3
XFILLER_0_14_65 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_30_53 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_28_41 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_1_3 vssd1 vccd1   sky130_ef_sc_hd__decap_12
Xinput4 vssd1 vccd1 input4/X data_in[12]   sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_44 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_2_53 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_22_65 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_8_41 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_17_21 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_28_53 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_14_77 vssd1 vccd1   sky130_fd_sc_hd__decap_4
XFILLER_0_30_65 vssd1 vccd1   sky130_ef_sc_hd__decap_12
Xinput5 vssd1 vccd1 _17_/A0 data_in[13]   sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_22 vccd1 vssd1   sky130_fd_sc_hd__decap_6
XFILLER_0_2_65 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_17_33 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_22_77 vssd1 vccd1   sky130_fd_sc_hd__decap_4
XFILLER_0_8_53 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_30_77 vssd1 vccd1   sky130_fd_sc_hd__decap_4
XFILLER_0_28_65 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_11_57 vssd1 vccd1   sky130_ef_sc_hd__decap_12
Xinput6 vssd1 vccd1 _19_/C data_in[14]   sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_77 vssd1 vccd1   sky130_fd_sc_hd__decap_4
XFILLER_0_8_65 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_17_45 vccd1 vssd1   sky130_fd_sc_hd__decap_8
Xinput20 vssd1 vccd1 _25_/A select[3]   sky130_fd_sc_hd__buf_1
XFILLER_0_28_77 vssd1 vccd1   sky130_fd_sc_hd__decap_4
XFILLER_0_28_3 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_12_6 vssd1 vccd1   sky130_ef_sc_hd__decap_12
Xinput7 vssd1 vccd1 _17_/A1 data_in[15]   sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_69 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_17_57 vssd1 vccd1   sky130_ef_sc_hd__decap_12
Xinput10 vssd1 vccd1 _22_/A1 data_in[3]   sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_77 vssd1 vccd1   sky130_fd_sc_hd__decap_4
XFILLER_0_5_12 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_25_57 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_25_24 vssd1 vccd1   sky130_ef_sc_hd__decap_12
Xinput8 vssd1 vccd1 _22_/A0 data_in[1]   sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_69 vssd1 vccd1   sky130_ef_sc_hd__decap_12
Xinput11 vssd1 vccd1 _23_/A2 data_in[4]   sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_15 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_5_24 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_5_57 vssd1 vccd1   sky130_ef_sc_hd__decap_12
Xinput9 vssd1 vccd1 _23_/A1 data_in[2]   sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_69 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_25_36 vssd1 vccd1   sky130_ef_sc_hd__decap_12
Xinput12 vssd1 vccd1 _22_/A2 data_in[5]   sky130_fd_sc_hd__clkbuf_1
XPHY_60 vccd1 vssd1   sky130_fd_sc_hd__decap_3
XFILLER_0_26_3 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_5_36 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_5_69 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_25_48 vccd1 vssd1   sky130_fd_sc_hd__decap_8
XPHY_61 vccd1 vssd1   sky130_fd_sc_hd__decap_3
XPHY_50 vccd1 vssd1   sky130_fd_sc_hd__decap_3
Xinput13 vssd1 vccd1 _23_/A3 data_in[6]   sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_15 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_8_14 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_19_3 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_5_48 vccd1 vssd1   sky130_fd_sc_hd__decap_8
XFILLER_0_8_3 vccd1 vssd1   sky130_fd_sc_hd__decap_3
Xinput14 vssd1 vccd1 _22_/A3 data_in[7]   sky130_fd_sc_hd__clkbuf_1
XPHY_40 vccd1 vssd1   sky130_fd_sc_hd__decap_3
XPHY_62 vccd1 vssd1   sky130_fd_sc_hd__decap_3
XPHY_51 vccd1 vssd1   sky130_fd_sc_hd__decap_3
X_19_   vssd1 vccd1 _19_/Y _20_/B _19_/C _24_/S sky130_fd_sc_hd__nand3b_1
XFILLER_0_14_29 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XPHY_30 vccd1 vssd1   sky130_fd_sc_hd__decap_3
XPHY_41 vccd1 vssd1   sky130_fd_sc_hd__decap_3
XFILLER_0_22_29 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XPHY_63 vccd1 vssd1   sky130_fd_sc_hd__decap_3
XPHY_52 vccd1 vssd1   sky130_fd_sc_hd__decap_3
Xinput15 vssd1 vccd1 _15_/C_N data_in[8]   sky130_fd_sc_hd__clkbuf_1
X_18_   vssd1 vccd1 _24_/S _18_/Y _18_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_30_29 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_30_18 vccd1 vssd1   sky130_fd_sc_hd__decap_8
XFILLER_0_31_61 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_2_18 vccd1 vssd1   sky130_fd_sc_hd__decap_8
XFILLER_0_2_29 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XPHY_20 vccd1 vssd1   sky130_fd_sc_hd__decap_3
XFILLER_0_12_41 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XPHY_31 vccd1 vssd1   sky130_fd_sc_hd__decap_3
XPHY_42 vccd1 vssd1   sky130_fd_sc_hd__decap_3
XPHY_53 vccd1 vssd1   sky130_fd_sc_hd__decap_3
X_17_ vssd1 vccd1   _18_/B _17_/A1 _20_/B _17_/A0 sky130_fd_sc_hd__mux2_1
Xinput16 vssd1 vccd1 _13_/A0 data_in[9]   sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_29 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_20_41 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XPHY_10 vccd1 vssd1   sky130_fd_sc_hd__decap_3
XPHY_21 vccd1 vssd1   sky130_fd_sc_hd__decap_3
XFILLER_0_15_30 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XPHY_32 vccd1 vssd1   sky130_fd_sc_hd__decap_3
XPHY_43 vccd1 vssd1   sky130_fd_sc_hd__decap_3
XFILLER_0_31_73 vssd1 vccd1   sky130_fd_sc_hd__decap_4
XPHY_54 vccd1 vssd1   sky130_fd_sc_hd__decap_3
XFILLER_0_3_51 vssd1 vccd1   sky130_fd_sc_hd__decap_4
XFILLER_0_12_53 vssd1 vccd1   sky130_ef_sc_hd__decap_12
Xinput17 vssd1 vccd1 select[0] _24_/S   sky130_fd_sc_hd__clkbuf_2
XFILLER_0_8_29 vssd1 vccd1   sky130_ef_sc_hd__decap_12
X_16_  vccd1 vssd1  _23_/S1 _15_/Y _14_/X _24_/S _16_/Y _13_/X sky130_fd_sc_hd__a2111oi_1
XFILLER_0_18_41 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_20_53 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_0_41 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_15_42 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_29_51 vssd1 vccd1   sky130_fd_sc_hd__decap_4
XPHY_11 vccd1 vssd1   sky130_fd_sc_hd__decap_3
XPHY_22 vccd1 vssd1   sky130_fd_sc_hd__decap_3
XFILLER_0_12_65 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XPHY_33 vccd1 vssd1   sky130_fd_sc_hd__decap_3
XPHY_44 vccd1 vssd1   sky130_fd_sc_hd__decap_3
XPHY_55 vccd1 vssd1   sky130_fd_sc_hd__decap_3
XFILLER_0_26_41 vssd1 vccd1   sky130_ef_sc_hd__decap_12
X_15_   vssd1 vccd1 _15_/C_N _20_/B _15_/Y _24_/S sky130_fd_sc_hd__nor3b_1
XFILLER_0_18_53 vssd1 vccd1   sky130_ef_sc_hd__decap_12
Xinput18 vccd1 vssd1 _20_/B select[1]   sky130_fd_sc_hd__buf_2
XFILLER_0_0_53 vccd1 vssd1   sky130_fd_sc_hd__decap_3
XFILLER_0_20_65 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_24_6 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XPHY_12 vccd1 vssd1   sky130_fd_sc_hd__decap_3
XFILLER_0_6_41 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_31_53 vccd1 vssd1   sky130_fd_sc_hd__decap_3
XFILLER_0_26_53 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XPHY_23 vccd1 vssd1   sky130_fd_sc_hd__decap_3
XFILLER_0_12_77 vssd1 vccd1   sky130_fd_sc_hd__decap_4
XPHY_34 vccd1 vssd1   sky130_fd_sc_hd__decap_3
XPHY_45 vccd1 vssd1   sky130_fd_sc_hd__decap_3
Xinput19 vssd1 vccd1 select[2] _23_/S1   sky130_fd_sc_hd__clkbuf_2
XPHY_56 vccd1 vssd1   sky130_fd_sc_hd__decap_3
X_14_ _24_/S _20_/B _14_/X _14_/C vssd1 vccd1   sky130_fd_sc_hd__and3b_1
XFILLER_0_18_65 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_0_21 vccd1 vssd1   sky130_fd_sc_hd__decap_6
XFILLER_0_9_30 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_17_6 vccd1 vssd1   sky130_fd_sc_hd__decap_8
XFILLER_0_20_77 vssd1 vccd1   sky130_fd_sc_hd__decap_4
XFILLER_0_6_53 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XPHY_13 vccd1 vssd1   sky130_fd_sc_hd__decap_3
XPHY_24 vccd1 vssd1   sky130_fd_sc_hd__decap_3
XPHY_35 vccd1 vssd1   sky130_fd_sc_hd__decap_3
XPHY_46 vccd1 vssd1   sky130_fd_sc_hd__decap_3
XPHY_57 vccd1 vssd1   sky130_fd_sc_hd__decap_3
XFILLER_0_26_65 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_9_42 vssd1 vccd1   sky130_ef_sc_hd__decap_12
X_13_ vssd1 vccd1   _13_/X _13_/A1 _20_/B _13_/A0 sky130_fd_sc_hd__mux2_1
XFILLER_0_18_77 vssd1 vccd1   sky130_fd_sc_hd__decap_4
XFILLER_0_6_10 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_31_33 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_26_77 vssd1 vccd1   sky130_fd_sc_hd__decap_4
XPHY_14 vccd1 vssd1   sky130_fd_sc_hd__decap_3
XFILLER_0_6_65 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XPHY_25 vccd1 vssd1   sky130_fd_sc_hd__decap_3
XPHY_36 vccd1 vssd1   sky130_fd_sc_hd__decap_3
XPHY_58 vccd1 vssd1   sky130_fd_sc_hd__decap_3
XPHY_47 vccd1 vssd1   sky130_fd_sc_hd__decap_3
XFILLER_0_15_57 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_22_6 vccd1 vssd1   sky130_fd_sc_hd__decap_6
XFILLER_0_31_45 vccd1 vssd1   sky130_fd_sc_hd__decap_8
XFILLER_0_6_22 vccd1 vssd1   sky130_fd_sc_hd__decap_6
XFILLER_0_6_77 vssd1 vccd1   sky130_fd_sc_hd__decap_4
XPHY_15 vccd1 vssd1   sky130_fd_sc_hd__decap_3
XPHY_26 vccd1 vssd1   sky130_fd_sc_hd__decap_3
XPHY_37 vccd1 vssd1   sky130_fd_sc_hd__decap_3
XPHY_59 vccd1 vssd1   sky130_fd_sc_hd__decap_3
XPHY_48 vccd1 vssd1   sky130_fd_sc_hd__decap_3
XFILLER_0_23_24 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_23_57 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_0_57 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_15_6 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_15_69 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_31_13 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_4_6 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XPHY_16 vccd1 vssd1   sky130_fd_sc_hd__decap_3
XPHY_27 vccd1 vssd1   sky130_fd_sc_hd__decap_3
XPHY_38 vccd1 vssd1   sky130_fd_sc_hd__decap_3
XPHY_49 vccd1 vssd1   sky130_fd_sc_hd__decap_3
XFILLER_0_3_57 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_23_36 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_23_69 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_0_69 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_31_25 vccd1 vssd1   sky130_fd_sc_hd__decap_3
XFILLER_0_29_57 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XPHY_17 vccd1 vssd1   sky130_fd_sc_hd__decap_3
XPHY_28 vccd1 vssd1   sky130_fd_sc_hd__decap_3
XPHY_39 vccd1 vssd1   sky130_fd_sc_hd__decap_3
XFILLER_0_3_69 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_23_48 vccd1 vssd1   sky130_fd_sc_hd__decap_8
XFILLER_0_29_69 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_9_57 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XPHY_18 vccd1 vssd1   sky130_fd_sc_hd__decap_3
XPHY_29 vccd1 vssd1   sky130_fd_sc_hd__decap_3
XFILLER_0_20_6 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_26_15 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_3_15 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_18_16 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_9_69 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_29_3 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_29_15 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XPHY_19 vccd1 vssd1   sky130_fd_sc_hd__decap_3
XFILLER_0_2_6 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_3_27 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_12_18 vccd1 vssd1   sky130_fd_sc_hd__decap_8
XFILLER_0_12_29 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_20_18 vccd1 vssd1   sky130_fd_sc_hd__decap_8
XFILLER_0_20_29 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_29_27 vssd1 vccd1   sky130_ef_sc_hd__decap_12
XFILLER_0_15_18 vssd1 vccd1   sky130_ef_sc_hd__decap_12
.ends

.subckt sky130_osu_sc_12T_hs__mux2_1 A1 A0 Y vssd1  vccd1 S0
X0 Y S0 A0 sky130_fd_pr__pfet_01v8 ad=0.1764 pd=1.54 as=0.3402 ps=3.06 w=1.26 l=0.15
X1 Y a_110_114# A0 vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0.077 pd=0.83 as=0.1485 ps=1.64 w=0.55 l=0.15
X2 A1 a_110_114# Y sky130_fd_pr__pfet_01v8 ad=0.3339 pd=3.05 as=0.1764 ps=1.54 w=1.26 l=0.15
X3 A1 S0 Y vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0.14575 pd=1.63 as=0.077 ps=0.83 w=0.55 l=0.15
X4 a_110_114# S0 vccd1 sky130_fd_pr__pfet_01v8 ad=0.3339 pd=3.05 as=0.3402 ps=3.06 w=1.26 l=0.15
X5 a_110_114# S0 vssd1  vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0.14575 pd=1.63 as=0.1485 ps=1.64 w=0.55 l=0.15
.ends

.subckt scs130hd_mpr2ca_8 A1 B1 R3 R1 R0 B0 A0 R2 vpwr  vgnd vgnd_uq0 
X0 a_772_910# B0 vgnd sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.234 ps=2.02 w=0.65 l=0.15
X1 a_178_822# A0 a_352_928# sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 a_296_52# a_108_92# a_208_310# sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1079 ps=1.36 w=0.42 l=0.15
X3 a_824_46# B1 a_752_46# sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 vgnd_uq0 a_844_910# R1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 vpwr A1 a_670_46# sky130_fd_pr__pfet_01v8_hvt ad=0.140425 pd=1.335 as=0.0672 ps=0.74 w=0.42 l=0.15
X6 R3 a_670_46# vpwr sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.140425 ps=1.335 w=1 l=0.15
X7 a_352_928# B0 vgnd sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1118 ps=1.04 w=0.42 l=0.15
X8 vpwr A1 a_208_310# sky130_fd_pr__pfet_01v8_hvt ad=0.140425 pd=1.335 as=0.07525 ps=0.82 w=0.42 l=0.15
X9 a_368_52# B1 a_296_52# sky130_fd_pr__nfet_01v8 ad=0.0525 pd=0.67 as=0.0441 ps=0.63 w=0.42 l=0.15
X10 vgnd_uq0 A1 a_824_46# sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X11 vpwr a_178_822# R0 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.47 ps=2.94 w=1 l=0.15
X12 a_208_310# B1 vpwr sky130_fd_pr__pfet_01v8_hvt ad=0.07525 pd=0.82 as=0.0567 ps=0.69 w=0.42 l=0.15
X13 vpwr a_844_910# a_1212_296# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X14 vpwr a_108_92# a_208_310# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1085 ps=1.36 w=0.42 l=0.15
X15 vpwr A1 a_760_590# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X16 a_670_46# B1 vpwr sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.0567 ps=0.69 w=0.42 l=0.15
X17 a_1212_296# R3 R1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X18 vpwr A0 a_178_822# sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X19 R2 a_208_310# vgnd_uq0 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1222 ps=1.08 w=0.65 l=0.15
X20 a_844_910# B1 a_760_590# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X21 vpwr R0 a_670_46# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X22 R3 a_670_46# vgnd_uq0 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X23 a_178_822# B0 vpwr sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.16655 ps=1.39 w=0.42 l=0.15
X24 a_760_590# B0 vpwr sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3 ps=2.6 w=1 l=0.15
X25 vgnd_uq0 A1 a_368_52# sky130_fd_pr__nfet_01v8 ad=0.1222 pd=1.08 as=0.0525 ps=0.67 w=0.42 l=0.15
X26 vgnd a_178_822# R0 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X27 a_1040_910# A0 a_844_910# sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X28 a_108_92# R3 vgnd_uq0 sky130_fd_pr__nfet_01v8 ad=0.1078 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X29 R1 R3 vgnd_uq0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X30 a_844_910# A1 a_772_910# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X31 a_108_92# R3 vpwr sky130_fd_pr__pfet_01v8_hvt ad=0.1087 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X32 R2 a_208_310# vpwr sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.140425 ps=1.335 w=1 l=0.15
X33 a_760_590# A0 a_844_910# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X34 a_752_46# R0 a_670_46# sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X35 vgnd B1 a_1040_910# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
.ends

.subckt sky130_osu_sc_12T_hs__inv_1 vssd1 A Y vccd1
X0 Y A vccd1 sky130_fd_pr__pfet_01v8 ad=0.3339 pd=3.05 as=0.3402 ps=3.06 w=1.26 l=0.15
X1 Y A vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0.14575 pd=1.63 as=0.1485 ps=1.64 w=0.55 l=0.15
.ends

.subckt sky130_osu_single_mpr2ca_8_b0r1 Y1 Y0 in sel scs130hd_mpr2ca_8_0/B1 vccd1
+ vssd1
Xsky130_osu_sc_12T_hs__mux2_1_0 scs130hd_mpr2ca_8_0/R1 in sky130_osu_sc_12T_hs__inv_1_1/A
+ vssd1 vccd1 sel sky130_osu_sc_12T_hs__mux2_1
Xsky130_osu_sc_12T_hs__mux2_1_1 in vssd1 scs130hd_mpr2ca_8_0/B1 vssd1 vccd1 sel sky130_osu_sc_12T_hs__mux2_1
Xscs130hd_mpr2ca_8_0 scs130hd_mpr2ca_8_0/B1 scs130hd_mpr2ca_8_0/B1 scs130hd_mpr2ca_8_0/R3
+ scs130hd_mpr2ca_8_0/R1 scs130hd_mpr2ca_8_0/R0 vssd1 scs130hd_mpr2ca_8_0/B1 scs130hd_mpr2ca_8_0/R2
+ vccd1  vssd1 vssd1  scs130hd_mpr2ca_8
Xsky130_osu_sc_12T_hs__mux2_1_2 in scs130hd_mpr2ca_8_0/R1 sky130_osu_sc_12T_hs__inv_1_4/A
+ vssd1 vccd1 sel sky130_osu_sc_12T_hs__mux2_1
Xsky130_osu_sc_12T_hs__inv_1_1 vssd1 sky130_osu_sc_12T_hs__inv_1_1/A sky130_osu_sc_12T_hs__inv_1_2/A
+ vccd1 sky130_osu_sc_12T_hs__inv_1
Xsky130_osu_sc_12T_hs__inv_1_2 vssd1 sky130_osu_sc_12T_hs__inv_1_2/A Y1 vccd1 sky130_osu_sc_12T_hs__inv_1
Xsky130_osu_sc_12T_hs__inv_1_3 vssd1 sky130_osu_sc_12T_hs__inv_1_4/Y Y0 vccd1 sky130_osu_sc_12T_hs__inv_1
Xsky130_osu_sc_12T_hs__inv_1_4 vssd1 sky130_osu_sc_12T_hs__inv_1_4/A sky130_osu_sc_12T_hs__inv_1_4/Y
+ vccd1 sky130_osu_sc_12T_hs__inv_1
.ends

.subckt sky130_osu_ring_oscillator_mpr2ca_8_b0r1 s4 s5 X5_Y1 X4_Y1 X3_Y1 X2_Y1 X1_Y1
+ start vccd1 s2 s3 s1 vssd1
Xsky130_osu_single_mpr2ca_8_b0r1_0 X5_Y1 sky130_osu_sc_12T_hs__mux2_1_0/A0 sky130_osu_single_mpr2ca_8_b0r1_4/Y0
+ s5 sky130_osu_single_mpr2ca_8_b0r1_0/scs130hd_mpr2ca_8_0/B1 vccd1 vssd1 sky130_osu_single_mpr2ca_8_b0r1
Xsky130_osu_single_mpr2ca_8_b0r1_1 X1_Y1 sky130_osu_single_mpr2ca_8_b0r1_2/in sky130_osu_sc_12T_hs__mux2_1_0/Y
+ s1 sky130_osu_single_mpr2ca_8_b0r1_1/scs130hd_mpr2ca_8_0/B1 vccd1 vssd1 sky130_osu_single_mpr2ca_8_b0r1
Xsky130_osu_single_mpr2ca_8_b0r1_2 X2_Y1 sky130_osu_single_mpr2ca_8_b0r1_3/in sky130_osu_single_mpr2ca_8_b0r1_2/in
+ s2 sky130_osu_single_mpr2ca_8_b0r1_2/scs130hd_mpr2ca_8_0/B1 vccd1 vssd1 sky130_osu_single_mpr2ca_8_b0r1
Xsky130_osu_sc_12T_hs__mux2_1_0 vccd1 sky130_osu_sc_12T_hs__mux2_1_0/A0 sky130_osu_sc_12T_hs__mux2_1_0/Y
+ vssd1 vccd1 start sky130_osu_sc_12T_hs__mux2_1
Xsky130_osu_single_mpr2ca_8_b0r1_3 X3_Y1 sky130_osu_single_mpr2ca_8_b0r1_4/in sky130_osu_single_mpr2ca_8_b0r1_3/in
+ s3 sky130_osu_single_mpr2ca_8_b0r1_3/scs130hd_mpr2ca_8_0/B1 vccd1 vssd1 sky130_osu_single_mpr2ca_8_b0r1
Xsky130_osu_single_mpr2ca_8_b0r1_4 X4_Y1 sky130_osu_single_mpr2ca_8_b0r1_4/Y0 sky130_osu_single_mpr2ca_8_b0r1_4/in
+ s4 sky130_osu_single_mpr2ca_8_b0r1_4/scs130hd_mpr2ca_8_0/B1 vccd1 vssd1 sky130_osu_single_mpr2ca_8_b0r1
.ends

.subckt scs130hd_mpr2xa_8   R0 R1 R2 R3 B1 B0 A0 vgnd vpwr A1
X0 R0 a_56_48# vpwr sky130_fd_pr__pfet_01v8 ad=0.27 pd=2.54 as=0.165 ps=1.33 w=1 l=0.15
X1 a_1294_296# a_676_198# R3 sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.27 ps=2.54 w=1 l=0.15
X2 vpwr a_56_48# a_1294_296# sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X3 a_1486_296# a_334_296# vpwr sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X4 R1 R3 a_1486_296# sky130_fd_pr__pfet_01v8 ad=0.27 pd=2.54 as=0.165 ps=1.33 w=1 l=0.15
X5 R2 a_676_198# vgnd sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X6 vgnd a_56_48# R3 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X7 vpwr B0 a_56_48# sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.27 ps=2.54 w=1 l=0.15
X8 a_334_296# A1 a_238_296# sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X9 a_238_296# B0 a_334_296# sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X10 a_676_198# B1 a_910_46# sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.10725 ps=0.98 w=0.65 l=0.15
X11 R3 a_676_198# vgnd sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X12 a_238_296# A0 vpwr sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X13 a_142_46# B0 a_56_48# sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.1802 ps=1.86 w=0.65 l=0.15
X14 vgnd a_56_48# R0 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.1755 ps=1.84 w=0.65 l=0.15
X15 vgnd R3 R1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.10725 ps=0.98 w=0.65 l=0.15
X16 a_334_296# B0 a_334_46# sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X17 R1 a_334_296# vgnd sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X18 a_334_46# A1 vgnd sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X19 vgnd A0 a_142_46# sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X20 vgnd A0 a_526_46# sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X21 a_526_46# B1 a_334_296# sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X22 a_910_46# A1 vgnd sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X23 a_56_48# A0 vpwr sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X24 a_676_198# A1 vpwr sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.27 ps=2.54 w=1 l=0.15
X25 vgnd R0 R2 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X26 vpwr B1 a_238_296# sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X27 R2 a_676_198# a_56_48# sky130_fd_pr__pfet_01v8 ad=0.27 pd=2.54 as=0.165 ps=1.33 w=1 l=0.15
X28 vpwr B1 a_676_198# sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
.ends

* Black-box entry subcircuit for sky130_osu_sc_12T_hs__fill_8 abstract view
.subckt sky130_osu_sc_12T_hs__fill_8
.ends

.subckt sky130_osu_single_mpr2xa_8_b0r2 Y0 Y1 sel vccd1 in vssd1
Xscs130hd_mpr2xa_8_0   scs130hd_mpr2xa_8_0/R0 scs130hd_mpr2xa_8_0/R1 scs130hd_mpr2xa_8_0/R2
+ scs130hd_mpr2xa_8_0/R3 scs130hd_mpr2xa_8_0/B1 vssd1 scs130hd_mpr2xa_8_0/B1 vssd1
+ vccd1 scs130hd_mpr2xa_8_0/B1 scs130hd_mpr2xa_8
Xsky130_osu_sc_12T_hs__mux2_1_0 scs130hd_mpr2xa_8_0/R2 in sky130_osu_sc_12T_hs__inv_1_1/A
+ vssd1 vccd1 sel sky130_osu_sc_12T_hs__mux2_1
Xsky130_osu_sc_12T_hs__mux2_1_1 in vssd1 scs130hd_mpr2xa_8_0/B1 vssd1 vccd1 sel sky130_osu_sc_12T_hs__mux2_1
Xsky130_osu_sc_12T_hs__mux2_1_2 in scs130hd_mpr2xa_8_0/R2 sky130_osu_sc_12T_hs__inv_1_4/A
+ vssd1 vccd1 sel sky130_osu_sc_12T_hs__mux2_1
Xsky130_osu_sc_12T_hs__inv_1_1 vssd1 sky130_osu_sc_12T_hs__inv_1_1/A sky130_osu_sc_12T_hs__inv_1_2/A
+ vccd1 sky130_osu_sc_12T_hs__inv_1
Xsky130_osu_sc_12T_hs__inv_1_2 vssd1 sky130_osu_sc_12T_hs__inv_1_2/A Y1 vccd1 sky130_osu_sc_12T_hs__inv_1
Xsky130_osu_sc_12T_hs__inv_1_3 vssd1 sky130_osu_sc_12T_hs__inv_1_4/Y Y0 vccd1 sky130_osu_sc_12T_hs__inv_1
Xsky130_osu_sc_12T_hs__inv_1_4 vssd1 sky130_osu_sc_12T_hs__inv_1_4/A sky130_osu_sc_12T_hs__inv_1_4/Y
+ vccd1 sky130_osu_sc_12T_hs__inv_1
.ends

.subckt sky130_osu_ring_oscillator_mpr2xa_8_b0r2 s1 s3 s4 s5 X1_Y1 X5_Y1 start vccd1
+ X4_Y1 X3_Y1 s2 X2_Y1 vssd1
Xsky130_osu_sc_12T_hs__mux2_1_0 vccd1 sky130_osu_sc_12T_hs__mux2_1_0/A0 sky130_osu_sc_12T_hs__mux2_1_0/Y
+ vssd1 vccd1 start sky130_osu_sc_12T_hs__mux2_1
Xsky130_osu_single_mpr2xa_8_b0r2_0 sky130_osu_sc_12T_hs__mux2_1_0/A0 X5_Y1 s5 vccd1
+ sky130_osu_single_mpr2xa_8_b0r2_4/Y0 vssd1 sky130_osu_single_mpr2xa_8_b0r2
Xsky130_osu_single_mpr2xa_8_b0r2_1 sky130_osu_single_mpr2xa_8_b0r2_2/in X1_Y1 s1 vccd1
+ sky130_osu_sc_12T_hs__mux2_1_0/Y vssd1 sky130_osu_single_mpr2xa_8_b0r2
Xsky130_osu_single_mpr2xa_8_b0r2_2 sky130_osu_single_mpr2xa_8_b0r2_3/in X2_Y1 s2 vccd1
+ sky130_osu_single_mpr2xa_8_b0r2_2/in vssd1 sky130_osu_single_mpr2xa_8_b0r2
Xsky130_osu_single_mpr2xa_8_b0r2_4 sky130_osu_single_mpr2xa_8_b0r2_4/Y0 X4_Y1 s4 vccd1
+ sky130_osu_single_mpr2xa_8_b0r2_4/in vssd1 sky130_osu_single_mpr2xa_8_b0r2
Xsky130_osu_single_mpr2xa_8_b0r2_3 sky130_osu_single_mpr2xa_8_b0r2_4/in X3_Y1 s3 vccd1
+ sky130_osu_single_mpr2xa_8_b0r2_3/in vssd1 sky130_osu_single_mpr2xa_8_b0r2
.ends

.subckt scs130hd_mpr2ct_8 A1 A0 B0 B1 R0 R1 R2 R3 vpwr  vgnd vgnd_uq0 
X0 vpwr B1 a_1131_911# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 vgnd_uq0 a_1131_911# a_1133_47# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 vpwr A1 a_665_591# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 vgnd_uq0 a_665_591# a_915_232# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_1131_911# A0 vpwr sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5 R3 a_443_21# a_401_297# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X6 a_945_297# a_665_591# vpwr sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7 a_665_591# B0 vpwr sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8 vpwr a_443_21# a_661_297# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X9 R0 a_81_21# vpwr sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15 M=2
X10 a_401_297# a_81_21# vpwr sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X11 R1 a_915_232# vgnd_uq0 sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.208 ps=1.94 w=0.65 l=0.15
X12 vgnd B1 a_937_911# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 vgnd B1 a_1213_911# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 a_443_21# A1 vpwr sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X15 vgnd_uq0 a_443_21# R3 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 a_661_297# R0 R2 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X17 vgnd_uq0 a_81_21# R0 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15 M=2
X18 a_665_591# A1 a_665_911# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 a_1213_911# A0 a_1131_911# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X20 a_665_911# B0 vgnd sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X21 vpwr A0 a_81_21# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X22 a_915_232# a_665_591# a_1301_297# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X23 R3 a_81_21# vgnd_uq0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X24 a_81_21# B0 vpwr sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X25 a_1301_297# a_1131_911# vpwr sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X26 a_937_911# A1 a_443_21# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X27 a_945_297# a_915_232# R1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3 ps=2.6 w=1 l=0.15
X28 R2 R0 vgnd_uq0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X29 a_1133_47# a_665_591# R1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25025 ps=1.42 w=0.65 l=0.15
X30 vpwr a_1131_911# a_945_297# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X31 a_915_232# a_1131_911# vgnd_uq0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X32 a_81_21# A0 a_205_911# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X33 a_205_911# B0 vgnd sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X34 vpwr B1 a_443_21# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X35 vgnd_uq0 a_443_21# R2 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_osu_single_mpr2ct_8_b0r1 Y0 Y1 in sel vccd1 vssd1
Xsky130_osu_sc_12T_hs__mux2_1_0 scs130hd_mpr2ct_8_1/R1 in sky130_osu_sc_12T_hs__inv_1_1/A
+ vssd1 vccd1 sel sky130_osu_sc_12T_hs__mux2_1
Xsky130_osu_sc_12T_hs__mux2_1_1 in vssd1 scs130hd_mpr2ct_8_1/B1 vssd1 vccd1 sel sky130_osu_sc_12T_hs__mux2_1
Xsky130_osu_sc_12T_hs__inv_1_0 vssd1 sky130_osu_sc_12T_hs__inv_1_1/Y Y1 vccd1 sky130_osu_sc_12T_hs__inv_1
Xsky130_osu_sc_12T_hs__mux2_1_2 in scs130hd_mpr2ct_8_1/R1 sky130_osu_sc_12T_hs__inv_1_4/A
+ vssd1 vccd1 sel sky130_osu_sc_12T_hs__mux2_1
Xsky130_osu_sc_12T_hs__inv_1_1 vssd1 sky130_osu_sc_12T_hs__inv_1_1/A sky130_osu_sc_12T_hs__inv_1_1/Y
+ vccd1 sky130_osu_sc_12T_hs__inv_1
Xsky130_osu_sc_12T_hs__inv_1_3 vssd1 sky130_osu_sc_12T_hs__inv_1_4/Y Y0 vccd1 sky130_osu_sc_12T_hs__inv_1
Xsky130_osu_sc_12T_hs__inv_1_4 vssd1 sky130_osu_sc_12T_hs__inv_1_4/A sky130_osu_sc_12T_hs__inv_1_4/Y
+ vccd1 sky130_osu_sc_12T_hs__inv_1
Xscs130hd_mpr2ct_8_1 scs130hd_mpr2ct_8_1/B1 scs130hd_mpr2ct_8_1/B1 vssd1 scs130hd_mpr2ct_8_1/B1
+ scs130hd_mpr2ct_8_1/R0 scs130hd_mpr2ct_8_1/R1 scs130hd_mpr2ct_8_1/R2 scs130hd_mpr2ct_8_1/R3
+ vccd1  vssd1 vssd1  scs130hd_mpr2ct_8
.ends

.subckt sky130_osu_ring_oscillator_mpr2ct_8_b0r1 s1 s2 s3 X5_Y1 X4_Y1 X3_Y1 X2_Y1
+ X1_Y1 s5 s4 start vccd1 vssd1
Xsky130_osu_sc_12T_hs__mux2_1_0 vccd1 sky130_osu_sc_12T_hs__mux2_1_0/A0 sky130_osu_sc_12T_hs__mux2_1_0/Y
+ vssd1 vccd1 start sky130_osu_sc_12T_hs__mux2_1
Xsky130_osu_single_mpr2ct_8_b0r1_0 sky130_osu_sc_12T_hs__mux2_1_0/A0 X5_Y1 sky130_osu_single_mpr2ct_8_b0r1_4/Y0
+ s5 vccd1 vssd1 sky130_osu_single_mpr2ct_8_b0r1
Xsky130_osu_single_mpr2ct_8_b0r1_2 sky130_osu_single_mpr2ct_8_b0r1_3/in X2_Y1 sky130_osu_single_mpr2ct_8_b0r1_2/in
+ s2 vccd1 vssd1 sky130_osu_single_mpr2ct_8_b0r1
Xsky130_osu_single_mpr2ct_8_b0r1_1 sky130_osu_single_mpr2ct_8_b0r1_2/in X1_Y1 sky130_osu_sc_12T_hs__mux2_1_0/Y
+ s1 vccd1 vssd1 sky130_osu_single_mpr2ct_8_b0r1
Xsky130_osu_single_mpr2ct_8_b0r1_3 sky130_osu_single_mpr2ct_8_b0r1_4/in X3_Y1 sky130_osu_single_mpr2ct_8_b0r1_3/in
+ s3 vccd1 vssd1 sky130_osu_single_mpr2ct_8_b0r1
Xsky130_osu_single_mpr2ct_8_b0r1_4 sky130_osu_single_mpr2ct_8_b0r1_4/Y0 X4_Y1 sky130_osu_single_mpr2ct_8_b0r1_4/in
+ s4 vccd1 vssd1 sky130_osu_single_mpr2ct_8_b0r1
.ends

* Black-box entry subcircuit for sky130_osu_sc_12T_hs__fill_2 abstract view
.subckt sky130_osu_sc_12T_hs__fill_2
.ends

.subckt scs130hd_mpr2ea_8   B0 A1 R2 A0 R0 R3 B1 R1 vpwr vgnd
X0 vgnd R0 R2 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1 a_826_46# A1 vgnd sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2 a_104_198# A1 vpwr sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X3 vpwr B1 a_104_198# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.165 ps=1.33 w=1 l=0.15
X4 R2 a_104_198# vgnd sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.1885 ps=1.88 w=0.65 l=0.15
X5 a_688_198# B0 a_1706_46# sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.10725 ps=0.98 w=0.65 l=0.15
X6 vpwr a_688_198# a_634_296# sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X7 vgnd R3 R1 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.10725 ps=0.98 w=0.65 l=0.15
X8 a_1706_46# A0 vgnd sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X9 a_634_296# a_104_198# R3 sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.29 ps=2.58 w=1 l=0.15
X10 a_1122_46# B1 a_296_198# sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.1885 ps=1.88 w=0.65 l=0.15
X11 R1 a_296_198# vgnd sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X12 a_296_198# B0 a_1314_46# sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.10725 ps=0.98 w=0.65 l=0.15
X13 vpwr B1 a_1034_296# sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.29 ps=2.58 w=1 l=0.15
X14 a_1034_296# B0 a_296_198# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.165 ps=1.33 w=1 l=0.15
X15 a_1034_296# A0 vpwr sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X16 a_296_198# A1 a_1034_296# sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X17 a_1314_46# A1 vgnd sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X18 vgnd a_688_198# R3 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X19 vgnd A0 a_1122_46# sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X20 R3 a_104_198# vgnd sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.1885 ps=1.88 w=0.65 l=0.15
X21 vpwr R0 a_146_296# sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X22 a_146_296# a_104_198# R2 sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.29 ps=2.58 w=1 l=0.15
X23 a_338_296# a_296_198# vpwr sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X24 R1 R3 a_338_296# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.165 ps=1.33 w=1 l=0.15
X25 vpwr a_688_198# R0 sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.29 ps=2.58 w=1 l=0.15
X26 vpwr B0 a_688_198# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.165 ps=1.33 w=1 l=0.15
X27 a_104_198# B1 a_826_46# sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.10725 ps=0.98 w=0.65 l=0.15
X28 vgnd a_688_198# R0 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.1885 ps=1.88 w=0.65 l=0.15
X29 a_688_198# A0 vpwr sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
.ends

.subckt sky130_osu_single_mpr2ea_8_b0r1 in Y0 Y1 sel vccd1 vssd1
Xsky130_osu_sc_12T_hs__mux2_1_0 scs130hd_mpr2ea_8_0/R1 in sky130_osu_sc_12T_hs__inv_1_1/A
+ vssd1 vccd1 sel sky130_osu_sc_12T_hs__mux2_1
Xsky130_osu_sc_12T_hs__mux2_1_1 in vssd1 scs130hd_mpr2ea_8_0/B1 vssd1 vccd1 sel sky130_osu_sc_12T_hs__mux2_1
Xsky130_osu_sc_12T_hs__inv_1_2 vssd1 sky130_osu_sc_12T_hs__inv_1_2/A Y1 vccd1 sky130_osu_sc_12T_hs__inv_1
Xsky130_osu_sc_12T_hs__inv_1_1 vssd1 sky130_osu_sc_12T_hs__inv_1_1/A sky130_osu_sc_12T_hs__inv_1_2/A
+ vccd1 sky130_osu_sc_12T_hs__inv_1
Xsky130_osu_sc_12T_hs__mux2_1_2 in scs130hd_mpr2ea_8_0/R1 sky130_osu_sc_12T_hs__inv_1_4/A
+ vssd1 vccd1 sel sky130_osu_sc_12T_hs__mux2_1
Xsky130_osu_sc_12T_hs__inv_1_3 vssd1 sky130_osu_sc_12T_hs__inv_1_4/Y Y0 vccd1 sky130_osu_sc_12T_hs__inv_1
Xsky130_osu_sc_12T_hs__inv_1_4 vssd1 sky130_osu_sc_12T_hs__inv_1_4/A sky130_osu_sc_12T_hs__inv_1_4/Y
+ vccd1 sky130_osu_sc_12T_hs__inv_1
Xscs130hd_mpr2ea_8_0   vssd1 scs130hd_mpr2ea_8_0/B1 scs130hd_mpr2ea_8_0/R2
+ scs130hd_mpr2ea_8_0/B1 scs130hd_mpr2ea_8_0/R0 scs130hd_mpr2ea_8_0/R3 scs130hd_mpr2ea_8_0/B1
+ scs130hd_mpr2ea_8_0/R1 vccd1 vssd1 scs130hd_mpr2ea_8
.ends

.subckt sky130_osu_ring_oscillator_mpr2ea_8_b0r1 s1 s2 s3 s4 s5 X2_Y1 X3_Y1 X4_Y1
+ X5_Y1 start vccd1 X1_Y1 vssd1
Xsky130_osu_single_mpr2ea_8_b0r1_2 sky130_osu_single_mpr2ea_8_b0r1_2/in sky130_osu_single_mpr2ea_8_b0r1_3/in
+ X2_Y1 s2 vccd1 vssd1 sky130_osu_single_mpr2ea_8_b0r1
Xsky130_osu_single_mpr2ea_8_b0r1_3 sky130_osu_single_mpr2ea_8_b0r1_3/in sky130_osu_single_mpr2ea_8_b0r1_4/in
+ X3_Y1 s3 vccd1 vssd1 sky130_osu_single_mpr2ea_8_b0r1
Xsky130_osu_single_mpr2ea_8_b0r1_4 sky130_osu_single_mpr2ea_8_b0r1_4/in sky130_osu_single_mpr2ea_8_b0r1_4/Y0
+ X4_Y1 s4 vccd1 vssd1 sky130_osu_single_mpr2ea_8_b0r1
Xsky130_osu_sc_12T_hs__mux2_1_0 vccd1 sky130_osu_sc_12T_hs__mux2_1_0/A0 sky130_osu_sc_12T_hs__mux2_1_0/Y
+ vssd1 vccd1 start sky130_osu_sc_12T_hs__mux2_1
Xsky130_osu_single_mpr2ea_8_b0r1_0 sky130_osu_single_mpr2ea_8_b0r1_4/Y0 sky130_osu_sc_12T_hs__mux2_1_0/A0
+ X5_Y1 s5 vccd1 vssd1 sky130_osu_single_mpr2ea_8_b0r1
Xsky130_osu_single_mpr2ea_8_b0r1_1 sky130_osu_sc_12T_hs__mux2_1_0/Y sky130_osu_single_mpr2ea_8_b0r1_2/in
+ X1_Y1 s1 vccd1 vssd1 sky130_osu_single_mpr2ea_8_b0r1
.ends

.subckt scs130hd_mpr2et_8   B0 A0 B1 R1 R2 R0 R3 A1 vpwr vgnd a_938_46#
X0 a_242_46# A0 vgnd sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1 vgnd A1 a_730_46# sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.10725 ps=0.98 w=0.65 l=0.15
X2 vgnd a_104_198# a_1176_198# sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.1885 ps=1.88 w=0.65 l=0.15
X3 a_450_296# A1 a_634_46# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.165 ps=1.33 w=1 l=0.15
X4 a_2098_296# a_104_198# vpwr sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X5 R3 a_938_46# a_2098_296# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.165 ps=1.33 w=1 l=0.15
X6 vgnd a_104_198# R0 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.1885 ps=1.88 w=0.65 l=0.15
X7 vgnd a_938_46# R3 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.10725 ps=0.98 w=0.65 l=0.15
X8 R3 a_104_198# vgnd sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X9 a_634_46# B0 a_450_296# sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X10 vgnd a_1664_198# R1 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.10725 ps=0.98 w=0.65 l=0.15
X11 vpwr A0 a_450_296# sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.29 ps=2.58 w=1 l=0.15
X12 a_450_296# B1 vpwr sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X13 vgnd A1 a_1026_46# sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X14 vpwr a_104_198# a_1906_296# sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X15 a_1906_296# a_938_46# a_1664_198# sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.29 ps=2.58 w=1 l=0.15
X16 a_104_198# B0 a_242_46# sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.10725 ps=0.98 w=0.65 l=0.15
X17 a_938_46# B1 vpwr sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.29 ps=2.58 w=1 l=0.15
X18 vpwr A1 a_938_46# sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X19 a_1026_46# B1 a_938_46# sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.1885 ps=1.88 w=0.65 l=0.15
X20 a_1218_296# a_1176_198# vpwr sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X21 R2 a_938_46# a_1218_296# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.165 ps=1.33 w=1 l=0.15
X22 vgnd a_938_46# R2 sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.10725 ps=0.98 w=0.65 l=0.15
X23 a_730_46# B0 a_634_46# sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X24 R2 a_1176_198# vgnd sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X25 vgnd a_104_198# a_1664_198# sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X26 a_634_46# B1 a_538_46# sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X27 a_1664_198# a_938_46# vgnd sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.1885 ps=1.88 w=0.65 l=0.15
X28 a_104_198# A0 vpwr sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X29 a_538_46# A0 vgnd sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.1885 ps=1.88 w=0.65 l=0.15
X30 vpwr a_104_198# R0 sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.29 ps=2.58 w=1 l=0.15
X31 vpwr B0 a_104_198# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.165 ps=1.33 w=1 l=0.15
X32 vpwr a_104_198# a_1176_198# sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.29 ps=2.58 w=1 l=0.15
X33 a_1610_296# a_634_46# vpwr sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X34 R1 a_634_46# vgnd sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X35 R1 a_1664_198# a_1610_296# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.165 ps=1.33 w=1 l=0.15
.ends

.subckt sky130_osu_single_mpr2et_8_b0r1 Y0 Y1 sky130_osu_sc_12T_hs__inv_1_2/A sel
+ in vccd1 vssd1
Xscs130hd_mpr2et_8_0   vssd1 scs130hd_mpr2et_8_0/B1 scs130hd_mpr2et_8_0/B1
+ scs130hd_mpr2et_8_0/R1 scs130hd_mpr2et_8_0/R2 scs130hd_mpr2et_8_0/R0 scs130hd_mpr2et_8_0/R3
+ scs130hd_mpr2et_8_0/B1 vccd1 vssd1 m3_1223_853# scs130hd_mpr2et_8
Xsky130_osu_sc_12T_hs__mux2_1_0 scs130hd_mpr2et_8_0/R1 in sky130_osu_sc_12T_hs__inv_1_1/A
+ vssd1 vccd1 sel sky130_osu_sc_12T_hs__mux2_1
Xsky130_osu_sc_12T_hs__mux2_1_1 in vssd1 scs130hd_mpr2et_8_0/B1 vssd1 vccd1 sel sky130_osu_sc_12T_hs__mux2_1
Xsky130_osu_sc_12T_hs__inv_1_1 vssd1 sky130_osu_sc_12T_hs__inv_1_1/A sky130_osu_sc_12T_hs__inv_1_2/A
+ vccd1 sky130_osu_sc_12T_hs__inv_1
Xsky130_osu_sc_12T_hs__inv_1_2 vssd1 sky130_osu_sc_12T_hs__inv_1_2/A Y1 vccd1 sky130_osu_sc_12T_hs__inv_1
Xsky130_osu_sc_12T_hs__mux2_1_2 in scs130hd_mpr2et_8_0/R1 sky130_osu_sc_12T_hs__inv_1_4/A
+ vssd1 vccd1 sel sky130_osu_sc_12T_hs__mux2_1
Xsky130_osu_sc_12T_hs__inv_1_3 vssd1 sky130_osu_sc_12T_hs__inv_1_4/Y Y0 vccd1 sky130_osu_sc_12T_hs__inv_1
Xsky130_osu_sc_12T_hs__inv_1_4 vssd1 sky130_osu_sc_12T_hs__inv_1_4/A sky130_osu_sc_12T_hs__inv_1_4/Y
+ vccd1 sky130_osu_sc_12T_hs__inv_1
.ends

.subckt sky130_osu_ring_oscillator_mpr2et_8_b0r1 s1 s4 s5 X2_Y1 X5_Y1 start vccd1
+ X4_Y1 X1_Y1 sky130_osu_single_mpr2et_8_b0r1_2/sky130_osu_sc_12T_hs__inv_1_2/A X3_Y1
+ s3 vssd1 s2
Xsky130_osu_single_mpr2et_8_b0r1_0 sky130_osu_sc_12T_hs__mux2_1_0/A0 X5_Y1 sky130_osu_single_mpr2et_8_b0r1_0/sky130_osu_sc_12T_hs__inv_1_2/A
+ s5 sky130_osu_single_mpr2et_8_b0r1_4/Y0 vccd1 vssd1 sky130_osu_single_mpr2et_8_b0r1
Xsky130_osu_single_mpr2et_8_b0r1_1 sky130_osu_single_mpr2et_8_b0r1_2/in X1_Y1 sky130_osu_single_mpr2et_8_b0r1_1/sky130_osu_sc_12T_hs__inv_1_2/A
+ s1 sky130_osu_sc_12T_hs__mux2_1_0/Y vccd1 vssd1 sky130_osu_single_mpr2et_8_b0r1
Xsky130_osu_single_mpr2et_8_b0r1_2 sky130_osu_single_mpr2et_8_b0r1_3/in X2_Y1 sky130_osu_single_mpr2et_8_b0r1_2/sky130_osu_sc_12T_hs__inv_1_2/A
+ s2 sky130_osu_single_mpr2et_8_b0r1_2/in vccd1 vssd1 sky130_osu_single_mpr2et_8_b0r1
Xsky130_osu_single_mpr2et_8_b0r1_3 sky130_osu_single_mpr2et_8_b0r1_4/in X3_Y1 sky130_osu_single_mpr2et_8_b0r1_3/sky130_osu_sc_12T_hs__inv_1_2/A
+ s3 sky130_osu_single_mpr2et_8_b0r1_3/in vccd1 vssd1 sky130_osu_single_mpr2et_8_b0r1
Xsky130_osu_single_mpr2et_8_b0r1_4 sky130_osu_single_mpr2et_8_b0r1_4/Y0 X4_Y1 sky130_osu_single_mpr2et_8_b0r1_4/sky130_osu_sc_12T_hs__inv_1_2/A
+ s4 sky130_osu_single_mpr2et_8_b0r1_4/in vccd1 vssd1 sky130_osu_single_mpr2et_8_b0r1
Xsky130_osu_sc_12T_hs__mux2_1_0 vccd1 sky130_osu_sc_12T_hs__mux2_1_0/A0 sky130_osu_sc_12T_hs__mux2_1_0/Y
+ vssd1 vccd1 start sky130_osu_sc_12T_hs__mux2_1
.ends

.subckt sky130_osu_single_mpr2xa_8_b0r1 Y0 Y1 in sel vccd1 vssd1
Xscs130hd_mpr2xa_8_0   scs130hd_mpr2xa_8_0/R0 scs130hd_mpr2xa_8_0/R1 scs130hd_mpr2xa_8_0/R2
+ scs130hd_mpr2xa_8_0/R3 scs130hd_mpr2xa_8_0/B1 vssd1 scs130hd_mpr2xa_8_0/B1 vssd1
+ vccd1 scs130hd_mpr2xa_8_0/B1 scs130hd_mpr2xa_8
Xsky130_osu_sc_12T_hs__mux2_1_0 scs130hd_mpr2xa_8_0/R1 in sky130_osu_sc_12T_hs__inv_1_1/A
+ vssd1 vccd1 sel sky130_osu_sc_12T_hs__mux2_1
Xsky130_osu_sc_12T_hs__mux2_1_1 in vssd1 scs130hd_mpr2xa_8_0/B1 vssd1 vccd1 sel sky130_osu_sc_12T_hs__mux2_1
Xsky130_osu_sc_12T_hs__mux2_1_2 in scs130hd_mpr2xa_8_0/R1 sky130_osu_sc_12T_hs__inv_1_4/A
+ vssd1 vccd1 sel sky130_osu_sc_12T_hs__mux2_1
Xsky130_osu_sc_12T_hs__inv_1_1 vssd1 sky130_osu_sc_12T_hs__inv_1_1/A sky130_osu_sc_12T_hs__inv_1_2/A
+ vccd1 sky130_osu_sc_12T_hs__inv_1
Xsky130_osu_sc_12T_hs__inv_1_2 vssd1 sky130_osu_sc_12T_hs__inv_1_2/A Y1 vccd1 sky130_osu_sc_12T_hs__inv_1
Xsky130_osu_sc_12T_hs__inv_1_3 vssd1 sky130_osu_sc_12T_hs__inv_1_4/Y Y0 vccd1 sky130_osu_sc_12T_hs__inv_1
Xsky130_osu_sc_12T_hs__inv_1_4 vssd1 sky130_osu_sc_12T_hs__inv_1_4/A sky130_osu_sc_12T_hs__inv_1_4/Y
+ vccd1 sky130_osu_sc_12T_hs__inv_1
.ends

.subckt sky130_osu_ring_oscillator_mpr2xa_8_b0r1 X1_Y1 X2_Y1 X3_Y1 X5_Y1 start vccd1
+ s1 s2 s3 s4 s5 X4_Y1 vssd1
Xsky130_osu_single_mpr2xa_8_b0r1_0 sky130_osu_sc_12T_hs__mux2_1_0/A0 X5_Y1 sky130_osu_single_mpr2xa_8_b0r1_4/Y0
+ s5 vccd1 vssd1 sky130_osu_single_mpr2xa_8_b0r1
Xsky130_osu_single_mpr2xa_8_b0r1_1 sky130_osu_single_mpr2xa_8_b0r1_2/in X1_Y1 sky130_osu_sc_12T_hs__mux2_1_0/Y
+ s1 vccd1 vssd1 sky130_osu_single_mpr2xa_8_b0r1
Xsky130_osu_single_mpr2xa_8_b0r1_2 sky130_osu_single_mpr2xa_8_b0r1_3/in X2_Y1 sky130_osu_single_mpr2xa_8_b0r1_2/in
+ s2 vccd1 vssd1 sky130_osu_single_mpr2xa_8_b0r1
Xsky130_osu_single_mpr2xa_8_b0r1_3 sky130_osu_single_mpr2xa_8_b0r1_4/in X3_Y1 sky130_osu_single_mpr2xa_8_b0r1_3/in
+ s3 vccd1 vssd1 sky130_osu_single_mpr2xa_8_b0r1
Xsky130_osu_single_mpr2xa_8_b0r1_4 sky130_osu_single_mpr2xa_8_b0r1_4/Y0 X4_Y1 sky130_osu_single_mpr2xa_8_b0r1_4/in
+ s4 vccd1 vssd1 sky130_osu_single_mpr2xa_8_b0r1
Xsky130_osu_sc_12T_hs__mux2_1_0 vccd1 sky130_osu_sc_12T_hs__mux2_1_0/A0 sky130_osu_sc_12T_hs__mux2_1_0/Y
+ vssd1 vccd1 start sky130_osu_sc_12T_hs__mux2_1
.ends

.subckt sky130_fd_sc_hd__conb_1 LO HI   VGND VPWR
R0 VPWR HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
R1 LO VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
.ends

.subckt sky130_osu_single_mpr2ca_8_b0r2 Y0 in Y1 sel vssd1 scs130hd_mpr2ca_8_0/B1
+ vccd1
Xsky130_osu_sc_12T_hs__mux2_1_0 scs130hd_mpr2ca_8_0/R2 in sky130_osu_sc_12T_hs__inv_1_1/A
+ vssd1 vccd1 sel sky130_osu_sc_12T_hs__mux2_1
Xsky130_osu_sc_12T_hs__mux2_1_1 in vssd1 scs130hd_mpr2ca_8_0/B1 vssd1 vccd1 sel sky130_osu_sc_12T_hs__mux2_1
Xscs130hd_mpr2ca_8_0 scs130hd_mpr2ca_8_0/B1 scs130hd_mpr2ca_8_0/B1 scs130hd_mpr2ca_8_0/R3
+ scs130hd_mpr2ca_8_0/R1 scs130hd_mpr2ca_8_0/R0 vssd1 scs130hd_mpr2ca_8_0/B1 scs130hd_mpr2ca_8_0/R2
+ vccd1  vssd1 vssd1  scs130hd_mpr2ca_8
Xsky130_osu_sc_12T_hs__mux2_1_2 in scs130hd_mpr2ca_8_0/R2 sky130_osu_sc_12T_hs__inv_1_4/A
+ vssd1 vccd1 sel sky130_osu_sc_12T_hs__mux2_1
Xsky130_osu_sc_12T_hs__inv_1_1 vssd1 sky130_osu_sc_12T_hs__inv_1_1/A sky130_osu_sc_12T_hs__inv_1_2/A
+ vccd1 sky130_osu_sc_12T_hs__inv_1
Xsky130_osu_sc_12T_hs__inv_1_2 vssd1 sky130_osu_sc_12T_hs__inv_1_2/A Y1 vccd1 sky130_osu_sc_12T_hs__inv_1
Xsky130_osu_sc_12T_hs__inv_1_3 vssd1 sky130_osu_sc_12T_hs__inv_1_4/Y Y0 vccd1 sky130_osu_sc_12T_hs__inv_1
Xsky130_osu_sc_12T_hs__inv_1_4 vssd1 sky130_osu_sc_12T_hs__inv_1_4/A sky130_osu_sc_12T_hs__inv_1_4/Y
+ vccd1 sky130_osu_sc_12T_hs__inv_1
.ends

.subckt sky130_osu_ring_oscillator_mpr2ca_8_b0r2 s1 s5 X5_Y1 X2_Y1 X1_Y1 start vccd1
+ X4_Y1 s4 X3_Y1 vssd1 s3 s2
Xsky130_osu_single_mpr2ca_8_b0r2_4 sky130_osu_single_mpr2ca_8_b0r2_4/Y0 sky130_osu_single_mpr2ca_8_b0r2_4/in
+ X4_Y1 s4 vssd1 sky130_osu_single_mpr2ca_8_b0r2_4/scs130hd_mpr2ca_8_0/B1 vccd1 sky130_osu_single_mpr2ca_8_b0r2
Xsky130_osu_sc_12T_hs__mux2_1_0 vccd1 sky130_osu_sc_12T_hs__mux2_1_0/A0 sky130_osu_sc_12T_hs__mux2_1_0/Y
+ vssd1 vccd1 start sky130_osu_sc_12T_hs__mux2_1
Xsky130_osu_single_mpr2ca_8_b0r2_0 sky130_osu_sc_12T_hs__mux2_1_0/A0 sky130_osu_single_mpr2ca_8_b0r2_4/Y0
+ X5_Y1 s5 vssd1 sky130_osu_single_mpr2ca_8_b0r2_0/scs130hd_mpr2ca_8_0/B1 vccd1 sky130_osu_single_mpr2ca_8_b0r2
Xsky130_osu_single_mpr2ca_8_b0r2_1 sky130_osu_single_mpr2ca_8_b0r2_2/in sky130_osu_sc_12T_hs__mux2_1_0/Y
+ X1_Y1 s1 vssd1 sky130_osu_single_mpr2ca_8_b0r2_1/scs130hd_mpr2ca_8_0/B1 vccd1 sky130_osu_single_mpr2ca_8_b0r2
Xsky130_osu_single_mpr2ca_8_b0r2_2 sky130_osu_single_mpr2ca_8_b0r2_3/in sky130_osu_single_mpr2ca_8_b0r2_2/in
+ X2_Y1 s2 vssd1 sky130_osu_single_mpr2ca_8_b0r2_2/scs130hd_mpr2ca_8_0/B1 vccd1 sky130_osu_single_mpr2ca_8_b0r2
Xsky130_osu_single_mpr2ca_8_b0r2_3 sky130_osu_single_mpr2ca_8_b0r2_4/in sky130_osu_single_mpr2ca_8_b0r2_3/in
+ X3_Y1 s3 vssd1 sky130_osu_single_mpr2ca_8_b0r2_3/scs130hd_mpr2ca_8_0/B1 vccd1 sky130_osu_single_mpr2ca_8_b0r2
.ends

.subckt sky130_osu_single_mpr2ct_8_b0r2 Y0 Y1 in sel vccd1 vssd1
Xsky130_osu_sc_12T_hs__mux2_1_0 scs130hd_mpr2ct_8_1/R2 in sky130_osu_sc_12T_hs__inv_1_1/A
+ vssd1 vccd1 sel sky130_osu_sc_12T_hs__mux2_1
Xsky130_osu_sc_12T_hs__mux2_1_1 in vssd1 scs130hd_mpr2ct_8_1/B1 vssd1 vccd1 sel sky130_osu_sc_12T_hs__mux2_1
Xsky130_osu_sc_12T_hs__mux2_1_2 in scs130hd_mpr2ct_8_1/R2 sky130_osu_sc_12T_hs__inv_1_4/A
+ vssd1 vccd1 sel sky130_osu_sc_12T_hs__mux2_1
Xsky130_osu_sc_12T_hs__inv_1_1 vssd1 sky130_osu_sc_12T_hs__inv_1_1/A sky130_osu_sc_12T_hs__inv_1_2/A
+ vccd1 sky130_osu_sc_12T_hs__inv_1
Xsky130_osu_sc_12T_hs__inv_1_2 vssd1 sky130_osu_sc_12T_hs__inv_1_2/A Y1 vccd1 sky130_osu_sc_12T_hs__inv_1
Xsky130_osu_sc_12T_hs__inv_1_3 vssd1 sky130_osu_sc_12T_hs__inv_1_4/Y Y0 vccd1 sky130_osu_sc_12T_hs__inv_1
Xsky130_osu_sc_12T_hs__inv_1_4 vssd1 sky130_osu_sc_12T_hs__inv_1_4/A sky130_osu_sc_12T_hs__inv_1_4/Y
+ vccd1 sky130_osu_sc_12T_hs__inv_1
Xscs130hd_mpr2ct_8_1 scs130hd_mpr2ct_8_1/B1 scs130hd_mpr2ct_8_1/B1 vssd1 scs130hd_mpr2ct_8_1/B1
+ scs130hd_mpr2ct_8_1/R0 scs130hd_mpr2ct_8_1/R1 scs130hd_mpr2ct_8_1/R2 scs130hd_mpr2ct_8_1/R3
+ vccd1  vssd1 vssd1  scs130hd_mpr2ct_8
.ends

.subckt sky130_osu_ring_oscillator_mpr2ct_8_b0r2 s1 s2 s3 X3_Y1 X2_Y1 X1_Y1 s5 s4
+ start vccd1 X4_Y1 X5_Y1 vssd1
Xsky130_osu_single_mpr2ct_8_b0r2_0 sky130_osu_sc_12T_hs__mux2_1_0/A0 X5_Y1 sky130_osu_single_mpr2ct_8_b0r2_4/Y0
+ s5 vccd1 vssd1 sky130_osu_single_mpr2ct_8_b0r2
Xsky130_osu_single_mpr2ct_8_b0r2_1 sky130_osu_single_mpr2ct_8_b0r2_2/in X1_Y1 sky130_osu_sc_12T_hs__mux2_1_0/Y
+ s1 vccd1 vssd1 sky130_osu_single_mpr2ct_8_b0r2
Xsky130_osu_single_mpr2ct_8_b0r2_2 sky130_osu_single_mpr2ct_8_b0r2_3/in X2_Y1 sky130_osu_single_mpr2ct_8_b0r2_2/in
+ s2 vccd1 vssd1 sky130_osu_single_mpr2ct_8_b0r2
Xsky130_osu_single_mpr2ct_8_b0r2_3 sky130_osu_single_mpr2ct_8_b0r2_4/in X3_Y1 sky130_osu_single_mpr2ct_8_b0r2_3/in
+ s3 vccd1 vssd1 sky130_osu_single_mpr2ct_8_b0r2
Xsky130_osu_single_mpr2ct_8_b0r2_4 sky130_osu_single_mpr2ct_8_b0r2_4/Y0 X4_Y1 sky130_osu_single_mpr2ct_8_b0r2_4/in
+ s4 vccd1 vssd1 sky130_osu_single_mpr2ct_8_b0r2
Xsky130_osu_sc_12T_hs__mux2_1_0 vccd1 sky130_osu_sc_12T_hs__mux2_1_0/A0 sky130_osu_sc_12T_hs__mux2_1_0/Y
+ vssd1 vccd1 start sky130_osu_sc_12T_hs__mux2_1
.ends

.subckt sky130_osu_single_mpr2ea_8_b0r2 in Y0 Y1 sky130_osu_sc_12T_hs__inv_1_2/A sel
+ sky130_osu_sc_12T_hs__inv_1_1/A vccd1 vssd1
Xsky130_osu_sc_12T_hs__mux2_1_0 scs130hd_mpr2ea_8_0/R2 in sky130_osu_sc_12T_hs__inv_1_1/A
+ vssd1 vccd1 sel sky130_osu_sc_12T_hs__mux2_1
Xsky130_osu_sc_12T_hs__mux2_1_1 in vssd1 scs130hd_mpr2ea_8_0/B1 vssd1 vccd1 sel sky130_osu_sc_12T_hs__mux2_1
Xsky130_osu_sc_12T_hs__inv_1_2 vssd1 sky130_osu_sc_12T_hs__inv_1_2/A Y1 vccd1 sky130_osu_sc_12T_hs__inv_1
Xsky130_osu_sc_12T_hs__inv_1_1 vssd1 sky130_osu_sc_12T_hs__inv_1_1/A sky130_osu_sc_12T_hs__inv_1_2/A
+ vccd1 sky130_osu_sc_12T_hs__inv_1
Xsky130_osu_sc_12T_hs__mux2_1_2 in scs130hd_mpr2ea_8_0/R2 sky130_osu_sc_12T_hs__inv_1_4/A
+ vssd1 vccd1 sel sky130_osu_sc_12T_hs__mux2_1
Xsky130_osu_sc_12T_hs__inv_1_3 vssd1 sky130_osu_sc_12T_hs__inv_1_4/Y Y0 vccd1 sky130_osu_sc_12T_hs__inv_1
Xsky130_osu_sc_12T_hs__inv_1_4 vssd1 sky130_osu_sc_12T_hs__inv_1_4/A sky130_osu_sc_12T_hs__inv_1_4/Y
+ vccd1 sky130_osu_sc_12T_hs__inv_1
Xscs130hd_mpr2ea_8_0   vssd1 scs130hd_mpr2ea_8_0/B1 scs130hd_mpr2ea_8_0/R2
+ scs130hd_mpr2ea_8_0/B1 scs130hd_mpr2ea_8_0/R0 scs130hd_mpr2ea_8_0/R3 scs130hd_mpr2ea_8_0/B1
+ scs130hd_mpr2ea_8_0/R1 vccd1 vssd1 scs130hd_mpr2ea_8
.ends

.subckt sky130_osu_ring_oscillator_mpr2ea_8_b0r2 s1 s3 s4 X1_Y1 X2_Y1 X4_Y1 X5_Y1
+ start vccd1 sky130_osu_single_mpr2ea_8_b0r2_0/sky130_osu_sc_12T_hs__inv_1_2/A X3_Y1
+ s5 sky130_osu_single_mpr2ea_8_b0r2_0/sky130_osu_sc_12T_hs__inv_1_1/A s2 vssd1
Xsky130_osu_single_mpr2ea_8_b0r2_1 sky130_osu_sc_12T_hs__mux2_1_0/Y sky130_osu_single_mpr2ea_8_b0r2_2/in
+ X1_Y1 sky130_osu_single_mpr2ea_8_b0r2_1/sky130_osu_sc_12T_hs__inv_1_2/A s1 sky130_osu_single_mpr2ea_8_b0r2_1/sky130_osu_sc_12T_hs__inv_1_1/A
+ vccd1 vssd1 sky130_osu_single_mpr2ea_8_b0r2
Xsky130_osu_single_mpr2ea_8_b0r2_0 sky130_osu_single_mpr2ea_8_b0r2_4/Y0 sky130_osu_sc_12T_hs__mux2_1_0/A0
+ X5_Y1 sky130_osu_single_mpr2ea_8_b0r2_0/sky130_osu_sc_12T_hs__inv_1_2/A s5 sky130_osu_single_mpr2ea_8_b0r2_0/sky130_osu_sc_12T_hs__inv_1_1/A
+ vccd1 vssd1 sky130_osu_single_mpr2ea_8_b0r2
Xsky130_osu_single_mpr2ea_8_b0r2_2 sky130_osu_single_mpr2ea_8_b0r2_2/in sky130_osu_single_mpr2ea_8_b0r2_3/in
+ X2_Y1 sky130_osu_single_mpr2ea_8_b0r2_2/sky130_osu_sc_12T_hs__inv_1_2/A s2 sky130_osu_single_mpr2ea_8_b0r2_2/sky130_osu_sc_12T_hs__inv_1_1/A
+ vccd1 vssd1 sky130_osu_single_mpr2ea_8_b0r2
Xsky130_osu_sc_12T_hs__mux2_1_0 vccd1 sky130_osu_sc_12T_hs__mux2_1_0/A0 sky130_osu_sc_12T_hs__mux2_1_0/Y
+ vssd1 vccd1 start sky130_osu_sc_12T_hs__mux2_1
Xsky130_osu_single_mpr2ea_8_b0r2_3 sky130_osu_single_mpr2ea_8_b0r2_3/in sky130_osu_single_mpr2ea_8_b0r2_4/in
+ X3_Y1 sky130_osu_single_mpr2ea_8_b0r2_3/sky130_osu_sc_12T_hs__inv_1_2/A s3 sky130_osu_single_mpr2ea_8_b0r2_3/sky130_osu_sc_12T_hs__inv_1_1/A
+ vccd1 vssd1 sky130_osu_single_mpr2ea_8_b0r2
Xsky130_osu_single_mpr2ea_8_b0r2_4 sky130_osu_single_mpr2ea_8_b0r2_4/in sky130_osu_single_mpr2ea_8_b0r2_4/Y0
+ X4_Y1 sky130_osu_single_mpr2ea_8_b0r2_4/sky130_osu_sc_12T_hs__inv_1_2/A s4 sky130_osu_single_mpr2ea_8_b0r2_4/sky130_osu_sc_12T_hs__inv_1_1/A
+ vccd1 vssd1 sky130_osu_single_mpr2ea_8_b0r2
.ends

.subckt sky130_osu_single_mpr2et_8_b0r2 Y0 Y1 sky130_osu_sc_12T_hs__inv_1_2/A sky130_osu_sc_12T_hs__inv_1_4/A
+ sel in sky130_osu_sc_12T_hs__inv_1_4/Y vccd1 vssd1
Xscs130hd_mpr2et_8_0   vssd1 scs130hd_mpr2et_8_0/B1 scs130hd_mpr2et_8_0/B1
+ scs130hd_mpr2et_8_0/R1 scs130hd_mpr2et_8_0/R2 scs130hd_mpr2et_8_0/R0 scs130hd_mpr2et_8_0/R3
+ scs130hd_mpr2et_8_0/B1 vccd1 vssd1 scs130hd_mpr2et_8_0/a_938_46# scs130hd_mpr2et_8
Xsky130_osu_sc_12T_hs__mux2_1_0 scs130hd_mpr2et_8_0/R2 in sky130_osu_sc_12T_hs__inv_1_1/A
+ vssd1 vccd1 sel sky130_osu_sc_12T_hs__mux2_1
Xsky130_osu_sc_12T_hs__mux2_1_1 in vssd1 scs130hd_mpr2et_8_0/B1 vssd1 vccd1 sel sky130_osu_sc_12T_hs__mux2_1
Xsky130_osu_sc_12T_hs__inv_1_1 vssd1 sky130_osu_sc_12T_hs__inv_1_1/A sky130_osu_sc_12T_hs__inv_1_2/A
+ vccd1 sky130_osu_sc_12T_hs__inv_1
Xsky130_osu_sc_12T_hs__inv_1_2 vssd1 sky130_osu_sc_12T_hs__inv_1_2/A Y1 vccd1 sky130_osu_sc_12T_hs__inv_1
Xsky130_osu_sc_12T_hs__mux2_1_2 in scs130hd_mpr2et_8_0/R2 sky130_osu_sc_12T_hs__inv_1_4/A
+ vssd1 vccd1 sel sky130_osu_sc_12T_hs__mux2_1
Xsky130_osu_sc_12T_hs__inv_1_3 vssd1 sky130_osu_sc_12T_hs__inv_1_4/Y Y0 vccd1 sky130_osu_sc_12T_hs__inv_1
Xsky130_osu_sc_12T_hs__inv_1_4 vssd1 sky130_osu_sc_12T_hs__inv_1_4/A sky130_osu_sc_12T_hs__inv_1_4/Y
+ vccd1 sky130_osu_sc_12T_hs__inv_1
.ends

.subckt sky130_osu_ring_oscillator_mpr2et_8_b0r2 s1 s2 s3 s5 X2_Y1 X5_Y1 start vccd1
+ sky130_osu_single_mpr2et_8_b0r2_1/sky130_osu_sc_12T_hs__inv_1_4/A sky130_osu_single_mpr2et_8_b0r2_2/sky130_osu_sc_12T_hs__inv_1_2/A
+ X4_Y1 X1_Y1 sky130_osu_single_mpr2et_8_b0r2_1/sky130_osu_sc_12T_hs__inv_1_4/Y X3_Y1
+ s4 vssd1
Xsky130_osu_sc_12T_hs__mux2_1_0 vccd1 sky130_osu_sc_12T_hs__mux2_1_0/A0 sky130_osu_sc_12T_hs__mux2_1_0/Y
+ vssd1 vccd1 start sky130_osu_sc_12T_hs__mux2_1
Xsky130_osu_single_mpr2et_8_b0r2_0 sky130_osu_sc_12T_hs__mux2_1_0/A0 X5_Y1 sky130_osu_single_mpr2et_8_b0r2_0/sky130_osu_sc_12T_hs__inv_1_2/A
+ sky130_osu_single_mpr2et_8_b0r2_0/sky130_osu_sc_12T_hs__inv_1_4/A s5 sky130_osu_single_mpr2et_8_b0r2_4/Y0
+ sky130_osu_single_mpr2et_8_b0r2_0/sky130_osu_sc_12T_hs__inv_1_4/Y vccd1 vssd1 sky130_osu_single_mpr2et_8_b0r2
Xsky130_osu_single_mpr2et_8_b0r2_2 sky130_osu_single_mpr2et_8_b0r2_3/in X2_Y1 sky130_osu_single_mpr2et_8_b0r2_2/sky130_osu_sc_12T_hs__inv_1_2/A
+ sky130_osu_single_mpr2et_8_b0r2_2/sky130_osu_sc_12T_hs__inv_1_4/A s2 sky130_osu_single_mpr2et_8_b0r2_2/in
+ sky130_osu_single_mpr2et_8_b0r2_2/sky130_osu_sc_12T_hs__inv_1_4/Y vccd1 vssd1 sky130_osu_single_mpr2et_8_b0r2
Xsky130_osu_single_mpr2et_8_b0r2_1 sky130_osu_single_mpr2et_8_b0r2_2/in X1_Y1 sky130_osu_single_mpr2et_8_b0r2_1/sky130_osu_sc_12T_hs__inv_1_2/A
+ sky130_osu_single_mpr2et_8_b0r2_1/sky130_osu_sc_12T_hs__inv_1_4/A s1 sky130_osu_sc_12T_hs__mux2_1_0/Y
+ sky130_osu_single_mpr2et_8_b0r2_1/sky130_osu_sc_12T_hs__inv_1_4/Y vccd1 vssd1 sky130_osu_single_mpr2et_8_b0r2
Xsky130_osu_single_mpr2et_8_b0r2_3 sky130_osu_single_mpr2et_8_b0r2_4/in X3_Y1 sky130_osu_single_mpr2et_8_b0r2_3/sky130_osu_sc_12T_hs__inv_1_2/A
+ sky130_osu_single_mpr2et_8_b0r2_3/sky130_osu_sc_12T_hs__inv_1_4/A s3 sky130_osu_single_mpr2et_8_b0r2_3/in
+ sky130_osu_single_mpr2et_8_b0r2_3/sky130_osu_sc_12T_hs__inv_1_4/Y vccd1 vssd1 sky130_osu_single_mpr2et_8_b0r2
Xsky130_osu_single_mpr2et_8_b0r2_4 sky130_osu_single_mpr2et_8_b0r2_4/Y0 X4_Y1 sky130_osu_single_mpr2et_8_b0r2_4/sky130_osu_sc_12T_hs__inv_1_2/A
+ sky130_osu_single_mpr2et_8_b0r2_4/sky130_osu_sc_12T_hs__inv_1_4/A s4 sky130_osu_single_mpr2et_8_b0r2_4/in
+ sky130_osu_single_mpr2et_8_b0r2_4/sky130_osu_sc_12T_hs__inv_1_4/Y vccd1 vssd1 sky130_osu_single_mpr2et_8_b0r2
.ends

.subckt user_project_wrapper    
+ io_in[0]        
+   io_in[1]      
+     io_in[2]    
+     io_in[3] io_in[4] io_in[5] io_in[6] io_in[7]
+ io_in[8] io_in[9]      
+ io_out[0]       
+   vccd1      vssd1  
Xmprj3 ro1/X3_Y1 mprj5/data_in[15] mprj5/data_in[15] mprj5/data_in[15] mprj5/data_in[15]
+ mprj5/data_in[15] mprj5/data_in[15] ro2/X3_Y1 ro3/X3_Y1 ro4/X3_Y1 ro5/X3_Y1 ro6/X3_Y1
+ ro7/X3_Y1 ro8/X3_Y1 ro9/X3_Y1 ro10/X3_Y1 io_in[6] io_in[7] io_in[8] io_in[9] io_out[0]
+ vssd1 vccd1 mux16x1_project
Xmprj4 ro1/X4_Y1 mprj5/data_in[15] mprj5/data_in[15] mprj5/data_in[15] mprj5/data_in[15]
+ mprj5/data_in[15] mprj5/data_in[15] ro2/X4_Y1 ro3/X4_Y1 ro4/X4_Y1 ro5/X4_Y1 ro6/X4_Y1
+ ro7/X4_Y1 ro8/X4_Y1 ro9/X4_Y1 ro10/X4_Y1 io_in[6] io_in[7] io_in[8] io_in[9] io_out[0]
+ vssd1 vccd1 mux16x1_project
Xmprj5 ro1/X5_Y1 mprj5/data_in[15] mprj5/data_in[15] mprj5/data_in[15] mprj5/data_in[15]
+ mprj5/data_in[15] mprj5/data_in[15] ro2/X5_Y1 ro3/X5_Y1 ro4/X5_Y1 ro5/X5_Y1 ro6/X5_Y1
+ ro7/X5_Y1 ro8/X5_Y1 ro9/X5_Y1 ro10/X5_Y1 io_in[6] io_in[7] io_in[8] io_in[9] io_out[0]
+ vssd1 vccd1 mux16x1_project
Xro1 io_in[3] io_in[4] ro1/X5_Y1 ro1/X4_Y1 ro1/X3_Y1 ro1/X2_Y1 ro1/X1_Y1 io_in[5]
+ vccd1 io_in[1] io_in[2] io_in[0] vssd1 sky130_osu_ring_oscillator_mpr2ca_8_b0r1
Xro10 io_in[0] io_in[2] io_in[3] io_in[4] ro10/X1_Y1 ro10/X5_Y1 io_in[5] vccd1 ro10/X4_Y1
+ ro10/X3_Y1 io_in[1] ro10/X2_Y1 vssd1 sky130_osu_ring_oscillator_mpr2xa_8_b0r2
Xro2 io_in[0] io_in[1] io_in[2] ro2/X5_Y1 ro2/X4_Y1 ro2/X3_Y1 ro2/X2_Y1 ro2/X1_Y1
+ io_in[4] io_in[3] io_in[5] vccd1 vssd1 sky130_osu_ring_oscillator_mpr2ct_8_b0r1
Xro3 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] ro3/X2_Y1 ro3/X3_Y1 ro3/X4_Y1 ro3/X5_Y1
+ io_in[5] vccd1 ro3/X1_Y1 vssd1 sky130_osu_ring_oscillator_mpr2ea_8_b0r1
Xro4 io_in[0] io_in[3] io_in[4] ro4/X2_Y1 ro4/X5_Y1 io_in[5] vccd1 ro4/X4_Y1 ro4/X1_Y1
+ ro4/X2_Y1 ro4/X3_Y1 io_in[2] vssd1 io_in[1] sky130_osu_ring_oscillator_mpr2et_8_b0r1
Xro5 ro5/X1_Y1 ro5/X2_Y1 ro5/X3_Y1 ro5/X5_Y1 io_in[5] vccd1 io_in[0] io_in[1] io_in[2]
+ io_in[3] io_in[4] ro5/X4_Y1 vssd1 sky130_osu_ring_oscillator_mpr2xa_8_b0r1
XTIE_ZERO_zero_ mprj5/data_in[15] TIE_ZERO_zero_/HI   TIE_ZERO_zero_/VGND
+ TIE_ZERO_zero_/VPWR sky130_fd_sc_hd__conb_1
Xro6 io_in[0] io_in[4] ro6/X5_Y1 ro6/X2_Y1 ro6/X1_Y1 io_in[5] vccd1 ro6/X4_Y1 io_in[3]
+ ro6/X3_Y1 vssd1 io_in[2] io_in[1] sky130_osu_ring_oscillator_mpr2ca_8_b0r2
Xro7 io_in[0] io_in[1] io_in[2] ro7/X3_Y1 ro7/X2_Y1 ro7/X1_Y1 io_in[4] io_in[3] io_in[5]
+ vccd1 ro7/X4_Y1 ro7/X5_Y1 vssd1 sky130_osu_ring_oscillator_mpr2ct_8_b0r2
Xro8 io_in[0] io_in[2] io_in[3] ro8/X1_Y1 ro8/X2_Y1 ro8/X4_Y1 ro8/X5_Y1 io_in[5] vccd1
+ io_in[4] ro8/X3_Y1 io_in[4] io_in[4] io_in[1] vssd1 sky130_osu_ring_oscillator_mpr2ea_8_b0r2
Xro9 io_in[0] io_in[1] io_in[2] io_in[4] ro9/X2_Y1 ro9/X5_Y1 io_in[5] vccd1 io_in[0]
+ ro9/X2_Y1 ro9/X4_Y1 ro9/X1_Y1 io_in[0] ro9/X3_Y1 io_in[3] vssd1 sky130_osu_ring_oscillator_mpr2et_8_b0r2
Xmprj1 ro1/X1_Y1 mprj5/data_in[15] mprj5/data_in[15] mprj5/data_in[15] mprj5/data_in[15]
+ mprj5/data_in[15] mprj5/data_in[15] ro2/X1_Y1 ro3/X1_Y1 ro4/X1_Y1 ro5/X1_Y1 ro6/X1_Y1
+ ro7/X1_Y1 ro8/X1_Y1 ro9/X1_Y1 ro10/X1_Y1 io_in[6] io_in[7] io_in[8] io_in[9] io_out[0]
+ vssd1 vccd1 mux16x1_project
Xmprj2 ro1/X2_Y1 mprj5/data_in[15] mprj5/data_in[15] mprj5/data_in[15] mprj5/data_in[15]
+ mprj5/data_in[15] mprj5/data_in[15] ro2/X2_Y1 ro3/X2_Y1 ro4/X2_Y1 ro5/X2_Y1 ro6/X2_Y1
+ ro7/X2_Y1 ro8/X2_Y1 ro9/X2_Y1 ro10/X2_Y1 io_in[6] io_in[7] io_in[8] io_in[9] io_out[0]
+ vssd1 vccd1 mux16x1_project
.ends

