magic
tech sky130A
magscale 1 2
timestamp 1699152421
<< viali >>
rect 2053 19465 2087 19499
rect 3985 19465 4019 19499
rect 1501 19397 1535 19431
rect 6561 19397 6595 19431
rect 1961 19329 1995 19363
rect 2237 19329 2271 19363
rect 3801 19329 3835 19363
rect 8493 19329 8527 19363
rect 1685 19261 1719 19295
rect 6377 19193 6411 19227
rect 1777 19125 1811 19159
rect 8309 19125 8343 19159
rect 1409 18717 1443 18751
rect 1593 18581 1627 18615
rect 1409 17153 1443 17187
rect 1593 16949 1627 16983
rect 1409 16065 1443 16099
rect 1593 16065 1627 16099
rect 2329 15997 2363 16031
rect 2446 15997 2480 16031
rect 2605 15997 2639 16031
rect 2053 15929 2087 15963
rect 3249 15861 3283 15895
rect 1593 15657 1627 15691
rect 1409 15453 1443 15487
rect 1409 14977 1443 15011
rect 1593 14977 1627 15011
rect 2605 14977 2639 15011
rect 2329 14909 2363 14943
rect 2446 14909 2480 14943
rect 2053 14841 2087 14875
rect 3249 14773 3283 14807
rect 1593 14569 1627 14603
rect 2789 14433 2823 14467
rect 2881 14433 2915 14467
rect 1409 14365 1443 14399
rect 2697 14297 2731 14331
rect 2329 14229 2363 14263
rect 1593 13481 1627 13515
rect 1409 13277 1443 13311
rect 2329 12189 2363 12223
rect 2513 12189 2547 12223
rect 2421 12053 2455 12087
rect 1593 11849 1627 11883
rect 1409 11713 1443 11747
rect 2421 11713 2455 11747
rect 2789 11713 2823 11747
rect 2973 11645 3007 11679
rect 2513 11577 2547 11611
rect 7113 11101 7147 11135
rect 8217 11033 8251 11067
rect 1409 10625 1443 10659
rect 1593 10421 1627 10455
rect 1593 9537 1627 9571
rect 1685 9537 1719 9571
rect 1501 9469 1535 9503
rect 1869 9333 1903 9367
rect 1409 8925 1443 8959
rect 1593 8789 1627 8823
rect 1777 8585 1811 8619
rect 2145 8585 2179 8619
rect 2329 8585 2363 8619
rect 2697 8585 2731 8619
rect 2421 8449 2455 8483
rect 2605 8449 2639 8483
rect 1593 8381 1627 8415
rect 1685 8381 1719 8415
rect 2697 8381 2731 8415
rect 2513 8245 2547 8279
rect 1777 8041 1811 8075
rect 1961 8041 1995 8075
rect 1409 7973 1443 8007
rect 1777 7701 1811 7735
rect 1593 7497 1627 7531
rect 1409 7361 1443 7395
rect 2053 6817 2087 6851
rect 1685 6749 1719 6783
rect 2145 6749 2179 6783
rect 1777 6613 1811 6647
rect 1869 6613 1903 6647
rect 2329 6613 2363 6647
rect 2237 6409 2271 6443
rect 1593 6273 1627 6307
rect 2421 6273 2455 6307
rect 2513 6273 2547 6307
rect 2605 6273 2639 6307
rect 1869 6205 1903 6239
rect 2145 6137 2179 6171
rect 1685 6069 1719 6103
rect 1593 5865 1627 5899
rect 1869 5865 1903 5899
rect 1409 5661 1443 5695
rect 1777 5661 1811 5695
rect 1961 5661 1995 5695
rect 2145 5321 2179 5355
rect 1777 5185 1811 5219
rect 1501 5117 1535 5151
rect 1685 5117 1719 5151
rect 1593 4777 1627 4811
rect 1409 4573 1443 4607
rect 1593 3689 1627 3723
rect 1409 3485 1443 3519
rect 1869 2601 1903 2635
rect 1593 2533 1627 2567
rect 1409 2397 1443 2431
rect 1685 2397 1719 2431
<< metal1 >>
rect 1104 19610 8992 19632
rect 1104 19558 2882 19610
rect 2934 19558 2946 19610
rect 2998 19558 3010 19610
rect 3062 19558 3074 19610
rect 3126 19558 3138 19610
rect 3190 19558 4814 19610
rect 4866 19558 4878 19610
rect 4930 19558 4942 19610
rect 4994 19558 5006 19610
rect 5058 19558 5070 19610
rect 5122 19558 6746 19610
rect 6798 19558 6810 19610
rect 6862 19558 6874 19610
rect 6926 19558 6938 19610
rect 6990 19558 7002 19610
rect 7054 19558 8678 19610
rect 8730 19558 8742 19610
rect 8794 19558 8806 19610
rect 8858 19558 8870 19610
rect 8922 19558 8934 19610
rect 8986 19558 8992 19610
rect 1104 19536 8992 19558
rect 1118 19456 1124 19508
rect 1176 19496 1182 19508
rect 1176 19468 1624 19496
rect 1176 19456 1182 19468
rect 1394 19388 1400 19440
rect 1452 19428 1458 19440
rect 1489 19431 1547 19437
rect 1489 19428 1501 19431
rect 1452 19400 1501 19428
rect 1452 19388 1458 19400
rect 1489 19397 1501 19400
rect 1535 19397 1547 19431
rect 1596 19428 1624 19468
rect 1762 19456 1768 19508
rect 1820 19496 1826 19508
rect 2041 19499 2099 19505
rect 2041 19496 2053 19499
rect 1820 19468 2053 19496
rect 1820 19456 1826 19468
rect 2041 19465 2053 19468
rect 2087 19465 2099 19499
rect 2041 19459 2099 19465
rect 2498 19456 2504 19508
rect 2556 19496 2562 19508
rect 3973 19499 4031 19505
rect 3973 19496 3985 19499
rect 2556 19468 3985 19496
rect 2556 19456 2562 19468
rect 3973 19465 3985 19468
rect 4019 19465 4031 19499
rect 3973 19459 4031 19465
rect 8570 19456 8576 19508
rect 8628 19456 8634 19508
rect 1596 19400 2268 19428
rect 1489 19391 1547 19397
rect 1026 19320 1032 19372
rect 1084 19360 1090 19372
rect 2240 19369 2268 19400
rect 6178 19388 6184 19440
rect 6236 19428 6242 19440
rect 6549 19431 6607 19437
rect 6549 19428 6561 19431
rect 6236 19400 6561 19428
rect 6236 19388 6242 19400
rect 6549 19397 6561 19400
rect 6595 19397 6607 19431
rect 6549 19391 6607 19397
rect 1949 19363 2007 19369
rect 1949 19360 1961 19363
rect 1084 19332 1961 19360
rect 1084 19320 1090 19332
rect 1949 19329 1961 19332
rect 1995 19329 2007 19363
rect 1949 19323 2007 19329
rect 2225 19363 2283 19369
rect 2225 19329 2237 19363
rect 2271 19329 2283 19363
rect 2225 19323 2283 19329
rect 3694 19320 3700 19372
rect 3752 19360 3758 19372
rect 3789 19363 3847 19369
rect 3789 19360 3801 19363
rect 3752 19332 3801 19360
rect 3752 19320 3758 19332
rect 3789 19329 3801 19332
rect 3835 19329 3847 19363
rect 3789 19323 3847 19329
rect 8481 19363 8539 19369
rect 8481 19329 8493 19363
rect 8527 19360 8539 19363
rect 8588 19360 8616 19456
rect 8527 19332 8616 19360
rect 8527 19329 8539 19332
rect 8481 19323 8539 19329
rect 1673 19295 1731 19301
rect 1673 19261 1685 19295
rect 1719 19292 1731 19295
rect 2314 19292 2320 19304
rect 1719 19264 2320 19292
rect 1719 19261 1731 19264
rect 1673 19255 1731 19261
rect 2314 19252 2320 19264
rect 2372 19252 2378 19304
rect 6362 19184 6368 19236
rect 6420 19184 6426 19236
rect 1670 19116 1676 19168
rect 1728 19156 1734 19168
rect 1765 19159 1823 19165
rect 1765 19156 1777 19159
rect 1728 19128 1777 19156
rect 1728 19116 1734 19128
rect 1765 19125 1777 19128
rect 1811 19125 1823 19159
rect 1765 19119 1823 19125
rect 8294 19116 8300 19168
rect 8352 19116 8358 19168
rect 1104 19066 8832 19088
rect 1104 19014 1916 19066
rect 1968 19014 1980 19066
rect 2032 19014 2044 19066
rect 2096 19014 2108 19066
rect 2160 19014 2172 19066
rect 2224 19014 3848 19066
rect 3900 19014 3912 19066
rect 3964 19014 3976 19066
rect 4028 19014 4040 19066
rect 4092 19014 4104 19066
rect 4156 19014 5780 19066
rect 5832 19014 5844 19066
rect 5896 19014 5908 19066
rect 5960 19014 5972 19066
rect 6024 19014 6036 19066
rect 6088 19014 7712 19066
rect 7764 19014 7776 19066
rect 7828 19014 7840 19066
rect 7892 19014 7904 19066
rect 7956 19014 7968 19066
rect 8020 19014 8832 19066
rect 1104 18992 8832 19014
rect 934 18708 940 18760
rect 992 18748 998 18760
rect 1397 18751 1455 18757
rect 1397 18748 1409 18751
rect 992 18720 1409 18748
rect 992 18708 998 18720
rect 1397 18717 1409 18720
rect 1443 18717 1455 18751
rect 1397 18711 1455 18717
rect 1578 18572 1584 18624
rect 1636 18572 1642 18624
rect 1104 18522 8992 18544
rect 1104 18470 2882 18522
rect 2934 18470 2946 18522
rect 2998 18470 3010 18522
rect 3062 18470 3074 18522
rect 3126 18470 3138 18522
rect 3190 18470 4814 18522
rect 4866 18470 4878 18522
rect 4930 18470 4942 18522
rect 4994 18470 5006 18522
rect 5058 18470 5070 18522
rect 5122 18470 6746 18522
rect 6798 18470 6810 18522
rect 6862 18470 6874 18522
rect 6926 18470 6938 18522
rect 6990 18470 7002 18522
rect 7054 18470 8678 18522
rect 8730 18470 8742 18522
rect 8794 18470 8806 18522
rect 8858 18470 8870 18522
rect 8922 18470 8934 18522
rect 8986 18470 8992 18522
rect 1104 18448 8992 18470
rect 1104 17978 8832 18000
rect 1104 17926 1916 17978
rect 1968 17926 1980 17978
rect 2032 17926 2044 17978
rect 2096 17926 2108 17978
rect 2160 17926 2172 17978
rect 2224 17926 3848 17978
rect 3900 17926 3912 17978
rect 3964 17926 3976 17978
rect 4028 17926 4040 17978
rect 4092 17926 4104 17978
rect 4156 17926 5780 17978
rect 5832 17926 5844 17978
rect 5896 17926 5908 17978
rect 5960 17926 5972 17978
rect 6024 17926 6036 17978
rect 6088 17926 7712 17978
rect 7764 17926 7776 17978
rect 7828 17926 7840 17978
rect 7892 17926 7904 17978
rect 7956 17926 7968 17978
rect 8020 17926 8832 17978
rect 1104 17904 8832 17926
rect 1104 17434 8992 17456
rect 1104 17382 2882 17434
rect 2934 17382 2946 17434
rect 2998 17382 3010 17434
rect 3062 17382 3074 17434
rect 3126 17382 3138 17434
rect 3190 17382 4814 17434
rect 4866 17382 4878 17434
rect 4930 17382 4942 17434
rect 4994 17382 5006 17434
rect 5058 17382 5070 17434
rect 5122 17382 6746 17434
rect 6798 17382 6810 17434
rect 6862 17382 6874 17434
rect 6926 17382 6938 17434
rect 6990 17382 7002 17434
rect 7054 17382 8678 17434
rect 8730 17382 8742 17434
rect 8794 17382 8806 17434
rect 8858 17382 8870 17434
rect 8922 17382 8934 17434
rect 8986 17382 8992 17434
rect 1104 17360 8992 17382
rect 934 17144 940 17196
rect 992 17184 998 17196
rect 1397 17187 1455 17193
rect 1397 17184 1409 17187
rect 992 17156 1409 17184
rect 992 17144 998 17156
rect 1397 17153 1409 17156
rect 1443 17153 1455 17187
rect 1397 17147 1455 17153
rect 1394 16940 1400 16992
rect 1452 16980 1458 16992
rect 1581 16983 1639 16989
rect 1581 16980 1593 16983
rect 1452 16952 1593 16980
rect 1452 16940 1458 16952
rect 1581 16949 1593 16952
rect 1627 16949 1639 16983
rect 1581 16943 1639 16949
rect 1104 16890 8832 16912
rect 1104 16838 1916 16890
rect 1968 16838 1980 16890
rect 2032 16838 2044 16890
rect 2096 16838 2108 16890
rect 2160 16838 2172 16890
rect 2224 16838 3848 16890
rect 3900 16838 3912 16890
rect 3964 16838 3976 16890
rect 4028 16838 4040 16890
rect 4092 16838 4104 16890
rect 4156 16838 5780 16890
rect 5832 16838 5844 16890
rect 5896 16838 5908 16890
rect 5960 16838 5972 16890
rect 6024 16838 6036 16890
rect 6088 16838 7712 16890
rect 7764 16838 7776 16890
rect 7828 16838 7840 16890
rect 7892 16838 7904 16890
rect 7956 16838 7968 16890
rect 8020 16838 8832 16890
rect 1104 16816 8832 16838
rect 1486 16600 1492 16652
rect 1544 16640 1550 16652
rect 1670 16640 1676 16652
rect 1544 16612 1676 16640
rect 1544 16600 1550 16612
rect 1670 16600 1676 16612
rect 1728 16600 1734 16652
rect 1104 16346 8992 16368
rect 1104 16294 2882 16346
rect 2934 16294 2946 16346
rect 2998 16294 3010 16346
rect 3062 16294 3074 16346
rect 3126 16294 3138 16346
rect 3190 16294 4814 16346
rect 4866 16294 4878 16346
rect 4930 16294 4942 16346
rect 4994 16294 5006 16346
rect 5058 16294 5070 16346
rect 5122 16294 6746 16346
rect 6798 16294 6810 16346
rect 6862 16294 6874 16346
rect 6926 16294 6938 16346
rect 6990 16294 7002 16346
rect 7054 16294 8678 16346
rect 8730 16294 8742 16346
rect 8794 16294 8806 16346
rect 8858 16294 8870 16346
rect 8922 16294 8934 16346
rect 8986 16294 8992 16346
rect 1104 16272 8992 16294
rect 1397 16099 1455 16105
rect 1397 16065 1409 16099
rect 1443 16096 1455 16099
rect 1486 16096 1492 16108
rect 1443 16068 1492 16096
rect 1443 16065 1455 16068
rect 1397 16059 1455 16065
rect 1486 16056 1492 16068
rect 1544 16056 1550 16108
rect 1578 16056 1584 16108
rect 1636 16056 1642 16108
rect 6362 16056 6368 16108
rect 6420 16056 6426 16108
rect 2317 16031 2375 16037
rect 2317 16028 2329 16031
rect 1504 16000 2329 16028
rect 1504 15972 1532 16000
rect 2317 15997 2329 16000
rect 2363 15997 2375 16031
rect 2317 15991 2375 15997
rect 2406 15988 2412 16040
rect 2464 16037 2470 16040
rect 2464 16031 2492 16037
rect 2480 15997 2492 16031
rect 2464 15991 2492 15997
rect 2464 15988 2470 15991
rect 2590 15988 2596 16040
rect 2648 16028 2654 16040
rect 6380 16028 6408 16056
rect 2648 16000 6408 16028
rect 2648 15988 2654 16000
rect 1486 15920 1492 15972
rect 1544 15920 1550 15972
rect 2041 15963 2099 15969
rect 2041 15929 2053 15963
rect 2087 15929 2099 15963
rect 2041 15923 2099 15929
rect 2056 15892 2084 15923
rect 2498 15892 2504 15904
rect 2056 15864 2504 15892
rect 2498 15852 2504 15864
rect 2556 15852 2562 15904
rect 2774 15852 2780 15904
rect 2832 15892 2838 15904
rect 3237 15895 3295 15901
rect 3237 15892 3249 15895
rect 2832 15864 3249 15892
rect 2832 15852 2838 15864
rect 3237 15861 3249 15864
rect 3283 15861 3295 15895
rect 3237 15855 3295 15861
rect 1104 15802 8832 15824
rect 1104 15750 1916 15802
rect 1968 15750 1980 15802
rect 2032 15750 2044 15802
rect 2096 15750 2108 15802
rect 2160 15750 2172 15802
rect 2224 15750 3848 15802
rect 3900 15750 3912 15802
rect 3964 15750 3976 15802
rect 4028 15750 4040 15802
rect 4092 15750 4104 15802
rect 4156 15750 5780 15802
rect 5832 15750 5844 15802
rect 5896 15750 5908 15802
rect 5960 15750 5972 15802
rect 6024 15750 6036 15802
rect 6088 15750 7712 15802
rect 7764 15750 7776 15802
rect 7828 15750 7840 15802
rect 7892 15750 7904 15802
rect 7956 15750 7968 15802
rect 8020 15750 8832 15802
rect 1104 15728 8832 15750
rect 1581 15691 1639 15697
rect 1581 15657 1593 15691
rect 1627 15688 1639 15691
rect 2406 15688 2412 15700
rect 1627 15660 2412 15688
rect 1627 15657 1639 15660
rect 1581 15651 1639 15657
rect 2406 15648 2412 15660
rect 2464 15648 2470 15700
rect 934 15444 940 15496
rect 992 15484 998 15496
rect 1397 15487 1455 15493
rect 1397 15484 1409 15487
rect 992 15456 1409 15484
rect 992 15444 998 15456
rect 1397 15453 1409 15456
rect 1443 15453 1455 15487
rect 1397 15447 1455 15453
rect 1104 15258 8992 15280
rect 1104 15206 2882 15258
rect 2934 15206 2946 15258
rect 2998 15206 3010 15258
rect 3062 15206 3074 15258
rect 3126 15206 3138 15258
rect 3190 15206 4814 15258
rect 4866 15206 4878 15258
rect 4930 15206 4942 15258
rect 4994 15206 5006 15258
rect 5058 15206 5070 15258
rect 5122 15206 6746 15258
rect 6798 15206 6810 15258
rect 6862 15206 6874 15258
rect 6926 15206 6938 15258
rect 6990 15206 7002 15258
rect 7054 15206 8678 15258
rect 8730 15206 8742 15258
rect 8794 15206 8806 15258
rect 8858 15206 8870 15258
rect 8922 15206 8934 15258
rect 8986 15206 8992 15258
rect 1104 15184 8992 15206
rect 1394 14968 1400 15020
rect 1452 14968 1458 15020
rect 1578 14968 1584 15020
rect 1636 14968 1642 15020
rect 2590 14968 2596 15020
rect 2648 14968 2654 15020
rect 1762 14900 1768 14952
rect 1820 14940 1826 14952
rect 2317 14943 2375 14949
rect 2317 14940 2329 14943
rect 1820 14912 2329 14940
rect 1820 14900 1826 14912
rect 2317 14909 2329 14912
rect 2363 14909 2375 14943
rect 2317 14903 2375 14909
rect 2406 14900 2412 14952
rect 2464 14949 2470 14952
rect 2464 14943 2492 14949
rect 2480 14909 2492 14943
rect 2464 14903 2492 14909
rect 2464 14900 2470 14903
rect 2041 14875 2099 14881
rect 2041 14841 2053 14875
rect 2087 14841 2099 14875
rect 2041 14835 2099 14841
rect 1670 14764 1676 14816
rect 1728 14804 1734 14816
rect 2056 14804 2084 14835
rect 2498 14804 2504 14816
rect 1728 14776 2504 14804
rect 1728 14764 1734 14776
rect 2498 14764 2504 14776
rect 2556 14764 2562 14816
rect 3234 14764 3240 14816
rect 3292 14764 3298 14816
rect 1104 14714 8832 14736
rect 1104 14662 1916 14714
rect 1968 14662 1980 14714
rect 2032 14662 2044 14714
rect 2096 14662 2108 14714
rect 2160 14662 2172 14714
rect 2224 14662 3848 14714
rect 3900 14662 3912 14714
rect 3964 14662 3976 14714
rect 4028 14662 4040 14714
rect 4092 14662 4104 14714
rect 4156 14662 5780 14714
rect 5832 14662 5844 14714
rect 5896 14662 5908 14714
rect 5960 14662 5972 14714
rect 6024 14662 6036 14714
rect 6088 14662 7712 14714
rect 7764 14662 7776 14714
rect 7828 14662 7840 14714
rect 7892 14662 7904 14714
rect 7956 14662 7968 14714
rect 8020 14662 8832 14714
rect 1104 14640 8832 14662
rect 1581 14603 1639 14609
rect 1581 14569 1593 14603
rect 1627 14600 1639 14603
rect 2406 14600 2412 14612
rect 1627 14572 2412 14600
rect 1627 14569 1639 14572
rect 1581 14563 1639 14569
rect 2406 14560 2412 14572
rect 2464 14560 2470 14612
rect 3234 14600 3240 14612
rect 2792 14572 3240 14600
rect 1578 14424 1584 14476
rect 1636 14464 1642 14476
rect 2314 14464 2320 14476
rect 1636 14436 2320 14464
rect 1636 14424 1642 14436
rect 2314 14424 2320 14436
rect 2372 14464 2378 14476
rect 2792 14473 2820 14572
rect 3234 14560 3240 14572
rect 3292 14560 3298 14612
rect 2777 14467 2835 14473
rect 2372 14436 2728 14464
rect 2372 14424 2378 14436
rect 934 14356 940 14408
rect 992 14396 998 14408
rect 1397 14399 1455 14405
rect 1397 14396 1409 14399
rect 992 14368 1409 14396
rect 992 14356 998 14368
rect 1397 14365 1409 14368
rect 1443 14365 1455 14399
rect 2700 14396 2728 14436
rect 2777 14433 2789 14467
rect 2823 14433 2835 14467
rect 2777 14427 2835 14433
rect 2869 14467 2927 14473
rect 2869 14433 2881 14467
rect 2915 14433 2927 14467
rect 2869 14427 2927 14433
rect 2884 14396 2912 14427
rect 2700 14368 2912 14396
rect 1397 14359 1455 14365
rect 2685 14331 2743 14337
rect 2685 14297 2697 14331
rect 2731 14328 2743 14331
rect 2774 14328 2780 14340
rect 2731 14300 2780 14328
rect 2731 14297 2743 14300
rect 2685 14291 2743 14297
rect 2774 14288 2780 14300
rect 2832 14288 2838 14340
rect 2314 14220 2320 14272
rect 2372 14220 2378 14272
rect 1104 14170 8992 14192
rect 1104 14118 2882 14170
rect 2934 14118 2946 14170
rect 2998 14118 3010 14170
rect 3062 14118 3074 14170
rect 3126 14118 3138 14170
rect 3190 14118 4814 14170
rect 4866 14118 4878 14170
rect 4930 14118 4942 14170
rect 4994 14118 5006 14170
rect 5058 14118 5070 14170
rect 5122 14118 6746 14170
rect 6798 14118 6810 14170
rect 6862 14118 6874 14170
rect 6926 14118 6938 14170
rect 6990 14118 7002 14170
rect 7054 14118 8678 14170
rect 8730 14118 8742 14170
rect 8794 14118 8806 14170
rect 8858 14118 8870 14170
rect 8922 14118 8934 14170
rect 8986 14118 8992 14170
rect 1104 14096 8992 14118
rect 1104 13626 8832 13648
rect 1104 13574 1916 13626
rect 1968 13574 1980 13626
rect 2032 13574 2044 13626
rect 2096 13574 2108 13626
rect 2160 13574 2172 13626
rect 2224 13574 3848 13626
rect 3900 13574 3912 13626
rect 3964 13574 3976 13626
rect 4028 13574 4040 13626
rect 4092 13574 4104 13626
rect 4156 13574 5780 13626
rect 5832 13574 5844 13626
rect 5896 13574 5908 13626
rect 5960 13574 5972 13626
rect 6024 13574 6036 13626
rect 6088 13574 7712 13626
rect 7764 13574 7776 13626
rect 7828 13574 7840 13626
rect 7892 13574 7904 13626
rect 7956 13574 7968 13626
rect 8020 13574 8832 13626
rect 1104 13552 8832 13574
rect 1486 13472 1492 13524
rect 1544 13512 1550 13524
rect 1581 13515 1639 13521
rect 1581 13512 1593 13515
rect 1544 13484 1593 13512
rect 1544 13472 1550 13484
rect 1581 13481 1593 13484
rect 1627 13481 1639 13515
rect 1581 13475 1639 13481
rect 934 13268 940 13320
rect 992 13308 998 13320
rect 1397 13311 1455 13317
rect 1397 13308 1409 13311
rect 992 13280 1409 13308
rect 992 13268 998 13280
rect 1397 13277 1409 13280
rect 1443 13277 1455 13311
rect 1397 13271 1455 13277
rect 1104 13082 8992 13104
rect 1104 13030 2882 13082
rect 2934 13030 2946 13082
rect 2998 13030 3010 13082
rect 3062 13030 3074 13082
rect 3126 13030 3138 13082
rect 3190 13030 4814 13082
rect 4866 13030 4878 13082
rect 4930 13030 4942 13082
rect 4994 13030 5006 13082
rect 5058 13030 5070 13082
rect 5122 13030 6746 13082
rect 6798 13030 6810 13082
rect 6862 13030 6874 13082
rect 6926 13030 6938 13082
rect 6990 13030 7002 13082
rect 7054 13030 8678 13082
rect 8730 13030 8742 13082
rect 8794 13030 8806 13082
rect 8858 13030 8870 13082
rect 8922 13030 8934 13082
rect 8986 13030 8992 13082
rect 1104 13008 8992 13030
rect 1104 12538 8832 12560
rect 1104 12486 1916 12538
rect 1968 12486 1980 12538
rect 2032 12486 2044 12538
rect 2096 12486 2108 12538
rect 2160 12486 2172 12538
rect 2224 12486 3848 12538
rect 3900 12486 3912 12538
rect 3964 12486 3976 12538
rect 4028 12486 4040 12538
rect 4092 12486 4104 12538
rect 4156 12486 5780 12538
rect 5832 12486 5844 12538
rect 5896 12486 5908 12538
rect 5960 12486 5972 12538
rect 6024 12486 6036 12538
rect 6088 12486 7712 12538
rect 7764 12486 7776 12538
rect 7828 12486 7840 12538
rect 7892 12486 7904 12538
rect 7956 12486 7968 12538
rect 8020 12486 8832 12538
rect 1104 12464 8832 12486
rect 2314 12180 2320 12232
rect 2372 12180 2378 12232
rect 2501 12223 2559 12229
rect 2501 12189 2513 12223
rect 2547 12220 2559 12223
rect 2774 12220 2780 12232
rect 2547 12192 2780 12220
rect 2547 12189 2559 12192
rect 2501 12183 2559 12189
rect 2774 12180 2780 12192
rect 2832 12220 2838 12232
rect 8294 12220 8300 12232
rect 2832 12192 8300 12220
rect 2832 12180 2838 12192
rect 8294 12180 8300 12192
rect 8352 12180 8358 12232
rect 2406 12044 2412 12096
rect 2464 12044 2470 12096
rect 1104 11994 8992 12016
rect 1104 11942 2882 11994
rect 2934 11942 2946 11994
rect 2998 11942 3010 11994
rect 3062 11942 3074 11994
rect 3126 11942 3138 11994
rect 3190 11942 4814 11994
rect 4866 11942 4878 11994
rect 4930 11942 4942 11994
rect 4994 11942 5006 11994
rect 5058 11942 5070 11994
rect 5122 11942 6746 11994
rect 6798 11942 6810 11994
rect 6862 11942 6874 11994
rect 6926 11942 6938 11994
rect 6990 11942 7002 11994
rect 7054 11942 8678 11994
rect 8730 11942 8742 11994
rect 8794 11942 8806 11994
rect 8858 11942 8870 11994
rect 8922 11942 8934 11994
rect 8986 11942 8992 11994
rect 1104 11920 8992 11942
rect 1581 11883 1639 11889
rect 1581 11849 1593 11883
rect 1627 11880 1639 11883
rect 1762 11880 1768 11892
rect 1627 11852 1768 11880
rect 1627 11849 1639 11852
rect 1581 11843 1639 11849
rect 1762 11840 1768 11852
rect 1820 11840 1826 11892
rect 2406 11840 2412 11892
rect 2464 11840 2470 11892
rect 2774 11840 2780 11892
rect 2832 11840 2838 11892
rect 934 11704 940 11756
rect 992 11744 998 11756
rect 2424 11753 2452 11840
rect 2792 11753 2820 11840
rect 1397 11747 1455 11753
rect 1397 11744 1409 11747
rect 992 11716 1409 11744
rect 992 11704 998 11716
rect 1397 11713 1409 11716
rect 1443 11713 1455 11747
rect 1397 11707 1455 11713
rect 2409 11747 2467 11753
rect 2409 11713 2421 11747
rect 2455 11713 2467 11747
rect 2409 11707 2467 11713
rect 2777 11747 2835 11753
rect 2777 11713 2789 11747
rect 2823 11713 2835 11747
rect 2777 11707 2835 11713
rect 2958 11636 2964 11688
rect 3016 11636 3022 11688
rect 2498 11568 2504 11620
rect 2556 11568 2562 11620
rect 1104 11450 8832 11472
rect 1104 11398 1916 11450
rect 1968 11398 1980 11450
rect 2032 11398 2044 11450
rect 2096 11398 2108 11450
rect 2160 11398 2172 11450
rect 2224 11398 3848 11450
rect 3900 11398 3912 11450
rect 3964 11398 3976 11450
rect 4028 11398 4040 11450
rect 4092 11398 4104 11450
rect 4156 11398 5780 11450
rect 5832 11398 5844 11450
rect 5896 11398 5908 11450
rect 5960 11398 5972 11450
rect 6024 11398 6036 11450
rect 6088 11398 7712 11450
rect 7764 11398 7776 11450
rect 7828 11398 7840 11450
rect 7892 11398 7904 11450
rect 7956 11398 7968 11450
rect 8020 11398 8832 11450
rect 1104 11376 8832 11398
rect 2498 11296 2504 11348
rect 2556 11336 2562 11348
rect 2556 11308 6914 11336
rect 2556 11296 2562 11308
rect 6886 11132 6914 11308
rect 7101 11135 7159 11141
rect 7101 11132 7113 11135
rect 6886 11104 7113 11132
rect 7101 11101 7113 11104
rect 7147 11101 7159 11135
rect 7101 11095 7159 11101
rect 8202 11024 8208 11076
rect 8260 11024 8266 11076
rect 1104 10906 8992 10928
rect 1104 10854 2882 10906
rect 2934 10854 2946 10906
rect 2998 10854 3010 10906
rect 3062 10854 3074 10906
rect 3126 10854 3138 10906
rect 3190 10854 4814 10906
rect 4866 10854 4878 10906
rect 4930 10854 4942 10906
rect 4994 10854 5006 10906
rect 5058 10854 5070 10906
rect 5122 10854 6746 10906
rect 6798 10854 6810 10906
rect 6862 10854 6874 10906
rect 6926 10854 6938 10906
rect 6990 10854 7002 10906
rect 7054 10854 8678 10906
rect 8730 10854 8742 10906
rect 8794 10854 8806 10906
rect 8858 10854 8870 10906
rect 8922 10854 8934 10906
rect 8986 10854 8992 10906
rect 1104 10832 8992 10854
rect 934 10616 940 10668
rect 992 10656 998 10668
rect 1397 10659 1455 10665
rect 1397 10656 1409 10659
rect 992 10628 1409 10656
rect 992 10616 998 10628
rect 1397 10625 1409 10628
rect 1443 10625 1455 10659
rect 1397 10619 1455 10625
rect 1486 10412 1492 10464
rect 1544 10452 1550 10464
rect 1581 10455 1639 10461
rect 1581 10452 1593 10455
rect 1544 10424 1593 10452
rect 1544 10412 1550 10424
rect 1581 10421 1593 10424
rect 1627 10421 1639 10455
rect 1581 10415 1639 10421
rect 1104 10362 8832 10384
rect 1104 10310 1916 10362
rect 1968 10310 1980 10362
rect 2032 10310 2044 10362
rect 2096 10310 2108 10362
rect 2160 10310 2172 10362
rect 2224 10310 3848 10362
rect 3900 10310 3912 10362
rect 3964 10310 3976 10362
rect 4028 10310 4040 10362
rect 4092 10310 4104 10362
rect 4156 10310 5780 10362
rect 5832 10310 5844 10362
rect 5896 10310 5908 10362
rect 5960 10310 5972 10362
rect 6024 10310 6036 10362
rect 6088 10310 7712 10362
rect 7764 10310 7776 10362
rect 7828 10310 7840 10362
rect 7892 10310 7904 10362
rect 7956 10310 7968 10362
rect 8020 10310 8832 10362
rect 1104 10288 8832 10310
rect 1104 9818 8992 9840
rect 1104 9766 2882 9818
rect 2934 9766 2946 9818
rect 2998 9766 3010 9818
rect 3062 9766 3074 9818
rect 3126 9766 3138 9818
rect 3190 9766 4814 9818
rect 4866 9766 4878 9818
rect 4930 9766 4942 9818
rect 4994 9766 5006 9818
rect 5058 9766 5070 9818
rect 5122 9766 6746 9818
rect 6798 9766 6810 9818
rect 6862 9766 6874 9818
rect 6926 9766 6938 9818
rect 6990 9766 7002 9818
rect 7054 9766 8678 9818
rect 8730 9766 8742 9818
rect 8794 9766 8806 9818
rect 8858 9766 8870 9818
rect 8922 9766 8934 9818
rect 8986 9766 8992 9818
rect 1104 9744 8992 9766
rect 1578 9528 1584 9580
rect 1636 9528 1642 9580
rect 1670 9528 1676 9580
rect 1728 9528 1734 9580
rect 1486 9460 1492 9512
rect 1544 9460 1550 9512
rect 1596 9500 1624 9528
rect 2406 9500 2412 9512
rect 1596 9472 2412 9500
rect 2406 9460 2412 9472
rect 2464 9460 2470 9512
rect 1857 9367 1915 9373
rect 1857 9333 1869 9367
rect 1903 9364 1915 9367
rect 2590 9364 2596 9376
rect 1903 9336 2596 9364
rect 1903 9333 1915 9336
rect 1857 9327 1915 9333
rect 2590 9324 2596 9336
rect 2648 9324 2654 9376
rect 1104 9274 8832 9296
rect 1104 9222 1916 9274
rect 1968 9222 1980 9274
rect 2032 9222 2044 9274
rect 2096 9222 2108 9274
rect 2160 9222 2172 9274
rect 2224 9222 3848 9274
rect 3900 9222 3912 9274
rect 3964 9222 3976 9274
rect 4028 9222 4040 9274
rect 4092 9222 4104 9274
rect 4156 9222 5780 9274
rect 5832 9222 5844 9274
rect 5896 9222 5908 9274
rect 5960 9222 5972 9274
rect 6024 9222 6036 9274
rect 6088 9222 7712 9274
rect 7764 9222 7776 9274
rect 7828 9222 7840 9274
rect 7892 9222 7904 9274
rect 7956 9222 7968 9274
rect 8020 9222 8832 9274
rect 1104 9200 8832 9222
rect 934 8916 940 8968
rect 992 8956 998 8968
rect 1397 8959 1455 8965
rect 1397 8956 1409 8959
rect 992 8928 1409 8956
rect 992 8916 998 8928
rect 1397 8925 1409 8928
rect 1443 8925 1455 8959
rect 1397 8919 1455 8925
rect 1578 8780 1584 8832
rect 1636 8780 1642 8832
rect 1104 8730 8992 8752
rect 1104 8678 2882 8730
rect 2934 8678 2946 8730
rect 2998 8678 3010 8730
rect 3062 8678 3074 8730
rect 3126 8678 3138 8730
rect 3190 8678 4814 8730
rect 4866 8678 4878 8730
rect 4930 8678 4942 8730
rect 4994 8678 5006 8730
rect 5058 8678 5070 8730
rect 5122 8678 6746 8730
rect 6798 8678 6810 8730
rect 6862 8678 6874 8730
rect 6926 8678 6938 8730
rect 6990 8678 7002 8730
rect 7054 8678 8678 8730
rect 8730 8678 8742 8730
rect 8794 8678 8806 8730
rect 8858 8678 8870 8730
rect 8922 8678 8934 8730
rect 8986 8678 8992 8730
rect 1104 8656 8992 8678
rect 1578 8576 1584 8628
rect 1636 8616 1642 8628
rect 1765 8619 1823 8625
rect 1765 8616 1777 8619
rect 1636 8588 1777 8616
rect 1636 8576 1642 8588
rect 1765 8585 1777 8588
rect 1811 8585 1823 8619
rect 1765 8579 1823 8585
rect 2133 8619 2191 8625
rect 2133 8585 2145 8619
rect 2179 8616 2191 8619
rect 2317 8619 2375 8625
rect 2317 8616 2329 8619
rect 2179 8588 2329 8616
rect 2179 8585 2191 8588
rect 2133 8579 2191 8585
rect 2317 8585 2329 8588
rect 2363 8585 2375 8619
rect 2317 8579 2375 8585
rect 2406 8576 2412 8628
rect 2464 8576 2470 8628
rect 2590 8576 2596 8628
rect 2648 8576 2654 8628
rect 2682 8576 2688 8628
rect 2740 8576 2746 8628
rect 1670 8548 1676 8560
rect 1596 8520 1676 8548
rect 1596 8421 1624 8520
rect 1670 8508 1676 8520
rect 1728 8508 1734 8560
rect 2424 8489 2452 8576
rect 2409 8483 2467 8489
rect 2409 8449 2421 8483
rect 2455 8449 2467 8483
rect 2409 8443 2467 8449
rect 2498 8440 2504 8492
rect 2556 8440 2562 8492
rect 2608 8489 2636 8576
rect 2593 8483 2651 8489
rect 2593 8449 2605 8483
rect 2639 8449 2651 8483
rect 2593 8443 2651 8449
rect 1581 8415 1639 8421
rect 1581 8381 1593 8415
rect 1627 8381 1639 8415
rect 1581 8375 1639 8381
rect 1670 8372 1676 8424
rect 1728 8372 1734 8424
rect 2516 8412 2544 8440
rect 2685 8415 2743 8421
rect 2685 8412 2697 8415
rect 2516 8384 2697 8412
rect 2685 8381 2697 8384
rect 2731 8381 2743 8415
rect 2685 8375 2743 8381
rect 2498 8236 2504 8288
rect 2556 8236 2562 8288
rect 1104 8186 8832 8208
rect 1104 8134 1916 8186
rect 1968 8134 1980 8186
rect 2032 8134 2044 8186
rect 2096 8134 2108 8186
rect 2160 8134 2172 8186
rect 2224 8134 3848 8186
rect 3900 8134 3912 8186
rect 3964 8134 3976 8186
rect 4028 8134 4040 8186
rect 4092 8134 4104 8186
rect 4156 8134 5780 8186
rect 5832 8134 5844 8186
rect 5896 8134 5908 8186
rect 5960 8134 5972 8186
rect 6024 8134 6036 8186
rect 6088 8134 7712 8186
rect 7764 8134 7776 8186
rect 7828 8134 7840 8186
rect 7892 8134 7904 8186
rect 7956 8134 7968 8186
rect 8020 8134 8832 8186
rect 1104 8112 8832 8134
rect 1762 8032 1768 8084
rect 1820 8032 1826 8084
rect 1949 8075 2007 8081
rect 1949 8041 1961 8075
rect 1995 8072 2007 8075
rect 2498 8072 2504 8084
rect 1995 8044 2504 8072
rect 1995 8041 2007 8044
rect 1949 8035 2007 8041
rect 2498 8032 2504 8044
rect 2556 8032 2562 8084
rect 1397 8007 1455 8013
rect 1397 7973 1409 8007
rect 1443 8004 1455 8007
rect 1486 8004 1492 8016
rect 1443 7976 1492 8004
rect 1443 7973 1455 7976
rect 1397 7967 1455 7973
rect 1486 7964 1492 7976
rect 1544 7964 1550 8016
rect 1780 8004 1808 8032
rect 2406 8004 2412 8016
rect 1780 7976 2412 8004
rect 2406 7964 2412 7976
rect 2464 7964 2470 8016
rect 1762 7692 1768 7744
rect 1820 7692 1826 7744
rect 1104 7642 8992 7664
rect 1104 7590 2882 7642
rect 2934 7590 2946 7642
rect 2998 7590 3010 7642
rect 3062 7590 3074 7642
rect 3126 7590 3138 7642
rect 3190 7590 4814 7642
rect 4866 7590 4878 7642
rect 4930 7590 4942 7642
rect 4994 7590 5006 7642
rect 5058 7590 5070 7642
rect 5122 7590 6746 7642
rect 6798 7590 6810 7642
rect 6862 7590 6874 7642
rect 6926 7590 6938 7642
rect 6990 7590 7002 7642
rect 7054 7590 8678 7642
rect 8730 7590 8742 7642
rect 8794 7590 8806 7642
rect 8858 7590 8870 7642
rect 8922 7590 8934 7642
rect 8986 7590 8992 7642
rect 1104 7568 8992 7590
rect 1581 7531 1639 7537
rect 1581 7497 1593 7531
rect 1627 7528 1639 7531
rect 1762 7528 1768 7540
rect 1627 7500 1768 7528
rect 1627 7497 1639 7500
rect 1581 7491 1639 7497
rect 1762 7488 1768 7500
rect 1820 7488 1826 7540
rect 934 7352 940 7404
rect 992 7392 998 7404
rect 1397 7395 1455 7401
rect 1397 7392 1409 7395
rect 992 7364 1409 7392
rect 992 7352 998 7364
rect 1397 7361 1409 7364
rect 1443 7361 1455 7395
rect 1397 7355 1455 7361
rect 1104 7098 8832 7120
rect 1104 7046 1916 7098
rect 1968 7046 1980 7098
rect 2032 7046 2044 7098
rect 2096 7046 2108 7098
rect 2160 7046 2172 7098
rect 2224 7046 3848 7098
rect 3900 7046 3912 7098
rect 3964 7046 3976 7098
rect 4028 7046 4040 7098
rect 4092 7046 4104 7098
rect 4156 7046 5780 7098
rect 5832 7046 5844 7098
rect 5896 7046 5908 7098
rect 5960 7046 5972 7098
rect 6024 7046 6036 7098
rect 6088 7046 7712 7098
rect 7764 7046 7776 7098
rect 7828 7046 7840 7098
rect 7892 7046 7904 7098
rect 7956 7046 7968 7098
rect 8020 7046 8832 7098
rect 1104 7024 8832 7046
rect 2041 6851 2099 6857
rect 2041 6817 2053 6851
rect 2087 6848 2099 6851
rect 2314 6848 2320 6860
rect 2087 6820 2320 6848
rect 2087 6817 2099 6820
rect 2041 6811 2099 6817
rect 2314 6808 2320 6820
rect 2372 6808 2378 6860
rect 1673 6783 1731 6789
rect 1673 6749 1685 6783
rect 1719 6780 1731 6783
rect 1946 6780 1952 6792
rect 1719 6752 1952 6780
rect 1719 6749 1731 6752
rect 1673 6743 1731 6749
rect 1946 6740 1952 6752
rect 2004 6740 2010 6792
rect 2133 6783 2191 6789
rect 2133 6749 2145 6783
rect 2179 6780 2191 6783
rect 2682 6780 2688 6792
rect 2179 6752 2688 6780
rect 2179 6749 2191 6752
rect 2133 6743 2191 6749
rect 2682 6740 2688 6752
rect 2740 6740 2746 6792
rect 1394 6672 1400 6724
rect 1452 6712 1458 6724
rect 2406 6712 2412 6724
rect 1452 6684 2412 6712
rect 1452 6672 1458 6684
rect 2406 6672 2412 6684
rect 2464 6672 2470 6724
rect 1762 6604 1768 6656
rect 1820 6604 1826 6656
rect 1854 6604 1860 6656
rect 1912 6604 1918 6656
rect 2317 6647 2375 6653
rect 2317 6613 2329 6647
rect 2363 6644 2375 6647
rect 2774 6644 2780 6656
rect 2363 6616 2780 6644
rect 2363 6613 2375 6616
rect 2317 6607 2375 6613
rect 2774 6604 2780 6616
rect 2832 6604 2838 6656
rect 1104 6554 8992 6576
rect 1104 6502 2882 6554
rect 2934 6502 2946 6554
rect 2998 6502 3010 6554
rect 3062 6502 3074 6554
rect 3126 6502 3138 6554
rect 3190 6502 4814 6554
rect 4866 6502 4878 6554
rect 4930 6502 4942 6554
rect 4994 6502 5006 6554
rect 5058 6502 5070 6554
rect 5122 6502 6746 6554
rect 6798 6502 6810 6554
rect 6862 6502 6874 6554
rect 6926 6502 6938 6554
rect 6990 6502 7002 6554
rect 7054 6502 8678 6554
rect 8730 6502 8742 6554
rect 8794 6502 8806 6554
rect 8858 6502 8870 6554
rect 8922 6502 8934 6554
rect 8986 6502 8992 6554
rect 1104 6480 8992 6502
rect 1762 6400 1768 6452
rect 1820 6440 1826 6452
rect 2225 6443 2283 6449
rect 2225 6440 2237 6443
rect 1820 6412 2237 6440
rect 1820 6400 1826 6412
rect 2225 6409 2237 6412
rect 2271 6409 2283 6443
rect 2225 6403 2283 6409
rect 1504 6344 1900 6372
rect 1504 6316 1532 6344
rect 1486 6264 1492 6316
rect 1544 6264 1550 6316
rect 1578 6264 1584 6316
rect 1636 6264 1642 6316
rect 1872 6245 1900 6344
rect 1946 6332 1952 6384
rect 2004 6372 2010 6384
rect 2004 6344 2176 6372
rect 2004 6332 2010 6344
rect 1857 6239 1915 6245
rect 1857 6205 1869 6239
rect 1903 6205 1915 6239
rect 1857 6199 1915 6205
rect 1394 6060 1400 6112
rect 1452 6100 1458 6112
rect 1673 6103 1731 6109
rect 1673 6100 1685 6103
rect 1452 6072 1685 6100
rect 1452 6060 1458 6072
rect 1673 6069 1685 6072
rect 1719 6069 1731 6103
rect 1872 6100 1900 6199
rect 2148 6177 2176 6344
rect 2406 6264 2412 6316
rect 2464 6264 2470 6316
rect 2498 6264 2504 6316
rect 2556 6264 2562 6316
rect 2593 6307 2651 6313
rect 2593 6273 2605 6307
rect 2639 6273 2651 6307
rect 2593 6267 2651 6273
rect 2608 6236 2636 6267
rect 2516 6208 2636 6236
rect 2133 6171 2191 6177
rect 2133 6137 2145 6171
rect 2179 6137 2191 6171
rect 2133 6131 2191 6137
rect 2516 6100 2544 6208
rect 1872 6072 2544 6100
rect 1673 6063 1731 6069
rect 1104 6010 8832 6032
rect 1104 5958 1916 6010
rect 1968 5958 1980 6010
rect 2032 5958 2044 6010
rect 2096 5958 2108 6010
rect 2160 5958 2172 6010
rect 2224 5958 3848 6010
rect 3900 5958 3912 6010
rect 3964 5958 3976 6010
rect 4028 5958 4040 6010
rect 4092 5958 4104 6010
rect 4156 5958 5780 6010
rect 5832 5958 5844 6010
rect 5896 5958 5908 6010
rect 5960 5958 5972 6010
rect 6024 5958 6036 6010
rect 6088 5958 7712 6010
rect 7764 5958 7776 6010
rect 7828 5958 7840 6010
rect 7892 5958 7904 6010
rect 7956 5958 7968 6010
rect 8020 5958 8832 6010
rect 1104 5936 8832 5958
rect 1581 5899 1639 5905
rect 1581 5865 1593 5899
rect 1627 5896 1639 5899
rect 1670 5896 1676 5908
rect 1627 5868 1676 5896
rect 1627 5865 1639 5868
rect 1581 5859 1639 5865
rect 1670 5856 1676 5868
rect 1728 5856 1734 5908
rect 1762 5856 1768 5908
rect 1820 5896 1826 5908
rect 1857 5899 1915 5905
rect 1857 5896 1869 5899
rect 1820 5868 1869 5896
rect 1820 5856 1826 5868
rect 1857 5865 1869 5868
rect 1903 5865 1915 5899
rect 1857 5859 1915 5865
rect 934 5652 940 5704
rect 992 5692 998 5704
rect 1397 5695 1455 5701
rect 1397 5692 1409 5695
rect 992 5664 1409 5692
rect 992 5652 998 5664
rect 1397 5661 1409 5664
rect 1443 5661 1455 5695
rect 1397 5655 1455 5661
rect 1486 5652 1492 5704
rect 1544 5692 1550 5704
rect 1765 5695 1823 5701
rect 1765 5692 1777 5695
rect 1544 5664 1777 5692
rect 1544 5652 1550 5664
rect 1765 5661 1777 5664
rect 1811 5661 1823 5695
rect 1765 5655 1823 5661
rect 1946 5652 1952 5704
rect 2004 5652 2010 5704
rect 1104 5466 8992 5488
rect 1104 5414 2882 5466
rect 2934 5414 2946 5466
rect 2998 5414 3010 5466
rect 3062 5414 3074 5466
rect 3126 5414 3138 5466
rect 3190 5414 4814 5466
rect 4866 5414 4878 5466
rect 4930 5414 4942 5466
rect 4994 5414 5006 5466
rect 5058 5414 5070 5466
rect 5122 5414 6746 5466
rect 6798 5414 6810 5466
rect 6862 5414 6874 5466
rect 6926 5414 6938 5466
rect 6990 5414 7002 5466
rect 7054 5414 8678 5466
rect 8730 5414 8742 5466
rect 8794 5414 8806 5466
rect 8858 5414 8870 5466
rect 8922 5414 8934 5466
rect 8986 5414 8992 5466
rect 1104 5392 8992 5414
rect 1946 5312 1952 5364
rect 2004 5352 2010 5364
rect 2133 5355 2191 5361
rect 2133 5352 2145 5355
rect 2004 5324 2145 5352
rect 2004 5312 2010 5324
rect 2133 5321 2145 5324
rect 2179 5321 2191 5355
rect 2133 5315 2191 5321
rect 1762 5176 1768 5228
rect 1820 5176 1826 5228
rect 1394 5108 1400 5160
rect 1452 5148 1458 5160
rect 1489 5151 1547 5157
rect 1489 5148 1501 5151
rect 1452 5120 1501 5148
rect 1452 5108 1458 5120
rect 1489 5117 1501 5120
rect 1535 5117 1547 5151
rect 1489 5111 1547 5117
rect 1670 5108 1676 5160
rect 1728 5108 1734 5160
rect 1104 4922 8832 4944
rect 1104 4870 1916 4922
rect 1968 4870 1980 4922
rect 2032 4870 2044 4922
rect 2096 4870 2108 4922
rect 2160 4870 2172 4922
rect 2224 4870 3848 4922
rect 3900 4870 3912 4922
rect 3964 4870 3976 4922
rect 4028 4870 4040 4922
rect 4092 4870 4104 4922
rect 4156 4870 5780 4922
rect 5832 4870 5844 4922
rect 5896 4870 5908 4922
rect 5960 4870 5972 4922
rect 6024 4870 6036 4922
rect 6088 4870 7712 4922
rect 7764 4870 7776 4922
rect 7828 4870 7840 4922
rect 7892 4870 7904 4922
rect 7956 4870 7968 4922
rect 8020 4870 8832 4922
rect 1104 4848 8832 4870
rect 1578 4768 1584 4820
rect 1636 4768 1642 4820
rect 934 4564 940 4616
rect 992 4604 998 4616
rect 1397 4607 1455 4613
rect 1397 4604 1409 4607
rect 992 4576 1409 4604
rect 992 4564 998 4576
rect 1397 4573 1409 4576
rect 1443 4573 1455 4607
rect 1397 4567 1455 4573
rect 1104 4378 8992 4400
rect 1104 4326 2882 4378
rect 2934 4326 2946 4378
rect 2998 4326 3010 4378
rect 3062 4326 3074 4378
rect 3126 4326 3138 4378
rect 3190 4326 4814 4378
rect 4866 4326 4878 4378
rect 4930 4326 4942 4378
rect 4994 4326 5006 4378
rect 5058 4326 5070 4378
rect 5122 4326 6746 4378
rect 6798 4326 6810 4378
rect 6862 4326 6874 4378
rect 6926 4326 6938 4378
rect 6990 4326 7002 4378
rect 7054 4326 8678 4378
rect 8730 4326 8742 4378
rect 8794 4326 8806 4378
rect 8858 4326 8870 4378
rect 8922 4326 8934 4378
rect 8986 4326 8992 4378
rect 1104 4304 8992 4326
rect 1104 3834 8832 3856
rect 1104 3782 1916 3834
rect 1968 3782 1980 3834
rect 2032 3782 2044 3834
rect 2096 3782 2108 3834
rect 2160 3782 2172 3834
rect 2224 3782 3848 3834
rect 3900 3782 3912 3834
rect 3964 3782 3976 3834
rect 4028 3782 4040 3834
rect 4092 3782 4104 3834
rect 4156 3782 5780 3834
rect 5832 3782 5844 3834
rect 5896 3782 5908 3834
rect 5960 3782 5972 3834
rect 6024 3782 6036 3834
rect 6088 3782 7712 3834
rect 7764 3782 7776 3834
rect 7828 3782 7840 3834
rect 7892 3782 7904 3834
rect 7956 3782 7968 3834
rect 8020 3782 8832 3834
rect 1104 3760 8832 3782
rect 1581 3723 1639 3729
rect 1581 3689 1593 3723
rect 1627 3720 1639 3723
rect 1762 3720 1768 3732
rect 1627 3692 1768 3720
rect 1627 3689 1639 3692
rect 1581 3683 1639 3689
rect 1762 3680 1768 3692
rect 1820 3680 1826 3732
rect 934 3476 940 3528
rect 992 3516 998 3528
rect 1397 3519 1455 3525
rect 1397 3516 1409 3519
rect 992 3488 1409 3516
rect 992 3476 998 3488
rect 1397 3485 1409 3488
rect 1443 3485 1455 3519
rect 1397 3479 1455 3485
rect 1104 3290 8992 3312
rect 1104 3238 2882 3290
rect 2934 3238 2946 3290
rect 2998 3238 3010 3290
rect 3062 3238 3074 3290
rect 3126 3238 3138 3290
rect 3190 3238 4814 3290
rect 4866 3238 4878 3290
rect 4930 3238 4942 3290
rect 4994 3238 5006 3290
rect 5058 3238 5070 3290
rect 5122 3238 6746 3290
rect 6798 3238 6810 3290
rect 6862 3238 6874 3290
rect 6926 3238 6938 3290
rect 6990 3238 7002 3290
rect 7054 3238 8678 3290
rect 8730 3238 8742 3290
rect 8794 3238 8806 3290
rect 8858 3238 8870 3290
rect 8922 3238 8934 3290
rect 8986 3238 8992 3290
rect 1104 3216 8992 3238
rect 1104 2746 8832 2768
rect 1104 2694 1916 2746
rect 1968 2694 1980 2746
rect 2032 2694 2044 2746
rect 2096 2694 2108 2746
rect 2160 2694 2172 2746
rect 2224 2694 3848 2746
rect 3900 2694 3912 2746
rect 3964 2694 3976 2746
rect 4028 2694 4040 2746
rect 4092 2694 4104 2746
rect 4156 2694 5780 2746
rect 5832 2694 5844 2746
rect 5896 2694 5908 2746
rect 5960 2694 5972 2746
rect 6024 2694 6036 2746
rect 6088 2694 7712 2746
rect 7764 2694 7776 2746
rect 7828 2694 7840 2746
rect 7892 2694 7904 2746
rect 7956 2694 7968 2746
rect 8020 2694 8832 2746
rect 1104 2672 8832 2694
rect 1670 2592 1676 2644
rect 1728 2632 1734 2644
rect 1857 2635 1915 2641
rect 1857 2632 1869 2635
rect 1728 2604 1869 2632
rect 1728 2592 1734 2604
rect 1857 2601 1869 2604
rect 1903 2601 1915 2635
rect 1857 2595 1915 2601
rect 2498 2592 2504 2644
rect 2556 2592 2562 2644
rect 1581 2567 1639 2573
rect 1581 2533 1593 2567
rect 1627 2564 1639 2567
rect 2516 2564 2544 2592
rect 1627 2536 2544 2564
rect 1627 2533 1639 2536
rect 1581 2527 1639 2533
rect 934 2388 940 2440
rect 992 2428 998 2440
rect 1397 2431 1455 2437
rect 1397 2428 1409 2431
rect 992 2400 1409 2428
rect 992 2388 998 2400
rect 1397 2397 1409 2400
rect 1443 2397 1455 2431
rect 1397 2391 1455 2397
rect 1670 2388 1676 2440
rect 1728 2388 1734 2440
rect 1104 2202 8992 2224
rect 1104 2150 2882 2202
rect 2934 2150 2946 2202
rect 2998 2150 3010 2202
rect 3062 2150 3074 2202
rect 3126 2150 3138 2202
rect 3190 2150 4814 2202
rect 4866 2150 4878 2202
rect 4930 2150 4942 2202
rect 4994 2150 5006 2202
rect 5058 2150 5070 2202
rect 5122 2150 6746 2202
rect 6798 2150 6810 2202
rect 6862 2150 6874 2202
rect 6926 2150 6938 2202
rect 6990 2150 7002 2202
rect 7054 2150 8678 2202
rect 8730 2150 8742 2202
rect 8794 2150 8806 2202
rect 8858 2150 8870 2202
rect 8922 2150 8934 2202
rect 8986 2150 8992 2202
rect 1104 2128 8992 2150
<< via1 >>
rect 2882 19558 2934 19610
rect 2946 19558 2998 19610
rect 3010 19558 3062 19610
rect 3074 19558 3126 19610
rect 3138 19558 3190 19610
rect 4814 19558 4866 19610
rect 4878 19558 4930 19610
rect 4942 19558 4994 19610
rect 5006 19558 5058 19610
rect 5070 19558 5122 19610
rect 6746 19558 6798 19610
rect 6810 19558 6862 19610
rect 6874 19558 6926 19610
rect 6938 19558 6990 19610
rect 7002 19558 7054 19610
rect 8678 19558 8730 19610
rect 8742 19558 8794 19610
rect 8806 19558 8858 19610
rect 8870 19558 8922 19610
rect 8934 19558 8986 19610
rect 1124 19456 1176 19508
rect 1400 19388 1452 19440
rect 1768 19456 1820 19508
rect 2504 19456 2556 19508
rect 8576 19456 8628 19508
rect 1032 19320 1084 19372
rect 6184 19388 6236 19440
rect 3700 19320 3752 19372
rect 2320 19252 2372 19304
rect 6368 19227 6420 19236
rect 6368 19193 6377 19227
rect 6377 19193 6411 19227
rect 6411 19193 6420 19227
rect 6368 19184 6420 19193
rect 1676 19116 1728 19168
rect 8300 19159 8352 19168
rect 8300 19125 8309 19159
rect 8309 19125 8343 19159
rect 8343 19125 8352 19159
rect 8300 19116 8352 19125
rect 1916 19014 1968 19066
rect 1980 19014 2032 19066
rect 2044 19014 2096 19066
rect 2108 19014 2160 19066
rect 2172 19014 2224 19066
rect 3848 19014 3900 19066
rect 3912 19014 3964 19066
rect 3976 19014 4028 19066
rect 4040 19014 4092 19066
rect 4104 19014 4156 19066
rect 5780 19014 5832 19066
rect 5844 19014 5896 19066
rect 5908 19014 5960 19066
rect 5972 19014 6024 19066
rect 6036 19014 6088 19066
rect 7712 19014 7764 19066
rect 7776 19014 7828 19066
rect 7840 19014 7892 19066
rect 7904 19014 7956 19066
rect 7968 19014 8020 19066
rect 940 18708 992 18760
rect 1584 18615 1636 18624
rect 1584 18581 1593 18615
rect 1593 18581 1627 18615
rect 1627 18581 1636 18615
rect 1584 18572 1636 18581
rect 2882 18470 2934 18522
rect 2946 18470 2998 18522
rect 3010 18470 3062 18522
rect 3074 18470 3126 18522
rect 3138 18470 3190 18522
rect 4814 18470 4866 18522
rect 4878 18470 4930 18522
rect 4942 18470 4994 18522
rect 5006 18470 5058 18522
rect 5070 18470 5122 18522
rect 6746 18470 6798 18522
rect 6810 18470 6862 18522
rect 6874 18470 6926 18522
rect 6938 18470 6990 18522
rect 7002 18470 7054 18522
rect 8678 18470 8730 18522
rect 8742 18470 8794 18522
rect 8806 18470 8858 18522
rect 8870 18470 8922 18522
rect 8934 18470 8986 18522
rect 1916 17926 1968 17978
rect 1980 17926 2032 17978
rect 2044 17926 2096 17978
rect 2108 17926 2160 17978
rect 2172 17926 2224 17978
rect 3848 17926 3900 17978
rect 3912 17926 3964 17978
rect 3976 17926 4028 17978
rect 4040 17926 4092 17978
rect 4104 17926 4156 17978
rect 5780 17926 5832 17978
rect 5844 17926 5896 17978
rect 5908 17926 5960 17978
rect 5972 17926 6024 17978
rect 6036 17926 6088 17978
rect 7712 17926 7764 17978
rect 7776 17926 7828 17978
rect 7840 17926 7892 17978
rect 7904 17926 7956 17978
rect 7968 17926 8020 17978
rect 2882 17382 2934 17434
rect 2946 17382 2998 17434
rect 3010 17382 3062 17434
rect 3074 17382 3126 17434
rect 3138 17382 3190 17434
rect 4814 17382 4866 17434
rect 4878 17382 4930 17434
rect 4942 17382 4994 17434
rect 5006 17382 5058 17434
rect 5070 17382 5122 17434
rect 6746 17382 6798 17434
rect 6810 17382 6862 17434
rect 6874 17382 6926 17434
rect 6938 17382 6990 17434
rect 7002 17382 7054 17434
rect 8678 17382 8730 17434
rect 8742 17382 8794 17434
rect 8806 17382 8858 17434
rect 8870 17382 8922 17434
rect 8934 17382 8986 17434
rect 940 17144 992 17196
rect 1400 16940 1452 16992
rect 1916 16838 1968 16890
rect 1980 16838 2032 16890
rect 2044 16838 2096 16890
rect 2108 16838 2160 16890
rect 2172 16838 2224 16890
rect 3848 16838 3900 16890
rect 3912 16838 3964 16890
rect 3976 16838 4028 16890
rect 4040 16838 4092 16890
rect 4104 16838 4156 16890
rect 5780 16838 5832 16890
rect 5844 16838 5896 16890
rect 5908 16838 5960 16890
rect 5972 16838 6024 16890
rect 6036 16838 6088 16890
rect 7712 16838 7764 16890
rect 7776 16838 7828 16890
rect 7840 16838 7892 16890
rect 7904 16838 7956 16890
rect 7968 16838 8020 16890
rect 1492 16600 1544 16652
rect 1676 16600 1728 16652
rect 2882 16294 2934 16346
rect 2946 16294 2998 16346
rect 3010 16294 3062 16346
rect 3074 16294 3126 16346
rect 3138 16294 3190 16346
rect 4814 16294 4866 16346
rect 4878 16294 4930 16346
rect 4942 16294 4994 16346
rect 5006 16294 5058 16346
rect 5070 16294 5122 16346
rect 6746 16294 6798 16346
rect 6810 16294 6862 16346
rect 6874 16294 6926 16346
rect 6938 16294 6990 16346
rect 7002 16294 7054 16346
rect 8678 16294 8730 16346
rect 8742 16294 8794 16346
rect 8806 16294 8858 16346
rect 8870 16294 8922 16346
rect 8934 16294 8986 16346
rect 1492 16056 1544 16108
rect 1584 16099 1636 16108
rect 1584 16065 1593 16099
rect 1593 16065 1627 16099
rect 1627 16065 1636 16099
rect 1584 16056 1636 16065
rect 6368 16056 6420 16108
rect 2412 16031 2464 16040
rect 2412 15997 2446 16031
rect 2446 15997 2464 16031
rect 2412 15988 2464 15997
rect 2596 16031 2648 16040
rect 2596 15997 2605 16031
rect 2605 15997 2639 16031
rect 2639 15997 2648 16031
rect 2596 15988 2648 15997
rect 1492 15920 1544 15972
rect 2504 15852 2556 15904
rect 2780 15852 2832 15904
rect 1916 15750 1968 15802
rect 1980 15750 2032 15802
rect 2044 15750 2096 15802
rect 2108 15750 2160 15802
rect 2172 15750 2224 15802
rect 3848 15750 3900 15802
rect 3912 15750 3964 15802
rect 3976 15750 4028 15802
rect 4040 15750 4092 15802
rect 4104 15750 4156 15802
rect 5780 15750 5832 15802
rect 5844 15750 5896 15802
rect 5908 15750 5960 15802
rect 5972 15750 6024 15802
rect 6036 15750 6088 15802
rect 7712 15750 7764 15802
rect 7776 15750 7828 15802
rect 7840 15750 7892 15802
rect 7904 15750 7956 15802
rect 7968 15750 8020 15802
rect 2412 15648 2464 15700
rect 940 15444 992 15496
rect 2882 15206 2934 15258
rect 2946 15206 2998 15258
rect 3010 15206 3062 15258
rect 3074 15206 3126 15258
rect 3138 15206 3190 15258
rect 4814 15206 4866 15258
rect 4878 15206 4930 15258
rect 4942 15206 4994 15258
rect 5006 15206 5058 15258
rect 5070 15206 5122 15258
rect 6746 15206 6798 15258
rect 6810 15206 6862 15258
rect 6874 15206 6926 15258
rect 6938 15206 6990 15258
rect 7002 15206 7054 15258
rect 8678 15206 8730 15258
rect 8742 15206 8794 15258
rect 8806 15206 8858 15258
rect 8870 15206 8922 15258
rect 8934 15206 8986 15258
rect 1400 15011 1452 15020
rect 1400 14977 1409 15011
rect 1409 14977 1443 15011
rect 1443 14977 1452 15011
rect 1400 14968 1452 14977
rect 1584 15011 1636 15020
rect 1584 14977 1593 15011
rect 1593 14977 1627 15011
rect 1627 14977 1636 15011
rect 1584 14968 1636 14977
rect 2596 15011 2648 15020
rect 2596 14977 2605 15011
rect 2605 14977 2639 15011
rect 2639 14977 2648 15011
rect 2596 14968 2648 14977
rect 1768 14900 1820 14952
rect 2412 14943 2464 14952
rect 2412 14909 2446 14943
rect 2446 14909 2464 14943
rect 2412 14900 2464 14909
rect 1676 14764 1728 14816
rect 2504 14764 2556 14816
rect 3240 14807 3292 14816
rect 3240 14773 3249 14807
rect 3249 14773 3283 14807
rect 3283 14773 3292 14807
rect 3240 14764 3292 14773
rect 1916 14662 1968 14714
rect 1980 14662 2032 14714
rect 2044 14662 2096 14714
rect 2108 14662 2160 14714
rect 2172 14662 2224 14714
rect 3848 14662 3900 14714
rect 3912 14662 3964 14714
rect 3976 14662 4028 14714
rect 4040 14662 4092 14714
rect 4104 14662 4156 14714
rect 5780 14662 5832 14714
rect 5844 14662 5896 14714
rect 5908 14662 5960 14714
rect 5972 14662 6024 14714
rect 6036 14662 6088 14714
rect 7712 14662 7764 14714
rect 7776 14662 7828 14714
rect 7840 14662 7892 14714
rect 7904 14662 7956 14714
rect 7968 14662 8020 14714
rect 2412 14560 2464 14612
rect 1584 14424 1636 14476
rect 2320 14424 2372 14476
rect 3240 14560 3292 14612
rect 940 14356 992 14408
rect 2780 14288 2832 14340
rect 2320 14263 2372 14272
rect 2320 14229 2329 14263
rect 2329 14229 2363 14263
rect 2363 14229 2372 14263
rect 2320 14220 2372 14229
rect 2882 14118 2934 14170
rect 2946 14118 2998 14170
rect 3010 14118 3062 14170
rect 3074 14118 3126 14170
rect 3138 14118 3190 14170
rect 4814 14118 4866 14170
rect 4878 14118 4930 14170
rect 4942 14118 4994 14170
rect 5006 14118 5058 14170
rect 5070 14118 5122 14170
rect 6746 14118 6798 14170
rect 6810 14118 6862 14170
rect 6874 14118 6926 14170
rect 6938 14118 6990 14170
rect 7002 14118 7054 14170
rect 8678 14118 8730 14170
rect 8742 14118 8794 14170
rect 8806 14118 8858 14170
rect 8870 14118 8922 14170
rect 8934 14118 8986 14170
rect 1916 13574 1968 13626
rect 1980 13574 2032 13626
rect 2044 13574 2096 13626
rect 2108 13574 2160 13626
rect 2172 13574 2224 13626
rect 3848 13574 3900 13626
rect 3912 13574 3964 13626
rect 3976 13574 4028 13626
rect 4040 13574 4092 13626
rect 4104 13574 4156 13626
rect 5780 13574 5832 13626
rect 5844 13574 5896 13626
rect 5908 13574 5960 13626
rect 5972 13574 6024 13626
rect 6036 13574 6088 13626
rect 7712 13574 7764 13626
rect 7776 13574 7828 13626
rect 7840 13574 7892 13626
rect 7904 13574 7956 13626
rect 7968 13574 8020 13626
rect 1492 13472 1544 13524
rect 940 13268 992 13320
rect 2882 13030 2934 13082
rect 2946 13030 2998 13082
rect 3010 13030 3062 13082
rect 3074 13030 3126 13082
rect 3138 13030 3190 13082
rect 4814 13030 4866 13082
rect 4878 13030 4930 13082
rect 4942 13030 4994 13082
rect 5006 13030 5058 13082
rect 5070 13030 5122 13082
rect 6746 13030 6798 13082
rect 6810 13030 6862 13082
rect 6874 13030 6926 13082
rect 6938 13030 6990 13082
rect 7002 13030 7054 13082
rect 8678 13030 8730 13082
rect 8742 13030 8794 13082
rect 8806 13030 8858 13082
rect 8870 13030 8922 13082
rect 8934 13030 8986 13082
rect 1916 12486 1968 12538
rect 1980 12486 2032 12538
rect 2044 12486 2096 12538
rect 2108 12486 2160 12538
rect 2172 12486 2224 12538
rect 3848 12486 3900 12538
rect 3912 12486 3964 12538
rect 3976 12486 4028 12538
rect 4040 12486 4092 12538
rect 4104 12486 4156 12538
rect 5780 12486 5832 12538
rect 5844 12486 5896 12538
rect 5908 12486 5960 12538
rect 5972 12486 6024 12538
rect 6036 12486 6088 12538
rect 7712 12486 7764 12538
rect 7776 12486 7828 12538
rect 7840 12486 7892 12538
rect 7904 12486 7956 12538
rect 7968 12486 8020 12538
rect 2320 12223 2372 12232
rect 2320 12189 2329 12223
rect 2329 12189 2363 12223
rect 2363 12189 2372 12223
rect 2320 12180 2372 12189
rect 2780 12180 2832 12232
rect 8300 12180 8352 12232
rect 2412 12087 2464 12096
rect 2412 12053 2421 12087
rect 2421 12053 2455 12087
rect 2455 12053 2464 12087
rect 2412 12044 2464 12053
rect 2882 11942 2934 11994
rect 2946 11942 2998 11994
rect 3010 11942 3062 11994
rect 3074 11942 3126 11994
rect 3138 11942 3190 11994
rect 4814 11942 4866 11994
rect 4878 11942 4930 11994
rect 4942 11942 4994 11994
rect 5006 11942 5058 11994
rect 5070 11942 5122 11994
rect 6746 11942 6798 11994
rect 6810 11942 6862 11994
rect 6874 11942 6926 11994
rect 6938 11942 6990 11994
rect 7002 11942 7054 11994
rect 8678 11942 8730 11994
rect 8742 11942 8794 11994
rect 8806 11942 8858 11994
rect 8870 11942 8922 11994
rect 8934 11942 8986 11994
rect 1768 11840 1820 11892
rect 2412 11840 2464 11892
rect 2780 11840 2832 11892
rect 940 11704 992 11756
rect 2964 11679 3016 11688
rect 2964 11645 2973 11679
rect 2973 11645 3007 11679
rect 3007 11645 3016 11679
rect 2964 11636 3016 11645
rect 2504 11611 2556 11620
rect 2504 11577 2513 11611
rect 2513 11577 2547 11611
rect 2547 11577 2556 11611
rect 2504 11568 2556 11577
rect 1916 11398 1968 11450
rect 1980 11398 2032 11450
rect 2044 11398 2096 11450
rect 2108 11398 2160 11450
rect 2172 11398 2224 11450
rect 3848 11398 3900 11450
rect 3912 11398 3964 11450
rect 3976 11398 4028 11450
rect 4040 11398 4092 11450
rect 4104 11398 4156 11450
rect 5780 11398 5832 11450
rect 5844 11398 5896 11450
rect 5908 11398 5960 11450
rect 5972 11398 6024 11450
rect 6036 11398 6088 11450
rect 7712 11398 7764 11450
rect 7776 11398 7828 11450
rect 7840 11398 7892 11450
rect 7904 11398 7956 11450
rect 7968 11398 8020 11450
rect 2504 11296 2556 11348
rect 8208 11067 8260 11076
rect 8208 11033 8217 11067
rect 8217 11033 8251 11067
rect 8251 11033 8260 11067
rect 8208 11024 8260 11033
rect 2882 10854 2934 10906
rect 2946 10854 2998 10906
rect 3010 10854 3062 10906
rect 3074 10854 3126 10906
rect 3138 10854 3190 10906
rect 4814 10854 4866 10906
rect 4878 10854 4930 10906
rect 4942 10854 4994 10906
rect 5006 10854 5058 10906
rect 5070 10854 5122 10906
rect 6746 10854 6798 10906
rect 6810 10854 6862 10906
rect 6874 10854 6926 10906
rect 6938 10854 6990 10906
rect 7002 10854 7054 10906
rect 8678 10854 8730 10906
rect 8742 10854 8794 10906
rect 8806 10854 8858 10906
rect 8870 10854 8922 10906
rect 8934 10854 8986 10906
rect 940 10616 992 10668
rect 1492 10412 1544 10464
rect 1916 10310 1968 10362
rect 1980 10310 2032 10362
rect 2044 10310 2096 10362
rect 2108 10310 2160 10362
rect 2172 10310 2224 10362
rect 3848 10310 3900 10362
rect 3912 10310 3964 10362
rect 3976 10310 4028 10362
rect 4040 10310 4092 10362
rect 4104 10310 4156 10362
rect 5780 10310 5832 10362
rect 5844 10310 5896 10362
rect 5908 10310 5960 10362
rect 5972 10310 6024 10362
rect 6036 10310 6088 10362
rect 7712 10310 7764 10362
rect 7776 10310 7828 10362
rect 7840 10310 7892 10362
rect 7904 10310 7956 10362
rect 7968 10310 8020 10362
rect 2882 9766 2934 9818
rect 2946 9766 2998 9818
rect 3010 9766 3062 9818
rect 3074 9766 3126 9818
rect 3138 9766 3190 9818
rect 4814 9766 4866 9818
rect 4878 9766 4930 9818
rect 4942 9766 4994 9818
rect 5006 9766 5058 9818
rect 5070 9766 5122 9818
rect 6746 9766 6798 9818
rect 6810 9766 6862 9818
rect 6874 9766 6926 9818
rect 6938 9766 6990 9818
rect 7002 9766 7054 9818
rect 8678 9766 8730 9818
rect 8742 9766 8794 9818
rect 8806 9766 8858 9818
rect 8870 9766 8922 9818
rect 8934 9766 8986 9818
rect 1584 9571 1636 9580
rect 1584 9537 1593 9571
rect 1593 9537 1627 9571
rect 1627 9537 1636 9571
rect 1584 9528 1636 9537
rect 1676 9571 1728 9580
rect 1676 9537 1685 9571
rect 1685 9537 1719 9571
rect 1719 9537 1728 9571
rect 1676 9528 1728 9537
rect 1492 9503 1544 9512
rect 1492 9469 1501 9503
rect 1501 9469 1535 9503
rect 1535 9469 1544 9503
rect 1492 9460 1544 9469
rect 2412 9460 2464 9512
rect 2596 9324 2648 9376
rect 1916 9222 1968 9274
rect 1980 9222 2032 9274
rect 2044 9222 2096 9274
rect 2108 9222 2160 9274
rect 2172 9222 2224 9274
rect 3848 9222 3900 9274
rect 3912 9222 3964 9274
rect 3976 9222 4028 9274
rect 4040 9222 4092 9274
rect 4104 9222 4156 9274
rect 5780 9222 5832 9274
rect 5844 9222 5896 9274
rect 5908 9222 5960 9274
rect 5972 9222 6024 9274
rect 6036 9222 6088 9274
rect 7712 9222 7764 9274
rect 7776 9222 7828 9274
rect 7840 9222 7892 9274
rect 7904 9222 7956 9274
rect 7968 9222 8020 9274
rect 940 8916 992 8968
rect 1584 8823 1636 8832
rect 1584 8789 1593 8823
rect 1593 8789 1627 8823
rect 1627 8789 1636 8823
rect 1584 8780 1636 8789
rect 2882 8678 2934 8730
rect 2946 8678 2998 8730
rect 3010 8678 3062 8730
rect 3074 8678 3126 8730
rect 3138 8678 3190 8730
rect 4814 8678 4866 8730
rect 4878 8678 4930 8730
rect 4942 8678 4994 8730
rect 5006 8678 5058 8730
rect 5070 8678 5122 8730
rect 6746 8678 6798 8730
rect 6810 8678 6862 8730
rect 6874 8678 6926 8730
rect 6938 8678 6990 8730
rect 7002 8678 7054 8730
rect 8678 8678 8730 8730
rect 8742 8678 8794 8730
rect 8806 8678 8858 8730
rect 8870 8678 8922 8730
rect 8934 8678 8986 8730
rect 1584 8576 1636 8628
rect 2412 8576 2464 8628
rect 2596 8576 2648 8628
rect 2688 8619 2740 8628
rect 2688 8585 2697 8619
rect 2697 8585 2731 8619
rect 2731 8585 2740 8619
rect 2688 8576 2740 8585
rect 1676 8508 1728 8560
rect 2504 8440 2556 8492
rect 1676 8415 1728 8424
rect 1676 8381 1685 8415
rect 1685 8381 1719 8415
rect 1719 8381 1728 8415
rect 1676 8372 1728 8381
rect 2504 8279 2556 8288
rect 2504 8245 2513 8279
rect 2513 8245 2547 8279
rect 2547 8245 2556 8279
rect 2504 8236 2556 8245
rect 1916 8134 1968 8186
rect 1980 8134 2032 8186
rect 2044 8134 2096 8186
rect 2108 8134 2160 8186
rect 2172 8134 2224 8186
rect 3848 8134 3900 8186
rect 3912 8134 3964 8186
rect 3976 8134 4028 8186
rect 4040 8134 4092 8186
rect 4104 8134 4156 8186
rect 5780 8134 5832 8186
rect 5844 8134 5896 8186
rect 5908 8134 5960 8186
rect 5972 8134 6024 8186
rect 6036 8134 6088 8186
rect 7712 8134 7764 8186
rect 7776 8134 7828 8186
rect 7840 8134 7892 8186
rect 7904 8134 7956 8186
rect 7968 8134 8020 8186
rect 1768 8075 1820 8084
rect 1768 8041 1777 8075
rect 1777 8041 1811 8075
rect 1811 8041 1820 8075
rect 1768 8032 1820 8041
rect 2504 8032 2556 8084
rect 1492 7964 1544 8016
rect 2412 7964 2464 8016
rect 1768 7735 1820 7744
rect 1768 7701 1777 7735
rect 1777 7701 1811 7735
rect 1811 7701 1820 7735
rect 1768 7692 1820 7701
rect 2882 7590 2934 7642
rect 2946 7590 2998 7642
rect 3010 7590 3062 7642
rect 3074 7590 3126 7642
rect 3138 7590 3190 7642
rect 4814 7590 4866 7642
rect 4878 7590 4930 7642
rect 4942 7590 4994 7642
rect 5006 7590 5058 7642
rect 5070 7590 5122 7642
rect 6746 7590 6798 7642
rect 6810 7590 6862 7642
rect 6874 7590 6926 7642
rect 6938 7590 6990 7642
rect 7002 7590 7054 7642
rect 8678 7590 8730 7642
rect 8742 7590 8794 7642
rect 8806 7590 8858 7642
rect 8870 7590 8922 7642
rect 8934 7590 8986 7642
rect 1768 7488 1820 7540
rect 940 7352 992 7404
rect 1916 7046 1968 7098
rect 1980 7046 2032 7098
rect 2044 7046 2096 7098
rect 2108 7046 2160 7098
rect 2172 7046 2224 7098
rect 3848 7046 3900 7098
rect 3912 7046 3964 7098
rect 3976 7046 4028 7098
rect 4040 7046 4092 7098
rect 4104 7046 4156 7098
rect 5780 7046 5832 7098
rect 5844 7046 5896 7098
rect 5908 7046 5960 7098
rect 5972 7046 6024 7098
rect 6036 7046 6088 7098
rect 7712 7046 7764 7098
rect 7776 7046 7828 7098
rect 7840 7046 7892 7098
rect 7904 7046 7956 7098
rect 7968 7046 8020 7098
rect 2320 6808 2372 6860
rect 1952 6740 2004 6792
rect 2688 6740 2740 6792
rect 1400 6672 1452 6724
rect 2412 6672 2464 6724
rect 1768 6647 1820 6656
rect 1768 6613 1777 6647
rect 1777 6613 1811 6647
rect 1811 6613 1820 6647
rect 1768 6604 1820 6613
rect 1860 6647 1912 6656
rect 1860 6613 1869 6647
rect 1869 6613 1903 6647
rect 1903 6613 1912 6647
rect 1860 6604 1912 6613
rect 2780 6604 2832 6656
rect 2882 6502 2934 6554
rect 2946 6502 2998 6554
rect 3010 6502 3062 6554
rect 3074 6502 3126 6554
rect 3138 6502 3190 6554
rect 4814 6502 4866 6554
rect 4878 6502 4930 6554
rect 4942 6502 4994 6554
rect 5006 6502 5058 6554
rect 5070 6502 5122 6554
rect 6746 6502 6798 6554
rect 6810 6502 6862 6554
rect 6874 6502 6926 6554
rect 6938 6502 6990 6554
rect 7002 6502 7054 6554
rect 8678 6502 8730 6554
rect 8742 6502 8794 6554
rect 8806 6502 8858 6554
rect 8870 6502 8922 6554
rect 8934 6502 8986 6554
rect 1768 6400 1820 6452
rect 1492 6264 1544 6316
rect 1584 6307 1636 6316
rect 1584 6273 1593 6307
rect 1593 6273 1627 6307
rect 1627 6273 1636 6307
rect 1584 6264 1636 6273
rect 1952 6332 2004 6384
rect 1400 6060 1452 6112
rect 2412 6307 2464 6316
rect 2412 6273 2421 6307
rect 2421 6273 2455 6307
rect 2455 6273 2464 6307
rect 2412 6264 2464 6273
rect 2504 6307 2556 6316
rect 2504 6273 2513 6307
rect 2513 6273 2547 6307
rect 2547 6273 2556 6307
rect 2504 6264 2556 6273
rect 1916 5958 1968 6010
rect 1980 5958 2032 6010
rect 2044 5958 2096 6010
rect 2108 5958 2160 6010
rect 2172 5958 2224 6010
rect 3848 5958 3900 6010
rect 3912 5958 3964 6010
rect 3976 5958 4028 6010
rect 4040 5958 4092 6010
rect 4104 5958 4156 6010
rect 5780 5958 5832 6010
rect 5844 5958 5896 6010
rect 5908 5958 5960 6010
rect 5972 5958 6024 6010
rect 6036 5958 6088 6010
rect 7712 5958 7764 6010
rect 7776 5958 7828 6010
rect 7840 5958 7892 6010
rect 7904 5958 7956 6010
rect 7968 5958 8020 6010
rect 1676 5856 1728 5908
rect 1768 5856 1820 5908
rect 940 5652 992 5704
rect 1492 5652 1544 5704
rect 1952 5695 2004 5704
rect 1952 5661 1961 5695
rect 1961 5661 1995 5695
rect 1995 5661 2004 5695
rect 1952 5652 2004 5661
rect 2882 5414 2934 5466
rect 2946 5414 2998 5466
rect 3010 5414 3062 5466
rect 3074 5414 3126 5466
rect 3138 5414 3190 5466
rect 4814 5414 4866 5466
rect 4878 5414 4930 5466
rect 4942 5414 4994 5466
rect 5006 5414 5058 5466
rect 5070 5414 5122 5466
rect 6746 5414 6798 5466
rect 6810 5414 6862 5466
rect 6874 5414 6926 5466
rect 6938 5414 6990 5466
rect 7002 5414 7054 5466
rect 8678 5414 8730 5466
rect 8742 5414 8794 5466
rect 8806 5414 8858 5466
rect 8870 5414 8922 5466
rect 8934 5414 8986 5466
rect 1952 5312 2004 5364
rect 1768 5219 1820 5228
rect 1768 5185 1777 5219
rect 1777 5185 1811 5219
rect 1811 5185 1820 5219
rect 1768 5176 1820 5185
rect 1400 5108 1452 5160
rect 1676 5151 1728 5160
rect 1676 5117 1685 5151
rect 1685 5117 1719 5151
rect 1719 5117 1728 5151
rect 1676 5108 1728 5117
rect 1916 4870 1968 4922
rect 1980 4870 2032 4922
rect 2044 4870 2096 4922
rect 2108 4870 2160 4922
rect 2172 4870 2224 4922
rect 3848 4870 3900 4922
rect 3912 4870 3964 4922
rect 3976 4870 4028 4922
rect 4040 4870 4092 4922
rect 4104 4870 4156 4922
rect 5780 4870 5832 4922
rect 5844 4870 5896 4922
rect 5908 4870 5960 4922
rect 5972 4870 6024 4922
rect 6036 4870 6088 4922
rect 7712 4870 7764 4922
rect 7776 4870 7828 4922
rect 7840 4870 7892 4922
rect 7904 4870 7956 4922
rect 7968 4870 8020 4922
rect 1584 4811 1636 4820
rect 1584 4777 1593 4811
rect 1593 4777 1627 4811
rect 1627 4777 1636 4811
rect 1584 4768 1636 4777
rect 940 4564 992 4616
rect 2882 4326 2934 4378
rect 2946 4326 2998 4378
rect 3010 4326 3062 4378
rect 3074 4326 3126 4378
rect 3138 4326 3190 4378
rect 4814 4326 4866 4378
rect 4878 4326 4930 4378
rect 4942 4326 4994 4378
rect 5006 4326 5058 4378
rect 5070 4326 5122 4378
rect 6746 4326 6798 4378
rect 6810 4326 6862 4378
rect 6874 4326 6926 4378
rect 6938 4326 6990 4378
rect 7002 4326 7054 4378
rect 8678 4326 8730 4378
rect 8742 4326 8794 4378
rect 8806 4326 8858 4378
rect 8870 4326 8922 4378
rect 8934 4326 8986 4378
rect 1916 3782 1968 3834
rect 1980 3782 2032 3834
rect 2044 3782 2096 3834
rect 2108 3782 2160 3834
rect 2172 3782 2224 3834
rect 3848 3782 3900 3834
rect 3912 3782 3964 3834
rect 3976 3782 4028 3834
rect 4040 3782 4092 3834
rect 4104 3782 4156 3834
rect 5780 3782 5832 3834
rect 5844 3782 5896 3834
rect 5908 3782 5960 3834
rect 5972 3782 6024 3834
rect 6036 3782 6088 3834
rect 7712 3782 7764 3834
rect 7776 3782 7828 3834
rect 7840 3782 7892 3834
rect 7904 3782 7956 3834
rect 7968 3782 8020 3834
rect 1768 3680 1820 3732
rect 940 3476 992 3528
rect 2882 3238 2934 3290
rect 2946 3238 2998 3290
rect 3010 3238 3062 3290
rect 3074 3238 3126 3290
rect 3138 3238 3190 3290
rect 4814 3238 4866 3290
rect 4878 3238 4930 3290
rect 4942 3238 4994 3290
rect 5006 3238 5058 3290
rect 5070 3238 5122 3290
rect 6746 3238 6798 3290
rect 6810 3238 6862 3290
rect 6874 3238 6926 3290
rect 6938 3238 6990 3290
rect 7002 3238 7054 3290
rect 8678 3238 8730 3290
rect 8742 3238 8794 3290
rect 8806 3238 8858 3290
rect 8870 3238 8922 3290
rect 8934 3238 8986 3290
rect 1916 2694 1968 2746
rect 1980 2694 2032 2746
rect 2044 2694 2096 2746
rect 2108 2694 2160 2746
rect 2172 2694 2224 2746
rect 3848 2694 3900 2746
rect 3912 2694 3964 2746
rect 3976 2694 4028 2746
rect 4040 2694 4092 2746
rect 4104 2694 4156 2746
rect 5780 2694 5832 2746
rect 5844 2694 5896 2746
rect 5908 2694 5960 2746
rect 5972 2694 6024 2746
rect 6036 2694 6088 2746
rect 7712 2694 7764 2746
rect 7776 2694 7828 2746
rect 7840 2694 7892 2746
rect 7904 2694 7956 2746
rect 7968 2694 8020 2746
rect 1676 2592 1728 2644
rect 2504 2592 2556 2644
rect 940 2388 992 2440
rect 1676 2431 1728 2440
rect 1676 2397 1685 2431
rect 1685 2397 1719 2431
rect 1719 2397 1728 2431
rect 1676 2388 1728 2397
rect 2882 2150 2934 2202
rect 2946 2150 2998 2202
rect 3010 2150 3062 2202
rect 3074 2150 3126 2202
rect 3138 2150 3190 2202
rect 4814 2150 4866 2202
rect 4878 2150 4930 2202
rect 4942 2150 4994 2202
rect 5006 2150 5058 2202
rect 5070 2150 5122 2202
rect 6746 2150 6798 2202
rect 6810 2150 6862 2202
rect 6874 2150 6926 2202
rect 6938 2150 6990 2202
rect 7002 2150 7054 2202
rect 8678 2150 8730 2202
rect 8742 2150 8794 2202
rect 8806 2150 8858 2202
rect 8870 2150 8922 2202
rect 8934 2150 8986 2202
<< metal2 >>
rect 1214 21298 1270 22000
rect 1214 21270 1440 21298
rect 1214 21200 1270 21270
rect 1030 21040 1086 21049
rect 1030 20975 1086 20984
rect 1044 19378 1072 20975
rect 1122 19680 1178 19689
rect 1122 19615 1178 19624
rect 1136 19514 1164 19615
rect 1124 19508 1176 19514
rect 1124 19450 1176 19456
rect 1412 19446 1440 21270
rect 3698 21200 3754 22000
rect 6182 21200 6238 22000
rect 8666 21298 8722 22000
rect 8588 21270 8722 21298
rect 2882 19612 3190 19621
rect 2882 19610 2888 19612
rect 2944 19610 2968 19612
rect 3024 19610 3048 19612
rect 3104 19610 3128 19612
rect 3184 19610 3190 19612
rect 2944 19558 2946 19610
rect 3126 19558 3128 19610
rect 2882 19556 2888 19558
rect 2944 19556 2968 19558
rect 3024 19556 3048 19558
rect 3104 19556 3128 19558
rect 3184 19556 3190 19558
rect 2882 19547 3190 19556
rect 1768 19508 1820 19514
rect 1768 19450 1820 19456
rect 2504 19508 2556 19514
rect 2504 19450 2556 19456
rect 1400 19440 1452 19446
rect 1400 19382 1452 19388
rect 1032 19372 1084 19378
rect 1032 19314 1084 19320
rect 1676 19168 1728 19174
rect 1676 19110 1728 19116
rect 940 18760 992 18766
rect 1688 18714 1716 19110
rect 940 18702 992 18708
rect 952 18329 980 18702
rect 1504 18686 1716 18714
rect 938 18320 994 18329
rect 938 18255 994 18264
rect 940 17196 992 17202
rect 940 17138 992 17144
rect 952 16969 980 17138
rect 1400 16992 1452 16998
rect 938 16960 994 16969
rect 1400 16934 1452 16940
rect 1504 16946 1532 18686
rect 1584 18624 1636 18630
rect 1584 18566 1636 18572
rect 1596 17082 1624 18566
rect 1596 17054 1716 17082
rect 938 16895 994 16904
rect 938 15600 994 15609
rect 938 15535 994 15544
rect 952 15502 980 15535
rect 940 15496 992 15502
rect 940 15438 992 15444
rect 1412 15026 1440 16934
rect 1504 16918 1624 16946
rect 1492 16652 1544 16658
rect 1492 16594 1544 16600
rect 1504 16114 1532 16594
rect 1596 16114 1624 16918
rect 1688 16658 1716 17054
rect 1676 16652 1728 16658
rect 1676 16594 1728 16600
rect 1492 16108 1544 16114
rect 1492 16050 1544 16056
rect 1584 16108 1636 16114
rect 1584 16050 1636 16056
rect 1492 15972 1544 15978
rect 1492 15914 1544 15920
rect 1400 15020 1452 15026
rect 1400 14962 1452 14968
rect 940 14408 992 14414
rect 940 14350 992 14356
rect 952 14249 980 14350
rect 938 14240 994 14249
rect 938 14175 994 14184
rect 1504 13530 1532 15914
rect 1780 15722 1808 19450
rect 2320 19304 2372 19310
rect 2320 19246 2372 19252
rect 1916 19068 2224 19077
rect 1916 19066 1922 19068
rect 1978 19066 2002 19068
rect 2058 19066 2082 19068
rect 2138 19066 2162 19068
rect 2218 19066 2224 19068
rect 1978 19014 1980 19066
rect 2160 19014 2162 19066
rect 1916 19012 1922 19014
rect 1978 19012 2002 19014
rect 2058 19012 2082 19014
rect 2138 19012 2162 19014
rect 2218 19012 2224 19014
rect 1916 19003 2224 19012
rect 1916 17980 2224 17989
rect 1916 17978 1922 17980
rect 1978 17978 2002 17980
rect 2058 17978 2082 17980
rect 2138 17978 2162 17980
rect 2218 17978 2224 17980
rect 1978 17926 1980 17978
rect 2160 17926 2162 17978
rect 1916 17924 1922 17926
rect 1978 17924 2002 17926
rect 2058 17924 2082 17926
rect 2138 17924 2162 17926
rect 2218 17924 2224 17926
rect 1916 17915 2224 17924
rect 1916 16892 2224 16901
rect 1916 16890 1922 16892
rect 1978 16890 2002 16892
rect 2058 16890 2082 16892
rect 2138 16890 2162 16892
rect 2218 16890 2224 16892
rect 1978 16838 1980 16890
rect 2160 16838 2162 16890
rect 1916 16836 1922 16838
rect 1978 16836 2002 16838
rect 2058 16836 2082 16838
rect 2138 16836 2162 16838
rect 2218 16836 2224 16838
rect 1916 16827 2224 16836
rect 1916 15804 2224 15813
rect 1916 15802 1922 15804
rect 1978 15802 2002 15804
rect 2058 15802 2082 15804
rect 2138 15802 2162 15804
rect 2218 15802 2224 15804
rect 1978 15750 1980 15802
rect 2160 15750 2162 15802
rect 1916 15748 1922 15750
rect 1978 15748 2002 15750
rect 2058 15748 2082 15750
rect 2138 15748 2162 15750
rect 2218 15748 2224 15750
rect 1916 15739 2224 15748
rect 1596 15694 1808 15722
rect 1596 15026 1624 15694
rect 1584 15020 1636 15026
rect 1584 14962 1636 14968
rect 1768 14952 1820 14958
rect 1768 14894 1820 14900
rect 1676 14816 1728 14822
rect 1676 14758 1728 14764
rect 1584 14476 1636 14482
rect 1584 14418 1636 14424
rect 1492 13524 1544 13530
rect 1492 13466 1544 13472
rect 940 13320 992 13326
rect 940 13262 992 13268
rect 952 12889 980 13262
rect 938 12880 994 12889
rect 938 12815 994 12824
rect 940 11756 992 11762
rect 940 11698 992 11704
rect 952 11529 980 11698
rect 938 11520 994 11529
rect 938 11455 994 11464
rect 940 10668 992 10674
rect 940 10610 992 10616
rect 952 10169 980 10610
rect 1492 10464 1544 10470
rect 1492 10406 1544 10412
rect 938 10160 994 10169
rect 938 10095 994 10104
rect 1504 9518 1532 10406
rect 1596 9586 1624 14418
rect 1688 9586 1716 14758
rect 1780 11898 1808 14894
rect 1916 14716 2224 14725
rect 1916 14714 1922 14716
rect 1978 14714 2002 14716
rect 2058 14714 2082 14716
rect 2138 14714 2162 14716
rect 2218 14714 2224 14716
rect 1978 14662 1980 14714
rect 2160 14662 2162 14714
rect 1916 14660 1922 14662
rect 1978 14660 2002 14662
rect 2058 14660 2082 14662
rect 2138 14660 2162 14662
rect 2218 14660 2224 14662
rect 1916 14651 2224 14660
rect 2332 14482 2360 19246
rect 2412 16040 2464 16046
rect 2412 15982 2464 15988
rect 2424 15706 2452 15982
rect 2516 15910 2544 19450
rect 3712 19378 3740 21200
rect 4814 19612 5122 19621
rect 4814 19610 4820 19612
rect 4876 19610 4900 19612
rect 4956 19610 4980 19612
rect 5036 19610 5060 19612
rect 5116 19610 5122 19612
rect 4876 19558 4878 19610
rect 5058 19558 5060 19610
rect 4814 19556 4820 19558
rect 4876 19556 4900 19558
rect 4956 19556 4980 19558
rect 5036 19556 5060 19558
rect 5116 19556 5122 19558
rect 4814 19547 5122 19556
rect 6196 19446 6224 21200
rect 6746 19612 7054 19621
rect 6746 19610 6752 19612
rect 6808 19610 6832 19612
rect 6888 19610 6912 19612
rect 6968 19610 6992 19612
rect 7048 19610 7054 19612
rect 6808 19558 6810 19610
rect 6990 19558 6992 19610
rect 6746 19556 6752 19558
rect 6808 19556 6832 19558
rect 6888 19556 6912 19558
rect 6968 19556 6992 19558
rect 7048 19556 7054 19558
rect 6746 19547 7054 19556
rect 8588 19514 8616 21270
rect 8666 21200 8722 21270
rect 8678 19612 8986 19621
rect 8678 19610 8684 19612
rect 8740 19610 8764 19612
rect 8820 19610 8844 19612
rect 8900 19610 8924 19612
rect 8980 19610 8986 19612
rect 8740 19558 8742 19610
rect 8922 19558 8924 19610
rect 8678 19556 8684 19558
rect 8740 19556 8764 19558
rect 8820 19556 8844 19558
rect 8900 19556 8924 19558
rect 8980 19556 8986 19558
rect 8678 19547 8986 19556
rect 8576 19508 8628 19514
rect 8576 19450 8628 19456
rect 6184 19440 6236 19446
rect 6184 19382 6236 19388
rect 3700 19372 3752 19378
rect 3700 19314 3752 19320
rect 6368 19236 6420 19242
rect 6368 19178 6420 19184
rect 3848 19068 4156 19077
rect 3848 19066 3854 19068
rect 3910 19066 3934 19068
rect 3990 19066 4014 19068
rect 4070 19066 4094 19068
rect 4150 19066 4156 19068
rect 3910 19014 3912 19066
rect 4092 19014 4094 19066
rect 3848 19012 3854 19014
rect 3910 19012 3934 19014
rect 3990 19012 4014 19014
rect 4070 19012 4094 19014
rect 4150 19012 4156 19014
rect 3848 19003 4156 19012
rect 5780 19068 6088 19077
rect 5780 19066 5786 19068
rect 5842 19066 5866 19068
rect 5922 19066 5946 19068
rect 6002 19066 6026 19068
rect 6082 19066 6088 19068
rect 5842 19014 5844 19066
rect 6024 19014 6026 19066
rect 5780 19012 5786 19014
rect 5842 19012 5866 19014
rect 5922 19012 5946 19014
rect 6002 19012 6026 19014
rect 6082 19012 6088 19014
rect 5780 19003 6088 19012
rect 2882 18524 3190 18533
rect 2882 18522 2888 18524
rect 2944 18522 2968 18524
rect 3024 18522 3048 18524
rect 3104 18522 3128 18524
rect 3184 18522 3190 18524
rect 2944 18470 2946 18522
rect 3126 18470 3128 18522
rect 2882 18468 2888 18470
rect 2944 18468 2968 18470
rect 3024 18468 3048 18470
rect 3104 18468 3128 18470
rect 3184 18468 3190 18470
rect 2882 18459 3190 18468
rect 4814 18524 5122 18533
rect 4814 18522 4820 18524
rect 4876 18522 4900 18524
rect 4956 18522 4980 18524
rect 5036 18522 5060 18524
rect 5116 18522 5122 18524
rect 4876 18470 4878 18522
rect 5058 18470 5060 18522
rect 4814 18468 4820 18470
rect 4876 18468 4900 18470
rect 4956 18468 4980 18470
rect 5036 18468 5060 18470
rect 5116 18468 5122 18470
rect 4814 18459 5122 18468
rect 3848 17980 4156 17989
rect 3848 17978 3854 17980
rect 3910 17978 3934 17980
rect 3990 17978 4014 17980
rect 4070 17978 4094 17980
rect 4150 17978 4156 17980
rect 3910 17926 3912 17978
rect 4092 17926 4094 17978
rect 3848 17924 3854 17926
rect 3910 17924 3934 17926
rect 3990 17924 4014 17926
rect 4070 17924 4094 17926
rect 4150 17924 4156 17926
rect 3848 17915 4156 17924
rect 5780 17980 6088 17989
rect 5780 17978 5786 17980
rect 5842 17978 5866 17980
rect 5922 17978 5946 17980
rect 6002 17978 6026 17980
rect 6082 17978 6088 17980
rect 5842 17926 5844 17978
rect 6024 17926 6026 17978
rect 5780 17924 5786 17926
rect 5842 17924 5866 17926
rect 5922 17924 5946 17926
rect 6002 17924 6026 17926
rect 6082 17924 6088 17926
rect 5780 17915 6088 17924
rect 2882 17436 3190 17445
rect 2882 17434 2888 17436
rect 2944 17434 2968 17436
rect 3024 17434 3048 17436
rect 3104 17434 3128 17436
rect 3184 17434 3190 17436
rect 2944 17382 2946 17434
rect 3126 17382 3128 17434
rect 2882 17380 2888 17382
rect 2944 17380 2968 17382
rect 3024 17380 3048 17382
rect 3104 17380 3128 17382
rect 3184 17380 3190 17382
rect 2882 17371 3190 17380
rect 4814 17436 5122 17445
rect 4814 17434 4820 17436
rect 4876 17434 4900 17436
rect 4956 17434 4980 17436
rect 5036 17434 5060 17436
rect 5116 17434 5122 17436
rect 4876 17382 4878 17434
rect 5058 17382 5060 17434
rect 4814 17380 4820 17382
rect 4876 17380 4900 17382
rect 4956 17380 4980 17382
rect 5036 17380 5060 17382
rect 5116 17380 5122 17382
rect 4814 17371 5122 17380
rect 3848 16892 4156 16901
rect 3848 16890 3854 16892
rect 3910 16890 3934 16892
rect 3990 16890 4014 16892
rect 4070 16890 4094 16892
rect 4150 16890 4156 16892
rect 3910 16838 3912 16890
rect 4092 16838 4094 16890
rect 3848 16836 3854 16838
rect 3910 16836 3934 16838
rect 3990 16836 4014 16838
rect 4070 16836 4094 16838
rect 4150 16836 4156 16838
rect 3848 16827 4156 16836
rect 5780 16892 6088 16901
rect 5780 16890 5786 16892
rect 5842 16890 5866 16892
rect 5922 16890 5946 16892
rect 6002 16890 6026 16892
rect 6082 16890 6088 16892
rect 5842 16838 5844 16890
rect 6024 16838 6026 16890
rect 5780 16836 5786 16838
rect 5842 16836 5866 16838
rect 5922 16836 5946 16838
rect 6002 16836 6026 16838
rect 6082 16836 6088 16838
rect 5780 16827 6088 16836
rect 2882 16348 3190 16357
rect 2882 16346 2888 16348
rect 2944 16346 2968 16348
rect 3024 16346 3048 16348
rect 3104 16346 3128 16348
rect 3184 16346 3190 16348
rect 2944 16294 2946 16346
rect 3126 16294 3128 16346
rect 2882 16292 2888 16294
rect 2944 16292 2968 16294
rect 3024 16292 3048 16294
rect 3104 16292 3128 16294
rect 3184 16292 3190 16294
rect 2882 16283 3190 16292
rect 4814 16348 5122 16357
rect 4814 16346 4820 16348
rect 4876 16346 4900 16348
rect 4956 16346 4980 16348
rect 5036 16346 5060 16348
rect 5116 16346 5122 16348
rect 4876 16294 4878 16346
rect 5058 16294 5060 16346
rect 4814 16292 4820 16294
rect 4876 16292 4900 16294
rect 4956 16292 4980 16294
rect 5036 16292 5060 16294
rect 5116 16292 5122 16294
rect 4814 16283 5122 16292
rect 6380 16114 6408 19178
rect 8300 19168 8352 19174
rect 8300 19110 8352 19116
rect 7712 19068 8020 19077
rect 7712 19066 7718 19068
rect 7774 19066 7798 19068
rect 7854 19066 7878 19068
rect 7934 19066 7958 19068
rect 8014 19066 8020 19068
rect 7774 19014 7776 19066
rect 7956 19014 7958 19066
rect 7712 19012 7718 19014
rect 7774 19012 7798 19014
rect 7854 19012 7878 19014
rect 7934 19012 7958 19014
rect 8014 19012 8020 19014
rect 7712 19003 8020 19012
rect 6746 18524 7054 18533
rect 6746 18522 6752 18524
rect 6808 18522 6832 18524
rect 6888 18522 6912 18524
rect 6968 18522 6992 18524
rect 7048 18522 7054 18524
rect 6808 18470 6810 18522
rect 6990 18470 6992 18522
rect 6746 18468 6752 18470
rect 6808 18468 6832 18470
rect 6888 18468 6912 18470
rect 6968 18468 6992 18470
rect 7048 18468 7054 18470
rect 6746 18459 7054 18468
rect 7712 17980 8020 17989
rect 7712 17978 7718 17980
rect 7774 17978 7798 17980
rect 7854 17978 7878 17980
rect 7934 17978 7958 17980
rect 8014 17978 8020 17980
rect 7774 17926 7776 17978
rect 7956 17926 7958 17978
rect 7712 17924 7718 17926
rect 7774 17924 7798 17926
rect 7854 17924 7878 17926
rect 7934 17924 7958 17926
rect 8014 17924 8020 17926
rect 7712 17915 8020 17924
rect 6746 17436 7054 17445
rect 6746 17434 6752 17436
rect 6808 17434 6832 17436
rect 6888 17434 6912 17436
rect 6968 17434 6992 17436
rect 7048 17434 7054 17436
rect 6808 17382 6810 17434
rect 6990 17382 6992 17434
rect 6746 17380 6752 17382
rect 6808 17380 6832 17382
rect 6888 17380 6912 17382
rect 6968 17380 6992 17382
rect 7048 17380 7054 17382
rect 6746 17371 7054 17380
rect 7712 16892 8020 16901
rect 7712 16890 7718 16892
rect 7774 16890 7798 16892
rect 7854 16890 7878 16892
rect 7934 16890 7958 16892
rect 8014 16890 8020 16892
rect 7774 16838 7776 16890
rect 7956 16838 7958 16890
rect 7712 16836 7718 16838
rect 7774 16836 7798 16838
rect 7854 16836 7878 16838
rect 7934 16836 7958 16838
rect 8014 16836 8020 16838
rect 7712 16827 8020 16836
rect 6746 16348 7054 16357
rect 6746 16346 6752 16348
rect 6808 16346 6832 16348
rect 6888 16346 6912 16348
rect 6968 16346 6992 16348
rect 7048 16346 7054 16348
rect 6808 16294 6810 16346
rect 6990 16294 6992 16346
rect 6746 16292 6752 16294
rect 6808 16292 6832 16294
rect 6888 16292 6912 16294
rect 6968 16292 6992 16294
rect 7048 16292 7054 16294
rect 6746 16283 7054 16292
rect 6368 16108 6420 16114
rect 6368 16050 6420 16056
rect 2596 16040 2648 16046
rect 2596 15982 2648 15988
rect 2504 15904 2556 15910
rect 2504 15846 2556 15852
rect 2412 15700 2464 15706
rect 2412 15642 2464 15648
rect 2412 14952 2464 14958
rect 2412 14894 2464 14900
rect 2424 14618 2452 14894
rect 2516 14822 2544 15846
rect 2608 15026 2636 15982
rect 2780 15904 2832 15910
rect 2780 15846 2832 15852
rect 2596 15020 2648 15026
rect 2596 14962 2648 14968
rect 2504 14816 2556 14822
rect 2504 14758 2556 14764
rect 2412 14612 2464 14618
rect 2412 14554 2464 14560
rect 2320 14476 2372 14482
rect 2320 14418 2372 14424
rect 2320 14272 2372 14278
rect 2320 14214 2372 14220
rect 1916 13628 2224 13637
rect 1916 13626 1922 13628
rect 1978 13626 2002 13628
rect 2058 13626 2082 13628
rect 2138 13626 2162 13628
rect 2218 13626 2224 13628
rect 1978 13574 1980 13626
rect 2160 13574 2162 13626
rect 1916 13572 1922 13574
rect 1978 13572 2002 13574
rect 2058 13572 2082 13574
rect 2138 13572 2162 13574
rect 2218 13572 2224 13574
rect 1916 13563 2224 13572
rect 1916 12540 2224 12549
rect 1916 12538 1922 12540
rect 1978 12538 2002 12540
rect 2058 12538 2082 12540
rect 2138 12538 2162 12540
rect 2218 12538 2224 12540
rect 1978 12486 1980 12538
rect 2160 12486 2162 12538
rect 1916 12484 1922 12486
rect 1978 12484 2002 12486
rect 2058 12484 2082 12486
rect 2138 12484 2162 12486
rect 2218 12484 2224 12486
rect 1916 12475 2224 12484
rect 2332 12238 2360 14214
rect 2320 12232 2372 12238
rect 2320 12174 2372 12180
rect 2412 12096 2464 12102
rect 2412 12038 2464 12044
rect 2424 11898 2452 12038
rect 1768 11892 1820 11898
rect 1768 11834 1820 11840
rect 2412 11892 2464 11898
rect 2412 11834 2464 11840
rect 2504 11620 2556 11626
rect 2504 11562 2556 11568
rect 1916 11452 2224 11461
rect 1916 11450 1922 11452
rect 1978 11450 2002 11452
rect 2058 11450 2082 11452
rect 2138 11450 2162 11452
rect 2218 11450 2224 11452
rect 1978 11398 1980 11450
rect 2160 11398 2162 11450
rect 1916 11396 1922 11398
rect 1978 11396 2002 11398
rect 2058 11396 2082 11398
rect 2138 11396 2162 11398
rect 2218 11396 2224 11398
rect 1916 11387 2224 11396
rect 2516 11354 2544 11562
rect 2504 11348 2556 11354
rect 2504 11290 2556 11296
rect 1916 10364 2224 10373
rect 1916 10362 1922 10364
rect 1978 10362 2002 10364
rect 2058 10362 2082 10364
rect 2138 10362 2162 10364
rect 2218 10362 2224 10364
rect 1978 10310 1980 10362
rect 2160 10310 2162 10362
rect 1916 10308 1922 10310
rect 1978 10308 2002 10310
rect 2058 10308 2082 10310
rect 2138 10308 2162 10310
rect 2218 10308 2224 10310
rect 1916 10299 2224 10308
rect 1584 9580 1636 9586
rect 1584 9522 1636 9528
rect 1676 9580 1728 9586
rect 1676 9522 1728 9528
rect 1492 9512 1544 9518
rect 1492 9454 1544 9460
rect 940 8968 992 8974
rect 1596 8922 1624 9522
rect 940 8910 992 8916
rect 952 8809 980 8910
rect 1504 8894 1624 8922
rect 938 8800 994 8809
rect 938 8735 994 8744
rect 1504 8022 1532 8894
rect 1584 8832 1636 8838
rect 1584 8774 1636 8780
rect 1596 8634 1624 8774
rect 1584 8628 1636 8634
rect 1584 8570 1636 8576
rect 1688 8566 1716 9522
rect 2412 9512 2464 9518
rect 2608 9466 2636 14962
rect 2792 14346 2820 15846
rect 3848 15804 4156 15813
rect 3848 15802 3854 15804
rect 3910 15802 3934 15804
rect 3990 15802 4014 15804
rect 4070 15802 4094 15804
rect 4150 15802 4156 15804
rect 3910 15750 3912 15802
rect 4092 15750 4094 15802
rect 3848 15748 3854 15750
rect 3910 15748 3934 15750
rect 3990 15748 4014 15750
rect 4070 15748 4094 15750
rect 4150 15748 4156 15750
rect 3848 15739 4156 15748
rect 5780 15804 6088 15813
rect 5780 15802 5786 15804
rect 5842 15802 5866 15804
rect 5922 15802 5946 15804
rect 6002 15802 6026 15804
rect 6082 15802 6088 15804
rect 5842 15750 5844 15802
rect 6024 15750 6026 15802
rect 5780 15748 5786 15750
rect 5842 15748 5866 15750
rect 5922 15748 5946 15750
rect 6002 15748 6026 15750
rect 6082 15748 6088 15750
rect 5780 15739 6088 15748
rect 7712 15804 8020 15813
rect 7712 15802 7718 15804
rect 7774 15802 7798 15804
rect 7854 15802 7878 15804
rect 7934 15802 7958 15804
rect 8014 15802 8020 15804
rect 7774 15750 7776 15802
rect 7956 15750 7958 15802
rect 7712 15748 7718 15750
rect 7774 15748 7798 15750
rect 7854 15748 7878 15750
rect 7934 15748 7958 15750
rect 8014 15748 8020 15750
rect 7712 15739 8020 15748
rect 2882 15260 3190 15269
rect 2882 15258 2888 15260
rect 2944 15258 2968 15260
rect 3024 15258 3048 15260
rect 3104 15258 3128 15260
rect 3184 15258 3190 15260
rect 2944 15206 2946 15258
rect 3126 15206 3128 15258
rect 2882 15204 2888 15206
rect 2944 15204 2968 15206
rect 3024 15204 3048 15206
rect 3104 15204 3128 15206
rect 3184 15204 3190 15206
rect 2882 15195 3190 15204
rect 4814 15260 5122 15269
rect 4814 15258 4820 15260
rect 4876 15258 4900 15260
rect 4956 15258 4980 15260
rect 5036 15258 5060 15260
rect 5116 15258 5122 15260
rect 4876 15206 4878 15258
rect 5058 15206 5060 15258
rect 4814 15204 4820 15206
rect 4876 15204 4900 15206
rect 4956 15204 4980 15206
rect 5036 15204 5060 15206
rect 5116 15204 5122 15206
rect 4814 15195 5122 15204
rect 6746 15260 7054 15269
rect 6746 15258 6752 15260
rect 6808 15258 6832 15260
rect 6888 15258 6912 15260
rect 6968 15258 6992 15260
rect 7048 15258 7054 15260
rect 6808 15206 6810 15258
rect 6990 15206 6992 15258
rect 6746 15204 6752 15206
rect 6808 15204 6832 15206
rect 6888 15204 6912 15206
rect 6968 15204 6992 15206
rect 7048 15204 7054 15206
rect 6746 15195 7054 15204
rect 3240 14816 3292 14822
rect 3240 14758 3292 14764
rect 3252 14618 3280 14758
rect 3848 14716 4156 14725
rect 3848 14714 3854 14716
rect 3910 14714 3934 14716
rect 3990 14714 4014 14716
rect 4070 14714 4094 14716
rect 4150 14714 4156 14716
rect 3910 14662 3912 14714
rect 4092 14662 4094 14714
rect 3848 14660 3854 14662
rect 3910 14660 3934 14662
rect 3990 14660 4014 14662
rect 4070 14660 4094 14662
rect 4150 14660 4156 14662
rect 3848 14651 4156 14660
rect 5780 14716 6088 14725
rect 5780 14714 5786 14716
rect 5842 14714 5866 14716
rect 5922 14714 5946 14716
rect 6002 14714 6026 14716
rect 6082 14714 6088 14716
rect 5842 14662 5844 14714
rect 6024 14662 6026 14714
rect 5780 14660 5786 14662
rect 5842 14660 5866 14662
rect 5922 14660 5946 14662
rect 6002 14660 6026 14662
rect 6082 14660 6088 14662
rect 5780 14651 6088 14660
rect 7712 14716 8020 14725
rect 7712 14714 7718 14716
rect 7774 14714 7798 14716
rect 7854 14714 7878 14716
rect 7934 14714 7958 14716
rect 8014 14714 8020 14716
rect 7774 14662 7776 14714
rect 7956 14662 7958 14714
rect 7712 14660 7718 14662
rect 7774 14660 7798 14662
rect 7854 14660 7878 14662
rect 7934 14660 7958 14662
rect 8014 14660 8020 14662
rect 7712 14651 8020 14660
rect 3240 14612 3292 14618
rect 3240 14554 3292 14560
rect 2780 14340 2832 14346
rect 2780 14282 2832 14288
rect 2882 14172 3190 14181
rect 2882 14170 2888 14172
rect 2944 14170 2968 14172
rect 3024 14170 3048 14172
rect 3104 14170 3128 14172
rect 3184 14170 3190 14172
rect 2944 14118 2946 14170
rect 3126 14118 3128 14170
rect 2882 14116 2888 14118
rect 2944 14116 2968 14118
rect 3024 14116 3048 14118
rect 3104 14116 3128 14118
rect 3184 14116 3190 14118
rect 2882 14107 3190 14116
rect 4814 14172 5122 14181
rect 4814 14170 4820 14172
rect 4876 14170 4900 14172
rect 4956 14170 4980 14172
rect 5036 14170 5060 14172
rect 5116 14170 5122 14172
rect 4876 14118 4878 14170
rect 5058 14118 5060 14170
rect 4814 14116 4820 14118
rect 4876 14116 4900 14118
rect 4956 14116 4980 14118
rect 5036 14116 5060 14118
rect 5116 14116 5122 14118
rect 4814 14107 5122 14116
rect 6746 14172 7054 14181
rect 6746 14170 6752 14172
rect 6808 14170 6832 14172
rect 6888 14170 6912 14172
rect 6968 14170 6992 14172
rect 7048 14170 7054 14172
rect 6808 14118 6810 14170
rect 6990 14118 6992 14170
rect 6746 14116 6752 14118
rect 6808 14116 6832 14118
rect 6888 14116 6912 14118
rect 6968 14116 6992 14118
rect 7048 14116 7054 14118
rect 6746 14107 7054 14116
rect 3848 13628 4156 13637
rect 3848 13626 3854 13628
rect 3910 13626 3934 13628
rect 3990 13626 4014 13628
rect 4070 13626 4094 13628
rect 4150 13626 4156 13628
rect 3910 13574 3912 13626
rect 4092 13574 4094 13626
rect 3848 13572 3854 13574
rect 3910 13572 3934 13574
rect 3990 13572 4014 13574
rect 4070 13572 4094 13574
rect 4150 13572 4156 13574
rect 3848 13563 4156 13572
rect 5780 13628 6088 13637
rect 5780 13626 5786 13628
rect 5842 13626 5866 13628
rect 5922 13626 5946 13628
rect 6002 13626 6026 13628
rect 6082 13626 6088 13628
rect 5842 13574 5844 13626
rect 6024 13574 6026 13626
rect 5780 13572 5786 13574
rect 5842 13572 5866 13574
rect 5922 13572 5946 13574
rect 6002 13572 6026 13574
rect 6082 13572 6088 13574
rect 5780 13563 6088 13572
rect 7712 13628 8020 13637
rect 7712 13626 7718 13628
rect 7774 13626 7798 13628
rect 7854 13626 7878 13628
rect 7934 13626 7958 13628
rect 8014 13626 8020 13628
rect 7774 13574 7776 13626
rect 7956 13574 7958 13626
rect 7712 13572 7718 13574
rect 7774 13572 7798 13574
rect 7854 13572 7878 13574
rect 7934 13572 7958 13574
rect 8014 13572 8020 13574
rect 7712 13563 8020 13572
rect 2882 13084 3190 13093
rect 2882 13082 2888 13084
rect 2944 13082 2968 13084
rect 3024 13082 3048 13084
rect 3104 13082 3128 13084
rect 3184 13082 3190 13084
rect 2944 13030 2946 13082
rect 3126 13030 3128 13082
rect 2882 13028 2888 13030
rect 2944 13028 2968 13030
rect 3024 13028 3048 13030
rect 3104 13028 3128 13030
rect 3184 13028 3190 13030
rect 2882 13019 3190 13028
rect 4814 13084 5122 13093
rect 4814 13082 4820 13084
rect 4876 13082 4900 13084
rect 4956 13082 4980 13084
rect 5036 13082 5060 13084
rect 5116 13082 5122 13084
rect 4876 13030 4878 13082
rect 5058 13030 5060 13082
rect 4814 13028 4820 13030
rect 4876 13028 4900 13030
rect 4956 13028 4980 13030
rect 5036 13028 5060 13030
rect 5116 13028 5122 13030
rect 4814 13019 5122 13028
rect 6746 13084 7054 13093
rect 6746 13082 6752 13084
rect 6808 13082 6832 13084
rect 6888 13082 6912 13084
rect 6968 13082 6992 13084
rect 7048 13082 7054 13084
rect 6808 13030 6810 13082
rect 6990 13030 6992 13082
rect 6746 13028 6752 13030
rect 6808 13028 6832 13030
rect 6888 13028 6912 13030
rect 6968 13028 6992 13030
rect 7048 13028 7054 13030
rect 6746 13019 7054 13028
rect 3848 12540 4156 12549
rect 3848 12538 3854 12540
rect 3910 12538 3934 12540
rect 3990 12538 4014 12540
rect 4070 12538 4094 12540
rect 4150 12538 4156 12540
rect 3910 12486 3912 12538
rect 4092 12486 4094 12538
rect 3848 12484 3854 12486
rect 3910 12484 3934 12486
rect 3990 12484 4014 12486
rect 4070 12484 4094 12486
rect 4150 12484 4156 12486
rect 3848 12475 4156 12484
rect 5780 12540 6088 12549
rect 5780 12538 5786 12540
rect 5842 12538 5866 12540
rect 5922 12538 5946 12540
rect 6002 12538 6026 12540
rect 6082 12538 6088 12540
rect 5842 12486 5844 12538
rect 6024 12486 6026 12538
rect 5780 12484 5786 12486
rect 5842 12484 5866 12486
rect 5922 12484 5946 12486
rect 6002 12484 6026 12486
rect 6082 12484 6088 12486
rect 5780 12475 6088 12484
rect 7712 12540 8020 12549
rect 7712 12538 7718 12540
rect 7774 12538 7798 12540
rect 7854 12538 7878 12540
rect 7934 12538 7958 12540
rect 8014 12538 8020 12540
rect 7774 12486 7776 12538
rect 7956 12486 7958 12538
rect 7712 12484 7718 12486
rect 7774 12484 7798 12486
rect 7854 12484 7878 12486
rect 7934 12484 7958 12486
rect 8014 12484 8020 12486
rect 7712 12475 8020 12484
rect 8312 12238 8340 19110
rect 8678 18524 8986 18533
rect 8678 18522 8684 18524
rect 8740 18522 8764 18524
rect 8820 18522 8844 18524
rect 8900 18522 8924 18524
rect 8980 18522 8986 18524
rect 8740 18470 8742 18522
rect 8922 18470 8924 18522
rect 8678 18468 8684 18470
rect 8740 18468 8764 18470
rect 8820 18468 8844 18470
rect 8900 18468 8924 18470
rect 8980 18468 8986 18470
rect 8678 18459 8986 18468
rect 8678 17436 8986 17445
rect 8678 17434 8684 17436
rect 8740 17434 8764 17436
rect 8820 17434 8844 17436
rect 8900 17434 8924 17436
rect 8980 17434 8986 17436
rect 8740 17382 8742 17434
rect 8922 17382 8924 17434
rect 8678 17380 8684 17382
rect 8740 17380 8764 17382
rect 8820 17380 8844 17382
rect 8900 17380 8924 17382
rect 8980 17380 8986 17382
rect 8678 17371 8986 17380
rect 8678 16348 8986 16357
rect 8678 16346 8684 16348
rect 8740 16346 8764 16348
rect 8820 16346 8844 16348
rect 8900 16346 8924 16348
rect 8980 16346 8986 16348
rect 8740 16294 8742 16346
rect 8922 16294 8924 16346
rect 8678 16292 8684 16294
rect 8740 16292 8764 16294
rect 8820 16292 8844 16294
rect 8900 16292 8924 16294
rect 8980 16292 8986 16294
rect 8678 16283 8986 16292
rect 8678 15260 8986 15269
rect 8678 15258 8684 15260
rect 8740 15258 8764 15260
rect 8820 15258 8844 15260
rect 8900 15258 8924 15260
rect 8980 15258 8986 15260
rect 8740 15206 8742 15258
rect 8922 15206 8924 15258
rect 8678 15204 8684 15206
rect 8740 15204 8764 15206
rect 8820 15204 8844 15206
rect 8900 15204 8924 15206
rect 8980 15204 8986 15206
rect 8678 15195 8986 15204
rect 8678 14172 8986 14181
rect 8678 14170 8684 14172
rect 8740 14170 8764 14172
rect 8820 14170 8844 14172
rect 8900 14170 8924 14172
rect 8980 14170 8986 14172
rect 8740 14118 8742 14170
rect 8922 14118 8924 14170
rect 8678 14116 8684 14118
rect 8740 14116 8764 14118
rect 8820 14116 8844 14118
rect 8900 14116 8924 14118
rect 8980 14116 8986 14118
rect 8678 14107 8986 14116
rect 8678 13084 8986 13093
rect 8678 13082 8684 13084
rect 8740 13082 8764 13084
rect 8820 13082 8844 13084
rect 8900 13082 8924 13084
rect 8980 13082 8986 13084
rect 8740 13030 8742 13082
rect 8922 13030 8924 13082
rect 8678 13028 8684 13030
rect 8740 13028 8764 13030
rect 8820 13028 8844 13030
rect 8900 13028 8924 13030
rect 8980 13028 8986 13030
rect 8678 13019 8986 13028
rect 2780 12232 2832 12238
rect 2780 12174 2832 12180
rect 8300 12232 8352 12238
rect 8300 12174 8352 12180
rect 2792 11898 2820 12174
rect 2882 11996 3190 12005
rect 2882 11994 2888 11996
rect 2944 11994 2968 11996
rect 3024 11994 3048 11996
rect 3104 11994 3128 11996
rect 3184 11994 3190 11996
rect 2944 11942 2946 11994
rect 3126 11942 3128 11994
rect 2882 11940 2888 11942
rect 2944 11940 2968 11942
rect 3024 11940 3048 11942
rect 3104 11940 3128 11942
rect 3184 11940 3190 11942
rect 2882 11931 3190 11940
rect 4814 11996 5122 12005
rect 4814 11994 4820 11996
rect 4876 11994 4900 11996
rect 4956 11994 4980 11996
rect 5036 11994 5060 11996
rect 5116 11994 5122 11996
rect 4876 11942 4878 11994
rect 5058 11942 5060 11994
rect 4814 11940 4820 11942
rect 4876 11940 4900 11942
rect 4956 11940 4980 11942
rect 5036 11940 5060 11942
rect 5116 11940 5122 11942
rect 4814 11931 5122 11940
rect 6746 11996 7054 12005
rect 6746 11994 6752 11996
rect 6808 11994 6832 11996
rect 6888 11994 6912 11996
rect 6968 11994 6992 11996
rect 7048 11994 7054 11996
rect 6808 11942 6810 11994
rect 6990 11942 6992 11994
rect 6746 11940 6752 11942
rect 6808 11940 6832 11942
rect 6888 11940 6912 11942
rect 6968 11940 6992 11942
rect 7048 11940 7054 11942
rect 6746 11931 7054 11940
rect 8678 11996 8986 12005
rect 8678 11994 8684 11996
rect 8740 11994 8764 11996
rect 8820 11994 8844 11996
rect 8900 11994 8924 11996
rect 8980 11994 8986 11996
rect 8740 11942 8742 11994
rect 8922 11942 8924 11994
rect 8678 11940 8684 11942
rect 8740 11940 8764 11942
rect 8820 11940 8844 11942
rect 8900 11940 8924 11942
rect 8980 11940 8986 11942
rect 8678 11931 8986 11940
rect 2780 11892 2832 11898
rect 2780 11834 2832 11840
rect 2964 11688 3016 11694
rect 2964 11630 3016 11636
rect 2976 11098 3004 11630
rect 3848 11452 4156 11461
rect 3848 11450 3854 11452
rect 3910 11450 3934 11452
rect 3990 11450 4014 11452
rect 4070 11450 4094 11452
rect 4150 11450 4156 11452
rect 3910 11398 3912 11450
rect 4092 11398 4094 11450
rect 3848 11396 3854 11398
rect 3910 11396 3934 11398
rect 3990 11396 4014 11398
rect 4070 11396 4094 11398
rect 4150 11396 4156 11398
rect 3848 11387 4156 11396
rect 5780 11452 6088 11461
rect 5780 11450 5786 11452
rect 5842 11450 5866 11452
rect 5922 11450 5946 11452
rect 6002 11450 6026 11452
rect 6082 11450 6088 11452
rect 5842 11398 5844 11450
rect 6024 11398 6026 11450
rect 5780 11396 5786 11398
rect 5842 11396 5866 11398
rect 5922 11396 5946 11398
rect 6002 11396 6026 11398
rect 6082 11396 6088 11398
rect 5780 11387 6088 11396
rect 7712 11452 8020 11461
rect 7712 11450 7718 11452
rect 7774 11450 7798 11452
rect 7854 11450 7878 11452
rect 7934 11450 7958 11452
rect 8014 11450 8020 11452
rect 7774 11398 7776 11450
rect 7956 11398 7958 11450
rect 7712 11396 7718 11398
rect 7774 11396 7798 11398
rect 7854 11396 7878 11398
rect 7934 11396 7958 11398
rect 8014 11396 8020 11398
rect 7712 11387 8020 11396
rect 2412 9454 2464 9460
rect 1916 9276 2224 9285
rect 1916 9274 1922 9276
rect 1978 9274 2002 9276
rect 2058 9274 2082 9276
rect 2138 9274 2162 9276
rect 2218 9274 2224 9276
rect 1978 9222 1980 9274
rect 2160 9222 2162 9274
rect 1916 9220 1922 9222
rect 1978 9220 2002 9222
rect 2058 9220 2082 9222
rect 2138 9220 2162 9222
rect 2218 9220 2224 9222
rect 1916 9211 2224 9220
rect 2424 8634 2452 9454
rect 2516 9438 2636 9466
rect 2792 11070 3004 11098
rect 8208 11076 8260 11082
rect 2412 8628 2464 8634
rect 2412 8570 2464 8576
rect 1676 8560 1728 8566
rect 1728 8508 1808 8514
rect 1676 8502 1808 8508
rect 1688 8486 1808 8502
rect 2516 8498 2544 9438
rect 2596 9376 2648 9382
rect 2596 9318 2648 9324
rect 2608 8634 2636 9318
rect 2596 8628 2648 8634
rect 2596 8570 2648 8576
rect 2688 8628 2740 8634
rect 2688 8570 2740 8576
rect 1676 8424 1728 8430
rect 1676 8366 1728 8372
rect 1492 8016 1544 8022
rect 1492 7958 1544 7964
rect 938 7440 994 7449
rect 938 7375 940 7384
rect 992 7375 994 7384
rect 940 7346 992 7352
rect 1400 6724 1452 6730
rect 1400 6666 1452 6672
rect 1412 6118 1440 6666
rect 1504 6322 1532 7958
rect 1492 6316 1544 6322
rect 1492 6258 1544 6264
rect 1584 6316 1636 6322
rect 1584 6258 1636 6264
rect 1400 6112 1452 6118
rect 938 6080 994 6089
rect 1400 6054 1452 6060
rect 938 6015 994 6024
rect 952 5710 980 6015
rect 940 5704 992 5710
rect 940 5646 992 5652
rect 1412 5166 1440 6054
rect 1504 5710 1532 6258
rect 1492 5704 1544 5710
rect 1492 5646 1544 5652
rect 1400 5160 1452 5166
rect 1400 5102 1452 5108
rect 1596 4826 1624 6258
rect 1688 5914 1716 8366
rect 1780 8090 1808 8486
rect 2504 8492 2556 8498
rect 2504 8434 2556 8440
rect 2516 8378 2544 8434
rect 2332 8350 2544 8378
rect 1916 8188 2224 8197
rect 1916 8186 1922 8188
rect 1978 8186 2002 8188
rect 2058 8186 2082 8188
rect 2138 8186 2162 8188
rect 2218 8186 2224 8188
rect 1978 8134 1980 8186
rect 2160 8134 2162 8186
rect 1916 8132 1922 8134
rect 1978 8132 2002 8134
rect 2058 8132 2082 8134
rect 2138 8132 2162 8134
rect 2218 8132 2224 8134
rect 1916 8123 2224 8132
rect 1768 8084 1820 8090
rect 1768 8026 1820 8032
rect 1768 7744 1820 7750
rect 1768 7686 1820 7692
rect 1780 7546 1808 7686
rect 1768 7540 1820 7546
rect 1768 7482 1820 7488
rect 1916 7100 2224 7109
rect 1916 7098 1922 7100
rect 1978 7098 2002 7100
rect 2058 7098 2082 7100
rect 2138 7098 2162 7100
rect 2218 7098 2224 7100
rect 1978 7046 1980 7098
rect 2160 7046 2162 7098
rect 1916 7044 1922 7046
rect 1978 7044 2002 7046
rect 2058 7044 2082 7046
rect 2138 7044 2162 7046
rect 2218 7044 2224 7046
rect 1916 7035 2224 7044
rect 2332 6866 2360 8350
rect 2504 8288 2556 8294
rect 2504 8230 2556 8236
rect 2516 8090 2544 8230
rect 2504 8084 2556 8090
rect 2504 8026 2556 8032
rect 2412 8016 2464 8022
rect 2412 7958 2464 7964
rect 2320 6860 2372 6866
rect 2320 6802 2372 6808
rect 1952 6792 2004 6798
rect 1952 6734 2004 6740
rect 1768 6656 1820 6662
rect 1768 6598 1820 6604
rect 1860 6656 1912 6662
rect 1860 6598 1912 6604
rect 1780 6458 1808 6598
rect 1768 6452 1820 6458
rect 1768 6394 1820 6400
rect 1872 6202 1900 6598
rect 1964 6390 1992 6734
rect 2424 6730 2452 7958
rect 2700 6798 2728 8570
rect 2688 6792 2740 6798
rect 2688 6734 2740 6740
rect 2412 6724 2464 6730
rect 2412 6666 2464 6672
rect 1952 6384 2004 6390
rect 1952 6326 2004 6332
rect 2424 6322 2452 6666
rect 2792 6662 2820 11070
rect 8208 11018 8260 11024
rect 2882 10908 3190 10917
rect 2882 10906 2888 10908
rect 2944 10906 2968 10908
rect 3024 10906 3048 10908
rect 3104 10906 3128 10908
rect 3184 10906 3190 10908
rect 2944 10854 2946 10906
rect 3126 10854 3128 10906
rect 2882 10852 2888 10854
rect 2944 10852 2968 10854
rect 3024 10852 3048 10854
rect 3104 10852 3128 10854
rect 3184 10852 3190 10854
rect 2882 10843 3190 10852
rect 4814 10908 5122 10917
rect 4814 10906 4820 10908
rect 4876 10906 4900 10908
rect 4956 10906 4980 10908
rect 5036 10906 5060 10908
rect 5116 10906 5122 10908
rect 4876 10854 4878 10906
rect 5058 10854 5060 10906
rect 4814 10852 4820 10854
rect 4876 10852 4900 10854
rect 4956 10852 4980 10854
rect 5036 10852 5060 10854
rect 5116 10852 5122 10854
rect 4814 10843 5122 10852
rect 6746 10908 7054 10917
rect 6746 10906 6752 10908
rect 6808 10906 6832 10908
rect 6888 10906 6912 10908
rect 6968 10906 6992 10908
rect 7048 10906 7054 10908
rect 6808 10854 6810 10906
rect 6990 10854 6992 10906
rect 6746 10852 6752 10854
rect 6808 10852 6832 10854
rect 6888 10852 6912 10854
rect 6968 10852 6992 10854
rect 7048 10852 7054 10854
rect 6746 10843 7054 10852
rect 8220 10713 8248 11018
rect 8678 10908 8986 10917
rect 8678 10906 8684 10908
rect 8740 10906 8764 10908
rect 8820 10906 8844 10908
rect 8900 10906 8924 10908
rect 8980 10906 8986 10908
rect 8740 10854 8742 10906
rect 8922 10854 8924 10906
rect 8678 10852 8684 10854
rect 8740 10852 8764 10854
rect 8820 10852 8844 10854
rect 8900 10852 8924 10854
rect 8980 10852 8986 10854
rect 8678 10843 8986 10852
rect 8206 10704 8262 10713
rect 8206 10639 8262 10648
rect 3848 10364 4156 10373
rect 3848 10362 3854 10364
rect 3910 10362 3934 10364
rect 3990 10362 4014 10364
rect 4070 10362 4094 10364
rect 4150 10362 4156 10364
rect 3910 10310 3912 10362
rect 4092 10310 4094 10362
rect 3848 10308 3854 10310
rect 3910 10308 3934 10310
rect 3990 10308 4014 10310
rect 4070 10308 4094 10310
rect 4150 10308 4156 10310
rect 3848 10299 4156 10308
rect 5780 10364 6088 10373
rect 5780 10362 5786 10364
rect 5842 10362 5866 10364
rect 5922 10362 5946 10364
rect 6002 10362 6026 10364
rect 6082 10362 6088 10364
rect 5842 10310 5844 10362
rect 6024 10310 6026 10362
rect 5780 10308 5786 10310
rect 5842 10308 5866 10310
rect 5922 10308 5946 10310
rect 6002 10308 6026 10310
rect 6082 10308 6088 10310
rect 5780 10299 6088 10308
rect 7712 10364 8020 10373
rect 7712 10362 7718 10364
rect 7774 10362 7798 10364
rect 7854 10362 7878 10364
rect 7934 10362 7958 10364
rect 8014 10362 8020 10364
rect 7774 10310 7776 10362
rect 7956 10310 7958 10362
rect 7712 10308 7718 10310
rect 7774 10308 7798 10310
rect 7854 10308 7878 10310
rect 7934 10308 7958 10310
rect 8014 10308 8020 10310
rect 7712 10299 8020 10308
rect 2882 9820 3190 9829
rect 2882 9818 2888 9820
rect 2944 9818 2968 9820
rect 3024 9818 3048 9820
rect 3104 9818 3128 9820
rect 3184 9818 3190 9820
rect 2944 9766 2946 9818
rect 3126 9766 3128 9818
rect 2882 9764 2888 9766
rect 2944 9764 2968 9766
rect 3024 9764 3048 9766
rect 3104 9764 3128 9766
rect 3184 9764 3190 9766
rect 2882 9755 3190 9764
rect 4814 9820 5122 9829
rect 4814 9818 4820 9820
rect 4876 9818 4900 9820
rect 4956 9818 4980 9820
rect 5036 9818 5060 9820
rect 5116 9818 5122 9820
rect 4876 9766 4878 9818
rect 5058 9766 5060 9818
rect 4814 9764 4820 9766
rect 4876 9764 4900 9766
rect 4956 9764 4980 9766
rect 5036 9764 5060 9766
rect 5116 9764 5122 9766
rect 4814 9755 5122 9764
rect 6746 9820 7054 9829
rect 6746 9818 6752 9820
rect 6808 9818 6832 9820
rect 6888 9818 6912 9820
rect 6968 9818 6992 9820
rect 7048 9818 7054 9820
rect 6808 9766 6810 9818
rect 6990 9766 6992 9818
rect 6746 9764 6752 9766
rect 6808 9764 6832 9766
rect 6888 9764 6912 9766
rect 6968 9764 6992 9766
rect 7048 9764 7054 9766
rect 6746 9755 7054 9764
rect 8678 9820 8986 9829
rect 8678 9818 8684 9820
rect 8740 9818 8764 9820
rect 8820 9818 8844 9820
rect 8900 9818 8924 9820
rect 8980 9818 8986 9820
rect 8740 9766 8742 9818
rect 8922 9766 8924 9818
rect 8678 9764 8684 9766
rect 8740 9764 8764 9766
rect 8820 9764 8844 9766
rect 8900 9764 8924 9766
rect 8980 9764 8986 9766
rect 8678 9755 8986 9764
rect 3848 9276 4156 9285
rect 3848 9274 3854 9276
rect 3910 9274 3934 9276
rect 3990 9274 4014 9276
rect 4070 9274 4094 9276
rect 4150 9274 4156 9276
rect 3910 9222 3912 9274
rect 4092 9222 4094 9274
rect 3848 9220 3854 9222
rect 3910 9220 3934 9222
rect 3990 9220 4014 9222
rect 4070 9220 4094 9222
rect 4150 9220 4156 9222
rect 3848 9211 4156 9220
rect 5780 9276 6088 9285
rect 5780 9274 5786 9276
rect 5842 9274 5866 9276
rect 5922 9274 5946 9276
rect 6002 9274 6026 9276
rect 6082 9274 6088 9276
rect 5842 9222 5844 9274
rect 6024 9222 6026 9274
rect 5780 9220 5786 9222
rect 5842 9220 5866 9222
rect 5922 9220 5946 9222
rect 6002 9220 6026 9222
rect 6082 9220 6088 9222
rect 5780 9211 6088 9220
rect 7712 9276 8020 9285
rect 7712 9274 7718 9276
rect 7774 9274 7798 9276
rect 7854 9274 7878 9276
rect 7934 9274 7958 9276
rect 8014 9274 8020 9276
rect 7774 9222 7776 9274
rect 7956 9222 7958 9274
rect 7712 9220 7718 9222
rect 7774 9220 7798 9222
rect 7854 9220 7878 9222
rect 7934 9220 7958 9222
rect 8014 9220 8020 9222
rect 7712 9211 8020 9220
rect 2882 8732 3190 8741
rect 2882 8730 2888 8732
rect 2944 8730 2968 8732
rect 3024 8730 3048 8732
rect 3104 8730 3128 8732
rect 3184 8730 3190 8732
rect 2944 8678 2946 8730
rect 3126 8678 3128 8730
rect 2882 8676 2888 8678
rect 2944 8676 2968 8678
rect 3024 8676 3048 8678
rect 3104 8676 3128 8678
rect 3184 8676 3190 8678
rect 2882 8667 3190 8676
rect 4814 8732 5122 8741
rect 4814 8730 4820 8732
rect 4876 8730 4900 8732
rect 4956 8730 4980 8732
rect 5036 8730 5060 8732
rect 5116 8730 5122 8732
rect 4876 8678 4878 8730
rect 5058 8678 5060 8730
rect 4814 8676 4820 8678
rect 4876 8676 4900 8678
rect 4956 8676 4980 8678
rect 5036 8676 5060 8678
rect 5116 8676 5122 8678
rect 4814 8667 5122 8676
rect 6746 8732 7054 8741
rect 6746 8730 6752 8732
rect 6808 8730 6832 8732
rect 6888 8730 6912 8732
rect 6968 8730 6992 8732
rect 7048 8730 7054 8732
rect 6808 8678 6810 8730
rect 6990 8678 6992 8730
rect 6746 8676 6752 8678
rect 6808 8676 6832 8678
rect 6888 8676 6912 8678
rect 6968 8676 6992 8678
rect 7048 8676 7054 8678
rect 6746 8667 7054 8676
rect 8678 8732 8986 8741
rect 8678 8730 8684 8732
rect 8740 8730 8764 8732
rect 8820 8730 8844 8732
rect 8900 8730 8924 8732
rect 8980 8730 8986 8732
rect 8740 8678 8742 8730
rect 8922 8678 8924 8730
rect 8678 8676 8684 8678
rect 8740 8676 8764 8678
rect 8820 8676 8844 8678
rect 8900 8676 8924 8678
rect 8980 8676 8986 8678
rect 8678 8667 8986 8676
rect 3848 8188 4156 8197
rect 3848 8186 3854 8188
rect 3910 8186 3934 8188
rect 3990 8186 4014 8188
rect 4070 8186 4094 8188
rect 4150 8186 4156 8188
rect 3910 8134 3912 8186
rect 4092 8134 4094 8186
rect 3848 8132 3854 8134
rect 3910 8132 3934 8134
rect 3990 8132 4014 8134
rect 4070 8132 4094 8134
rect 4150 8132 4156 8134
rect 3848 8123 4156 8132
rect 5780 8188 6088 8197
rect 5780 8186 5786 8188
rect 5842 8186 5866 8188
rect 5922 8186 5946 8188
rect 6002 8186 6026 8188
rect 6082 8186 6088 8188
rect 5842 8134 5844 8186
rect 6024 8134 6026 8186
rect 5780 8132 5786 8134
rect 5842 8132 5866 8134
rect 5922 8132 5946 8134
rect 6002 8132 6026 8134
rect 6082 8132 6088 8134
rect 5780 8123 6088 8132
rect 7712 8188 8020 8197
rect 7712 8186 7718 8188
rect 7774 8186 7798 8188
rect 7854 8186 7878 8188
rect 7934 8186 7958 8188
rect 8014 8186 8020 8188
rect 7774 8134 7776 8186
rect 7956 8134 7958 8186
rect 7712 8132 7718 8134
rect 7774 8132 7798 8134
rect 7854 8132 7878 8134
rect 7934 8132 7958 8134
rect 8014 8132 8020 8134
rect 7712 8123 8020 8132
rect 2882 7644 3190 7653
rect 2882 7642 2888 7644
rect 2944 7642 2968 7644
rect 3024 7642 3048 7644
rect 3104 7642 3128 7644
rect 3184 7642 3190 7644
rect 2944 7590 2946 7642
rect 3126 7590 3128 7642
rect 2882 7588 2888 7590
rect 2944 7588 2968 7590
rect 3024 7588 3048 7590
rect 3104 7588 3128 7590
rect 3184 7588 3190 7590
rect 2882 7579 3190 7588
rect 4814 7644 5122 7653
rect 4814 7642 4820 7644
rect 4876 7642 4900 7644
rect 4956 7642 4980 7644
rect 5036 7642 5060 7644
rect 5116 7642 5122 7644
rect 4876 7590 4878 7642
rect 5058 7590 5060 7642
rect 4814 7588 4820 7590
rect 4876 7588 4900 7590
rect 4956 7588 4980 7590
rect 5036 7588 5060 7590
rect 5116 7588 5122 7590
rect 4814 7579 5122 7588
rect 6746 7644 7054 7653
rect 6746 7642 6752 7644
rect 6808 7642 6832 7644
rect 6888 7642 6912 7644
rect 6968 7642 6992 7644
rect 7048 7642 7054 7644
rect 6808 7590 6810 7642
rect 6990 7590 6992 7642
rect 6746 7588 6752 7590
rect 6808 7588 6832 7590
rect 6888 7588 6912 7590
rect 6968 7588 6992 7590
rect 7048 7588 7054 7590
rect 6746 7579 7054 7588
rect 8678 7644 8986 7653
rect 8678 7642 8684 7644
rect 8740 7642 8764 7644
rect 8820 7642 8844 7644
rect 8900 7642 8924 7644
rect 8980 7642 8986 7644
rect 8740 7590 8742 7642
rect 8922 7590 8924 7642
rect 8678 7588 8684 7590
rect 8740 7588 8764 7590
rect 8820 7588 8844 7590
rect 8900 7588 8924 7590
rect 8980 7588 8986 7590
rect 8678 7579 8986 7588
rect 3848 7100 4156 7109
rect 3848 7098 3854 7100
rect 3910 7098 3934 7100
rect 3990 7098 4014 7100
rect 4070 7098 4094 7100
rect 4150 7098 4156 7100
rect 3910 7046 3912 7098
rect 4092 7046 4094 7098
rect 3848 7044 3854 7046
rect 3910 7044 3934 7046
rect 3990 7044 4014 7046
rect 4070 7044 4094 7046
rect 4150 7044 4156 7046
rect 3848 7035 4156 7044
rect 5780 7100 6088 7109
rect 5780 7098 5786 7100
rect 5842 7098 5866 7100
rect 5922 7098 5946 7100
rect 6002 7098 6026 7100
rect 6082 7098 6088 7100
rect 5842 7046 5844 7098
rect 6024 7046 6026 7098
rect 5780 7044 5786 7046
rect 5842 7044 5866 7046
rect 5922 7044 5946 7046
rect 6002 7044 6026 7046
rect 6082 7044 6088 7046
rect 5780 7035 6088 7044
rect 7712 7100 8020 7109
rect 7712 7098 7718 7100
rect 7774 7098 7798 7100
rect 7854 7098 7878 7100
rect 7934 7098 7958 7100
rect 8014 7098 8020 7100
rect 7774 7046 7776 7098
rect 7956 7046 7958 7098
rect 7712 7044 7718 7046
rect 7774 7044 7798 7046
rect 7854 7044 7878 7046
rect 7934 7044 7958 7046
rect 8014 7044 8020 7046
rect 7712 7035 8020 7044
rect 2780 6656 2832 6662
rect 2780 6598 2832 6604
rect 2882 6556 3190 6565
rect 2882 6554 2888 6556
rect 2944 6554 2968 6556
rect 3024 6554 3048 6556
rect 3104 6554 3128 6556
rect 3184 6554 3190 6556
rect 2944 6502 2946 6554
rect 3126 6502 3128 6554
rect 2882 6500 2888 6502
rect 2944 6500 2968 6502
rect 3024 6500 3048 6502
rect 3104 6500 3128 6502
rect 3184 6500 3190 6502
rect 2882 6491 3190 6500
rect 4814 6556 5122 6565
rect 4814 6554 4820 6556
rect 4876 6554 4900 6556
rect 4956 6554 4980 6556
rect 5036 6554 5060 6556
rect 5116 6554 5122 6556
rect 4876 6502 4878 6554
rect 5058 6502 5060 6554
rect 4814 6500 4820 6502
rect 4876 6500 4900 6502
rect 4956 6500 4980 6502
rect 5036 6500 5060 6502
rect 5116 6500 5122 6502
rect 4814 6491 5122 6500
rect 6746 6556 7054 6565
rect 6746 6554 6752 6556
rect 6808 6554 6832 6556
rect 6888 6554 6912 6556
rect 6968 6554 6992 6556
rect 7048 6554 7054 6556
rect 6808 6502 6810 6554
rect 6990 6502 6992 6554
rect 6746 6500 6752 6502
rect 6808 6500 6832 6502
rect 6888 6500 6912 6502
rect 6968 6500 6992 6502
rect 7048 6500 7054 6502
rect 6746 6491 7054 6500
rect 8678 6556 8986 6565
rect 8678 6554 8684 6556
rect 8740 6554 8764 6556
rect 8820 6554 8844 6556
rect 8900 6554 8924 6556
rect 8980 6554 8986 6556
rect 8740 6502 8742 6554
rect 8922 6502 8924 6554
rect 8678 6500 8684 6502
rect 8740 6500 8764 6502
rect 8820 6500 8844 6502
rect 8900 6500 8924 6502
rect 8980 6500 8986 6502
rect 8678 6491 8986 6500
rect 2412 6316 2464 6322
rect 2412 6258 2464 6264
rect 2504 6316 2556 6322
rect 2504 6258 2556 6264
rect 1780 6174 1900 6202
rect 1780 5914 1808 6174
rect 1916 6012 2224 6021
rect 1916 6010 1922 6012
rect 1978 6010 2002 6012
rect 2058 6010 2082 6012
rect 2138 6010 2162 6012
rect 2218 6010 2224 6012
rect 1978 5958 1980 6010
rect 2160 5958 2162 6010
rect 1916 5956 1922 5958
rect 1978 5956 2002 5958
rect 2058 5956 2082 5958
rect 2138 5956 2162 5958
rect 2218 5956 2224 5958
rect 1916 5947 2224 5956
rect 1676 5908 1728 5914
rect 1676 5850 1728 5856
rect 1768 5908 1820 5914
rect 1768 5850 1820 5856
rect 1952 5704 2004 5710
rect 1952 5646 2004 5652
rect 1964 5370 1992 5646
rect 1952 5364 2004 5370
rect 1952 5306 2004 5312
rect 1768 5228 1820 5234
rect 1768 5170 1820 5176
rect 1676 5160 1728 5166
rect 1676 5102 1728 5108
rect 1584 4820 1636 4826
rect 1584 4762 1636 4768
rect 938 4720 994 4729
rect 938 4655 994 4664
rect 952 4622 980 4655
rect 940 4616 992 4622
rect 940 4558 992 4564
rect 940 3528 992 3534
rect 940 3470 992 3476
rect 952 3369 980 3470
rect 938 3360 994 3369
rect 938 3295 994 3304
rect 1688 2650 1716 5102
rect 1780 3738 1808 5170
rect 1916 4924 2224 4933
rect 1916 4922 1922 4924
rect 1978 4922 2002 4924
rect 2058 4922 2082 4924
rect 2138 4922 2162 4924
rect 2218 4922 2224 4924
rect 1978 4870 1980 4922
rect 2160 4870 2162 4922
rect 1916 4868 1922 4870
rect 1978 4868 2002 4870
rect 2058 4868 2082 4870
rect 2138 4868 2162 4870
rect 2218 4868 2224 4870
rect 1916 4859 2224 4868
rect 1916 3836 2224 3845
rect 1916 3834 1922 3836
rect 1978 3834 2002 3836
rect 2058 3834 2082 3836
rect 2138 3834 2162 3836
rect 2218 3834 2224 3836
rect 1978 3782 1980 3834
rect 2160 3782 2162 3834
rect 1916 3780 1922 3782
rect 1978 3780 2002 3782
rect 2058 3780 2082 3782
rect 2138 3780 2162 3782
rect 2218 3780 2224 3782
rect 1916 3771 2224 3780
rect 1768 3732 1820 3738
rect 1768 3674 1820 3680
rect 1916 2748 2224 2757
rect 1916 2746 1922 2748
rect 1978 2746 2002 2748
rect 2058 2746 2082 2748
rect 2138 2746 2162 2748
rect 2218 2746 2224 2748
rect 1978 2694 1980 2746
rect 2160 2694 2162 2746
rect 1916 2692 1922 2694
rect 1978 2692 2002 2694
rect 2058 2692 2082 2694
rect 2138 2692 2162 2694
rect 2218 2692 2224 2694
rect 1916 2683 2224 2692
rect 2516 2650 2544 6258
rect 3848 6012 4156 6021
rect 3848 6010 3854 6012
rect 3910 6010 3934 6012
rect 3990 6010 4014 6012
rect 4070 6010 4094 6012
rect 4150 6010 4156 6012
rect 3910 5958 3912 6010
rect 4092 5958 4094 6010
rect 3848 5956 3854 5958
rect 3910 5956 3934 5958
rect 3990 5956 4014 5958
rect 4070 5956 4094 5958
rect 4150 5956 4156 5958
rect 3848 5947 4156 5956
rect 5780 6012 6088 6021
rect 5780 6010 5786 6012
rect 5842 6010 5866 6012
rect 5922 6010 5946 6012
rect 6002 6010 6026 6012
rect 6082 6010 6088 6012
rect 5842 5958 5844 6010
rect 6024 5958 6026 6010
rect 5780 5956 5786 5958
rect 5842 5956 5866 5958
rect 5922 5956 5946 5958
rect 6002 5956 6026 5958
rect 6082 5956 6088 5958
rect 5780 5947 6088 5956
rect 7712 6012 8020 6021
rect 7712 6010 7718 6012
rect 7774 6010 7798 6012
rect 7854 6010 7878 6012
rect 7934 6010 7958 6012
rect 8014 6010 8020 6012
rect 7774 5958 7776 6010
rect 7956 5958 7958 6010
rect 7712 5956 7718 5958
rect 7774 5956 7798 5958
rect 7854 5956 7878 5958
rect 7934 5956 7958 5958
rect 8014 5956 8020 5958
rect 7712 5947 8020 5956
rect 2882 5468 3190 5477
rect 2882 5466 2888 5468
rect 2944 5466 2968 5468
rect 3024 5466 3048 5468
rect 3104 5466 3128 5468
rect 3184 5466 3190 5468
rect 2944 5414 2946 5466
rect 3126 5414 3128 5466
rect 2882 5412 2888 5414
rect 2944 5412 2968 5414
rect 3024 5412 3048 5414
rect 3104 5412 3128 5414
rect 3184 5412 3190 5414
rect 2882 5403 3190 5412
rect 4814 5468 5122 5477
rect 4814 5466 4820 5468
rect 4876 5466 4900 5468
rect 4956 5466 4980 5468
rect 5036 5466 5060 5468
rect 5116 5466 5122 5468
rect 4876 5414 4878 5466
rect 5058 5414 5060 5466
rect 4814 5412 4820 5414
rect 4876 5412 4900 5414
rect 4956 5412 4980 5414
rect 5036 5412 5060 5414
rect 5116 5412 5122 5414
rect 4814 5403 5122 5412
rect 6746 5468 7054 5477
rect 6746 5466 6752 5468
rect 6808 5466 6832 5468
rect 6888 5466 6912 5468
rect 6968 5466 6992 5468
rect 7048 5466 7054 5468
rect 6808 5414 6810 5466
rect 6990 5414 6992 5466
rect 6746 5412 6752 5414
rect 6808 5412 6832 5414
rect 6888 5412 6912 5414
rect 6968 5412 6992 5414
rect 7048 5412 7054 5414
rect 6746 5403 7054 5412
rect 8678 5468 8986 5477
rect 8678 5466 8684 5468
rect 8740 5466 8764 5468
rect 8820 5466 8844 5468
rect 8900 5466 8924 5468
rect 8980 5466 8986 5468
rect 8740 5414 8742 5466
rect 8922 5414 8924 5466
rect 8678 5412 8684 5414
rect 8740 5412 8764 5414
rect 8820 5412 8844 5414
rect 8900 5412 8924 5414
rect 8980 5412 8986 5414
rect 8678 5403 8986 5412
rect 3848 4924 4156 4933
rect 3848 4922 3854 4924
rect 3910 4922 3934 4924
rect 3990 4922 4014 4924
rect 4070 4922 4094 4924
rect 4150 4922 4156 4924
rect 3910 4870 3912 4922
rect 4092 4870 4094 4922
rect 3848 4868 3854 4870
rect 3910 4868 3934 4870
rect 3990 4868 4014 4870
rect 4070 4868 4094 4870
rect 4150 4868 4156 4870
rect 3848 4859 4156 4868
rect 5780 4924 6088 4933
rect 5780 4922 5786 4924
rect 5842 4922 5866 4924
rect 5922 4922 5946 4924
rect 6002 4922 6026 4924
rect 6082 4922 6088 4924
rect 5842 4870 5844 4922
rect 6024 4870 6026 4922
rect 5780 4868 5786 4870
rect 5842 4868 5866 4870
rect 5922 4868 5946 4870
rect 6002 4868 6026 4870
rect 6082 4868 6088 4870
rect 5780 4859 6088 4868
rect 7712 4924 8020 4933
rect 7712 4922 7718 4924
rect 7774 4922 7798 4924
rect 7854 4922 7878 4924
rect 7934 4922 7958 4924
rect 8014 4922 8020 4924
rect 7774 4870 7776 4922
rect 7956 4870 7958 4922
rect 7712 4868 7718 4870
rect 7774 4868 7798 4870
rect 7854 4868 7878 4870
rect 7934 4868 7958 4870
rect 8014 4868 8020 4870
rect 7712 4859 8020 4868
rect 2882 4380 3190 4389
rect 2882 4378 2888 4380
rect 2944 4378 2968 4380
rect 3024 4378 3048 4380
rect 3104 4378 3128 4380
rect 3184 4378 3190 4380
rect 2944 4326 2946 4378
rect 3126 4326 3128 4378
rect 2882 4324 2888 4326
rect 2944 4324 2968 4326
rect 3024 4324 3048 4326
rect 3104 4324 3128 4326
rect 3184 4324 3190 4326
rect 2882 4315 3190 4324
rect 4814 4380 5122 4389
rect 4814 4378 4820 4380
rect 4876 4378 4900 4380
rect 4956 4378 4980 4380
rect 5036 4378 5060 4380
rect 5116 4378 5122 4380
rect 4876 4326 4878 4378
rect 5058 4326 5060 4378
rect 4814 4324 4820 4326
rect 4876 4324 4900 4326
rect 4956 4324 4980 4326
rect 5036 4324 5060 4326
rect 5116 4324 5122 4326
rect 4814 4315 5122 4324
rect 6746 4380 7054 4389
rect 6746 4378 6752 4380
rect 6808 4378 6832 4380
rect 6888 4378 6912 4380
rect 6968 4378 6992 4380
rect 7048 4378 7054 4380
rect 6808 4326 6810 4378
rect 6990 4326 6992 4378
rect 6746 4324 6752 4326
rect 6808 4324 6832 4326
rect 6888 4324 6912 4326
rect 6968 4324 6992 4326
rect 7048 4324 7054 4326
rect 6746 4315 7054 4324
rect 8678 4380 8986 4389
rect 8678 4378 8684 4380
rect 8740 4378 8764 4380
rect 8820 4378 8844 4380
rect 8900 4378 8924 4380
rect 8980 4378 8986 4380
rect 8740 4326 8742 4378
rect 8922 4326 8924 4378
rect 8678 4324 8684 4326
rect 8740 4324 8764 4326
rect 8820 4324 8844 4326
rect 8900 4324 8924 4326
rect 8980 4324 8986 4326
rect 8678 4315 8986 4324
rect 3848 3836 4156 3845
rect 3848 3834 3854 3836
rect 3910 3834 3934 3836
rect 3990 3834 4014 3836
rect 4070 3834 4094 3836
rect 4150 3834 4156 3836
rect 3910 3782 3912 3834
rect 4092 3782 4094 3834
rect 3848 3780 3854 3782
rect 3910 3780 3934 3782
rect 3990 3780 4014 3782
rect 4070 3780 4094 3782
rect 4150 3780 4156 3782
rect 3848 3771 4156 3780
rect 5780 3836 6088 3845
rect 5780 3834 5786 3836
rect 5842 3834 5866 3836
rect 5922 3834 5946 3836
rect 6002 3834 6026 3836
rect 6082 3834 6088 3836
rect 5842 3782 5844 3834
rect 6024 3782 6026 3834
rect 5780 3780 5786 3782
rect 5842 3780 5866 3782
rect 5922 3780 5946 3782
rect 6002 3780 6026 3782
rect 6082 3780 6088 3782
rect 5780 3771 6088 3780
rect 7712 3836 8020 3845
rect 7712 3834 7718 3836
rect 7774 3834 7798 3836
rect 7854 3834 7878 3836
rect 7934 3834 7958 3836
rect 8014 3834 8020 3836
rect 7774 3782 7776 3834
rect 7956 3782 7958 3834
rect 7712 3780 7718 3782
rect 7774 3780 7798 3782
rect 7854 3780 7878 3782
rect 7934 3780 7958 3782
rect 8014 3780 8020 3782
rect 7712 3771 8020 3780
rect 2882 3292 3190 3301
rect 2882 3290 2888 3292
rect 2944 3290 2968 3292
rect 3024 3290 3048 3292
rect 3104 3290 3128 3292
rect 3184 3290 3190 3292
rect 2944 3238 2946 3290
rect 3126 3238 3128 3290
rect 2882 3236 2888 3238
rect 2944 3236 2968 3238
rect 3024 3236 3048 3238
rect 3104 3236 3128 3238
rect 3184 3236 3190 3238
rect 2882 3227 3190 3236
rect 4814 3292 5122 3301
rect 4814 3290 4820 3292
rect 4876 3290 4900 3292
rect 4956 3290 4980 3292
rect 5036 3290 5060 3292
rect 5116 3290 5122 3292
rect 4876 3238 4878 3290
rect 5058 3238 5060 3290
rect 4814 3236 4820 3238
rect 4876 3236 4900 3238
rect 4956 3236 4980 3238
rect 5036 3236 5060 3238
rect 5116 3236 5122 3238
rect 4814 3227 5122 3236
rect 6746 3292 7054 3301
rect 6746 3290 6752 3292
rect 6808 3290 6832 3292
rect 6888 3290 6912 3292
rect 6968 3290 6992 3292
rect 7048 3290 7054 3292
rect 6808 3238 6810 3290
rect 6990 3238 6992 3290
rect 6746 3236 6752 3238
rect 6808 3236 6832 3238
rect 6888 3236 6912 3238
rect 6968 3236 6992 3238
rect 7048 3236 7054 3238
rect 6746 3227 7054 3236
rect 8678 3292 8986 3301
rect 8678 3290 8684 3292
rect 8740 3290 8764 3292
rect 8820 3290 8844 3292
rect 8900 3290 8924 3292
rect 8980 3290 8986 3292
rect 8740 3238 8742 3290
rect 8922 3238 8924 3290
rect 8678 3236 8684 3238
rect 8740 3236 8764 3238
rect 8820 3236 8844 3238
rect 8900 3236 8924 3238
rect 8980 3236 8986 3238
rect 8678 3227 8986 3236
rect 3848 2748 4156 2757
rect 3848 2746 3854 2748
rect 3910 2746 3934 2748
rect 3990 2746 4014 2748
rect 4070 2746 4094 2748
rect 4150 2746 4156 2748
rect 3910 2694 3912 2746
rect 4092 2694 4094 2746
rect 3848 2692 3854 2694
rect 3910 2692 3934 2694
rect 3990 2692 4014 2694
rect 4070 2692 4094 2694
rect 4150 2692 4156 2694
rect 3848 2683 4156 2692
rect 5780 2748 6088 2757
rect 5780 2746 5786 2748
rect 5842 2746 5866 2748
rect 5922 2746 5946 2748
rect 6002 2746 6026 2748
rect 6082 2746 6088 2748
rect 5842 2694 5844 2746
rect 6024 2694 6026 2746
rect 5780 2692 5786 2694
rect 5842 2692 5866 2694
rect 5922 2692 5946 2694
rect 6002 2692 6026 2694
rect 6082 2692 6088 2694
rect 5780 2683 6088 2692
rect 7712 2748 8020 2757
rect 7712 2746 7718 2748
rect 7774 2746 7798 2748
rect 7854 2746 7878 2748
rect 7934 2746 7958 2748
rect 8014 2746 8020 2748
rect 7774 2694 7776 2746
rect 7956 2694 7958 2746
rect 7712 2692 7718 2694
rect 7774 2692 7798 2694
rect 7854 2692 7878 2694
rect 7934 2692 7958 2694
rect 8014 2692 8020 2694
rect 7712 2683 8020 2692
rect 1676 2644 1728 2650
rect 1676 2586 1728 2592
rect 2504 2644 2556 2650
rect 2504 2586 2556 2592
rect 940 2440 992 2446
rect 940 2382 992 2388
rect 1676 2440 1728 2446
rect 1676 2382 1728 2388
rect 952 2009 980 2382
rect 938 2000 994 2009
rect 938 1935 994 1944
rect 1688 785 1716 2382
rect 2882 2204 3190 2213
rect 2882 2202 2888 2204
rect 2944 2202 2968 2204
rect 3024 2202 3048 2204
rect 3104 2202 3128 2204
rect 3184 2202 3190 2204
rect 2944 2150 2946 2202
rect 3126 2150 3128 2202
rect 2882 2148 2888 2150
rect 2944 2148 2968 2150
rect 3024 2148 3048 2150
rect 3104 2148 3128 2150
rect 3184 2148 3190 2150
rect 2882 2139 3190 2148
rect 4814 2204 5122 2213
rect 4814 2202 4820 2204
rect 4876 2202 4900 2204
rect 4956 2202 4980 2204
rect 5036 2202 5060 2204
rect 5116 2202 5122 2204
rect 4876 2150 4878 2202
rect 5058 2150 5060 2202
rect 4814 2148 4820 2150
rect 4876 2148 4900 2150
rect 4956 2148 4980 2150
rect 5036 2148 5060 2150
rect 5116 2148 5122 2150
rect 4814 2139 5122 2148
rect 6746 2204 7054 2213
rect 6746 2202 6752 2204
rect 6808 2202 6832 2204
rect 6888 2202 6912 2204
rect 6968 2202 6992 2204
rect 7048 2202 7054 2204
rect 6808 2150 6810 2202
rect 6990 2150 6992 2202
rect 6746 2148 6752 2150
rect 6808 2148 6832 2150
rect 6888 2148 6912 2150
rect 6968 2148 6992 2150
rect 7048 2148 7054 2150
rect 6746 2139 7054 2148
rect 8678 2204 8986 2213
rect 8678 2202 8684 2204
rect 8740 2202 8764 2204
rect 8820 2202 8844 2204
rect 8900 2202 8924 2204
rect 8980 2202 8986 2204
rect 8740 2150 8742 2202
rect 8922 2150 8924 2202
rect 8678 2148 8684 2150
rect 8740 2148 8764 2150
rect 8820 2148 8844 2150
rect 8900 2148 8924 2150
rect 8980 2148 8986 2150
rect 8678 2139 8986 2148
rect 1674 776 1730 785
rect 1674 711 1730 720
<< via2 >>
rect 1030 20984 1086 21040
rect 1122 19624 1178 19680
rect 2888 19610 2944 19612
rect 2968 19610 3024 19612
rect 3048 19610 3104 19612
rect 3128 19610 3184 19612
rect 2888 19558 2934 19610
rect 2934 19558 2944 19610
rect 2968 19558 2998 19610
rect 2998 19558 3010 19610
rect 3010 19558 3024 19610
rect 3048 19558 3062 19610
rect 3062 19558 3074 19610
rect 3074 19558 3104 19610
rect 3128 19558 3138 19610
rect 3138 19558 3184 19610
rect 2888 19556 2944 19558
rect 2968 19556 3024 19558
rect 3048 19556 3104 19558
rect 3128 19556 3184 19558
rect 938 18264 994 18320
rect 938 16904 994 16960
rect 938 15544 994 15600
rect 938 14184 994 14240
rect 1922 19066 1978 19068
rect 2002 19066 2058 19068
rect 2082 19066 2138 19068
rect 2162 19066 2218 19068
rect 1922 19014 1968 19066
rect 1968 19014 1978 19066
rect 2002 19014 2032 19066
rect 2032 19014 2044 19066
rect 2044 19014 2058 19066
rect 2082 19014 2096 19066
rect 2096 19014 2108 19066
rect 2108 19014 2138 19066
rect 2162 19014 2172 19066
rect 2172 19014 2218 19066
rect 1922 19012 1978 19014
rect 2002 19012 2058 19014
rect 2082 19012 2138 19014
rect 2162 19012 2218 19014
rect 1922 17978 1978 17980
rect 2002 17978 2058 17980
rect 2082 17978 2138 17980
rect 2162 17978 2218 17980
rect 1922 17926 1968 17978
rect 1968 17926 1978 17978
rect 2002 17926 2032 17978
rect 2032 17926 2044 17978
rect 2044 17926 2058 17978
rect 2082 17926 2096 17978
rect 2096 17926 2108 17978
rect 2108 17926 2138 17978
rect 2162 17926 2172 17978
rect 2172 17926 2218 17978
rect 1922 17924 1978 17926
rect 2002 17924 2058 17926
rect 2082 17924 2138 17926
rect 2162 17924 2218 17926
rect 1922 16890 1978 16892
rect 2002 16890 2058 16892
rect 2082 16890 2138 16892
rect 2162 16890 2218 16892
rect 1922 16838 1968 16890
rect 1968 16838 1978 16890
rect 2002 16838 2032 16890
rect 2032 16838 2044 16890
rect 2044 16838 2058 16890
rect 2082 16838 2096 16890
rect 2096 16838 2108 16890
rect 2108 16838 2138 16890
rect 2162 16838 2172 16890
rect 2172 16838 2218 16890
rect 1922 16836 1978 16838
rect 2002 16836 2058 16838
rect 2082 16836 2138 16838
rect 2162 16836 2218 16838
rect 1922 15802 1978 15804
rect 2002 15802 2058 15804
rect 2082 15802 2138 15804
rect 2162 15802 2218 15804
rect 1922 15750 1968 15802
rect 1968 15750 1978 15802
rect 2002 15750 2032 15802
rect 2032 15750 2044 15802
rect 2044 15750 2058 15802
rect 2082 15750 2096 15802
rect 2096 15750 2108 15802
rect 2108 15750 2138 15802
rect 2162 15750 2172 15802
rect 2172 15750 2218 15802
rect 1922 15748 1978 15750
rect 2002 15748 2058 15750
rect 2082 15748 2138 15750
rect 2162 15748 2218 15750
rect 938 12824 994 12880
rect 938 11464 994 11520
rect 938 10104 994 10160
rect 1922 14714 1978 14716
rect 2002 14714 2058 14716
rect 2082 14714 2138 14716
rect 2162 14714 2218 14716
rect 1922 14662 1968 14714
rect 1968 14662 1978 14714
rect 2002 14662 2032 14714
rect 2032 14662 2044 14714
rect 2044 14662 2058 14714
rect 2082 14662 2096 14714
rect 2096 14662 2108 14714
rect 2108 14662 2138 14714
rect 2162 14662 2172 14714
rect 2172 14662 2218 14714
rect 1922 14660 1978 14662
rect 2002 14660 2058 14662
rect 2082 14660 2138 14662
rect 2162 14660 2218 14662
rect 4820 19610 4876 19612
rect 4900 19610 4956 19612
rect 4980 19610 5036 19612
rect 5060 19610 5116 19612
rect 4820 19558 4866 19610
rect 4866 19558 4876 19610
rect 4900 19558 4930 19610
rect 4930 19558 4942 19610
rect 4942 19558 4956 19610
rect 4980 19558 4994 19610
rect 4994 19558 5006 19610
rect 5006 19558 5036 19610
rect 5060 19558 5070 19610
rect 5070 19558 5116 19610
rect 4820 19556 4876 19558
rect 4900 19556 4956 19558
rect 4980 19556 5036 19558
rect 5060 19556 5116 19558
rect 6752 19610 6808 19612
rect 6832 19610 6888 19612
rect 6912 19610 6968 19612
rect 6992 19610 7048 19612
rect 6752 19558 6798 19610
rect 6798 19558 6808 19610
rect 6832 19558 6862 19610
rect 6862 19558 6874 19610
rect 6874 19558 6888 19610
rect 6912 19558 6926 19610
rect 6926 19558 6938 19610
rect 6938 19558 6968 19610
rect 6992 19558 7002 19610
rect 7002 19558 7048 19610
rect 6752 19556 6808 19558
rect 6832 19556 6888 19558
rect 6912 19556 6968 19558
rect 6992 19556 7048 19558
rect 8684 19610 8740 19612
rect 8764 19610 8820 19612
rect 8844 19610 8900 19612
rect 8924 19610 8980 19612
rect 8684 19558 8730 19610
rect 8730 19558 8740 19610
rect 8764 19558 8794 19610
rect 8794 19558 8806 19610
rect 8806 19558 8820 19610
rect 8844 19558 8858 19610
rect 8858 19558 8870 19610
rect 8870 19558 8900 19610
rect 8924 19558 8934 19610
rect 8934 19558 8980 19610
rect 8684 19556 8740 19558
rect 8764 19556 8820 19558
rect 8844 19556 8900 19558
rect 8924 19556 8980 19558
rect 3854 19066 3910 19068
rect 3934 19066 3990 19068
rect 4014 19066 4070 19068
rect 4094 19066 4150 19068
rect 3854 19014 3900 19066
rect 3900 19014 3910 19066
rect 3934 19014 3964 19066
rect 3964 19014 3976 19066
rect 3976 19014 3990 19066
rect 4014 19014 4028 19066
rect 4028 19014 4040 19066
rect 4040 19014 4070 19066
rect 4094 19014 4104 19066
rect 4104 19014 4150 19066
rect 3854 19012 3910 19014
rect 3934 19012 3990 19014
rect 4014 19012 4070 19014
rect 4094 19012 4150 19014
rect 5786 19066 5842 19068
rect 5866 19066 5922 19068
rect 5946 19066 6002 19068
rect 6026 19066 6082 19068
rect 5786 19014 5832 19066
rect 5832 19014 5842 19066
rect 5866 19014 5896 19066
rect 5896 19014 5908 19066
rect 5908 19014 5922 19066
rect 5946 19014 5960 19066
rect 5960 19014 5972 19066
rect 5972 19014 6002 19066
rect 6026 19014 6036 19066
rect 6036 19014 6082 19066
rect 5786 19012 5842 19014
rect 5866 19012 5922 19014
rect 5946 19012 6002 19014
rect 6026 19012 6082 19014
rect 2888 18522 2944 18524
rect 2968 18522 3024 18524
rect 3048 18522 3104 18524
rect 3128 18522 3184 18524
rect 2888 18470 2934 18522
rect 2934 18470 2944 18522
rect 2968 18470 2998 18522
rect 2998 18470 3010 18522
rect 3010 18470 3024 18522
rect 3048 18470 3062 18522
rect 3062 18470 3074 18522
rect 3074 18470 3104 18522
rect 3128 18470 3138 18522
rect 3138 18470 3184 18522
rect 2888 18468 2944 18470
rect 2968 18468 3024 18470
rect 3048 18468 3104 18470
rect 3128 18468 3184 18470
rect 4820 18522 4876 18524
rect 4900 18522 4956 18524
rect 4980 18522 5036 18524
rect 5060 18522 5116 18524
rect 4820 18470 4866 18522
rect 4866 18470 4876 18522
rect 4900 18470 4930 18522
rect 4930 18470 4942 18522
rect 4942 18470 4956 18522
rect 4980 18470 4994 18522
rect 4994 18470 5006 18522
rect 5006 18470 5036 18522
rect 5060 18470 5070 18522
rect 5070 18470 5116 18522
rect 4820 18468 4876 18470
rect 4900 18468 4956 18470
rect 4980 18468 5036 18470
rect 5060 18468 5116 18470
rect 3854 17978 3910 17980
rect 3934 17978 3990 17980
rect 4014 17978 4070 17980
rect 4094 17978 4150 17980
rect 3854 17926 3900 17978
rect 3900 17926 3910 17978
rect 3934 17926 3964 17978
rect 3964 17926 3976 17978
rect 3976 17926 3990 17978
rect 4014 17926 4028 17978
rect 4028 17926 4040 17978
rect 4040 17926 4070 17978
rect 4094 17926 4104 17978
rect 4104 17926 4150 17978
rect 3854 17924 3910 17926
rect 3934 17924 3990 17926
rect 4014 17924 4070 17926
rect 4094 17924 4150 17926
rect 5786 17978 5842 17980
rect 5866 17978 5922 17980
rect 5946 17978 6002 17980
rect 6026 17978 6082 17980
rect 5786 17926 5832 17978
rect 5832 17926 5842 17978
rect 5866 17926 5896 17978
rect 5896 17926 5908 17978
rect 5908 17926 5922 17978
rect 5946 17926 5960 17978
rect 5960 17926 5972 17978
rect 5972 17926 6002 17978
rect 6026 17926 6036 17978
rect 6036 17926 6082 17978
rect 5786 17924 5842 17926
rect 5866 17924 5922 17926
rect 5946 17924 6002 17926
rect 6026 17924 6082 17926
rect 2888 17434 2944 17436
rect 2968 17434 3024 17436
rect 3048 17434 3104 17436
rect 3128 17434 3184 17436
rect 2888 17382 2934 17434
rect 2934 17382 2944 17434
rect 2968 17382 2998 17434
rect 2998 17382 3010 17434
rect 3010 17382 3024 17434
rect 3048 17382 3062 17434
rect 3062 17382 3074 17434
rect 3074 17382 3104 17434
rect 3128 17382 3138 17434
rect 3138 17382 3184 17434
rect 2888 17380 2944 17382
rect 2968 17380 3024 17382
rect 3048 17380 3104 17382
rect 3128 17380 3184 17382
rect 4820 17434 4876 17436
rect 4900 17434 4956 17436
rect 4980 17434 5036 17436
rect 5060 17434 5116 17436
rect 4820 17382 4866 17434
rect 4866 17382 4876 17434
rect 4900 17382 4930 17434
rect 4930 17382 4942 17434
rect 4942 17382 4956 17434
rect 4980 17382 4994 17434
rect 4994 17382 5006 17434
rect 5006 17382 5036 17434
rect 5060 17382 5070 17434
rect 5070 17382 5116 17434
rect 4820 17380 4876 17382
rect 4900 17380 4956 17382
rect 4980 17380 5036 17382
rect 5060 17380 5116 17382
rect 3854 16890 3910 16892
rect 3934 16890 3990 16892
rect 4014 16890 4070 16892
rect 4094 16890 4150 16892
rect 3854 16838 3900 16890
rect 3900 16838 3910 16890
rect 3934 16838 3964 16890
rect 3964 16838 3976 16890
rect 3976 16838 3990 16890
rect 4014 16838 4028 16890
rect 4028 16838 4040 16890
rect 4040 16838 4070 16890
rect 4094 16838 4104 16890
rect 4104 16838 4150 16890
rect 3854 16836 3910 16838
rect 3934 16836 3990 16838
rect 4014 16836 4070 16838
rect 4094 16836 4150 16838
rect 5786 16890 5842 16892
rect 5866 16890 5922 16892
rect 5946 16890 6002 16892
rect 6026 16890 6082 16892
rect 5786 16838 5832 16890
rect 5832 16838 5842 16890
rect 5866 16838 5896 16890
rect 5896 16838 5908 16890
rect 5908 16838 5922 16890
rect 5946 16838 5960 16890
rect 5960 16838 5972 16890
rect 5972 16838 6002 16890
rect 6026 16838 6036 16890
rect 6036 16838 6082 16890
rect 5786 16836 5842 16838
rect 5866 16836 5922 16838
rect 5946 16836 6002 16838
rect 6026 16836 6082 16838
rect 2888 16346 2944 16348
rect 2968 16346 3024 16348
rect 3048 16346 3104 16348
rect 3128 16346 3184 16348
rect 2888 16294 2934 16346
rect 2934 16294 2944 16346
rect 2968 16294 2998 16346
rect 2998 16294 3010 16346
rect 3010 16294 3024 16346
rect 3048 16294 3062 16346
rect 3062 16294 3074 16346
rect 3074 16294 3104 16346
rect 3128 16294 3138 16346
rect 3138 16294 3184 16346
rect 2888 16292 2944 16294
rect 2968 16292 3024 16294
rect 3048 16292 3104 16294
rect 3128 16292 3184 16294
rect 4820 16346 4876 16348
rect 4900 16346 4956 16348
rect 4980 16346 5036 16348
rect 5060 16346 5116 16348
rect 4820 16294 4866 16346
rect 4866 16294 4876 16346
rect 4900 16294 4930 16346
rect 4930 16294 4942 16346
rect 4942 16294 4956 16346
rect 4980 16294 4994 16346
rect 4994 16294 5006 16346
rect 5006 16294 5036 16346
rect 5060 16294 5070 16346
rect 5070 16294 5116 16346
rect 4820 16292 4876 16294
rect 4900 16292 4956 16294
rect 4980 16292 5036 16294
rect 5060 16292 5116 16294
rect 7718 19066 7774 19068
rect 7798 19066 7854 19068
rect 7878 19066 7934 19068
rect 7958 19066 8014 19068
rect 7718 19014 7764 19066
rect 7764 19014 7774 19066
rect 7798 19014 7828 19066
rect 7828 19014 7840 19066
rect 7840 19014 7854 19066
rect 7878 19014 7892 19066
rect 7892 19014 7904 19066
rect 7904 19014 7934 19066
rect 7958 19014 7968 19066
rect 7968 19014 8014 19066
rect 7718 19012 7774 19014
rect 7798 19012 7854 19014
rect 7878 19012 7934 19014
rect 7958 19012 8014 19014
rect 6752 18522 6808 18524
rect 6832 18522 6888 18524
rect 6912 18522 6968 18524
rect 6992 18522 7048 18524
rect 6752 18470 6798 18522
rect 6798 18470 6808 18522
rect 6832 18470 6862 18522
rect 6862 18470 6874 18522
rect 6874 18470 6888 18522
rect 6912 18470 6926 18522
rect 6926 18470 6938 18522
rect 6938 18470 6968 18522
rect 6992 18470 7002 18522
rect 7002 18470 7048 18522
rect 6752 18468 6808 18470
rect 6832 18468 6888 18470
rect 6912 18468 6968 18470
rect 6992 18468 7048 18470
rect 7718 17978 7774 17980
rect 7798 17978 7854 17980
rect 7878 17978 7934 17980
rect 7958 17978 8014 17980
rect 7718 17926 7764 17978
rect 7764 17926 7774 17978
rect 7798 17926 7828 17978
rect 7828 17926 7840 17978
rect 7840 17926 7854 17978
rect 7878 17926 7892 17978
rect 7892 17926 7904 17978
rect 7904 17926 7934 17978
rect 7958 17926 7968 17978
rect 7968 17926 8014 17978
rect 7718 17924 7774 17926
rect 7798 17924 7854 17926
rect 7878 17924 7934 17926
rect 7958 17924 8014 17926
rect 6752 17434 6808 17436
rect 6832 17434 6888 17436
rect 6912 17434 6968 17436
rect 6992 17434 7048 17436
rect 6752 17382 6798 17434
rect 6798 17382 6808 17434
rect 6832 17382 6862 17434
rect 6862 17382 6874 17434
rect 6874 17382 6888 17434
rect 6912 17382 6926 17434
rect 6926 17382 6938 17434
rect 6938 17382 6968 17434
rect 6992 17382 7002 17434
rect 7002 17382 7048 17434
rect 6752 17380 6808 17382
rect 6832 17380 6888 17382
rect 6912 17380 6968 17382
rect 6992 17380 7048 17382
rect 7718 16890 7774 16892
rect 7798 16890 7854 16892
rect 7878 16890 7934 16892
rect 7958 16890 8014 16892
rect 7718 16838 7764 16890
rect 7764 16838 7774 16890
rect 7798 16838 7828 16890
rect 7828 16838 7840 16890
rect 7840 16838 7854 16890
rect 7878 16838 7892 16890
rect 7892 16838 7904 16890
rect 7904 16838 7934 16890
rect 7958 16838 7968 16890
rect 7968 16838 8014 16890
rect 7718 16836 7774 16838
rect 7798 16836 7854 16838
rect 7878 16836 7934 16838
rect 7958 16836 8014 16838
rect 6752 16346 6808 16348
rect 6832 16346 6888 16348
rect 6912 16346 6968 16348
rect 6992 16346 7048 16348
rect 6752 16294 6798 16346
rect 6798 16294 6808 16346
rect 6832 16294 6862 16346
rect 6862 16294 6874 16346
rect 6874 16294 6888 16346
rect 6912 16294 6926 16346
rect 6926 16294 6938 16346
rect 6938 16294 6968 16346
rect 6992 16294 7002 16346
rect 7002 16294 7048 16346
rect 6752 16292 6808 16294
rect 6832 16292 6888 16294
rect 6912 16292 6968 16294
rect 6992 16292 7048 16294
rect 1922 13626 1978 13628
rect 2002 13626 2058 13628
rect 2082 13626 2138 13628
rect 2162 13626 2218 13628
rect 1922 13574 1968 13626
rect 1968 13574 1978 13626
rect 2002 13574 2032 13626
rect 2032 13574 2044 13626
rect 2044 13574 2058 13626
rect 2082 13574 2096 13626
rect 2096 13574 2108 13626
rect 2108 13574 2138 13626
rect 2162 13574 2172 13626
rect 2172 13574 2218 13626
rect 1922 13572 1978 13574
rect 2002 13572 2058 13574
rect 2082 13572 2138 13574
rect 2162 13572 2218 13574
rect 1922 12538 1978 12540
rect 2002 12538 2058 12540
rect 2082 12538 2138 12540
rect 2162 12538 2218 12540
rect 1922 12486 1968 12538
rect 1968 12486 1978 12538
rect 2002 12486 2032 12538
rect 2032 12486 2044 12538
rect 2044 12486 2058 12538
rect 2082 12486 2096 12538
rect 2096 12486 2108 12538
rect 2108 12486 2138 12538
rect 2162 12486 2172 12538
rect 2172 12486 2218 12538
rect 1922 12484 1978 12486
rect 2002 12484 2058 12486
rect 2082 12484 2138 12486
rect 2162 12484 2218 12486
rect 1922 11450 1978 11452
rect 2002 11450 2058 11452
rect 2082 11450 2138 11452
rect 2162 11450 2218 11452
rect 1922 11398 1968 11450
rect 1968 11398 1978 11450
rect 2002 11398 2032 11450
rect 2032 11398 2044 11450
rect 2044 11398 2058 11450
rect 2082 11398 2096 11450
rect 2096 11398 2108 11450
rect 2108 11398 2138 11450
rect 2162 11398 2172 11450
rect 2172 11398 2218 11450
rect 1922 11396 1978 11398
rect 2002 11396 2058 11398
rect 2082 11396 2138 11398
rect 2162 11396 2218 11398
rect 1922 10362 1978 10364
rect 2002 10362 2058 10364
rect 2082 10362 2138 10364
rect 2162 10362 2218 10364
rect 1922 10310 1968 10362
rect 1968 10310 1978 10362
rect 2002 10310 2032 10362
rect 2032 10310 2044 10362
rect 2044 10310 2058 10362
rect 2082 10310 2096 10362
rect 2096 10310 2108 10362
rect 2108 10310 2138 10362
rect 2162 10310 2172 10362
rect 2172 10310 2218 10362
rect 1922 10308 1978 10310
rect 2002 10308 2058 10310
rect 2082 10308 2138 10310
rect 2162 10308 2218 10310
rect 938 8744 994 8800
rect 3854 15802 3910 15804
rect 3934 15802 3990 15804
rect 4014 15802 4070 15804
rect 4094 15802 4150 15804
rect 3854 15750 3900 15802
rect 3900 15750 3910 15802
rect 3934 15750 3964 15802
rect 3964 15750 3976 15802
rect 3976 15750 3990 15802
rect 4014 15750 4028 15802
rect 4028 15750 4040 15802
rect 4040 15750 4070 15802
rect 4094 15750 4104 15802
rect 4104 15750 4150 15802
rect 3854 15748 3910 15750
rect 3934 15748 3990 15750
rect 4014 15748 4070 15750
rect 4094 15748 4150 15750
rect 5786 15802 5842 15804
rect 5866 15802 5922 15804
rect 5946 15802 6002 15804
rect 6026 15802 6082 15804
rect 5786 15750 5832 15802
rect 5832 15750 5842 15802
rect 5866 15750 5896 15802
rect 5896 15750 5908 15802
rect 5908 15750 5922 15802
rect 5946 15750 5960 15802
rect 5960 15750 5972 15802
rect 5972 15750 6002 15802
rect 6026 15750 6036 15802
rect 6036 15750 6082 15802
rect 5786 15748 5842 15750
rect 5866 15748 5922 15750
rect 5946 15748 6002 15750
rect 6026 15748 6082 15750
rect 7718 15802 7774 15804
rect 7798 15802 7854 15804
rect 7878 15802 7934 15804
rect 7958 15802 8014 15804
rect 7718 15750 7764 15802
rect 7764 15750 7774 15802
rect 7798 15750 7828 15802
rect 7828 15750 7840 15802
rect 7840 15750 7854 15802
rect 7878 15750 7892 15802
rect 7892 15750 7904 15802
rect 7904 15750 7934 15802
rect 7958 15750 7968 15802
rect 7968 15750 8014 15802
rect 7718 15748 7774 15750
rect 7798 15748 7854 15750
rect 7878 15748 7934 15750
rect 7958 15748 8014 15750
rect 2888 15258 2944 15260
rect 2968 15258 3024 15260
rect 3048 15258 3104 15260
rect 3128 15258 3184 15260
rect 2888 15206 2934 15258
rect 2934 15206 2944 15258
rect 2968 15206 2998 15258
rect 2998 15206 3010 15258
rect 3010 15206 3024 15258
rect 3048 15206 3062 15258
rect 3062 15206 3074 15258
rect 3074 15206 3104 15258
rect 3128 15206 3138 15258
rect 3138 15206 3184 15258
rect 2888 15204 2944 15206
rect 2968 15204 3024 15206
rect 3048 15204 3104 15206
rect 3128 15204 3184 15206
rect 4820 15258 4876 15260
rect 4900 15258 4956 15260
rect 4980 15258 5036 15260
rect 5060 15258 5116 15260
rect 4820 15206 4866 15258
rect 4866 15206 4876 15258
rect 4900 15206 4930 15258
rect 4930 15206 4942 15258
rect 4942 15206 4956 15258
rect 4980 15206 4994 15258
rect 4994 15206 5006 15258
rect 5006 15206 5036 15258
rect 5060 15206 5070 15258
rect 5070 15206 5116 15258
rect 4820 15204 4876 15206
rect 4900 15204 4956 15206
rect 4980 15204 5036 15206
rect 5060 15204 5116 15206
rect 6752 15258 6808 15260
rect 6832 15258 6888 15260
rect 6912 15258 6968 15260
rect 6992 15258 7048 15260
rect 6752 15206 6798 15258
rect 6798 15206 6808 15258
rect 6832 15206 6862 15258
rect 6862 15206 6874 15258
rect 6874 15206 6888 15258
rect 6912 15206 6926 15258
rect 6926 15206 6938 15258
rect 6938 15206 6968 15258
rect 6992 15206 7002 15258
rect 7002 15206 7048 15258
rect 6752 15204 6808 15206
rect 6832 15204 6888 15206
rect 6912 15204 6968 15206
rect 6992 15204 7048 15206
rect 3854 14714 3910 14716
rect 3934 14714 3990 14716
rect 4014 14714 4070 14716
rect 4094 14714 4150 14716
rect 3854 14662 3900 14714
rect 3900 14662 3910 14714
rect 3934 14662 3964 14714
rect 3964 14662 3976 14714
rect 3976 14662 3990 14714
rect 4014 14662 4028 14714
rect 4028 14662 4040 14714
rect 4040 14662 4070 14714
rect 4094 14662 4104 14714
rect 4104 14662 4150 14714
rect 3854 14660 3910 14662
rect 3934 14660 3990 14662
rect 4014 14660 4070 14662
rect 4094 14660 4150 14662
rect 5786 14714 5842 14716
rect 5866 14714 5922 14716
rect 5946 14714 6002 14716
rect 6026 14714 6082 14716
rect 5786 14662 5832 14714
rect 5832 14662 5842 14714
rect 5866 14662 5896 14714
rect 5896 14662 5908 14714
rect 5908 14662 5922 14714
rect 5946 14662 5960 14714
rect 5960 14662 5972 14714
rect 5972 14662 6002 14714
rect 6026 14662 6036 14714
rect 6036 14662 6082 14714
rect 5786 14660 5842 14662
rect 5866 14660 5922 14662
rect 5946 14660 6002 14662
rect 6026 14660 6082 14662
rect 7718 14714 7774 14716
rect 7798 14714 7854 14716
rect 7878 14714 7934 14716
rect 7958 14714 8014 14716
rect 7718 14662 7764 14714
rect 7764 14662 7774 14714
rect 7798 14662 7828 14714
rect 7828 14662 7840 14714
rect 7840 14662 7854 14714
rect 7878 14662 7892 14714
rect 7892 14662 7904 14714
rect 7904 14662 7934 14714
rect 7958 14662 7968 14714
rect 7968 14662 8014 14714
rect 7718 14660 7774 14662
rect 7798 14660 7854 14662
rect 7878 14660 7934 14662
rect 7958 14660 8014 14662
rect 2888 14170 2944 14172
rect 2968 14170 3024 14172
rect 3048 14170 3104 14172
rect 3128 14170 3184 14172
rect 2888 14118 2934 14170
rect 2934 14118 2944 14170
rect 2968 14118 2998 14170
rect 2998 14118 3010 14170
rect 3010 14118 3024 14170
rect 3048 14118 3062 14170
rect 3062 14118 3074 14170
rect 3074 14118 3104 14170
rect 3128 14118 3138 14170
rect 3138 14118 3184 14170
rect 2888 14116 2944 14118
rect 2968 14116 3024 14118
rect 3048 14116 3104 14118
rect 3128 14116 3184 14118
rect 4820 14170 4876 14172
rect 4900 14170 4956 14172
rect 4980 14170 5036 14172
rect 5060 14170 5116 14172
rect 4820 14118 4866 14170
rect 4866 14118 4876 14170
rect 4900 14118 4930 14170
rect 4930 14118 4942 14170
rect 4942 14118 4956 14170
rect 4980 14118 4994 14170
rect 4994 14118 5006 14170
rect 5006 14118 5036 14170
rect 5060 14118 5070 14170
rect 5070 14118 5116 14170
rect 4820 14116 4876 14118
rect 4900 14116 4956 14118
rect 4980 14116 5036 14118
rect 5060 14116 5116 14118
rect 6752 14170 6808 14172
rect 6832 14170 6888 14172
rect 6912 14170 6968 14172
rect 6992 14170 7048 14172
rect 6752 14118 6798 14170
rect 6798 14118 6808 14170
rect 6832 14118 6862 14170
rect 6862 14118 6874 14170
rect 6874 14118 6888 14170
rect 6912 14118 6926 14170
rect 6926 14118 6938 14170
rect 6938 14118 6968 14170
rect 6992 14118 7002 14170
rect 7002 14118 7048 14170
rect 6752 14116 6808 14118
rect 6832 14116 6888 14118
rect 6912 14116 6968 14118
rect 6992 14116 7048 14118
rect 3854 13626 3910 13628
rect 3934 13626 3990 13628
rect 4014 13626 4070 13628
rect 4094 13626 4150 13628
rect 3854 13574 3900 13626
rect 3900 13574 3910 13626
rect 3934 13574 3964 13626
rect 3964 13574 3976 13626
rect 3976 13574 3990 13626
rect 4014 13574 4028 13626
rect 4028 13574 4040 13626
rect 4040 13574 4070 13626
rect 4094 13574 4104 13626
rect 4104 13574 4150 13626
rect 3854 13572 3910 13574
rect 3934 13572 3990 13574
rect 4014 13572 4070 13574
rect 4094 13572 4150 13574
rect 5786 13626 5842 13628
rect 5866 13626 5922 13628
rect 5946 13626 6002 13628
rect 6026 13626 6082 13628
rect 5786 13574 5832 13626
rect 5832 13574 5842 13626
rect 5866 13574 5896 13626
rect 5896 13574 5908 13626
rect 5908 13574 5922 13626
rect 5946 13574 5960 13626
rect 5960 13574 5972 13626
rect 5972 13574 6002 13626
rect 6026 13574 6036 13626
rect 6036 13574 6082 13626
rect 5786 13572 5842 13574
rect 5866 13572 5922 13574
rect 5946 13572 6002 13574
rect 6026 13572 6082 13574
rect 7718 13626 7774 13628
rect 7798 13626 7854 13628
rect 7878 13626 7934 13628
rect 7958 13626 8014 13628
rect 7718 13574 7764 13626
rect 7764 13574 7774 13626
rect 7798 13574 7828 13626
rect 7828 13574 7840 13626
rect 7840 13574 7854 13626
rect 7878 13574 7892 13626
rect 7892 13574 7904 13626
rect 7904 13574 7934 13626
rect 7958 13574 7968 13626
rect 7968 13574 8014 13626
rect 7718 13572 7774 13574
rect 7798 13572 7854 13574
rect 7878 13572 7934 13574
rect 7958 13572 8014 13574
rect 2888 13082 2944 13084
rect 2968 13082 3024 13084
rect 3048 13082 3104 13084
rect 3128 13082 3184 13084
rect 2888 13030 2934 13082
rect 2934 13030 2944 13082
rect 2968 13030 2998 13082
rect 2998 13030 3010 13082
rect 3010 13030 3024 13082
rect 3048 13030 3062 13082
rect 3062 13030 3074 13082
rect 3074 13030 3104 13082
rect 3128 13030 3138 13082
rect 3138 13030 3184 13082
rect 2888 13028 2944 13030
rect 2968 13028 3024 13030
rect 3048 13028 3104 13030
rect 3128 13028 3184 13030
rect 4820 13082 4876 13084
rect 4900 13082 4956 13084
rect 4980 13082 5036 13084
rect 5060 13082 5116 13084
rect 4820 13030 4866 13082
rect 4866 13030 4876 13082
rect 4900 13030 4930 13082
rect 4930 13030 4942 13082
rect 4942 13030 4956 13082
rect 4980 13030 4994 13082
rect 4994 13030 5006 13082
rect 5006 13030 5036 13082
rect 5060 13030 5070 13082
rect 5070 13030 5116 13082
rect 4820 13028 4876 13030
rect 4900 13028 4956 13030
rect 4980 13028 5036 13030
rect 5060 13028 5116 13030
rect 6752 13082 6808 13084
rect 6832 13082 6888 13084
rect 6912 13082 6968 13084
rect 6992 13082 7048 13084
rect 6752 13030 6798 13082
rect 6798 13030 6808 13082
rect 6832 13030 6862 13082
rect 6862 13030 6874 13082
rect 6874 13030 6888 13082
rect 6912 13030 6926 13082
rect 6926 13030 6938 13082
rect 6938 13030 6968 13082
rect 6992 13030 7002 13082
rect 7002 13030 7048 13082
rect 6752 13028 6808 13030
rect 6832 13028 6888 13030
rect 6912 13028 6968 13030
rect 6992 13028 7048 13030
rect 3854 12538 3910 12540
rect 3934 12538 3990 12540
rect 4014 12538 4070 12540
rect 4094 12538 4150 12540
rect 3854 12486 3900 12538
rect 3900 12486 3910 12538
rect 3934 12486 3964 12538
rect 3964 12486 3976 12538
rect 3976 12486 3990 12538
rect 4014 12486 4028 12538
rect 4028 12486 4040 12538
rect 4040 12486 4070 12538
rect 4094 12486 4104 12538
rect 4104 12486 4150 12538
rect 3854 12484 3910 12486
rect 3934 12484 3990 12486
rect 4014 12484 4070 12486
rect 4094 12484 4150 12486
rect 5786 12538 5842 12540
rect 5866 12538 5922 12540
rect 5946 12538 6002 12540
rect 6026 12538 6082 12540
rect 5786 12486 5832 12538
rect 5832 12486 5842 12538
rect 5866 12486 5896 12538
rect 5896 12486 5908 12538
rect 5908 12486 5922 12538
rect 5946 12486 5960 12538
rect 5960 12486 5972 12538
rect 5972 12486 6002 12538
rect 6026 12486 6036 12538
rect 6036 12486 6082 12538
rect 5786 12484 5842 12486
rect 5866 12484 5922 12486
rect 5946 12484 6002 12486
rect 6026 12484 6082 12486
rect 7718 12538 7774 12540
rect 7798 12538 7854 12540
rect 7878 12538 7934 12540
rect 7958 12538 8014 12540
rect 7718 12486 7764 12538
rect 7764 12486 7774 12538
rect 7798 12486 7828 12538
rect 7828 12486 7840 12538
rect 7840 12486 7854 12538
rect 7878 12486 7892 12538
rect 7892 12486 7904 12538
rect 7904 12486 7934 12538
rect 7958 12486 7968 12538
rect 7968 12486 8014 12538
rect 7718 12484 7774 12486
rect 7798 12484 7854 12486
rect 7878 12484 7934 12486
rect 7958 12484 8014 12486
rect 8684 18522 8740 18524
rect 8764 18522 8820 18524
rect 8844 18522 8900 18524
rect 8924 18522 8980 18524
rect 8684 18470 8730 18522
rect 8730 18470 8740 18522
rect 8764 18470 8794 18522
rect 8794 18470 8806 18522
rect 8806 18470 8820 18522
rect 8844 18470 8858 18522
rect 8858 18470 8870 18522
rect 8870 18470 8900 18522
rect 8924 18470 8934 18522
rect 8934 18470 8980 18522
rect 8684 18468 8740 18470
rect 8764 18468 8820 18470
rect 8844 18468 8900 18470
rect 8924 18468 8980 18470
rect 8684 17434 8740 17436
rect 8764 17434 8820 17436
rect 8844 17434 8900 17436
rect 8924 17434 8980 17436
rect 8684 17382 8730 17434
rect 8730 17382 8740 17434
rect 8764 17382 8794 17434
rect 8794 17382 8806 17434
rect 8806 17382 8820 17434
rect 8844 17382 8858 17434
rect 8858 17382 8870 17434
rect 8870 17382 8900 17434
rect 8924 17382 8934 17434
rect 8934 17382 8980 17434
rect 8684 17380 8740 17382
rect 8764 17380 8820 17382
rect 8844 17380 8900 17382
rect 8924 17380 8980 17382
rect 8684 16346 8740 16348
rect 8764 16346 8820 16348
rect 8844 16346 8900 16348
rect 8924 16346 8980 16348
rect 8684 16294 8730 16346
rect 8730 16294 8740 16346
rect 8764 16294 8794 16346
rect 8794 16294 8806 16346
rect 8806 16294 8820 16346
rect 8844 16294 8858 16346
rect 8858 16294 8870 16346
rect 8870 16294 8900 16346
rect 8924 16294 8934 16346
rect 8934 16294 8980 16346
rect 8684 16292 8740 16294
rect 8764 16292 8820 16294
rect 8844 16292 8900 16294
rect 8924 16292 8980 16294
rect 8684 15258 8740 15260
rect 8764 15258 8820 15260
rect 8844 15258 8900 15260
rect 8924 15258 8980 15260
rect 8684 15206 8730 15258
rect 8730 15206 8740 15258
rect 8764 15206 8794 15258
rect 8794 15206 8806 15258
rect 8806 15206 8820 15258
rect 8844 15206 8858 15258
rect 8858 15206 8870 15258
rect 8870 15206 8900 15258
rect 8924 15206 8934 15258
rect 8934 15206 8980 15258
rect 8684 15204 8740 15206
rect 8764 15204 8820 15206
rect 8844 15204 8900 15206
rect 8924 15204 8980 15206
rect 8684 14170 8740 14172
rect 8764 14170 8820 14172
rect 8844 14170 8900 14172
rect 8924 14170 8980 14172
rect 8684 14118 8730 14170
rect 8730 14118 8740 14170
rect 8764 14118 8794 14170
rect 8794 14118 8806 14170
rect 8806 14118 8820 14170
rect 8844 14118 8858 14170
rect 8858 14118 8870 14170
rect 8870 14118 8900 14170
rect 8924 14118 8934 14170
rect 8934 14118 8980 14170
rect 8684 14116 8740 14118
rect 8764 14116 8820 14118
rect 8844 14116 8900 14118
rect 8924 14116 8980 14118
rect 8684 13082 8740 13084
rect 8764 13082 8820 13084
rect 8844 13082 8900 13084
rect 8924 13082 8980 13084
rect 8684 13030 8730 13082
rect 8730 13030 8740 13082
rect 8764 13030 8794 13082
rect 8794 13030 8806 13082
rect 8806 13030 8820 13082
rect 8844 13030 8858 13082
rect 8858 13030 8870 13082
rect 8870 13030 8900 13082
rect 8924 13030 8934 13082
rect 8934 13030 8980 13082
rect 8684 13028 8740 13030
rect 8764 13028 8820 13030
rect 8844 13028 8900 13030
rect 8924 13028 8980 13030
rect 2888 11994 2944 11996
rect 2968 11994 3024 11996
rect 3048 11994 3104 11996
rect 3128 11994 3184 11996
rect 2888 11942 2934 11994
rect 2934 11942 2944 11994
rect 2968 11942 2998 11994
rect 2998 11942 3010 11994
rect 3010 11942 3024 11994
rect 3048 11942 3062 11994
rect 3062 11942 3074 11994
rect 3074 11942 3104 11994
rect 3128 11942 3138 11994
rect 3138 11942 3184 11994
rect 2888 11940 2944 11942
rect 2968 11940 3024 11942
rect 3048 11940 3104 11942
rect 3128 11940 3184 11942
rect 4820 11994 4876 11996
rect 4900 11994 4956 11996
rect 4980 11994 5036 11996
rect 5060 11994 5116 11996
rect 4820 11942 4866 11994
rect 4866 11942 4876 11994
rect 4900 11942 4930 11994
rect 4930 11942 4942 11994
rect 4942 11942 4956 11994
rect 4980 11942 4994 11994
rect 4994 11942 5006 11994
rect 5006 11942 5036 11994
rect 5060 11942 5070 11994
rect 5070 11942 5116 11994
rect 4820 11940 4876 11942
rect 4900 11940 4956 11942
rect 4980 11940 5036 11942
rect 5060 11940 5116 11942
rect 6752 11994 6808 11996
rect 6832 11994 6888 11996
rect 6912 11994 6968 11996
rect 6992 11994 7048 11996
rect 6752 11942 6798 11994
rect 6798 11942 6808 11994
rect 6832 11942 6862 11994
rect 6862 11942 6874 11994
rect 6874 11942 6888 11994
rect 6912 11942 6926 11994
rect 6926 11942 6938 11994
rect 6938 11942 6968 11994
rect 6992 11942 7002 11994
rect 7002 11942 7048 11994
rect 6752 11940 6808 11942
rect 6832 11940 6888 11942
rect 6912 11940 6968 11942
rect 6992 11940 7048 11942
rect 8684 11994 8740 11996
rect 8764 11994 8820 11996
rect 8844 11994 8900 11996
rect 8924 11994 8980 11996
rect 8684 11942 8730 11994
rect 8730 11942 8740 11994
rect 8764 11942 8794 11994
rect 8794 11942 8806 11994
rect 8806 11942 8820 11994
rect 8844 11942 8858 11994
rect 8858 11942 8870 11994
rect 8870 11942 8900 11994
rect 8924 11942 8934 11994
rect 8934 11942 8980 11994
rect 8684 11940 8740 11942
rect 8764 11940 8820 11942
rect 8844 11940 8900 11942
rect 8924 11940 8980 11942
rect 3854 11450 3910 11452
rect 3934 11450 3990 11452
rect 4014 11450 4070 11452
rect 4094 11450 4150 11452
rect 3854 11398 3900 11450
rect 3900 11398 3910 11450
rect 3934 11398 3964 11450
rect 3964 11398 3976 11450
rect 3976 11398 3990 11450
rect 4014 11398 4028 11450
rect 4028 11398 4040 11450
rect 4040 11398 4070 11450
rect 4094 11398 4104 11450
rect 4104 11398 4150 11450
rect 3854 11396 3910 11398
rect 3934 11396 3990 11398
rect 4014 11396 4070 11398
rect 4094 11396 4150 11398
rect 5786 11450 5842 11452
rect 5866 11450 5922 11452
rect 5946 11450 6002 11452
rect 6026 11450 6082 11452
rect 5786 11398 5832 11450
rect 5832 11398 5842 11450
rect 5866 11398 5896 11450
rect 5896 11398 5908 11450
rect 5908 11398 5922 11450
rect 5946 11398 5960 11450
rect 5960 11398 5972 11450
rect 5972 11398 6002 11450
rect 6026 11398 6036 11450
rect 6036 11398 6082 11450
rect 5786 11396 5842 11398
rect 5866 11396 5922 11398
rect 5946 11396 6002 11398
rect 6026 11396 6082 11398
rect 7718 11450 7774 11452
rect 7798 11450 7854 11452
rect 7878 11450 7934 11452
rect 7958 11450 8014 11452
rect 7718 11398 7764 11450
rect 7764 11398 7774 11450
rect 7798 11398 7828 11450
rect 7828 11398 7840 11450
rect 7840 11398 7854 11450
rect 7878 11398 7892 11450
rect 7892 11398 7904 11450
rect 7904 11398 7934 11450
rect 7958 11398 7968 11450
rect 7968 11398 8014 11450
rect 7718 11396 7774 11398
rect 7798 11396 7854 11398
rect 7878 11396 7934 11398
rect 7958 11396 8014 11398
rect 1922 9274 1978 9276
rect 2002 9274 2058 9276
rect 2082 9274 2138 9276
rect 2162 9274 2218 9276
rect 1922 9222 1968 9274
rect 1968 9222 1978 9274
rect 2002 9222 2032 9274
rect 2032 9222 2044 9274
rect 2044 9222 2058 9274
rect 2082 9222 2096 9274
rect 2096 9222 2108 9274
rect 2108 9222 2138 9274
rect 2162 9222 2172 9274
rect 2172 9222 2218 9274
rect 1922 9220 1978 9222
rect 2002 9220 2058 9222
rect 2082 9220 2138 9222
rect 2162 9220 2218 9222
rect 938 7404 994 7440
rect 938 7384 940 7404
rect 940 7384 992 7404
rect 992 7384 994 7404
rect 938 6024 994 6080
rect 1922 8186 1978 8188
rect 2002 8186 2058 8188
rect 2082 8186 2138 8188
rect 2162 8186 2218 8188
rect 1922 8134 1968 8186
rect 1968 8134 1978 8186
rect 2002 8134 2032 8186
rect 2032 8134 2044 8186
rect 2044 8134 2058 8186
rect 2082 8134 2096 8186
rect 2096 8134 2108 8186
rect 2108 8134 2138 8186
rect 2162 8134 2172 8186
rect 2172 8134 2218 8186
rect 1922 8132 1978 8134
rect 2002 8132 2058 8134
rect 2082 8132 2138 8134
rect 2162 8132 2218 8134
rect 1922 7098 1978 7100
rect 2002 7098 2058 7100
rect 2082 7098 2138 7100
rect 2162 7098 2218 7100
rect 1922 7046 1968 7098
rect 1968 7046 1978 7098
rect 2002 7046 2032 7098
rect 2032 7046 2044 7098
rect 2044 7046 2058 7098
rect 2082 7046 2096 7098
rect 2096 7046 2108 7098
rect 2108 7046 2138 7098
rect 2162 7046 2172 7098
rect 2172 7046 2218 7098
rect 1922 7044 1978 7046
rect 2002 7044 2058 7046
rect 2082 7044 2138 7046
rect 2162 7044 2218 7046
rect 2888 10906 2944 10908
rect 2968 10906 3024 10908
rect 3048 10906 3104 10908
rect 3128 10906 3184 10908
rect 2888 10854 2934 10906
rect 2934 10854 2944 10906
rect 2968 10854 2998 10906
rect 2998 10854 3010 10906
rect 3010 10854 3024 10906
rect 3048 10854 3062 10906
rect 3062 10854 3074 10906
rect 3074 10854 3104 10906
rect 3128 10854 3138 10906
rect 3138 10854 3184 10906
rect 2888 10852 2944 10854
rect 2968 10852 3024 10854
rect 3048 10852 3104 10854
rect 3128 10852 3184 10854
rect 4820 10906 4876 10908
rect 4900 10906 4956 10908
rect 4980 10906 5036 10908
rect 5060 10906 5116 10908
rect 4820 10854 4866 10906
rect 4866 10854 4876 10906
rect 4900 10854 4930 10906
rect 4930 10854 4942 10906
rect 4942 10854 4956 10906
rect 4980 10854 4994 10906
rect 4994 10854 5006 10906
rect 5006 10854 5036 10906
rect 5060 10854 5070 10906
rect 5070 10854 5116 10906
rect 4820 10852 4876 10854
rect 4900 10852 4956 10854
rect 4980 10852 5036 10854
rect 5060 10852 5116 10854
rect 6752 10906 6808 10908
rect 6832 10906 6888 10908
rect 6912 10906 6968 10908
rect 6992 10906 7048 10908
rect 6752 10854 6798 10906
rect 6798 10854 6808 10906
rect 6832 10854 6862 10906
rect 6862 10854 6874 10906
rect 6874 10854 6888 10906
rect 6912 10854 6926 10906
rect 6926 10854 6938 10906
rect 6938 10854 6968 10906
rect 6992 10854 7002 10906
rect 7002 10854 7048 10906
rect 6752 10852 6808 10854
rect 6832 10852 6888 10854
rect 6912 10852 6968 10854
rect 6992 10852 7048 10854
rect 8684 10906 8740 10908
rect 8764 10906 8820 10908
rect 8844 10906 8900 10908
rect 8924 10906 8980 10908
rect 8684 10854 8730 10906
rect 8730 10854 8740 10906
rect 8764 10854 8794 10906
rect 8794 10854 8806 10906
rect 8806 10854 8820 10906
rect 8844 10854 8858 10906
rect 8858 10854 8870 10906
rect 8870 10854 8900 10906
rect 8924 10854 8934 10906
rect 8934 10854 8980 10906
rect 8684 10852 8740 10854
rect 8764 10852 8820 10854
rect 8844 10852 8900 10854
rect 8924 10852 8980 10854
rect 8206 10648 8262 10704
rect 3854 10362 3910 10364
rect 3934 10362 3990 10364
rect 4014 10362 4070 10364
rect 4094 10362 4150 10364
rect 3854 10310 3900 10362
rect 3900 10310 3910 10362
rect 3934 10310 3964 10362
rect 3964 10310 3976 10362
rect 3976 10310 3990 10362
rect 4014 10310 4028 10362
rect 4028 10310 4040 10362
rect 4040 10310 4070 10362
rect 4094 10310 4104 10362
rect 4104 10310 4150 10362
rect 3854 10308 3910 10310
rect 3934 10308 3990 10310
rect 4014 10308 4070 10310
rect 4094 10308 4150 10310
rect 5786 10362 5842 10364
rect 5866 10362 5922 10364
rect 5946 10362 6002 10364
rect 6026 10362 6082 10364
rect 5786 10310 5832 10362
rect 5832 10310 5842 10362
rect 5866 10310 5896 10362
rect 5896 10310 5908 10362
rect 5908 10310 5922 10362
rect 5946 10310 5960 10362
rect 5960 10310 5972 10362
rect 5972 10310 6002 10362
rect 6026 10310 6036 10362
rect 6036 10310 6082 10362
rect 5786 10308 5842 10310
rect 5866 10308 5922 10310
rect 5946 10308 6002 10310
rect 6026 10308 6082 10310
rect 7718 10362 7774 10364
rect 7798 10362 7854 10364
rect 7878 10362 7934 10364
rect 7958 10362 8014 10364
rect 7718 10310 7764 10362
rect 7764 10310 7774 10362
rect 7798 10310 7828 10362
rect 7828 10310 7840 10362
rect 7840 10310 7854 10362
rect 7878 10310 7892 10362
rect 7892 10310 7904 10362
rect 7904 10310 7934 10362
rect 7958 10310 7968 10362
rect 7968 10310 8014 10362
rect 7718 10308 7774 10310
rect 7798 10308 7854 10310
rect 7878 10308 7934 10310
rect 7958 10308 8014 10310
rect 2888 9818 2944 9820
rect 2968 9818 3024 9820
rect 3048 9818 3104 9820
rect 3128 9818 3184 9820
rect 2888 9766 2934 9818
rect 2934 9766 2944 9818
rect 2968 9766 2998 9818
rect 2998 9766 3010 9818
rect 3010 9766 3024 9818
rect 3048 9766 3062 9818
rect 3062 9766 3074 9818
rect 3074 9766 3104 9818
rect 3128 9766 3138 9818
rect 3138 9766 3184 9818
rect 2888 9764 2944 9766
rect 2968 9764 3024 9766
rect 3048 9764 3104 9766
rect 3128 9764 3184 9766
rect 4820 9818 4876 9820
rect 4900 9818 4956 9820
rect 4980 9818 5036 9820
rect 5060 9818 5116 9820
rect 4820 9766 4866 9818
rect 4866 9766 4876 9818
rect 4900 9766 4930 9818
rect 4930 9766 4942 9818
rect 4942 9766 4956 9818
rect 4980 9766 4994 9818
rect 4994 9766 5006 9818
rect 5006 9766 5036 9818
rect 5060 9766 5070 9818
rect 5070 9766 5116 9818
rect 4820 9764 4876 9766
rect 4900 9764 4956 9766
rect 4980 9764 5036 9766
rect 5060 9764 5116 9766
rect 6752 9818 6808 9820
rect 6832 9818 6888 9820
rect 6912 9818 6968 9820
rect 6992 9818 7048 9820
rect 6752 9766 6798 9818
rect 6798 9766 6808 9818
rect 6832 9766 6862 9818
rect 6862 9766 6874 9818
rect 6874 9766 6888 9818
rect 6912 9766 6926 9818
rect 6926 9766 6938 9818
rect 6938 9766 6968 9818
rect 6992 9766 7002 9818
rect 7002 9766 7048 9818
rect 6752 9764 6808 9766
rect 6832 9764 6888 9766
rect 6912 9764 6968 9766
rect 6992 9764 7048 9766
rect 8684 9818 8740 9820
rect 8764 9818 8820 9820
rect 8844 9818 8900 9820
rect 8924 9818 8980 9820
rect 8684 9766 8730 9818
rect 8730 9766 8740 9818
rect 8764 9766 8794 9818
rect 8794 9766 8806 9818
rect 8806 9766 8820 9818
rect 8844 9766 8858 9818
rect 8858 9766 8870 9818
rect 8870 9766 8900 9818
rect 8924 9766 8934 9818
rect 8934 9766 8980 9818
rect 8684 9764 8740 9766
rect 8764 9764 8820 9766
rect 8844 9764 8900 9766
rect 8924 9764 8980 9766
rect 3854 9274 3910 9276
rect 3934 9274 3990 9276
rect 4014 9274 4070 9276
rect 4094 9274 4150 9276
rect 3854 9222 3900 9274
rect 3900 9222 3910 9274
rect 3934 9222 3964 9274
rect 3964 9222 3976 9274
rect 3976 9222 3990 9274
rect 4014 9222 4028 9274
rect 4028 9222 4040 9274
rect 4040 9222 4070 9274
rect 4094 9222 4104 9274
rect 4104 9222 4150 9274
rect 3854 9220 3910 9222
rect 3934 9220 3990 9222
rect 4014 9220 4070 9222
rect 4094 9220 4150 9222
rect 5786 9274 5842 9276
rect 5866 9274 5922 9276
rect 5946 9274 6002 9276
rect 6026 9274 6082 9276
rect 5786 9222 5832 9274
rect 5832 9222 5842 9274
rect 5866 9222 5896 9274
rect 5896 9222 5908 9274
rect 5908 9222 5922 9274
rect 5946 9222 5960 9274
rect 5960 9222 5972 9274
rect 5972 9222 6002 9274
rect 6026 9222 6036 9274
rect 6036 9222 6082 9274
rect 5786 9220 5842 9222
rect 5866 9220 5922 9222
rect 5946 9220 6002 9222
rect 6026 9220 6082 9222
rect 7718 9274 7774 9276
rect 7798 9274 7854 9276
rect 7878 9274 7934 9276
rect 7958 9274 8014 9276
rect 7718 9222 7764 9274
rect 7764 9222 7774 9274
rect 7798 9222 7828 9274
rect 7828 9222 7840 9274
rect 7840 9222 7854 9274
rect 7878 9222 7892 9274
rect 7892 9222 7904 9274
rect 7904 9222 7934 9274
rect 7958 9222 7968 9274
rect 7968 9222 8014 9274
rect 7718 9220 7774 9222
rect 7798 9220 7854 9222
rect 7878 9220 7934 9222
rect 7958 9220 8014 9222
rect 2888 8730 2944 8732
rect 2968 8730 3024 8732
rect 3048 8730 3104 8732
rect 3128 8730 3184 8732
rect 2888 8678 2934 8730
rect 2934 8678 2944 8730
rect 2968 8678 2998 8730
rect 2998 8678 3010 8730
rect 3010 8678 3024 8730
rect 3048 8678 3062 8730
rect 3062 8678 3074 8730
rect 3074 8678 3104 8730
rect 3128 8678 3138 8730
rect 3138 8678 3184 8730
rect 2888 8676 2944 8678
rect 2968 8676 3024 8678
rect 3048 8676 3104 8678
rect 3128 8676 3184 8678
rect 4820 8730 4876 8732
rect 4900 8730 4956 8732
rect 4980 8730 5036 8732
rect 5060 8730 5116 8732
rect 4820 8678 4866 8730
rect 4866 8678 4876 8730
rect 4900 8678 4930 8730
rect 4930 8678 4942 8730
rect 4942 8678 4956 8730
rect 4980 8678 4994 8730
rect 4994 8678 5006 8730
rect 5006 8678 5036 8730
rect 5060 8678 5070 8730
rect 5070 8678 5116 8730
rect 4820 8676 4876 8678
rect 4900 8676 4956 8678
rect 4980 8676 5036 8678
rect 5060 8676 5116 8678
rect 6752 8730 6808 8732
rect 6832 8730 6888 8732
rect 6912 8730 6968 8732
rect 6992 8730 7048 8732
rect 6752 8678 6798 8730
rect 6798 8678 6808 8730
rect 6832 8678 6862 8730
rect 6862 8678 6874 8730
rect 6874 8678 6888 8730
rect 6912 8678 6926 8730
rect 6926 8678 6938 8730
rect 6938 8678 6968 8730
rect 6992 8678 7002 8730
rect 7002 8678 7048 8730
rect 6752 8676 6808 8678
rect 6832 8676 6888 8678
rect 6912 8676 6968 8678
rect 6992 8676 7048 8678
rect 8684 8730 8740 8732
rect 8764 8730 8820 8732
rect 8844 8730 8900 8732
rect 8924 8730 8980 8732
rect 8684 8678 8730 8730
rect 8730 8678 8740 8730
rect 8764 8678 8794 8730
rect 8794 8678 8806 8730
rect 8806 8678 8820 8730
rect 8844 8678 8858 8730
rect 8858 8678 8870 8730
rect 8870 8678 8900 8730
rect 8924 8678 8934 8730
rect 8934 8678 8980 8730
rect 8684 8676 8740 8678
rect 8764 8676 8820 8678
rect 8844 8676 8900 8678
rect 8924 8676 8980 8678
rect 3854 8186 3910 8188
rect 3934 8186 3990 8188
rect 4014 8186 4070 8188
rect 4094 8186 4150 8188
rect 3854 8134 3900 8186
rect 3900 8134 3910 8186
rect 3934 8134 3964 8186
rect 3964 8134 3976 8186
rect 3976 8134 3990 8186
rect 4014 8134 4028 8186
rect 4028 8134 4040 8186
rect 4040 8134 4070 8186
rect 4094 8134 4104 8186
rect 4104 8134 4150 8186
rect 3854 8132 3910 8134
rect 3934 8132 3990 8134
rect 4014 8132 4070 8134
rect 4094 8132 4150 8134
rect 5786 8186 5842 8188
rect 5866 8186 5922 8188
rect 5946 8186 6002 8188
rect 6026 8186 6082 8188
rect 5786 8134 5832 8186
rect 5832 8134 5842 8186
rect 5866 8134 5896 8186
rect 5896 8134 5908 8186
rect 5908 8134 5922 8186
rect 5946 8134 5960 8186
rect 5960 8134 5972 8186
rect 5972 8134 6002 8186
rect 6026 8134 6036 8186
rect 6036 8134 6082 8186
rect 5786 8132 5842 8134
rect 5866 8132 5922 8134
rect 5946 8132 6002 8134
rect 6026 8132 6082 8134
rect 7718 8186 7774 8188
rect 7798 8186 7854 8188
rect 7878 8186 7934 8188
rect 7958 8186 8014 8188
rect 7718 8134 7764 8186
rect 7764 8134 7774 8186
rect 7798 8134 7828 8186
rect 7828 8134 7840 8186
rect 7840 8134 7854 8186
rect 7878 8134 7892 8186
rect 7892 8134 7904 8186
rect 7904 8134 7934 8186
rect 7958 8134 7968 8186
rect 7968 8134 8014 8186
rect 7718 8132 7774 8134
rect 7798 8132 7854 8134
rect 7878 8132 7934 8134
rect 7958 8132 8014 8134
rect 2888 7642 2944 7644
rect 2968 7642 3024 7644
rect 3048 7642 3104 7644
rect 3128 7642 3184 7644
rect 2888 7590 2934 7642
rect 2934 7590 2944 7642
rect 2968 7590 2998 7642
rect 2998 7590 3010 7642
rect 3010 7590 3024 7642
rect 3048 7590 3062 7642
rect 3062 7590 3074 7642
rect 3074 7590 3104 7642
rect 3128 7590 3138 7642
rect 3138 7590 3184 7642
rect 2888 7588 2944 7590
rect 2968 7588 3024 7590
rect 3048 7588 3104 7590
rect 3128 7588 3184 7590
rect 4820 7642 4876 7644
rect 4900 7642 4956 7644
rect 4980 7642 5036 7644
rect 5060 7642 5116 7644
rect 4820 7590 4866 7642
rect 4866 7590 4876 7642
rect 4900 7590 4930 7642
rect 4930 7590 4942 7642
rect 4942 7590 4956 7642
rect 4980 7590 4994 7642
rect 4994 7590 5006 7642
rect 5006 7590 5036 7642
rect 5060 7590 5070 7642
rect 5070 7590 5116 7642
rect 4820 7588 4876 7590
rect 4900 7588 4956 7590
rect 4980 7588 5036 7590
rect 5060 7588 5116 7590
rect 6752 7642 6808 7644
rect 6832 7642 6888 7644
rect 6912 7642 6968 7644
rect 6992 7642 7048 7644
rect 6752 7590 6798 7642
rect 6798 7590 6808 7642
rect 6832 7590 6862 7642
rect 6862 7590 6874 7642
rect 6874 7590 6888 7642
rect 6912 7590 6926 7642
rect 6926 7590 6938 7642
rect 6938 7590 6968 7642
rect 6992 7590 7002 7642
rect 7002 7590 7048 7642
rect 6752 7588 6808 7590
rect 6832 7588 6888 7590
rect 6912 7588 6968 7590
rect 6992 7588 7048 7590
rect 8684 7642 8740 7644
rect 8764 7642 8820 7644
rect 8844 7642 8900 7644
rect 8924 7642 8980 7644
rect 8684 7590 8730 7642
rect 8730 7590 8740 7642
rect 8764 7590 8794 7642
rect 8794 7590 8806 7642
rect 8806 7590 8820 7642
rect 8844 7590 8858 7642
rect 8858 7590 8870 7642
rect 8870 7590 8900 7642
rect 8924 7590 8934 7642
rect 8934 7590 8980 7642
rect 8684 7588 8740 7590
rect 8764 7588 8820 7590
rect 8844 7588 8900 7590
rect 8924 7588 8980 7590
rect 3854 7098 3910 7100
rect 3934 7098 3990 7100
rect 4014 7098 4070 7100
rect 4094 7098 4150 7100
rect 3854 7046 3900 7098
rect 3900 7046 3910 7098
rect 3934 7046 3964 7098
rect 3964 7046 3976 7098
rect 3976 7046 3990 7098
rect 4014 7046 4028 7098
rect 4028 7046 4040 7098
rect 4040 7046 4070 7098
rect 4094 7046 4104 7098
rect 4104 7046 4150 7098
rect 3854 7044 3910 7046
rect 3934 7044 3990 7046
rect 4014 7044 4070 7046
rect 4094 7044 4150 7046
rect 5786 7098 5842 7100
rect 5866 7098 5922 7100
rect 5946 7098 6002 7100
rect 6026 7098 6082 7100
rect 5786 7046 5832 7098
rect 5832 7046 5842 7098
rect 5866 7046 5896 7098
rect 5896 7046 5908 7098
rect 5908 7046 5922 7098
rect 5946 7046 5960 7098
rect 5960 7046 5972 7098
rect 5972 7046 6002 7098
rect 6026 7046 6036 7098
rect 6036 7046 6082 7098
rect 5786 7044 5842 7046
rect 5866 7044 5922 7046
rect 5946 7044 6002 7046
rect 6026 7044 6082 7046
rect 7718 7098 7774 7100
rect 7798 7098 7854 7100
rect 7878 7098 7934 7100
rect 7958 7098 8014 7100
rect 7718 7046 7764 7098
rect 7764 7046 7774 7098
rect 7798 7046 7828 7098
rect 7828 7046 7840 7098
rect 7840 7046 7854 7098
rect 7878 7046 7892 7098
rect 7892 7046 7904 7098
rect 7904 7046 7934 7098
rect 7958 7046 7968 7098
rect 7968 7046 8014 7098
rect 7718 7044 7774 7046
rect 7798 7044 7854 7046
rect 7878 7044 7934 7046
rect 7958 7044 8014 7046
rect 2888 6554 2944 6556
rect 2968 6554 3024 6556
rect 3048 6554 3104 6556
rect 3128 6554 3184 6556
rect 2888 6502 2934 6554
rect 2934 6502 2944 6554
rect 2968 6502 2998 6554
rect 2998 6502 3010 6554
rect 3010 6502 3024 6554
rect 3048 6502 3062 6554
rect 3062 6502 3074 6554
rect 3074 6502 3104 6554
rect 3128 6502 3138 6554
rect 3138 6502 3184 6554
rect 2888 6500 2944 6502
rect 2968 6500 3024 6502
rect 3048 6500 3104 6502
rect 3128 6500 3184 6502
rect 4820 6554 4876 6556
rect 4900 6554 4956 6556
rect 4980 6554 5036 6556
rect 5060 6554 5116 6556
rect 4820 6502 4866 6554
rect 4866 6502 4876 6554
rect 4900 6502 4930 6554
rect 4930 6502 4942 6554
rect 4942 6502 4956 6554
rect 4980 6502 4994 6554
rect 4994 6502 5006 6554
rect 5006 6502 5036 6554
rect 5060 6502 5070 6554
rect 5070 6502 5116 6554
rect 4820 6500 4876 6502
rect 4900 6500 4956 6502
rect 4980 6500 5036 6502
rect 5060 6500 5116 6502
rect 6752 6554 6808 6556
rect 6832 6554 6888 6556
rect 6912 6554 6968 6556
rect 6992 6554 7048 6556
rect 6752 6502 6798 6554
rect 6798 6502 6808 6554
rect 6832 6502 6862 6554
rect 6862 6502 6874 6554
rect 6874 6502 6888 6554
rect 6912 6502 6926 6554
rect 6926 6502 6938 6554
rect 6938 6502 6968 6554
rect 6992 6502 7002 6554
rect 7002 6502 7048 6554
rect 6752 6500 6808 6502
rect 6832 6500 6888 6502
rect 6912 6500 6968 6502
rect 6992 6500 7048 6502
rect 8684 6554 8740 6556
rect 8764 6554 8820 6556
rect 8844 6554 8900 6556
rect 8924 6554 8980 6556
rect 8684 6502 8730 6554
rect 8730 6502 8740 6554
rect 8764 6502 8794 6554
rect 8794 6502 8806 6554
rect 8806 6502 8820 6554
rect 8844 6502 8858 6554
rect 8858 6502 8870 6554
rect 8870 6502 8900 6554
rect 8924 6502 8934 6554
rect 8934 6502 8980 6554
rect 8684 6500 8740 6502
rect 8764 6500 8820 6502
rect 8844 6500 8900 6502
rect 8924 6500 8980 6502
rect 1922 6010 1978 6012
rect 2002 6010 2058 6012
rect 2082 6010 2138 6012
rect 2162 6010 2218 6012
rect 1922 5958 1968 6010
rect 1968 5958 1978 6010
rect 2002 5958 2032 6010
rect 2032 5958 2044 6010
rect 2044 5958 2058 6010
rect 2082 5958 2096 6010
rect 2096 5958 2108 6010
rect 2108 5958 2138 6010
rect 2162 5958 2172 6010
rect 2172 5958 2218 6010
rect 1922 5956 1978 5958
rect 2002 5956 2058 5958
rect 2082 5956 2138 5958
rect 2162 5956 2218 5958
rect 938 4664 994 4720
rect 938 3304 994 3360
rect 1922 4922 1978 4924
rect 2002 4922 2058 4924
rect 2082 4922 2138 4924
rect 2162 4922 2218 4924
rect 1922 4870 1968 4922
rect 1968 4870 1978 4922
rect 2002 4870 2032 4922
rect 2032 4870 2044 4922
rect 2044 4870 2058 4922
rect 2082 4870 2096 4922
rect 2096 4870 2108 4922
rect 2108 4870 2138 4922
rect 2162 4870 2172 4922
rect 2172 4870 2218 4922
rect 1922 4868 1978 4870
rect 2002 4868 2058 4870
rect 2082 4868 2138 4870
rect 2162 4868 2218 4870
rect 1922 3834 1978 3836
rect 2002 3834 2058 3836
rect 2082 3834 2138 3836
rect 2162 3834 2218 3836
rect 1922 3782 1968 3834
rect 1968 3782 1978 3834
rect 2002 3782 2032 3834
rect 2032 3782 2044 3834
rect 2044 3782 2058 3834
rect 2082 3782 2096 3834
rect 2096 3782 2108 3834
rect 2108 3782 2138 3834
rect 2162 3782 2172 3834
rect 2172 3782 2218 3834
rect 1922 3780 1978 3782
rect 2002 3780 2058 3782
rect 2082 3780 2138 3782
rect 2162 3780 2218 3782
rect 1922 2746 1978 2748
rect 2002 2746 2058 2748
rect 2082 2746 2138 2748
rect 2162 2746 2218 2748
rect 1922 2694 1968 2746
rect 1968 2694 1978 2746
rect 2002 2694 2032 2746
rect 2032 2694 2044 2746
rect 2044 2694 2058 2746
rect 2082 2694 2096 2746
rect 2096 2694 2108 2746
rect 2108 2694 2138 2746
rect 2162 2694 2172 2746
rect 2172 2694 2218 2746
rect 1922 2692 1978 2694
rect 2002 2692 2058 2694
rect 2082 2692 2138 2694
rect 2162 2692 2218 2694
rect 3854 6010 3910 6012
rect 3934 6010 3990 6012
rect 4014 6010 4070 6012
rect 4094 6010 4150 6012
rect 3854 5958 3900 6010
rect 3900 5958 3910 6010
rect 3934 5958 3964 6010
rect 3964 5958 3976 6010
rect 3976 5958 3990 6010
rect 4014 5958 4028 6010
rect 4028 5958 4040 6010
rect 4040 5958 4070 6010
rect 4094 5958 4104 6010
rect 4104 5958 4150 6010
rect 3854 5956 3910 5958
rect 3934 5956 3990 5958
rect 4014 5956 4070 5958
rect 4094 5956 4150 5958
rect 5786 6010 5842 6012
rect 5866 6010 5922 6012
rect 5946 6010 6002 6012
rect 6026 6010 6082 6012
rect 5786 5958 5832 6010
rect 5832 5958 5842 6010
rect 5866 5958 5896 6010
rect 5896 5958 5908 6010
rect 5908 5958 5922 6010
rect 5946 5958 5960 6010
rect 5960 5958 5972 6010
rect 5972 5958 6002 6010
rect 6026 5958 6036 6010
rect 6036 5958 6082 6010
rect 5786 5956 5842 5958
rect 5866 5956 5922 5958
rect 5946 5956 6002 5958
rect 6026 5956 6082 5958
rect 7718 6010 7774 6012
rect 7798 6010 7854 6012
rect 7878 6010 7934 6012
rect 7958 6010 8014 6012
rect 7718 5958 7764 6010
rect 7764 5958 7774 6010
rect 7798 5958 7828 6010
rect 7828 5958 7840 6010
rect 7840 5958 7854 6010
rect 7878 5958 7892 6010
rect 7892 5958 7904 6010
rect 7904 5958 7934 6010
rect 7958 5958 7968 6010
rect 7968 5958 8014 6010
rect 7718 5956 7774 5958
rect 7798 5956 7854 5958
rect 7878 5956 7934 5958
rect 7958 5956 8014 5958
rect 2888 5466 2944 5468
rect 2968 5466 3024 5468
rect 3048 5466 3104 5468
rect 3128 5466 3184 5468
rect 2888 5414 2934 5466
rect 2934 5414 2944 5466
rect 2968 5414 2998 5466
rect 2998 5414 3010 5466
rect 3010 5414 3024 5466
rect 3048 5414 3062 5466
rect 3062 5414 3074 5466
rect 3074 5414 3104 5466
rect 3128 5414 3138 5466
rect 3138 5414 3184 5466
rect 2888 5412 2944 5414
rect 2968 5412 3024 5414
rect 3048 5412 3104 5414
rect 3128 5412 3184 5414
rect 4820 5466 4876 5468
rect 4900 5466 4956 5468
rect 4980 5466 5036 5468
rect 5060 5466 5116 5468
rect 4820 5414 4866 5466
rect 4866 5414 4876 5466
rect 4900 5414 4930 5466
rect 4930 5414 4942 5466
rect 4942 5414 4956 5466
rect 4980 5414 4994 5466
rect 4994 5414 5006 5466
rect 5006 5414 5036 5466
rect 5060 5414 5070 5466
rect 5070 5414 5116 5466
rect 4820 5412 4876 5414
rect 4900 5412 4956 5414
rect 4980 5412 5036 5414
rect 5060 5412 5116 5414
rect 6752 5466 6808 5468
rect 6832 5466 6888 5468
rect 6912 5466 6968 5468
rect 6992 5466 7048 5468
rect 6752 5414 6798 5466
rect 6798 5414 6808 5466
rect 6832 5414 6862 5466
rect 6862 5414 6874 5466
rect 6874 5414 6888 5466
rect 6912 5414 6926 5466
rect 6926 5414 6938 5466
rect 6938 5414 6968 5466
rect 6992 5414 7002 5466
rect 7002 5414 7048 5466
rect 6752 5412 6808 5414
rect 6832 5412 6888 5414
rect 6912 5412 6968 5414
rect 6992 5412 7048 5414
rect 8684 5466 8740 5468
rect 8764 5466 8820 5468
rect 8844 5466 8900 5468
rect 8924 5466 8980 5468
rect 8684 5414 8730 5466
rect 8730 5414 8740 5466
rect 8764 5414 8794 5466
rect 8794 5414 8806 5466
rect 8806 5414 8820 5466
rect 8844 5414 8858 5466
rect 8858 5414 8870 5466
rect 8870 5414 8900 5466
rect 8924 5414 8934 5466
rect 8934 5414 8980 5466
rect 8684 5412 8740 5414
rect 8764 5412 8820 5414
rect 8844 5412 8900 5414
rect 8924 5412 8980 5414
rect 3854 4922 3910 4924
rect 3934 4922 3990 4924
rect 4014 4922 4070 4924
rect 4094 4922 4150 4924
rect 3854 4870 3900 4922
rect 3900 4870 3910 4922
rect 3934 4870 3964 4922
rect 3964 4870 3976 4922
rect 3976 4870 3990 4922
rect 4014 4870 4028 4922
rect 4028 4870 4040 4922
rect 4040 4870 4070 4922
rect 4094 4870 4104 4922
rect 4104 4870 4150 4922
rect 3854 4868 3910 4870
rect 3934 4868 3990 4870
rect 4014 4868 4070 4870
rect 4094 4868 4150 4870
rect 5786 4922 5842 4924
rect 5866 4922 5922 4924
rect 5946 4922 6002 4924
rect 6026 4922 6082 4924
rect 5786 4870 5832 4922
rect 5832 4870 5842 4922
rect 5866 4870 5896 4922
rect 5896 4870 5908 4922
rect 5908 4870 5922 4922
rect 5946 4870 5960 4922
rect 5960 4870 5972 4922
rect 5972 4870 6002 4922
rect 6026 4870 6036 4922
rect 6036 4870 6082 4922
rect 5786 4868 5842 4870
rect 5866 4868 5922 4870
rect 5946 4868 6002 4870
rect 6026 4868 6082 4870
rect 7718 4922 7774 4924
rect 7798 4922 7854 4924
rect 7878 4922 7934 4924
rect 7958 4922 8014 4924
rect 7718 4870 7764 4922
rect 7764 4870 7774 4922
rect 7798 4870 7828 4922
rect 7828 4870 7840 4922
rect 7840 4870 7854 4922
rect 7878 4870 7892 4922
rect 7892 4870 7904 4922
rect 7904 4870 7934 4922
rect 7958 4870 7968 4922
rect 7968 4870 8014 4922
rect 7718 4868 7774 4870
rect 7798 4868 7854 4870
rect 7878 4868 7934 4870
rect 7958 4868 8014 4870
rect 2888 4378 2944 4380
rect 2968 4378 3024 4380
rect 3048 4378 3104 4380
rect 3128 4378 3184 4380
rect 2888 4326 2934 4378
rect 2934 4326 2944 4378
rect 2968 4326 2998 4378
rect 2998 4326 3010 4378
rect 3010 4326 3024 4378
rect 3048 4326 3062 4378
rect 3062 4326 3074 4378
rect 3074 4326 3104 4378
rect 3128 4326 3138 4378
rect 3138 4326 3184 4378
rect 2888 4324 2944 4326
rect 2968 4324 3024 4326
rect 3048 4324 3104 4326
rect 3128 4324 3184 4326
rect 4820 4378 4876 4380
rect 4900 4378 4956 4380
rect 4980 4378 5036 4380
rect 5060 4378 5116 4380
rect 4820 4326 4866 4378
rect 4866 4326 4876 4378
rect 4900 4326 4930 4378
rect 4930 4326 4942 4378
rect 4942 4326 4956 4378
rect 4980 4326 4994 4378
rect 4994 4326 5006 4378
rect 5006 4326 5036 4378
rect 5060 4326 5070 4378
rect 5070 4326 5116 4378
rect 4820 4324 4876 4326
rect 4900 4324 4956 4326
rect 4980 4324 5036 4326
rect 5060 4324 5116 4326
rect 6752 4378 6808 4380
rect 6832 4378 6888 4380
rect 6912 4378 6968 4380
rect 6992 4378 7048 4380
rect 6752 4326 6798 4378
rect 6798 4326 6808 4378
rect 6832 4326 6862 4378
rect 6862 4326 6874 4378
rect 6874 4326 6888 4378
rect 6912 4326 6926 4378
rect 6926 4326 6938 4378
rect 6938 4326 6968 4378
rect 6992 4326 7002 4378
rect 7002 4326 7048 4378
rect 6752 4324 6808 4326
rect 6832 4324 6888 4326
rect 6912 4324 6968 4326
rect 6992 4324 7048 4326
rect 8684 4378 8740 4380
rect 8764 4378 8820 4380
rect 8844 4378 8900 4380
rect 8924 4378 8980 4380
rect 8684 4326 8730 4378
rect 8730 4326 8740 4378
rect 8764 4326 8794 4378
rect 8794 4326 8806 4378
rect 8806 4326 8820 4378
rect 8844 4326 8858 4378
rect 8858 4326 8870 4378
rect 8870 4326 8900 4378
rect 8924 4326 8934 4378
rect 8934 4326 8980 4378
rect 8684 4324 8740 4326
rect 8764 4324 8820 4326
rect 8844 4324 8900 4326
rect 8924 4324 8980 4326
rect 3854 3834 3910 3836
rect 3934 3834 3990 3836
rect 4014 3834 4070 3836
rect 4094 3834 4150 3836
rect 3854 3782 3900 3834
rect 3900 3782 3910 3834
rect 3934 3782 3964 3834
rect 3964 3782 3976 3834
rect 3976 3782 3990 3834
rect 4014 3782 4028 3834
rect 4028 3782 4040 3834
rect 4040 3782 4070 3834
rect 4094 3782 4104 3834
rect 4104 3782 4150 3834
rect 3854 3780 3910 3782
rect 3934 3780 3990 3782
rect 4014 3780 4070 3782
rect 4094 3780 4150 3782
rect 5786 3834 5842 3836
rect 5866 3834 5922 3836
rect 5946 3834 6002 3836
rect 6026 3834 6082 3836
rect 5786 3782 5832 3834
rect 5832 3782 5842 3834
rect 5866 3782 5896 3834
rect 5896 3782 5908 3834
rect 5908 3782 5922 3834
rect 5946 3782 5960 3834
rect 5960 3782 5972 3834
rect 5972 3782 6002 3834
rect 6026 3782 6036 3834
rect 6036 3782 6082 3834
rect 5786 3780 5842 3782
rect 5866 3780 5922 3782
rect 5946 3780 6002 3782
rect 6026 3780 6082 3782
rect 7718 3834 7774 3836
rect 7798 3834 7854 3836
rect 7878 3834 7934 3836
rect 7958 3834 8014 3836
rect 7718 3782 7764 3834
rect 7764 3782 7774 3834
rect 7798 3782 7828 3834
rect 7828 3782 7840 3834
rect 7840 3782 7854 3834
rect 7878 3782 7892 3834
rect 7892 3782 7904 3834
rect 7904 3782 7934 3834
rect 7958 3782 7968 3834
rect 7968 3782 8014 3834
rect 7718 3780 7774 3782
rect 7798 3780 7854 3782
rect 7878 3780 7934 3782
rect 7958 3780 8014 3782
rect 2888 3290 2944 3292
rect 2968 3290 3024 3292
rect 3048 3290 3104 3292
rect 3128 3290 3184 3292
rect 2888 3238 2934 3290
rect 2934 3238 2944 3290
rect 2968 3238 2998 3290
rect 2998 3238 3010 3290
rect 3010 3238 3024 3290
rect 3048 3238 3062 3290
rect 3062 3238 3074 3290
rect 3074 3238 3104 3290
rect 3128 3238 3138 3290
rect 3138 3238 3184 3290
rect 2888 3236 2944 3238
rect 2968 3236 3024 3238
rect 3048 3236 3104 3238
rect 3128 3236 3184 3238
rect 4820 3290 4876 3292
rect 4900 3290 4956 3292
rect 4980 3290 5036 3292
rect 5060 3290 5116 3292
rect 4820 3238 4866 3290
rect 4866 3238 4876 3290
rect 4900 3238 4930 3290
rect 4930 3238 4942 3290
rect 4942 3238 4956 3290
rect 4980 3238 4994 3290
rect 4994 3238 5006 3290
rect 5006 3238 5036 3290
rect 5060 3238 5070 3290
rect 5070 3238 5116 3290
rect 4820 3236 4876 3238
rect 4900 3236 4956 3238
rect 4980 3236 5036 3238
rect 5060 3236 5116 3238
rect 6752 3290 6808 3292
rect 6832 3290 6888 3292
rect 6912 3290 6968 3292
rect 6992 3290 7048 3292
rect 6752 3238 6798 3290
rect 6798 3238 6808 3290
rect 6832 3238 6862 3290
rect 6862 3238 6874 3290
rect 6874 3238 6888 3290
rect 6912 3238 6926 3290
rect 6926 3238 6938 3290
rect 6938 3238 6968 3290
rect 6992 3238 7002 3290
rect 7002 3238 7048 3290
rect 6752 3236 6808 3238
rect 6832 3236 6888 3238
rect 6912 3236 6968 3238
rect 6992 3236 7048 3238
rect 8684 3290 8740 3292
rect 8764 3290 8820 3292
rect 8844 3290 8900 3292
rect 8924 3290 8980 3292
rect 8684 3238 8730 3290
rect 8730 3238 8740 3290
rect 8764 3238 8794 3290
rect 8794 3238 8806 3290
rect 8806 3238 8820 3290
rect 8844 3238 8858 3290
rect 8858 3238 8870 3290
rect 8870 3238 8900 3290
rect 8924 3238 8934 3290
rect 8934 3238 8980 3290
rect 8684 3236 8740 3238
rect 8764 3236 8820 3238
rect 8844 3236 8900 3238
rect 8924 3236 8980 3238
rect 3854 2746 3910 2748
rect 3934 2746 3990 2748
rect 4014 2746 4070 2748
rect 4094 2746 4150 2748
rect 3854 2694 3900 2746
rect 3900 2694 3910 2746
rect 3934 2694 3964 2746
rect 3964 2694 3976 2746
rect 3976 2694 3990 2746
rect 4014 2694 4028 2746
rect 4028 2694 4040 2746
rect 4040 2694 4070 2746
rect 4094 2694 4104 2746
rect 4104 2694 4150 2746
rect 3854 2692 3910 2694
rect 3934 2692 3990 2694
rect 4014 2692 4070 2694
rect 4094 2692 4150 2694
rect 5786 2746 5842 2748
rect 5866 2746 5922 2748
rect 5946 2746 6002 2748
rect 6026 2746 6082 2748
rect 5786 2694 5832 2746
rect 5832 2694 5842 2746
rect 5866 2694 5896 2746
rect 5896 2694 5908 2746
rect 5908 2694 5922 2746
rect 5946 2694 5960 2746
rect 5960 2694 5972 2746
rect 5972 2694 6002 2746
rect 6026 2694 6036 2746
rect 6036 2694 6082 2746
rect 5786 2692 5842 2694
rect 5866 2692 5922 2694
rect 5946 2692 6002 2694
rect 6026 2692 6082 2694
rect 7718 2746 7774 2748
rect 7798 2746 7854 2748
rect 7878 2746 7934 2748
rect 7958 2746 8014 2748
rect 7718 2694 7764 2746
rect 7764 2694 7774 2746
rect 7798 2694 7828 2746
rect 7828 2694 7840 2746
rect 7840 2694 7854 2746
rect 7878 2694 7892 2746
rect 7892 2694 7904 2746
rect 7904 2694 7934 2746
rect 7958 2694 7968 2746
rect 7968 2694 8014 2746
rect 7718 2692 7774 2694
rect 7798 2692 7854 2694
rect 7878 2692 7934 2694
rect 7958 2692 8014 2694
rect 938 1944 994 2000
rect 2888 2202 2944 2204
rect 2968 2202 3024 2204
rect 3048 2202 3104 2204
rect 3128 2202 3184 2204
rect 2888 2150 2934 2202
rect 2934 2150 2944 2202
rect 2968 2150 2998 2202
rect 2998 2150 3010 2202
rect 3010 2150 3024 2202
rect 3048 2150 3062 2202
rect 3062 2150 3074 2202
rect 3074 2150 3104 2202
rect 3128 2150 3138 2202
rect 3138 2150 3184 2202
rect 2888 2148 2944 2150
rect 2968 2148 3024 2150
rect 3048 2148 3104 2150
rect 3128 2148 3184 2150
rect 4820 2202 4876 2204
rect 4900 2202 4956 2204
rect 4980 2202 5036 2204
rect 5060 2202 5116 2204
rect 4820 2150 4866 2202
rect 4866 2150 4876 2202
rect 4900 2150 4930 2202
rect 4930 2150 4942 2202
rect 4942 2150 4956 2202
rect 4980 2150 4994 2202
rect 4994 2150 5006 2202
rect 5006 2150 5036 2202
rect 5060 2150 5070 2202
rect 5070 2150 5116 2202
rect 4820 2148 4876 2150
rect 4900 2148 4956 2150
rect 4980 2148 5036 2150
rect 5060 2148 5116 2150
rect 6752 2202 6808 2204
rect 6832 2202 6888 2204
rect 6912 2202 6968 2204
rect 6992 2202 7048 2204
rect 6752 2150 6798 2202
rect 6798 2150 6808 2202
rect 6832 2150 6862 2202
rect 6862 2150 6874 2202
rect 6874 2150 6888 2202
rect 6912 2150 6926 2202
rect 6926 2150 6938 2202
rect 6938 2150 6968 2202
rect 6992 2150 7002 2202
rect 7002 2150 7048 2202
rect 6752 2148 6808 2150
rect 6832 2148 6888 2150
rect 6912 2148 6968 2150
rect 6992 2148 7048 2150
rect 8684 2202 8740 2204
rect 8764 2202 8820 2204
rect 8844 2202 8900 2204
rect 8924 2202 8980 2204
rect 8684 2150 8730 2202
rect 8730 2150 8740 2202
rect 8764 2150 8794 2202
rect 8794 2150 8806 2202
rect 8806 2150 8820 2202
rect 8844 2150 8858 2202
rect 8858 2150 8870 2202
rect 8870 2150 8900 2202
rect 8924 2150 8934 2202
rect 8934 2150 8980 2202
rect 8684 2148 8740 2150
rect 8764 2148 8820 2150
rect 8844 2148 8900 2150
rect 8924 2148 8980 2150
rect 1674 720 1730 776
<< metal3 >>
rect 0 21042 800 21072
rect 1025 21042 1091 21045
rect 0 21040 1091 21042
rect 0 20984 1030 21040
rect 1086 20984 1091 21040
rect 0 20982 1091 20984
rect 0 20952 800 20982
rect 1025 20979 1091 20982
rect 0 19682 800 19712
rect 1117 19682 1183 19685
rect 0 19680 1183 19682
rect 0 19624 1122 19680
rect 1178 19624 1183 19680
rect 0 19622 1183 19624
rect 0 19592 800 19622
rect 1117 19619 1183 19622
rect 2878 19616 3194 19617
rect 2878 19552 2884 19616
rect 2948 19552 2964 19616
rect 3028 19552 3044 19616
rect 3108 19552 3124 19616
rect 3188 19552 3194 19616
rect 2878 19551 3194 19552
rect 4810 19616 5126 19617
rect 4810 19552 4816 19616
rect 4880 19552 4896 19616
rect 4960 19552 4976 19616
rect 5040 19552 5056 19616
rect 5120 19552 5126 19616
rect 4810 19551 5126 19552
rect 6742 19616 7058 19617
rect 6742 19552 6748 19616
rect 6812 19552 6828 19616
rect 6892 19552 6908 19616
rect 6972 19552 6988 19616
rect 7052 19552 7058 19616
rect 6742 19551 7058 19552
rect 8674 19616 8990 19617
rect 8674 19552 8680 19616
rect 8744 19552 8760 19616
rect 8824 19552 8840 19616
rect 8904 19552 8920 19616
rect 8984 19552 8990 19616
rect 8674 19551 8990 19552
rect 1912 19072 2228 19073
rect 1912 19008 1918 19072
rect 1982 19008 1998 19072
rect 2062 19008 2078 19072
rect 2142 19008 2158 19072
rect 2222 19008 2228 19072
rect 1912 19007 2228 19008
rect 3844 19072 4160 19073
rect 3844 19008 3850 19072
rect 3914 19008 3930 19072
rect 3994 19008 4010 19072
rect 4074 19008 4090 19072
rect 4154 19008 4160 19072
rect 3844 19007 4160 19008
rect 5776 19072 6092 19073
rect 5776 19008 5782 19072
rect 5846 19008 5862 19072
rect 5926 19008 5942 19072
rect 6006 19008 6022 19072
rect 6086 19008 6092 19072
rect 5776 19007 6092 19008
rect 7708 19072 8024 19073
rect 7708 19008 7714 19072
rect 7778 19008 7794 19072
rect 7858 19008 7874 19072
rect 7938 19008 7954 19072
rect 8018 19008 8024 19072
rect 7708 19007 8024 19008
rect 2878 18528 3194 18529
rect 2878 18464 2884 18528
rect 2948 18464 2964 18528
rect 3028 18464 3044 18528
rect 3108 18464 3124 18528
rect 3188 18464 3194 18528
rect 2878 18463 3194 18464
rect 4810 18528 5126 18529
rect 4810 18464 4816 18528
rect 4880 18464 4896 18528
rect 4960 18464 4976 18528
rect 5040 18464 5056 18528
rect 5120 18464 5126 18528
rect 4810 18463 5126 18464
rect 6742 18528 7058 18529
rect 6742 18464 6748 18528
rect 6812 18464 6828 18528
rect 6892 18464 6908 18528
rect 6972 18464 6988 18528
rect 7052 18464 7058 18528
rect 6742 18463 7058 18464
rect 8674 18528 8990 18529
rect 8674 18464 8680 18528
rect 8744 18464 8760 18528
rect 8824 18464 8840 18528
rect 8904 18464 8920 18528
rect 8984 18464 8990 18528
rect 8674 18463 8990 18464
rect 0 18322 800 18352
rect 933 18322 999 18325
rect 0 18320 999 18322
rect 0 18264 938 18320
rect 994 18264 999 18320
rect 0 18262 999 18264
rect 0 18232 800 18262
rect 933 18259 999 18262
rect 1912 17984 2228 17985
rect 1912 17920 1918 17984
rect 1982 17920 1998 17984
rect 2062 17920 2078 17984
rect 2142 17920 2158 17984
rect 2222 17920 2228 17984
rect 1912 17919 2228 17920
rect 3844 17984 4160 17985
rect 3844 17920 3850 17984
rect 3914 17920 3930 17984
rect 3994 17920 4010 17984
rect 4074 17920 4090 17984
rect 4154 17920 4160 17984
rect 3844 17919 4160 17920
rect 5776 17984 6092 17985
rect 5776 17920 5782 17984
rect 5846 17920 5862 17984
rect 5926 17920 5942 17984
rect 6006 17920 6022 17984
rect 6086 17920 6092 17984
rect 5776 17919 6092 17920
rect 7708 17984 8024 17985
rect 7708 17920 7714 17984
rect 7778 17920 7794 17984
rect 7858 17920 7874 17984
rect 7938 17920 7954 17984
rect 8018 17920 8024 17984
rect 7708 17919 8024 17920
rect 2878 17440 3194 17441
rect 2878 17376 2884 17440
rect 2948 17376 2964 17440
rect 3028 17376 3044 17440
rect 3108 17376 3124 17440
rect 3188 17376 3194 17440
rect 2878 17375 3194 17376
rect 4810 17440 5126 17441
rect 4810 17376 4816 17440
rect 4880 17376 4896 17440
rect 4960 17376 4976 17440
rect 5040 17376 5056 17440
rect 5120 17376 5126 17440
rect 4810 17375 5126 17376
rect 6742 17440 7058 17441
rect 6742 17376 6748 17440
rect 6812 17376 6828 17440
rect 6892 17376 6908 17440
rect 6972 17376 6988 17440
rect 7052 17376 7058 17440
rect 6742 17375 7058 17376
rect 8674 17440 8990 17441
rect 8674 17376 8680 17440
rect 8744 17376 8760 17440
rect 8824 17376 8840 17440
rect 8904 17376 8920 17440
rect 8984 17376 8990 17440
rect 8674 17375 8990 17376
rect 0 16962 800 16992
rect 933 16962 999 16965
rect 0 16960 999 16962
rect 0 16904 938 16960
rect 994 16904 999 16960
rect 0 16902 999 16904
rect 0 16872 800 16902
rect 933 16899 999 16902
rect 1912 16896 2228 16897
rect 1912 16832 1918 16896
rect 1982 16832 1998 16896
rect 2062 16832 2078 16896
rect 2142 16832 2158 16896
rect 2222 16832 2228 16896
rect 1912 16831 2228 16832
rect 3844 16896 4160 16897
rect 3844 16832 3850 16896
rect 3914 16832 3930 16896
rect 3994 16832 4010 16896
rect 4074 16832 4090 16896
rect 4154 16832 4160 16896
rect 3844 16831 4160 16832
rect 5776 16896 6092 16897
rect 5776 16832 5782 16896
rect 5846 16832 5862 16896
rect 5926 16832 5942 16896
rect 6006 16832 6022 16896
rect 6086 16832 6092 16896
rect 5776 16831 6092 16832
rect 7708 16896 8024 16897
rect 7708 16832 7714 16896
rect 7778 16832 7794 16896
rect 7858 16832 7874 16896
rect 7938 16832 7954 16896
rect 8018 16832 8024 16896
rect 7708 16831 8024 16832
rect 2878 16352 3194 16353
rect 2878 16288 2884 16352
rect 2948 16288 2964 16352
rect 3028 16288 3044 16352
rect 3108 16288 3124 16352
rect 3188 16288 3194 16352
rect 2878 16287 3194 16288
rect 4810 16352 5126 16353
rect 4810 16288 4816 16352
rect 4880 16288 4896 16352
rect 4960 16288 4976 16352
rect 5040 16288 5056 16352
rect 5120 16288 5126 16352
rect 4810 16287 5126 16288
rect 6742 16352 7058 16353
rect 6742 16288 6748 16352
rect 6812 16288 6828 16352
rect 6892 16288 6908 16352
rect 6972 16288 6988 16352
rect 7052 16288 7058 16352
rect 6742 16287 7058 16288
rect 8674 16352 8990 16353
rect 8674 16288 8680 16352
rect 8744 16288 8760 16352
rect 8824 16288 8840 16352
rect 8904 16288 8920 16352
rect 8984 16288 8990 16352
rect 8674 16287 8990 16288
rect 1912 15808 2228 15809
rect 1912 15744 1918 15808
rect 1982 15744 1998 15808
rect 2062 15744 2078 15808
rect 2142 15744 2158 15808
rect 2222 15744 2228 15808
rect 1912 15743 2228 15744
rect 3844 15808 4160 15809
rect 3844 15744 3850 15808
rect 3914 15744 3930 15808
rect 3994 15744 4010 15808
rect 4074 15744 4090 15808
rect 4154 15744 4160 15808
rect 3844 15743 4160 15744
rect 5776 15808 6092 15809
rect 5776 15744 5782 15808
rect 5846 15744 5862 15808
rect 5926 15744 5942 15808
rect 6006 15744 6022 15808
rect 6086 15744 6092 15808
rect 5776 15743 6092 15744
rect 7708 15808 8024 15809
rect 7708 15744 7714 15808
rect 7778 15744 7794 15808
rect 7858 15744 7874 15808
rect 7938 15744 7954 15808
rect 8018 15744 8024 15808
rect 7708 15743 8024 15744
rect 0 15602 800 15632
rect 933 15602 999 15605
rect 0 15600 999 15602
rect 0 15544 938 15600
rect 994 15544 999 15600
rect 0 15542 999 15544
rect 0 15512 800 15542
rect 933 15539 999 15542
rect 2878 15264 3194 15265
rect 2878 15200 2884 15264
rect 2948 15200 2964 15264
rect 3028 15200 3044 15264
rect 3108 15200 3124 15264
rect 3188 15200 3194 15264
rect 2878 15199 3194 15200
rect 4810 15264 5126 15265
rect 4810 15200 4816 15264
rect 4880 15200 4896 15264
rect 4960 15200 4976 15264
rect 5040 15200 5056 15264
rect 5120 15200 5126 15264
rect 4810 15199 5126 15200
rect 6742 15264 7058 15265
rect 6742 15200 6748 15264
rect 6812 15200 6828 15264
rect 6892 15200 6908 15264
rect 6972 15200 6988 15264
rect 7052 15200 7058 15264
rect 6742 15199 7058 15200
rect 8674 15264 8990 15265
rect 8674 15200 8680 15264
rect 8744 15200 8760 15264
rect 8824 15200 8840 15264
rect 8904 15200 8920 15264
rect 8984 15200 8990 15264
rect 8674 15199 8990 15200
rect 1912 14720 2228 14721
rect 1912 14656 1918 14720
rect 1982 14656 1998 14720
rect 2062 14656 2078 14720
rect 2142 14656 2158 14720
rect 2222 14656 2228 14720
rect 1912 14655 2228 14656
rect 3844 14720 4160 14721
rect 3844 14656 3850 14720
rect 3914 14656 3930 14720
rect 3994 14656 4010 14720
rect 4074 14656 4090 14720
rect 4154 14656 4160 14720
rect 3844 14655 4160 14656
rect 5776 14720 6092 14721
rect 5776 14656 5782 14720
rect 5846 14656 5862 14720
rect 5926 14656 5942 14720
rect 6006 14656 6022 14720
rect 6086 14656 6092 14720
rect 5776 14655 6092 14656
rect 7708 14720 8024 14721
rect 7708 14656 7714 14720
rect 7778 14656 7794 14720
rect 7858 14656 7874 14720
rect 7938 14656 7954 14720
rect 8018 14656 8024 14720
rect 7708 14655 8024 14656
rect 0 14242 800 14272
rect 933 14242 999 14245
rect 0 14240 999 14242
rect 0 14184 938 14240
rect 994 14184 999 14240
rect 0 14182 999 14184
rect 0 14152 800 14182
rect 933 14179 999 14182
rect 2878 14176 3194 14177
rect 2878 14112 2884 14176
rect 2948 14112 2964 14176
rect 3028 14112 3044 14176
rect 3108 14112 3124 14176
rect 3188 14112 3194 14176
rect 2878 14111 3194 14112
rect 4810 14176 5126 14177
rect 4810 14112 4816 14176
rect 4880 14112 4896 14176
rect 4960 14112 4976 14176
rect 5040 14112 5056 14176
rect 5120 14112 5126 14176
rect 4810 14111 5126 14112
rect 6742 14176 7058 14177
rect 6742 14112 6748 14176
rect 6812 14112 6828 14176
rect 6892 14112 6908 14176
rect 6972 14112 6988 14176
rect 7052 14112 7058 14176
rect 6742 14111 7058 14112
rect 8674 14176 8990 14177
rect 8674 14112 8680 14176
rect 8744 14112 8760 14176
rect 8824 14112 8840 14176
rect 8904 14112 8920 14176
rect 8984 14112 8990 14176
rect 8674 14111 8990 14112
rect 1912 13632 2228 13633
rect 1912 13568 1918 13632
rect 1982 13568 1998 13632
rect 2062 13568 2078 13632
rect 2142 13568 2158 13632
rect 2222 13568 2228 13632
rect 1912 13567 2228 13568
rect 3844 13632 4160 13633
rect 3844 13568 3850 13632
rect 3914 13568 3930 13632
rect 3994 13568 4010 13632
rect 4074 13568 4090 13632
rect 4154 13568 4160 13632
rect 3844 13567 4160 13568
rect 5776 13632 6092 13633
rect 5776 13568 5782 13632
rect 5846 13568 5862 13632
rect 5926 13568 5942 13632
rect 6006 13568 6022 13632
rect 6086 13568 6092 13632
rect 5776 13567 6092 13568
rect 7708 13632 8024 13633
rect 7708 13568 7714 13632
rect 7778 13568 7794 13632
rect 7858 13568 7874 13632
rect 7938 13568 7954 13632
rect 8018 13568 8024 13632
rect 7708 13567 8024 13568
rect 2878 13088 3194 13089
rect 2878 13024 2884 13088
rect 2948 13024 2964 13088
rect 3028 13024 3044 13088
rect 3108 13024 3124 13088
rect 3188 13024 3194 13088
rect 2878 13023 3194 13024
rect 4810 13088 5126 13089
rect 4810 13024 4816 13088
rect 4880 13024 4896 13088
rect 4960 13024 4976 13088
rect 5040 13024 5056 13088
rect 5120 13024 5126 13088
rect 4810 13023 5126 13024
rect 6742 13088 7058 13089
rect 6742 13024 6748 13088
rect 6812 13024 6828 13088
rect 6892 13024 6908 13088
rect 6972 13024 6988 13088
rect 7052 13024 7058 13088
rect 6742 13023 7058 13024
rect 8674 13088 8990 13089
rect 8674 13024 8680 13088
rect 8744 13024 8760 13088
rect 8824 13024 8840 13088
rect 8904 13024 8920 13088
rect 8984 13024 8990 13088
rect 8674 13023 8990 13024
rect 0 12882 800 12912
rect 933 12882 999 12885
rect 0 12880 999 12882
rect 0 12824 938 12880
rect 994 12824 999 12880
rect 0 12822 999 12824
rect 0 12792 800 12822
rect 933 12819 999 12822
rect 1912 12544 2228 12545
rect 1912 12480 1918 12544
rect 1982 12480 1998 12544
rect 2062 12480 2078 12544
rect 2142 12480 2158 12544
rect 2222 12480 2228 12544
rect 1912 12479 2228 12480
rect 3844 12544 4160 12545
rect 3844 12480 3850 12544
rect 3914 12480 3930 12544
rect 3994 12480 4010 12544
rect 4074 12480 4090 12544
rect 4154 12480 4160 12544
rect 3844 12479 4160 12480
rect 5776 12544 6092 12545
rect 5776 12480 5782 12544
rect 5846 12480 5862 12544
rect 5926 12480 5942 12544
rect 6006 12480 6022 12544
rect 6086 12480 6092 12544
rect 5776 12479 6092 12480
rect 7708 12544 8024 12545
rect 7708 12480 7714 12544
rect 7778 12480 7794 12544
rect 7858 12480 7874 12544
rect 7938 12480 7954 12544
rect 8018 12480 8024 12544
rect 7708 12479 8024 12480
rect 2878 12000 3194 12001
rect 2878 11936 2884 12000
rect 2948 11936 2964 12000
rect 3028 11936 3044 12000
rect 3108 11936 3124 12000
rect 3188 11936 3194 12000
rect 2878 11935 3194 11936
rect 4810 12000 5126 12001
rect 4810 11936 4816 12000
rect 4880 11936 4896 12000
rect 4960 11936 4976 12000
rect 5040 11936 5056 12000
rect 5120 11936 5126 12000
rect 4810 11935 5126 11936
rect 6742 12000 7058 12001
rect 6742 11936 6748 12000
rect 6812 11936 6828 12000
rect 6892 11936 6908 12000
rect 6972 11936 6988 12000
rect 7052 11936 7058 12000
rect 6742 11935 7058 11936
rect 8674 12000 8990 12001
rect 8674 11936 8680 12000
rect 8744 11936 8760 12000
rect 8824 11936 8840 12000
rect 8904 11936 8920 12000
rect 8984 11936 8990 12000
rect 8674 11935 8990 11936
rect 0 11522 800 11552
rect 933 11522 999 11525
rect 0 11520 999 11522
rect 0 11464 938 11520
rect 994 11464 999 11520
rect 0 11462 999 11464
rect 0 11432 800 11462
rect 933 11459 999 11462
rect 1912 11456 2228 11457
rect 1912 11392 1918 11456
rect 1982 11392 1998 11456
rect 2062 11392 2078 11456
rect 2142 11392 2158 11456
rect 2222 11392 2228 11456
rect 1912 11391 2228 11392
rect 3844 11456 4160 11457
rect 3844 11392 3850 11456
rect 3914 11392 3930 11456
rect 3994 11392 4010 11456
rect 4074 11392 4090 11456
rect 4154 11392 4160 11456
rect 3844 11391 4160 11392
rect 5776 11456 6092 11457
rect 5776 11392 5782 11456
rect 5846 11392 5862 11456
rect 5926 11392 5942 11456
rect 6006 11392 6022 11456
rect 6086 11392 6092 11456
rect 5776 11391 6092 11392
rect 7708 11456 8024 11457
rect 7708 11392 7714 11456
rect 7778 11392 7794 11456
rect 7858 11392 7874 11456
rect 7938 11392 7954 11456
rect 8018 11392 8024 11456
rect 7708 11391 8024 11392
rect 9200 10978 10000 11008
rect 9078 10918 10000 10978
rect 2878 10912 3194 10913
rect 2878 10848 2884 10912
rect 2948 10848 2964 10912
rect 3028 10848 3044 10912
rect 3108 10848 3124 10912
rect 3188 10848 3194 10912
rect 2878 10847 3194 10848
rect 4810 10912 5126 10913
rect 4810 10848 4816 10912
rect 4880 10848 4896 10912
rect 4960 10848 4976 10912
rect 5040 10848 5056 10912
rect 5120 10848 5126 10912
rect 4810 10847 5126 10848
rect 6742 10912 7058 10913
rect 6742 10848 6748 10912
rect 6812 10848 6828 10912
rect 6892 10848 6908 10912
rect 6972 10848 6988 10912
rect 7052 10848 7058 10912
rect 6742 10847 7058 10848
rect 8674 10912 8990 10913
rect 8674 10848 8680 10912
rect 8744 10848 8760 10912
rect 8824 10848 8840 10912
rect 8904 10848 8920 10912
rect 8984 10848 8990 10912
rect 8674 10847 8990 10848
rect 8201 10706 8267 10709
rect 9078 10706 9138 10918
rect 9200 10888 10000 10918
rect 8201 10704 9138 10706
rect 8201 10648 8206 10704
rect 8262 10648 9138 10704
rect 8201 10646 9138 10648
rect 8201 10643 8267 10646
rect 1912 10368 2228 10369
rect 1912 10304 1918 10368
rect 1982 10304 1998 10368
rect 2062 10304 2078 10368
rect 2142 10304 2158 10368
rect 2222 10304 2228 10368
rect 1912 10303 2228 10304
rect 3844 10368 4160 10369
rect 3844 10304 3850 10368
rect 3914 10304 3930 10368
rect 3994 10304 4010 10368
rect 4074 10304 4090 10368
rect 4154 10304 4160 10368
rect 3844 10303 4160 10304
rect 5776 10368 6092 10369
rect 5776 10304 5782 10368
rect 5846 10304 5862 10368
rect 5926 10304 5942 10368
rect 6006 10304 6022 10368
rect 6086 10304 6092 10368
rect 5776 10303 6092 10304
rect 7708 10368 8024 10369
rect 7708 10304 7714 10368
rect 7778 10304 7794 10368
rect 7858 10304 7874 10368
rect 7938 10304 7954 10368
rect 8018 10304 8024 10368
rect 7708 10303 8024 10304
rect 0 10162 800 10192
rect 933 10162 999 10165
rect 0 10160 999 10162
rect 0 10104 938 10160
rect 994 10104 999 10160
rect 0 10102 999 10104
rect 0 10072 800 10102
rect 933 10099 999 10102
rect 2878 9824 3194 9825
rect 2878 9760 2884 9824
rect 2948 9760 2964 9824
rect 3028 9760 3044 9824
rect 3108 9760 3124 9824
rect 3188 9760 3194 9824
rect 2878 9759 3194 9760
rect 4810 9824 5126 9825
rect 4810 9760 4816 9824
rect 4880 9760 4896 9824
rect 4960 9760 4976 9824
rect 5040 9760 5056 9824
rect 5120 9760 5126 9824
rect 4810 9759 5126 9760
rect 6742 9824 7058 9825
rect 6742 9760 6748 9824
rect 6812 9760 6828 9824
rect 6892 9760 6908 9824
rect 6972 9760 6988 9824
rect 7052 9760 7058 9824
rect 6742 9759 7058 9760
rect 8674 9824 8990 9825
rect 8674 9760 8680 9824
rect 8744 9760 8760 9824
rect 8824 9760 8840 9824
rect 8904 9760 8920 9824
rect 8984 9760 8990 9824
rect 8674 9759 8990 9760
rect 1912 9280 2228 9281
rect 1912 9216 1918 9280
rect 1982 9216 1998 9280
rect 2062 9216 2078 9280
rect 2142 9216 2158 9280
rect 2222 9216 2228 9280
rect 1912 9215 2228 9216
rect 3844 9280 4160 9281
rect 3844 9216 3850 9280
rect 3914 9216 3930 9280
rect 3994 9216 4010 9280
rect 4074 9216 4090 9280
rect 4154 9216 4160 9280
rect 3844 9215 4160 9216
rect 5776 9280 6092 9281
rect 5776 9216 5782 9280
rect 5846 9216 5862 9280
rect 5926 9216 5942 9280
rect 6006 9216 6022 9280
rect 6086 9216 6092 9280
rect 5776 9215 6092 9216
rect 7708 9280 8024 9281
rect 7708 9216 7714 9280
rect 7778 9216 7794 9280
rect 7858 9216 7874 9280
rect 7938 9216 7954 9280
rect 8018 9216 8024 9280
rect 7708 9215 8024 9216
rect 0 8802 800 8832
rect 933 8802 999 8805
rect 0 8800 999 8802
rect 0 8744 938 8800
rect 994 8744 999 8800
rect 0 8742 999 8744
rect 0 8712 800 8742
rect 933 8739 999 8742
rect 2878 8736 3194 8737
rect 2878 8672 2884 8736
rect 2948 8672 2964 8736
rect 3028 8672 3044 8736
rect 3108 8672 3124 8736
rect 3188 8672 3194 8736
rect 2878 8671 3194 8672
rect 4810 8736 5126 8737
rect 4810 8672 4816 8736
rect 4880 8672 4896 8736
rect 4960 8672 4976 8736
rect 5040 8672 5056 8736
rect 5120 8672 5126 8736
rect 4810 8671 5126 8672
rect 6742 8736 7058 8737
rect 6742 8672 6748 8736
rect 6812 8672 6828 8736
rect 6892 8672 6908 8736
rect 6972 8672 6988 8736
rect 7052 8672 7058 8736
rect 6742 8671 7058 8672
rect 8674 8736 8990 8737
rect 8674 8672 8680 8736
rect 8744 8672 8760 8736
rect 8824 8672 8840 8736
rect 8904 8672 8920 8736
rect 8984 8672 8990 8736
rect 8674 8671 8990 8672
rect 1912 8192 2228 8193
rect 1912 8128 1918 8192
rect 1982 8128 1998 8192
rect 2062 8128 2078 8192
rect 2142 8128 2158 8192
rect 2222 8128 2228 8192
rect 1912 8127 2228 8128
rect 3844 8192 4160 8193
rect 3844 8128 3850 8192
rect 3914 8128 3930 8192
rect 3994 8128 4010 8192
rect 4074 8128 4090 8192
rect 4154 8128 4160 8192
rect 3844 8127 4160 8128
rect 5776 8192 6092 8193
rect 5776 8128 5782 8192
rect 5846 8128 5862 8192
rect 5926 8128 5942 8192
rect 6006 8128 6022 8192
rect 6086 8128 6092 8192
rect 5776 8127 6092 8128
rect 7708 8192 8024 8193
rect 7708 8128 7714 8192
rect 7778 8128 7794 8192
rect 7858 8128 7874 8192
rect 7938 8128 7954 8192
rect 8018 8128 8024 8192
rect 7708 8127 8024 8128
rect 2878 7648 3194 7649
rect 2878 7584 2884 7648
rect 2948 7584 2964 7648
rect 3028 7584 3044 7648
rect 3108 7584 3124 7648
rect 3188 7584 3194 7648
rect 2878 7583 3194 7584
rect 4810 7648 5126 7649
rect 4810 7584 4816 7648
rect 4880 7584 4896 7648
rect 4960 7584 4976 7648
rect 5040 7584 5056 7648
rect 5120 7584 5126 7648
rect 4810 7583 5126 7584
rect 6742 7648 7058 7649
rect 6742 7584 6748 7648
rect 6812 7584 6828 7648
rect 6892 7584 6908 7648
rect 6972 7584 6988 7648
rect 7052 7584 7058 7648
rect 6742 7583 7058 7584
rect 8674 7648 8990 7649
rect 8674 7584 8680 7648
rect 8744 7584 8760 7648
rect 8824 7584 8840 7648
rect 8904 7584 8920 7648
rect 8984 7584 8990 7648
rect 8674 7583 8990 7584
rect 0 7442 800 7472
rect 933 7442 999 7445
rect 0 7440 999 7442
rect 0 7384 938 7440
rect 994 7384 999 7440
rect 0 7382 999 7384
rect 0 7352 800 7382
rect 933 7379 999 7382
rect 1912 7104 2228 7105
rect 1912 7040 1918 7104
rect 1982 7040 1998 7104
rect 2062 7040 2078 7104
rect 2142 7040 2158 7104
rect 2222 7040 2228 7104
rect 1912 7039 2228 7040
rect 3844 7104 4160 7105
rect 3844 7040 3850 7104
rect 3914 7040 3930 7104
rect 3994 7040 4010 7104
rect 4074 7040 4090 7104
rect 4154 7040 4160 7104
rect 3844 7039 4160 7040
rect 5776 7104 6092 7105
rect 5776 7040 5782 7104
rect 5846 7040 5862 7104
rect 5926 7040 5942 7104
rect 6006 7040 6022 7104
rect 6086 7040 6092 7104
rect 5776 7039 6092 7040
rect 7708 7104 8024 7105
rect 7708 7040 7714 7104
rect 7778 7040 7794 7104
rect 7858 7040 7874 7104
rect 7938 7040 7954 7104
rect 8018 7040 8024 7104
rect 7708 7039 8024 7040
rect 2878 6560 3194 6561
rect 2878 6496 2884 6560
rect 2948 6496 2964 6560
rect 3028 6496 3044 6560
rect 3108 6496 3124 6560
rect 3188 6496 3194 6560
rect 2878 6495 3194 6496
rect 4810 6560 5126 6561
rect 4810 6496 4816 6560
rect 4880 6496 4896 6560
rect 4960 6496 4976 6560
rect 5040 6496 5056 6560
rect 5120 6496 5126 6560
rect 4810 6495 5126 6496
rect 6742 6560 7058 6561
rect 6742 6496 6748 6560
rect 6812 6496 6828 6560
rect 6892 6496 6908 6560
rect 6972 6496 6988 6560
rect 7052 6496 7058 6560
rect 6742 6495 7058 6496
rect 8674 6560 8990 6561
rect 8674 6496 8680 6560
rect 8744 6496 8760 6560
rect 8824 6496 8840 6560
rect 8904 6496 8920 6560
rect 8984 6496 8990 6560
rect 8674 6495 8990 6496
rect 0 6082 800 6112
rect 933 6082 999 6085
rect 0 6080 999 6082
rect 0 6024 938 6080
rect 994 6024 999 6080
rect 0 6022 999 6024
rect 0 5992 800 6022
rect 933 6019 999 6022
rect 1912 6016 2228 6017
rect 1912 5952 1918 6016
rect 1982 5952 1998 6016
rect 2062 5952 2078 6016
rect 2142 5952 2158 6016
rect 2222 5952 2228 6016
rect 1912 5951 2228 5952
rect 3844 6016 4160 6017
rect 3844 5952 3850 6016
rect 3914 5952 3930 6016
rect 3994 5952 4010 6016
rect 4074 5952 4090 6016
rect 4154 5952 4160 6016
rect 3844 5951 4160 5952
rect 5776 6016 6092 6017
rect 5776 5952 5782 6016
rect 5846 5952 5862 6016
rect 5926 5952 5942 6016
rect 6006 5952 6022 6016
rect 6086 5952 6092 6016
rect 5776 5951 6092 5952
rect 7708 6016 8024 6017
rect 7708 5952 7714 6016
rect 7778 5952 7794 6016
rect 7858 5952 7874 6016
rect 7938 5952 7954 6016
rect 8018 5952 8024 6016
rect 7708 5951 8024 5952
rect 2878 5472 3194 5473
rect 2878 5408 2884 5472
rect 2948 5408 2964 5472
rect 3028 5408 3044 5472
rect 3108 5408 3124 5472
rect 3188 5408 3194 5472
rect 2878 5407 3194 5408
rect 4810 5472 5126 5473
rect 4810 5408 4816 5472
rect 4880 5408 4896 5472
rect 4960 5408 4976 5472
rect 5040 5408 5056 5472
rect 5120 5408 5126 5472
rect 4810 5407 5126 5408
rect 6742 5472 7058 5473
rect 6742 5408 6748 5472
rect 6812 5408 6828 5472
rect 6892 5408 6908 5472
rect 6972 5408 6988 5472
rect 7052 5408 7058 5472
rect 6742 5407 7058 5408
rect 8674 5472 8990 5473
rect 8674 5408 8680 5472
rect 8744 5408 8760 5472
rect 8824 5408 8840 5472
rect 8904 5408 8920 5472
rect 8984 5408 8990 5472
rect 8674 5407 8990 5408
rect 1912 4928 2228 4929
rect 1912 4864 1918 4928
rect 1982 4864 1998 4928
rect 2062 4864 2078 4928
rect 2142 4864 2158 4928
rect 2222 4864 2228 4928
rect 1912 4863 2228 4864
rect 3844 4928 4160 4929
rect 3844 4864 3850 4928
rect 3914 4864 3930 4928
rect 3994 4864 4010 4928
rect 4074 4864 4090 4928
rect 4154 4864 4160 4928
rect 3844 4863 4160 4864
rect 5776 4928 6092 4929
rect 5776 4864 5782 4928
rect 5846 4864 5862 4928
rect 5926 4864 5942 4928
rect 6006 4864 6022 4928
rect 6086 4864 6092 4928
rect 5776 4863 6092 4864
rect 7708 4928 8024 4929
rect 7708 4864 7714 4928
rect 7778 4864 7794 4928
rect 7858 4864 7874 4928
rect 7938 4864 7954 4928
rect 8018 4864 8024 4928
rect 7708 4863 8024 4864
rect 0 4722 800 4752
rect 933 4722 999 4725
rect 0 4720 999 4722
rect 0 4664 938 4720
rect 994 4664 999 4720
rect 0 4662 999 4664
rect 0 4632 800 4662
rect 933 4659 999 4662
rect 2878 4384 3194 4385
rect 2878 4320 2884 4384
rect 2948 4320 2964 4384
rect 3028 4320 3044 4384
rect 3108 4320 3124 4384
rect 3188 4320 3194 4384
rect 2878 4319 3194 4320
rect 4810 4384 5126 4385
rect 4810 4320 4816 4384
rect 4880 4320 4896 4384
rect 4960 4320 4976 4384
rect 5040 4320 5056 4384
rect 5120 4320 5126 4384
rect 4810 4319 5126 4320
rect 6742 4384 7058 4385
rect 6742 4320 6748 4384
rect 6812 4320 6828 4384
rect 6892 4320 6908 4384
rect 6972 4320 6988 4384
rect 7052 4320 7058 4384
rect 6742 4319 7058 4320
rect 8674 4384 8990 4385
rect 8674 4320 8680 4384
rect 8744 4320 8760 4384
rect 8824 4320 8840 4384
rect 8904 4320 8920 4384
rect 8984 4320 8990 4384
rect 8674 4319 8990 4320
rect 1912 3840 2228 3841
rect 1912 3776 1918 3840
rect 1982 3776 1998 3840
rect 2062 3776 2078 3840
rect 2142 3776 2158 3840
rect 2222 3776 2228 3840
rect 1912 3775 2228 3776
rect 3844 3840 4160 3841
rect 3844 3776 3850 3840
rect 3914 3776 3930 3840
rect 3994 3776 4010 3840
rect 4074 3776 4090 3840
rect 4154 3776 4160 3840
rect 3844 3775 4160 3776
rect 5776 3840 6092 3841
rect 5776 3776 5782 3840
rect 5846 3776 5862 3840
rect 5926 3776 5942 3840
rect 6006 3776 6022 3840
rect 6086 3776 6092 3840
rect 5776 3775 6092 3776
rect 7708 3840 8024 3841
rect 7708 3776 7714 3840
rect 7778 3776 7794 3840
rect 7858 3776 7874 3840
rect 7938 3776 7954 3840
rect 8018 3776 8024 3840
rect 7708 3775 8024 3776
rect 0 3362 800 3392
rect 933 3362 999 3365
rect 0 3360 999 3362
rect 0 3304 938 3360
rect 994 3304 999 3360
rect 0 3302 999 3304
rect 0 3272 800 3302
rect 933 3299 999 3302
rect 2878 3296 3194 3297
rect 2878 3232 2884 3296
rect 2948 3232 2964 3296
rect 3028 3232 3044 3296
rect 3108 3232 3124 3296
rect 3188 3232 3194 3296
rect 2878 3231 3194 3232
rect 4810 3296 5126 3297
rect 4810 3232 4816 3296
rect 4880 3232 4896 3296
rect 4960 3232 4976 3296
rect 5040 3232 5056 3296
rect 5120 3232 5126 3296
rect 4810 3231 5126 3232
rect 6742 3296 7058 3297
rect 6742 3232 6748 3296
rect 6812 3232 6828 3296
rect 6892 3232 6908 3296
rect 6972 3232 6988 3296
rect 7052 3232 7058 3296
rect 6742 3231 7058 3232
rect 8674 3296 8990 3297
rect 8674 3232 8680 3296
rect 8744 3232 8760 3296
rect 8824 3232 8840 3296
rect 8904 3232 8920 3296
rect 8984 3232 8990 3296
rect 8674 3231 8990 3232
rect 1912 2752 2228 2753
rect 1912 2688 1918 2752
rect 1982 2688 1998 2752
rect 2062 2688 2078 2752
rect 2142 2688 2158 2752
rect 2222 2688 2228 2752
rect 1912 2687 2228 2688
rect 3844 2752 4160 2753
rect 3844 2688 3850 2752
rect 3914 2688 3930 2752
rect 3994 2688 4010 2752
rect 4074 2688 4090 2752
rect 4154 2688 4160 2752
rect 3844 2687 4160 2688
rect 5776 2752 6092 2753
rect 5776 2688 5782 2752
rect 5846 2688 5862 2752
rect 5926 2688 5942 2752
rect 6006 2688 6022 2752
rect 6086 2688 6092 2752
rect 5776 2687 6092 2688
rect 7708 2752 8024 2753
rect 7708 2688 7714 2752
rect 7778 2688 7794 2752
rect 7858 2688 7874 2752
rect 7938 2688 7954 2752
rect 8018 2688 8024 2752
rect 7708 2687 8024 2688
rect 2878 2208 3194 2209
rect 2878 2144 2884 2208
rect 2948 2144 2964 2208
rect 3028 2144 3044 2208
rect 3108 2144 3124 2208
rect 3188 2144 3194 2208
rect 2878 2143 3194 2144
rect 4810 2208 5126 2209
rect 4810 2144 4816 2208
rect 4880 2144 4896 2208
rect 4960 2144 4976 2208
rect 5040 2144 5056 2208
rect 5120 2144 5126 2208
rect 4810 2143 5126 2144
rect 6742 2208 7058 2209
rect 6742 2144 6748 2208
rect 6812 2144 6828 2208
rect 6892 2144 6908 2208
rect 6972 2144 6988 2208
rect 7052 2144 7058 2208
rect 6742 2143 7058 2144
rect 8674 2208 8990 2209
rect 8674 2144 8680 2208
rect 8744 2144 8760 2208
rect 8824 2144 8840 2208
rect 8904 2144 8920 2208
rect 8984 2144 8990 2208
rect 8674 2143 8990 2144
rect 0 2002 800 2032
rect 933 2002 999 2005
rect 0 2000 999 2002
rect 0 1944 938 2000
rect 994 1944 999 2000
rect 0 1942 999 1944
rect 0 1912 800 1942
rect 933 1939 999 1942
rect 1669 778 1735 781
rect 982 776 1735 778
rect 982 720 1674 776
rect 1730 720 1735 776
rect 982 718 1735 720
rect 0 642 800 672
rect 982 642 1042 718
rect 1669 715 1735 718
rect 0 582 1042 642
rect 0 552 800 582
<< via3 >>
rect 2884 19612 2948 19616
rect 2884 19556 2888 19612
rect 2888 19556 2944 19612
rect 2944 19556 2948 19612
rect 2884 19552 2948 19556
rect 2964 19612 3028 19616
rect 2964 19556 2968 19612
rect 2968 19556 3024 19612
rect 3024 19556 3028 19612
rect 2964 19552 3028 19556
rect 3044 19612 3108 19616
rect 3044 19556 3048 19612
rect 3048 19556 3104 19612
rect 3104 19556 3108 19612
rect 3044 19552 3108 19556
rect 3124 19612 3188 19616
rect 3124 19556 3128 19612
rect 3128 19556 3184 19612
rect 3184 19556 3188 19612
rect 3124 19552 3188 19556
rect 4816 19612 4880 19616
rect 4816 19556 4820 19612
rect 4820 19556 4876 19612
rect 4876 19556 4880 19612
rect 4816 19552 4880 19556
rect 4896 19612 4960 19616
rect 4896 19556 4900 19612
rect 4900 19556 4956 19612
rect 4956 19556 4960 19612
rect 4896 19552 4960 19556
rect 4976 19612 5040 19616
rect 4976 19556 4980 19612
rect 4980 19556 5036 19612
rect 5036 19556 5040 19612
rect 4976 19552 5040 19556
rect 5056 19612 5120 19616
rect 5056 19556 5060 19612
rect 5060 19556 5116 19612
rect 5116 19556 5120 19612
rect 5056 19552 5120 19556
rect 6748 19612 6812 19616
rect 6748 19556 6752 19612
rect 6752 19556 6808 19612
rect 6808 19556 6812 19612
rect 6748 19552 6812 19556
rect 6828 19612 6892 19616
rect 6828 19556 6832 19612
rect 6832 19556 6888 19612
rect 6888 19556 6892 19612
rect 6828 19552 6892 19556
rect 6908 19612 6972 19616
rect 6908 19556 6912 19612
rect 6912 19556 6968 19612
rect 6968 19556 6972 19612
rect 6908 19552 6972 19556
rect 6988 19612 7052 19616
rect 6988 19556 6992 19612
rect 6992 19556 7048 19612
rect 7048 19556 7052 19612
rect 6988 19552 7052 19556
rect 8680 19612 8744 19616
rect 8680 19556 8684 19612
rect 8684 19556 8740 19612
rect 8740 19556 8744 19612
rect 8680 19552 8744 19556
rect 8760 19612 8824 19616
rect 8760 19556 8764 19612
rect 8764 19556 8820 19612
rect 8820 19556 8824 19612
rect 8760 19552 8824 19556
rect 8840 19612 8904 19616
rect 8840 19556 8844 19612
rect 8844 19556 8900 19612
rect 8900 19556 8904 19612
rect 8840 19552 8904 19556
rect 8920 19612 8984 19616
rect 8920 19556 8924 19612
rect 8924 19556 8980 19612
rect 8980 19556 8984 19612
rect 8920 19552 8984 19556
rect 1918 19068 1982 19072
rect 1918 19012 1922 19068
rect 1922 19012 1978 19068
rect 1978 19012 1982 19068
rect 1918 19008 1982 19012
rect 1998 19068 2062 19072
rect 1998 19012 2002 19068
rect 2002 19012 2058 19068
rect 2058 19012 2062 19068
rect 1998 19008 2062 19012
rect 2078 19068 2142 19072
rect 2078 19012 2082 19068
rect 2082 19012 2138 19068
rect 2138 19012 2142 19068
rect 2078 19008 2142 19012
rect 2158 19068 2222 19072
rect 2158 19012 2162 19068
rect 2162 19012 2218 19068
rect 2218 19012 2222 19068
rect 2158 19008 2222 19012
rect 3850 19068 3914 19072
rect 3850 19012 3854 19068
rect 3854 19012 3910 19068
rect 3910 19012 3914 19068
rect 3850 19008 3914 19012
rect 3930 19068 3994 19072
rect 3930 19012 3934 19068
rect 3934 19012 3990 19068
rect 3990 19012 3994 19068
rect 3930 19008 3994 19012
rect 4010 19068 4074 19072
rect 4010 19012 4014 19068
rect 4014 19012 4070 19068
rect 4070 19012 4074 19068
rect 4010 19008 4074 19012
rect 4090 19068 4154 19072
rect 4090 19012 4094 19068
rect 4094 19012 4150 19068
rect 4150 19012 4154 19068
rect 4090 19008 4154 19012
rect 5782 19068 5846 19072
rect 5782 19012 5786 19068
rect 5786 19012 5842 19068
rect 5842 19012 5846 19068
rect 5782 19008 5846 19012
rect 5862 19068 5926 19072
rect 5862 19012 5866 19068
rect 5866 19012 5922 19068
rect 5922 19012 5926 19068
rect 5862 19008 5926 19012
rect 5942 19068 6006 19072
rect 5942 19012 5946 19068
rect 5946 19012 6002 19068
rect 6002 19012 6006 19068
rect 5942 19008 6006 19012
rect 6022 19068 6086 19072
rect 6022 19012 6026 19068
rect 6026 19012 6082 19068
rect 6082 19012 6086 19068
rect 6022 19008 6086 19012
rect 7714 19068 7778 19072
rect 7714 19012 7718 19068
rect 7718 19012 7774 19068
rect 7774 19012 7778 19068
rect 7714 19008 7778 19012
rect 7794 19068 7858 19072
rect 7794 19012 7798 19068
rect 7798 19012 7854 19068
rect 7854 19012 7858 19068
rect 7794 19008 7858 19012
rect 7874 19068 7938 19072
rect 7874 19012 7878 19068
rect 7878 19012 7934 19068
rect 7934 19012 7938 19068
rect 7874 19008 7938 19012
rect 7954 19068 8018 19072
rect 7954 19012 7958 19068
rect 7958 19012 8014 19068
rect 8014 19012 8018 19068
rect 7954 19008 8018 19012
rect 2884 18524 2948 18528
rect 2884 18468 2888 18524
rect 2888 18468 2944 18524
rect 2944 18468 2948 18524
rect 2884 18464 2948 18468
rect 2964 18524 3028 18528
rect 2964 18468 2968 18524
rect 2968 18468 3024 18524
rect 3024 18468 3028 18524
rect 2964 18464 3028 18468
rect 3044 18524 3108 18528
rect 3044 18468 3048 18524
rect 3048 18468 3104 18524
rect 3104 18468 3108 18524
rect 3044 18464 3108 18468
rect 3124 18524 3188 18528
rect 3124 18468 3128 18524
rect 3128 18468 3184 18524
rect 3184 18468 3188 18524
rect 3124 18464 3188 18468
rect 4816 18524 4880 18528
rect 4816 18468 4820 18524
rect 4820 18468 4876 18524
rect 4876 18468 4880 18524
rect 4816 18464 4880 18468
rect 4896 18524 4960 18528
rect 4896 18468 4900 18524
rect 4900 18468 4956 18524
rect 4956 18468 4960 18524
rect 4896 18464 4960 18468
rect 4976 18524 5040 18528
rect 4976 18468 4980 18524
rect 4980 18468 5036 18524
rect 5036 18468 5040 18524
rect 4976 18464 5040 18468
rect 5056 18524 5120 18528
rect 5056 18468 5060 18524
rect 5060 18468 5116 18524
rect 5116 18468 5120 18524
rect 5056 18464 5120 18468
rect 6748 18524 6812 18528
rect 6748 18468 6752 18524
rect 6752 18468 6808 18524
rect 6808 18468 6812 18524
rect 6748 18464 6812 18468
rect 6828 18524 6892 18528
rect 6828 18468 6832 18524
rect 6832 18468 6888 18524
rect 6888 18468 6892 18524
rect 6828 18464 6892 18468
rect 6908 18524 6972 18528
rect 6908 18468 6912 18524
rect 6912 18468 6968 18524
rect 6968 18468 6972 18524
rect 6908 18464 6972 18468
rect 6988 18524 7052 18528
rect 6988 18468 6992 18524
rect 6992 18468 7048 18524
rect 7048 18468 7052 18524
rect 6988 18464 7052 18468
rect 8680 18524 8744 18528
rect 8680 18468 8684 18524
rect 8684 18468 8740 18524
rect 8740 18468 8744 18524
rect 8680 18464 8744 18468
rect 8760 18524 8824 18528
rect 8760 18468 8764 18524
rect 8764 18468 8820 18524
rect 8820 18468 8824 18524
rect 8760 18464 8824 18468
rect 8840 18524 8904 18528
rect 8840 18468 8844 18524
rect 8844 18468 8900 18524
rect 8900 18468 8904 18524
rect 8840 18464 8904 18468
rect 8920 18524 8984 18528
rect 8920 18468 8924 18524
rect 8924 18468 8980 18524
rect 8980 18468 8984 18524
rect 8920 18464 8984 18468
rect 1918 17980 1982 17984
rect 1918 17924 1922 17980
rect 1922 17924 1978 17980
rect 1978 17924 1982 17980
rect 1918 17920 1982 17924
rect 1998 17980 2062 17984
rect 1998 17924 2002 17980
rect 2002 17924 2058 17980
rect 2058 17924 2062 17980
rect 1998 17920 2062 17924
rect 2078 17980 2142 17984
rect 2078 17924 2082 17980
rect 2082 17924 2138 17980
rect 2138 17924 2142 17980
rect 2078 17920 2142 17924
rect 2158 17980 2222 17984
rect 2158 17924 2162 17980
rect 2162 17924 2218 17980
rect 2218 17924 2222 17980
rect 2158 17920 2222 17924
rect 3850 17980 3914 17984
rect 3850 17924 3854 17980
rect 3854 17924 3910 17980
rect 3910 17924 3914 17980
rect 3850 17920 3914 17924
rect 3930 17980 3994 17984
rect 3930 17924 3934 17980
rect 3934 17924 3990 17980
rect 3990 17924 3994 17980
rect 3930 17920 3994 17924
rect 4010 17980 4074 17984
rect 4010 17924 4014 17980
rect 4014 17924 4070 17980
rect 4070 17924 4074 17980
rect 4010 17920 4074 17924
rect 4090 17980 4154 17984
rect 4090 17924 4094 17980
rect 4094 17924 4150 17980
rect 4150 17924 4154 17980
rect 4090 17920 4154 17924
rect 5782 17980 5846 17984
rect 5782 17924 5786 17980
rect 5786 17924 5842 17980
rect 5842 17924 5846 17980
rect 5782 17920 5846 17924
rect 5862 17980 5926 17984
rect 5862 17924 5866 17980
rect 5866 17924 5922 17980
rect 5922 17924 5926 17980
rect 5862 17920 5926 17924
rect 5942 17980 6006 17984
rect 5942 17924 5946 17980
rect 5946 17924 6002 17980
rect 6002 17924 6006 17980
rect 5942 17920 6006 17924
rect 6022 17980 6086 17984
rect 6022 17924 6026 17980
rect 6026 17924 6082 17980
rect 6082 17924 6086 17980
rect 6022 17920 6086 17924
rect 7714 17980 7778 17984
rect 7714 17924 7718 17980
rect 7718 17924 7774 17980
rect 7774 17924 7778 17980
rect 7714 17920 7778 17924
rect 7794 17980 7858 17984
rect 7794 17924 7798 17980
rect 7798 17924 7854 17980
rect 7854 17924 7858 17980
rect 7794 17920 7858 17924
rect 7874 17980 7938 17984
rect 7874 17924 7878 17980
rect 7878 17924 7934 17980
rect 7934 17924 7938 17980
rect 7874 17920 7938 17924
rect 7954 17980 8018 17984
rect 7954 17924 7958 17980
rect 7958 17924 8014 17980
rect 8014 17924 8018 17980
rect 7954 17920 8018 17924
rect 2884 17436 2948 17440
rect 2884 17380 2888 17436
rect 2888 17380 2944 17436
rect 2944 17380 2948 17436
rect 2884 17376 2948 17380
rect 2964 17436 3028 17440
rect 2964 17380 2968 17436
rect 2968 17380 3024 17436
rect 3024 17380 3028 17436
rect 2964 17376 3028 17380
rect 3044 17436 3108 17440
rect 3044 17380 3048 17436
rect 3048 17380 3104 17436
rect 3104 17380 3108 17436
rect 3044 17376 3108 17380
rect 3124 17436 3188 17440
rect 3124 17380 3128 17436
rect 3128 17380 3184 17436
rect 3184 17380 3188 17436
rect 3124 17376 3188 17380
rect 4816 17436 4880 17440
rect 4816 17380 4820 17436
rect 4820 17380 4876 17436
rect 4876 17380 4880 17436
rect 4816 17376 4880 17380
rect 4896 17436 4960 17440
rect 4896 17380 4900 17436
rect 4900 17380 4956 17436
rect 4956 17380 4960 17436
rect 4896 17376 4960 17380
rect 4976 17436 5040 17440
rect 4976 17380 4980 17436
rect 4980 17380 5036 17436
rect 5036 17380 5040 17436
rect 4976 17376 5040 17380
rect 5056 17436 5120 17440
rect 5056 17380 5060 17436
rect 5060 17380 5116 17436
rect 5116 17380 5120 17436
rect 5056 17376 5120 17380
rect 6748 17436 6812 17440
rect 6748 17380 6752 17436
rect 6752 17380 6808 17436
rect 6808 17380 6812 17436
rect 6748 17376 6812 17380
rect 6828 17436 6892 17440
rect 6828 17380 6832 17436
rect 6832 17380 6888 17436
rect 6888 17380 6892 17436
rect 6828 17376 6892 17380
rect 6908 17436 6972 17440
rect 6908 17380 6912 17436
rect 6912 17380 6968 17436
rect 6968 17380 6972 17436
rect 6908 17376 6972 17380
rect 6988 17436 7052 17440
rect 6988 17380 6992 17436
rect 6992 17380 7048 17436
rect 7048 17380 7052 17436
rect 6988 17376 7052 17380
rect 8680 17436 8744 17440
rect 8680 17380 8684 17436
rect 8684 17380 8740 17436
rect 8740 17380 8744 17436
rect 8680 17376 8744 17380
rect 8760 17436 8824 17440
rect 8760 17380 8764 17436
rect 8764 17380 8820 17436
rect 8820 17380 8824 17436
rect 8760 17376 8824 17380
rect 8840 17436 8904 17440
rect 8840 17380 8844 17436
rect 8844 17380 8900 17436
rect 8900 17380 8904 17436
rect 8840 17376 8904 17380
rect 8920 17436 8984 17440
rect 8920 17380 8924 17436
rect 8924 17380 8980 17436
rect 8980 17380 8984 17436
rect 8920 17376 8984 17380
rect 1918 16892 1982 16896
rect 1918 16836 1922 16892
rect 1922 16836 1978 16892
rect 1978 16836 1982 16892
rect 1918 16832 1982 16836
rect 1998 16892 2062 16896
rect 1998 16836 2002 16892
rect 2002 16836 2058 16892
rect 2058 16836 2062 16892
rect 1998 16832 2062 16836
rect 2078 16892 2142 16896
rect 2078 16836 2082 16892
rect 2082 16836 2138 16892
rect 2138 16836 2142 16892
rect 2078 16832 2142 16836
rect 2158 16892 2222 16896
rect 2158 16836 2162 16892
rect 2162 16836 2218 16892
rect 2218 16836 2222 16892
rect 2158 16832 2222 16836
rect 3850 16892 3914 16896
rect 3850 16836 3854 16892
rect 3854 16836 3910 16892
rect 3910 16836 3914 16892
rect 3850 16832 3914 16836
rect 3930 16892 3994 16896
rect 3930 16836 3934 16892
rect 3934 16836 3990 16892
rect 3990 16836 3994 16892
rect 3930 16832 3994 16836
rect 4010 16892 4074 16896
rect 4010 16836 4014 16892
rect 4014 16836 4070 16892
rect 4070 16836 4074 16892
rect 4010 16832 4074 16836
rect 4090 16892 4154 16896
rect 4090 16836 4094 16892
rect 4094 16836 4150 16892
rect 4150 16836 4154 16892
rect 4090 16832 4154 16836
rect 5782 16892 5846 16896
rect 5782 16836 5786 16892
rect 5786 16836 5842 16892
rect 5842 16836 5846 16892
rect 5782 16832 5846 16836
rect 5862 16892 5926 16896
rect 5862 16836 5866 16892
rect 5866 16836 5922 16892
rect 5922 16836 5926 16892
rect 5862 16832 5926 16836
rect 5942 16892 6006 16896
rect 5942 16836 5946 16892
rect 5946 16836 6002 16892
rect 6002 16836 6006 16892
rect 5942 16832 6006 16836
rect 6022 16892 6086 16896
rect 6022 16836 6026 16892
rect 6026 16836 6082 16892
rect 6082 16836 6086 16892
rect 6022 16832 6086 16836
rect 7714 16892 7778 16896
rect 7714 16836 7718 16892
rect 7718 16836 7774 16892
rect 7774 16836 7778 16892
rect 7714 16832 7778 16836
rect 7794 16892 7858 16896
rect 7794 16836 7798 16892
rect 7798 16836 7854 16892
rect 7854 16836 7858 16892
rect 7794 16832 7858 16836
rect 7874 16892 7938 16896
rect 7874 16836 7878 16892
rect 7878 16836 7934 16892
rect 7934 16836 7938 16892
rect 7874 16832 7938 16836
rect 7954 16892 8018 16896
rect 7954 16836 7958 16892
rect 7958 16836 8014 16892
rect 8014 16836 8018 16892
rect 7954 16832 8018 16836
rect 2884 16348 2948 16352
rect 2884 16292 2888 16348
rect 2888 16292 2944 16348
rect 2944 16292 2948 16348
rect 2884 16288 2948 16292
rect 2964 16348 3028 16352
rect 2964 16292 2968 16348
rect 2968 16292 3024 16348
rect 3024 16292 3028 16348
rect 2964 16288 3028 16292
rect 3044 16348 3108 16352
rect 3044 16292 3048 16348
rect 3048 16292 3104 16348
rect 3104 16292 3108 16348
rect 3044 16288 3108 16292
rect 3124 16348 3188 16352
rect 3124 16292 3128 16348
rect 3128 16292 3184 16348
rect 3184 16292 3188 16348
rect 3124 16288 3188 16292
rect 4816 16348 4880 16352
rect 4816 16292 4820 16348
rect 4820 16292 4876 16348
rect 4876 16292 4880 16348
rect 4816 16288 4880 16292
rect 4896 16348 4960 16352
rect 4896 16292 4900 16348
rect 4900 16292 4956 16348
rect 4956 16292 4960 16348
rect 4896 16288 4960 16292
rect 4976 16348 5040 16352
rect 4976 16292 4980 16348
rect 4980 16292 5036 16348
rect 5036 16292 5040 16348
rect 4976 16288 5040 16292
rect 5056 16348 5120 16352
rect 5056 16292 5060 16348
rect 5060 16292 5116 16348
rect 5116 16292 5120 16348
rect 5056 16288 5120 16292
rect 6748 16348 6812 16352
rect 6748 16292 6752 16348
rect 6752 16292 6808 16348
rect 6808 16292 6812 16348
rect 6748 16288 6812 16292
rect 6828 16348 6892 16352
rect 6828 16292 6832 16348
rect 6832 16292 6888 16348
rect 6888 16292 6892 16348
rect 6828 16288 6892 16292
rect 6908 16348 6972 16352
rect 6908 16292 6912 16348
rect 6912 16292 6968 16348
rect 6968 16292 6972 16348
rect 6908 16288 6972 16292
rect 6988 16348 7052 16352
rect 6988 16292 6992 16348
rect 6992 16292 7048 16348
rect 7048 16292 7052 16348
rect 6988 16288 7052 16292
rect 8680 16348 8744 16352
rect 8680 16292 8684 16348
rect 8684 16292 8740 16348
rect 8740 16292 8744 16348
rect 8680 16288 8744 16292
rect 8760 16348 8824 16352
rect 8760 16292 8764 16348
rect 8764 16292 8820 16348
rect 8820 16292 8824 16348
rect 8760 16288 8824 16292
rect 8840 16348 8904 16352
rect 8840 16292 8844 16348
rect 8844 16292 8900 16348
rect 8900 16292 8904 16348
rect 8840 16288 8904 16292
rect 8920 16348 8984 16352
rect 8920 16292 8924 16348
rect 8924 16292 8980 16348
rect 8980 16292 8984 16348
rect 8920 16288 8984 16292
rect 1918 15804 1982 15808
rect 1918 15748 1922 15804
rect 1922 15748 1978 15804
rect 1978 15748 1982 15804
rect 1918 15744 1982 15748
rect 1998 15804 2062 15808
rect 1998 15748 2002 15804
rect 2002 15748 2058 15804
rect 2058 15748 2062 15804
rect 1998 15744 2062 15748
rect 2078 15804 2142 15808
rect 2078 15748 2082 15804
rect 2082 15748 2138 15804
rect 2138 15748 2142 15804
rect 2078 15744 2142 15748
rect 2158 15804 2222 15808
rect 2158 15748 2162 15804
rect 2162 15748 2218 15804
rect 2218 15748 2222 15804
rect 2158 15744 2222 15748
rect 3850 15804 3914 15808
rect 3850 15748 3854 15804
rect 3854 15748 3910 15804
rect 3910 15748 3914 15804
rect 3850 15744 3914 15748
rect 3930 15804 3994 15808
rect 3930 15748 3934 15804
rect 3934 15748 3990 15804
rect 3990 15748 3994 15804
rect 3930 15744 3994 15748
rect 4010 15804 4074 15808
rect 4010 15748 4014 15804
rect 4014 15748 4070 15804
rect 4070 15748 4074 15804
rect 4010 15744 4074 15748
rect 4090 15804 4154 15808
rect 4090 15748 4094 15804
rect 4094 15748 4150 15804
rect 4150 15748 4154 15804
rect 4090 15744 4154 15748
rect 5782 15804 5846 15808
rect 5782 15748 5786 15804
rect 5786 15748 5842 15804
rect 5842 15748 5846 15804
rect 5782 15744 5846 15748
rect 5862 15804 5926 15808
rect 5862 15748 5866 15804
rect 5866 15748 5922 15804
rect 5922 15748 5926 15804
rect 5862 15744 5926 15748
rect 5942 15804 6006 15808
rect 5942 15748 5946 15804
rect 5946 15748 6002 15804
rect 6002 15748 6006 15804
rect 5942 15744 6006 15748
rect 6022 15804 6086 15808
rect 6022 15748 6026 15804
rect 6026 15748 6082 15804
rect 6082 15748 6086 15804
rect 6022 15744 6086 15748
rect 7714 15804 7778 15808
rect 7714 15748 7718 15804
rect 7718 15748 7774 15804
rect 7774 15748 7778 15804
rect 7714 15744 7778 15748
rect 7794 15804 7858 15808
rect 7794 15748 7798 15804
rect 7798 15748 7854 15804
rect 7854 15748 7858 15804
rect 7794 15744 7858 15748
rect 7874 15804 7938 15808
rect 7874 15748 7878 15804
rect 7878 15748 7934 15804
rect 7934 15748 7938 15804
rect 7874 15744 7938 15748
rect 7954 15804 8018 15808
rect 7954 15748 7958 15804
rect 7958 15748 8014 15804
rect 8014 15748 8018 15804
rect 7954 15744 8018 15748
rect 2884 15260 2948 15264
rect 2884 15204 2888 15260
rect 2888 15204 2944 15260
rect 2944 15204 2948 15260
rect 2884 15200 2948 15204
rect 2964 15260 3028 15264
rect 2964 15204 2968 15260
rect 2968 15204 3024 15260
rect 3024 15204 3028 15260
rect 2964 15200 3028 15204
rect 3044 15260 3108 15264
rect 3044 15204 3048 15260
rect 3048 15204 3104 15260
rect 3104 15204 3108 15260
rect 3044 15200 3108 15204
rect 3124 15260 3188 15264
rect 3124 15204 3128 15260
rect 3128 15204 3184 15260
rect 3184 15204 3188 15260
rect 3124 15200 3188 15204
rect 4816 15260 4880 15264
rect 4816 15204 4820 15260
rect 4820 15204 4876 15260
rect 4876 15204 4880 15260
rect 4816 15200 4880 15204
rect 4896 15260 4960 15264
rect 4896 15204 4900 15260
rect 4900 15204 4956 15260
rect 4956 15204 4960 15260
rect 4896 15200 4960 15204
rect 4976 15260 5040 15264
rect 4976 15204 4980 15260
rect 4980 15204 5036 15260
rect 5036 15204 5040 15260
rect 4976 15200 5040 15204
rect 5056 15260 5120 15264
rect 5056 15204 5060 15260
rect 5060 15204 5116 15260
rect 5116 15204 5120 15260
rect 5056 15200 5120 15204
rect 6748 15260 6812 15264
rect 6748 15204 6752 15260
rect 6752 15204 6808 15260
rect 6808 15204 6812 15260
rect 6748 15200 6812 15204
rect 6828 15260 6892 15264
rect 6828 15204 6832 15260
rect 6832 15204 6888 15260
rect 6888 15204 6892 15260
rect 6828 15200 6892 15204
rect 6908 15260 6972 15264
rect 6908 15204 6912 15260
rect 6912 15204 6968 15260
rect 6968 15204 6972 15260
rect 6908 15200 6972 15204
rect 6988 15260 7052 15264
rect 6988 15204 6992 15260
rect 6992 15204 7048 15260
rect 7048 15204 7052 15260
rect 6988 15200 7052 15204
rect 8680 15260 8744 15264
rect 8680 15204 8684 15260
rect 8684 15204 8740 15260
rect 8740 15204 8744 15260
rect 8680 15200 8744 15204
rect 8760 15260 8824 15264
rect 8760 15204 8764 15260
rect 8764 15204 8820 15260
rect 8820 15204 8824 15260
rect 8760 15200 8824 15204
rect 8840 15260 8904 15264
rect 8840 15204 8844 15260
rect 8844 15204 8900 15260
rect 8900 15204 8904 15260
rect 8840 15200 8904 15204
rect 8920 15260 8984 15264
rect 8920 15204 8924 15260
rect 8924 15204 8980 15260
rect 8980 15204 8984 15260
rect 8920 15200 8984 15204
rect 1918 14716 1982 14720
rect 1918 14660 1922 14716
rect 1922 14660 1978 14716
rect 1978 14660 1982 14716
rect 1918 14656 1982 14660
rect 1998 14716 2062 14720
rect 1998 14660 2002 14716
rect 2002 14660 2058 14716
rect 2058 14660 2062 14716
rect 1998 14656 2062 14660
rect 2078 14716 2142 14720
rect 2078 14660 2082 14716
rect 2082 14660 2138 14716
rect 2138 14660 2142 14716
rect 2078 14656 2142 14660
rect 2158 14716 2222 14720
rect 2158 14660 2162 14716
rect 2162 14660 2218 14716
rect 2218 14660 2222 14716
rect 2158 14656 2222 14660
rect 3850 14716 3914 14720
rect 3850 14660 3854 14716
rect 3854 14660 3910 14716
rect 3910 14660 3914 14716
rect 3850 14656 3914 14660
rect 3930 14716 3994 14720
rect 3930 14660 3934 14716
rect 3934 14660 3990 14716
rect 3990 14660 3994 14716
rect 3930 14656 3994 14660
rect 4010 14716 4074 14720
rect 4010 14660 4014 14716
rect 4014 14660 4070 14716
rect 4070 14660 4074 14716
rect 4010 14656 4074 14660
rect 4090 14716 4154 14720
rect 4090 14660 4094 14716
rect 4094 14660 4150 14716
rect 4150 14660 4154 14716
rect 4090 14656 4154 14660
rect 5782 14716 5846 14720
rect 5782 14660 5786 14716
rect 5786 14660 5842 14716
rect 5842 14660 5846 14716
rect 5782 14656 5846 14660
rect 5862 14716 5926 14720
rect 5862 14660 5866 14716
rect 5866 14660 5922 14716
rect 5922 14660 5926 14716
rect 5862 14656 5926 14660
rect 5942 14716 6006 14720
rect 5942 14660 5946 14716
rect 5946 14660 6002 14716
rect 6002 14660 6006 14716
rect 5942 14656 6006 14660
rect 6022 14716 6086 14720
rect 6022 14660 6026 14716
rect 6026 14660 6082 14716
rect 6082 14660 6086 14716
rect 6022 14656 6086 14660
rect 7714 14716 7778 14720
rect 7714 14660 7718 14716
rect 7718 14660 7774 14716
rect 7774 14660 7778 14716
rect 7714 14656 7778 14660
rect 7794 14716 7858 14720
rect 7794 14660 7798 14716
rect 7798 14660 7854 14716
rect 7854 14660 7858 14716
rect 7794 14656 7858 14660
rect 7874 14716 7938 14720
rect 7874 14660 7878 14716
rect 7878 14660 7934 14716
rect 7934 14660 7938 14716
rect 7874 14656 7938 14660
rect 7954 14716 8018 14720
rect 7954 14660 7958 14716
rect 7958 14660 8014 14716
rect 8014 14660 8018 14716
rect 7954 14656 8018 14660
rect 2884 14172 2948 14176
rect 2884 14116 2888 14172
rect 2888 14116 2944 14172
rect 2944 14116 2948 14172
rect 2884 14112 2948 14116
rect 2964 14172 3028 14176
rect 2964 14116 2968 14172
rect 2968 14116 3024 14172
rect 3024 14116 3028 14172
rect 2964 14112 3028 14116
rect 3044 14172 3108 14176
rect 3044 14116 3048 14172
rect 3048 14116 3104 14172
rect 3104 14116 3108 14172
rect 3044 14112 3108 14116
rect 3124 14172 3188 14176
rect 3124 14116 3128 14172
rect 3128 14116 3184 14172
rect 3184 14116 3188 14172
rect 3124 14112 3188 14116
rect 4816 14172 4880 14176
rect 4816 14116 4820 14172
rect 4820 14116 4876 14172
rect 4876 14116 4880 14172
rect 4816 14112 4880 14116
rect 4896 14172 4960 14176
rect 4896 14116 4900 14172
rect 4900 14116 4956 14172
rect 4956 14116 4960 14172
rect 4896 14112 4960 14116
rect 4976 14172 5040 14176
rect 4976 14116 4980 14172
rect 4980 14116 5036 14172
rect 5036 14116 5040 14172
rect 4976 14112 5040 14116
rect 5056 14172 5120 14176
rect 5056 14116 5060 14172
rect 5060 14116 5116 14172
rect 5116 14116 5120 14172
rect 5056 14112 5120 14116
rect 6748 14172 6812 14176
rect 6748 14116 6752 14172
rect 6752 14116 6808 14172
rect 6808 14116 6812 14172
rect 6748 14112 6812 14116
rect 6828 14172 6892 14176
rect 6828 14116 6832 14172
rect 6832 14116 6888 14172
rect 6888 14116 6892 14172
rect 6828 14112 6892 14116
rect 6908 14172 6972 14176
rect 6908 14116 6912 14172
rect 6912 14116 6968 14172
rect 6968 14116 6972 14172
rect 6908 14112 6972 14116
rect 6988 14172 7052 14176
rect 6988 14116 6992 14172
rect 6992 14116 7048 14172
rect 7048 14116 7052 14172
rect 6988 14112 7052 14116
rect 8680 14172 8744 14176
rect 8680 14116 8684 14172
rect 8684 14116 8740 14172
rect 8740 14116 8744 14172
rect 8680 14112 8744 14116
rect 8760 14172 8824 14176
rect 8760 14116 8764 14172
rect 8764 14116 8820 14172
rect 8820 14116 8824 14172
rect 8760 14112 8824 14116
rect 8840 14172 8904 14176
rect 8840 14116 8844 14172
rect 8844 14116 8900 14172
rect 8900 14116 8904 14172
rect 8840 14112 8904 14116
rect 8920 14172 8984 14176
rect 8920 14116 8924 14172
rect 8924 14116 8980 14172
rect 8980 14116 8984 14172
rect 8920 14112 8984 14116
rect 1918 13628 1982 13632
rect 1918 13572 1922 13628
rect 1922 13572 1978 13628
rect 1978 13572 1982 13628
rect 1918 13568 1982 13572
rect 1998 13628 2062 13632
rect 1998 13572 2002 13628
rect 2002 13572 2058 13628
rect 2058 13572 2062 13628
rect 1998 13568 2062 13572
rect 2078 13628 2142 13632
rect 2078 13572 2082 13628
rect 2082 13572 2138 13628
rect 2138 13572 2142 13628
rect 2078 13568 2142 13572
rect 2158 13628 2222 13632
rect 2158 13572 2162 13628
rect 2162 13572 2218 13628
rect 2218 13572 2222 13628
rect 2158 13568 2222 13572
rect 3850 13628 3914 13632
rect 3850 13572 3854 13628
rect 3854 13572 3910 13628
rect 3910 13572 3914 13628
rect 3850 13568 3914 13572
rect 3930 13628 3994 13632
rect 3930 13572 3934 13628
rect 3934 13572 3990 13628
rect 3990 13572 3994 13628
rect 3930 13568 3994 13572
rect 4010 13628 4074 13632
rect 4010 13572 4014 13628
rect 4014 13572 4070 13628
rect 4070 13572 4074 13628
rect 4010 13568 4074 13572
rect 4090 13628 4154 13632
rect 4090 13572 4094 13628
rect 4094 13572 4150 13628
rect 4150 13572 4154 13628
rect 4090 13568 4154 13572
rect 5782 13628 5846 13632
rect 5782 13572 5786 13628
rect 5786 13572 5842 13628
rect 5842 13572 5846 13628
rect 5782 13568 5846 13572
rect 5862 13628 5926 13632
rect 5862 13572 5866 13628
rect 5866 13572 5922 13628
rect 5922 13572 5926 13628
rect 5862 13568 5926 13572
rect 5942 13628 6006 13632
rect 5942 13572 5946 13628
rect 5946 13572 6002 13628
rect 6002 13572 6006 13628
rect 5942 13568 6006 13572
rect 6022 13628 6086 13632
rect 6022 13572 6026 13628
rect 6026 13572 6082 13628
rect 6082 13572 6086 13628
rect 6022 13568 6086 13572
rect 7714 13628 7778 13632
rect 7714 13572 7718 13628
rect 7718 13572 7774 13628
rect 7774 13572 7778 13628
rect 7714 13568 7778 13572
rect 7794 13628 7858 13632
rect 7794 13572 7798 13628
rect 7798 13572 7854 13628
rect 7854 13572 7858 13628
rect 7794 13568 7858 13572
rect 7874 13628 7938 13632
rect 7874 13572 7878 13628
rect 7878 13572 7934 13628
rect 7934 13572 7938 13628
rect 7874 13568 7938 13572
rect 7954 13628 8018 13632
rect 7954 13572 7958 13628
rect 7958 13572 8014 13628
rect 8014 13572 8018 13628
rect 7954 13568 8018 13572
rect 2884 13084 2948 13088
rect 2884 13028 2888 13084
rect 2888 13028 2944 13084
rect 2944 13028 2948 13084
rect 2884 13024 2948 13028
rect 2964 13084 3028 13088
rect 2964 13028 2968 13084
rect 2968 13028 3024 13084
rect 3024 13028 3028 13084
rect 2964 13024 3028 13028
rect 3044 13084 3108 13088
rect 3044 13028 3048 13084
rect 3048 13028 3104 13084
rect 3104 13028 3108 13084
rect 3044 13024 3108 13028
rect 3124 13084 3188 13088
rect 3124 13028 3128 13084
rect 3128 13028 3184 13084
rect 3184 13028 3188 13084
rect 3124 13024 3188 13028
rect 4816 13084 4880 13088
rect 4816 13028 4820 13084
rect 4820 13028 4876 13084
rect 4876 13028 4880 13084
rect 4816 13024 4880 13028
rect 4896 13084 4960 13088
rect 4896 13028 4900 13084
rect 4900 13028 4956 13084
rect 4956 13028 4960 13084
rect 4896 13024 4960 13028
rect 4976 13084 5040 13088
rect 4976 13028 4980 13084
rect 4980 13028 5036 13084
rect 5036 13028 5040 13084
rect 4976 13024 5040 13028
rect 5056 13084 5120 13088
rect 5056 13028 5060 13084
rect 5060 13028 5116 13084
rect 5116 13028 5120 13084
rect 5056 13024 5120 13028
rect 6748 13084 6812 13088
rect 6748 13028 6752 13084
rect 6752 13028 6808 13084
rect 6808 13028 6812 13084
rect 6748 13024 6812 13028
rect 6828 13084 6892 13088
rect 6828 13028 6832 13084
rect 6832 13028 6888 13084
rect 6888 13028 6892 13084
rect 6828 13024 6892 13028
rect 6908 13084 6972 13088
rect 6908 13028 6912 13084
rect 6912 13028 6968 13084
rect 6968 13028 6972 13084
rect 6908 13024 6972 13028
rect 6988 13084 7052 13088
rect 6988 13028 6992 13084
rect 6992 13028 7048 13084
rect 7048 13028 7052 13084
rect 6988 13024 7052 13028
rect 8680 13084 8744 13088
rect 8680 13028 8684 13084
rect 8684 13028 8740 13084
rect 8740 13028 8744 13084
rect 8680 13024 8744 13028
rect 8760 13084 8824 13088
rect 8760 13028 8764 13084
rect 8764 13028 8820 13084
rect 8820 13028 8824 13084
rect 8760 13024 8824 13028
rect 8840 13084 8904 13088
rect 8840 13028 8844 13084
rect 8844 13028 8900 13084
rect 8900 13028 8904 13084
rect 8840 13024 8904 13028
rect 8920 13084 8984 13088
rect 8920 13028 8924 13084
rect 8924 13028 8980 13084
rect 8980 13028 8984 13084
rect 8920 13024 8984 13028
rect 1918 12540 1982 12544
rect 1918 12484 1922 12540
rect 1922 12484 1978 12540
rect 1978 12484 1982 12540
rect 1918 12480 1982 12484
rect 1998 12540 2062 12544
rect 1998 12484 2002 12540
rect 2002 12484 2058 12540
rect 2058 12484 2062 12540
rect 1998 12480 2062 12484
rect 2078 12540 2142 12544
rect 2078 12484 2082 12540
rect 2082 12484 2138 12540
rect 2138 12484 2142 12540
rect 2078 12480 2142 12484
rect 2158 12540 2222 12544
rect 2158 12484 2162 12540
rect 2162 12484 2218 12540
rect 2218 12484 2222 12540
rect 2158 12480 2222 12484
rect 3850 12540 3914 12544
rect 3850 12484 3854 12540
rect 3854 12484 3910 12540
rect 3910 12484 3914 12540
rect 3850 12480 3914 12484
rect 3930 12540 3994 12544
rect 3930 12484 3934 12540
rect 3934 12484 3990 12540
rect 3990 12484 3994 12540
rect 3930 12480 3994 12484
rect 4010 12540 4074 12544
rect 4010 12484 4014 12540
rect 4014 12484 4070 12540
rect 4070 12484 4074 12540
rect 4010 12480 4074 12484
rect 4090 12540 4154 12544
rect 4090 12484 4094 12540
rect 4094 12484 4150 12540
rect 4150 12484 4154 12540
rect 4090 12480 4154 12484
rect 5782 12540 5846 12544
rect 5782 12484 5786 12540
rect 5786 12484 5842 12540
rect 5842 12484 5846 12540
rect 5782 12480 5846 12484
rect 5862 12540 5926 12544
rect 5862 12484 5866 12540
rect 5866 12484 5922 12540
rect 5922 12484 5926 12540
rect 5862 12480 5926 12484
rect 5942 12540 6006 12544
rect 5942 12484 5946 12540
rect 5946 12484 6002 12540
rect 6002 12484 6006 12540
rect 5942 12480 6006 12484
rect 6022 12540 6086 12544
rect 6022 12484 6026 12540
rect 6026 12484 6082 12540
rect 6082 12484 6086 12540
rect 6022 12480 6086 12484
rect 7714 12540 7778 12544
rect 7714 12484 7718 12540
rect 7718 12484 7774 12540
rect 7774 12484 7778 12540
rect 7714 12480 7778 12484
rect 7794 12540 7858 12544
rect 7794 12484 7798 12540
rect 7798 12484 7854 12540
rect 7854 12484 7858 12540
rect 7794 12480 7858 12484
rect 7874 12540 7938 12544
rect 7874 12484 7878 12540
rect 7878 12484 7934 12540
rect 7934 12484 7938 12540
rect 7874 12480 7938 12484
rect 7954 12540 8018 12544
rect 7954 12484 7958 12540
rect 7958 12484 8014 12540
rect 8014 12484 8018 12540
rect 7954 12480 8018 12484
rect 2884 11996 2948 12000
rect 2884 11940 2888 11996
rect 2888 11940 2944 11996
rect 2944 11940 2948 11996
rect 2884 11936 2948 11940
rect 2964 11996 3028 12000
rect 2964 11940 2968 11996
rect 2968 11940 3024 11996
rect 3024 11940 3028 11996
rect 2964 11936 3028 11940
rect 3044 11996 3108 12000
rect 3044 11940 3048 11996
rect 3048 11940 3104 11996
rect 3104 11940 3108 11996
rect 3044 11936 3108 11940
rect 3124 11996 3188 12000
rect 3124 11940 3128 11996
rect 3128 11940 3184 11996
rect 3184 11940 3188 11996
rect 3124 11936 3188 11940
rect 4816 11996 4880 12000
rect 4816 11940 4820 11996
rect 4820 11940 4876 11996
rect 4876 11940 4880 11996
rect 4816 11936 4880 11940
rect 4896 11996 4960 12000
rect 4896 11940 4900 11996
rect 4900 11940 4956 11996
rect 4956 11940 4960 11996
rect 4896 11936 4960 11940
rect 4976 11996 5040 12000
rect 4976 11940 4980 11996
rect 4980 11940 5036 11996
rect 5036 11940 5040 11996
rect 4976 11936 5040 11940
rect 5056 11996 5120 12000
rect 5056 11940 5060 11996
rect 5060 11940 5116 11996
rect 5116 11940 5120 11996
rect 5056 11936 5120 11940
rect 6748 11996 6812 12000
rect 6748 11940 6752 11996
rect 6752 11940 6808 11996
rect 6808 11940 6812 11996
rect 6748 11936 6812 11940
rect 6828 11996 6892 12000
rect 6828 11940 6832 11996
rect 6832 11940 6888 11996
rect 6888 11940 6892 11996
rect 6828 11936 6892 11940
rect 6908 11996 6972 12000
rect 6908 11940 6912 11996
rect 6912 11940 6968 11996
rect 6968 11940 6972 11996
rect 6908 11936 6972 11940
rect 6988 11996 7052 12000
rect 6988 11940 6992 11996
rect 6992 11940 7048 11996
rect 7048 11940 7052 11996
rect 6988 11936 7052 11940
rect 8680 11996 8744 12000
rect 8680 11940 8684 11996
rect 8684 11940 8740 11996
rect 8740 11940 8744 11996
rect 8680 11936 8744 11940
rect 8760 11996 8824 12000
rect 8760 11940 8764 11996
rect 8764 11940 8820 11996
rect 8820 11940 8824 11996
rect 8760 11936 8824 11940
rect 8840 11996 8904 12000
rect 8840 11940 8844 11996
rect 8844 11940 8900 11996
rect 8900 11940 8904 11996
rect 8840 11936 8904 11940
rect 8920 11996 8984 12000
rect 8920 11940 8924 11996
rect 8924 11940 8980 11996
rect 8980 11940 8984 11996
rect 8920 11936 8984 11940
rect 1918 11452 1982 11456
rect 1918 11396 1922 11452
rect 1922 11396 1978 11452
rect 1978 11396 1982 11452
rect 1918 11392 1982 11396
rect 1998 11452 2062 11456
rect 1998 11396 2002 11452
rect 2002 11396 2058 11452
rect 2058 11396 2062 11452
rect 1998 11392 2062 11396
rect 2078 11452 2142 11456
rect 2078 11396 2082 11452
rect 2082 11396 2138 11452
rect 2138 11396 2142 11452
rect 2078 11392 2142 11396
rect 2158 11452 2222 11456
rect 2158 11396 2162 11452
rect 2162 11396 2218 11452
rect 2218 11396 2222 11452
rect 2158 11392 2222 11396
rect 3850 11452 3914 11456
rect 3850 11396 3854 11452
rect 3854 11396 3910 11452
rect 3910 11396 3914 11452
rect 3850 11392 3914 11396
rect 3930 11452 3994 11456
rect 3930 11396 3934 11452
rect 3934 11396 3990 11452
rect 3990 11396 3994 11452
rect 3930 11392 3994 11396
rect 4010 11452 4074 11456
rect 4010 11396 4014 11452
rect 4014 11396 4070 11452
rect 4070 11396 4074 11452
rect 4010 11392 4074 11396
rect 4090 11452 4154 11456
rect 4090 11396 4094 11452
rect 4094 11396 4150 11452
rect 4150 11396 4154 11452
rect 4090 11392 4154 11396
rect 5782 11452 5846 11456
rect 5782 11396 5786 11452
rect 5786 11396 5842 11452
rect 5842 11396 5846 11452
rect 5782 11392 5846 11396
rect 5862 11452 5926 11456
rect 5862 11396 5866 11452
rect 5866 11396 5922 11452
rect 5922 11396 5926 11452
rect 5862 11392 5926 11396
rect 5942 11452 6006 11456
rect 5942 11396 5946 11452
rect 5946 11396 6002 11452
rect 6002 11396 6006 11452
rect 5942 11392 6006 11396
rect 6022 11452 6086 11456
rect 6022 11396 6026 11452
rect 6026 11396 6082 11452
rect 6082 11396 6086 11452
rect 6022 11392 6086 11396
rect 7714 11452 7778 11456
rect 7714 11396 7718 11452
rect 7718 11396 7774 11452
rect 7774 11396 7778 11452
rect 7714 11392 7778 11396
rect 7794 11452 7858 11456
rect 7794 11396 7798 11452
rect 7798 11396 7854 11452
rect 7854 11396 7858 11452
rect 7794 11392 7858 11396
rect 7874 11452 7938 11456
rect 7874 11396 7878 11452
rect 7878 11396 7934 11452
rect 7934 11396 7938 11452
rect 7874 11392 7938 11396
rect 7954 11452 8018 11456
rect 7954 11396 7958 11452
rect 7958 11396 8014 11452
rect 8014 11396 8018 11452
rect 7954 11392 8018 11396
rect 2884 10908 2948 10912
rect 2884 10852 2888 10908
rect 2888 10852 2944 10908
rect 2944 10852 2948 10908
rect 2884 10848 2948 10852
rect 2964 10908 3028 10912
rect 2964 10852 2968 10908
rect 2968 10852 3024 10908
rect 3024 10852 3028 10908
rect 2964 10848 3028 10852
rect 3044 10908 3108 10912
rect 3044 10852 3048 10908
rect 3048 10852 3104 10908
rect 3104 10852 3108 10908
rect 3044 10848 3108 10852
rect 3124 10908 3188 10912
rect 3124 10852 3128 10908
rect 3128 10852 3184 10908
rect 3184 10852 3188 10908
rect 3124 10848 3188 10852
rect 4816 10908 4880 10912
rect 4816 10852 4820 10908
rect 4820 10852 4876 10908
rect 4876 10852 4880 10908
rect 4816 10848 4880 10852
rect 4896 10908 4960 10912
rect 4896 10852 4900 10908
rect 4900 10852 4956 10908
rect 4956 10852 4960 10908
rect 4896 10848 4960 10852
rect 4976 10908 5040 10912
rect 4976 10852 4980 10908
rect 4980 10852 5036 10908
rect 5036 10852 5040 10908
rect 4976 10848 5040 10852
rect 5056 10908 5120 10912
rect 5056 10852 5060 10908
rect 5060 10852 5116 10908
rect 5116 10852 5120 10908
rect 5056 10848 5120 10852
rect 6748 10908 6812 10912
rect 6748 10852 6752 10908
rect 6752 10852 6808 10908
rect 6808 10852 6812 10908
rect 6748 10848 6812 10852
rect 6828 10908 6892 10912
rect 6828 10852 6832 10908
rect 6832 10852 6888 10908
rect 6888 10852 6892 10908
rect 6828 10848 6892 10852
rect 6908 10908 6972 10912
rect 6908 10852 6912 10908
rect 6912 10852 6968 10908
rect 6968 10852 6972 10908
rect 6908 10848 6972 10852
rect 6988 10908 7052 10912
rect 6988 10852 6992 10908
rect 6992 10852 7048 10908
rect 7048 10852 7052 10908
rect 6988 10848 7052 10852
rect 8680 10908 8744 10912
rect 8680 10852 8684 10908
rect 8684 10852 8740 10908
rect 8740 10852 8744 10908
rect 8680 10848 8744 10852
rect 8760 10908 8824 10912
rect 8760 10852 8764 10908
rect 8764 10852 8820 10908
rect 8820 10852 8824 10908
rect 8760 10848 8824 10852
rect 8840 10908 8904 10912
rect 8840 10852 8844 10908
rect 8844 10852 8900 10908
rect 8900 10852 8904 10908
rect 8840 10848 8904 10852
rect 8920 10908 8984 10912
rect 8920 10852 8924 10908
rect 8924 10852 8980 10908
rect 8980 10852 8984 10908
rect 8920 10848 8984 10852
rect 1918 10364 1982 10368
rect 1918 10308 1922 10364
rect 1922 10308 1978 10364
rect 1978 10308 1982 10364
rect 1918 10304 1982 10308
rect 1998 10364 2062 10368
rect 1998 10308 2002 10364
rect 2002 10308 2058 10364
rect 2058 10308 2062 10364
rect 1998 10304 2062 10308
rect 2078 10364 2142 10368
rect 2078 10308 2082 10364
rect 2082 10308 2138 10364
rect 2138 10308 2142 10364
rect 2078 10304 2142 10308
rect 2158 10364 2222 10368
rect 2158 10308 2162 10364
rect 2162 10308 2218 10364
rect 2218 10308 2222 10364
rect 2158 10304 2222 10308
rect 3850 10364 3914 10368
rect 3850 10308 3854 10364
rect 3854 10308 3910 10364
rect 3910 10308 3914 10364
rect 3850 10304 3914 10308
rect 3930 10364 3994 10368
rect 3930 10308 3934 10364
rect 3934 10308 3990 10364
rect 3990 10308 3994 10364
rect 3930 10304 3994 10308
rect 4010 10364 4074 10368
rect 4010 10308 4014 10364
rect 4014 10308 4070 10364
rect 4070 10308 4074 10364
rect 4010 10304 4074 10308
rect 4090 10364 4154 10368
rect 4090 10308 4094 10364
rect 4094 10308 4150 10364
rect 4150 10308 4154 10364
rect 4090 10304 4154 10308
rect 5782 10364 5846 10368
rect 5782 10308 5786 10364
rect 5786 10308 5842 10364
rect 5842 10308 5846 10364
rect 5782 10304 5846 10308
rect 5862 10364 5926 10368
rect 5862 10308 5866 10364
rect 5866 10308 5922 10364
rect 5922 10308 5926 10364
rect 5862 10304 5926 10308
rect 5942 10364 6006 10368
rect 5942 10308 5946 10364
rect 5946 10308 6002 10364
rect 6002 10308 6006 10364
rect 5942 10304 6006 10308
rect 6022 10364 6086 10368
rect 6022 10308 6026 10364
rect 6026 10308 6082 10364
rect 6082 10308 6086 10364
rect 6022 10304 6086 10308
rect 7714 10364 7778 10368
rect 7714 10308 7718 10364
rect 7718 10308 7774 10364
rect 7774 10308 7778 10364
rect 7714 10304 7778 10308
rect 7794 10364 7858 10368
rect 7794 10308 7798 10364
rect 7798 10308 7854 10364
rect 7854 10308 7858 10364
rect 7794 10304 7858 10308
rect 7874 10364 7938 10368
rect 7874 10308 7878 10364
rect 7878 10308 7934 10364
rect 7934 10308 7938 10364
rect 7874 10304 7938 10308
rect 7954 10364 8018 10368
rect 7954 10308 7958 10364
rect 7958 10308 8014 10364
rect 8014 10308 8018 10364
rect 7954 10304 8018 10308
rect 2884 9820 2948 9824
rect 2884 9764 2888 9820
rect 2888 9764 2944 9820
rect 2944 9764 2948 9820
rect 2884 9760 2948 9764
rect 2964 9820 3028 9824
rect 2964 9764 2968 9820
rect 2968 9764 3024 9820
rect 3024 9764 3028 9820
rect 2964 9760 3028 9764
rect 3044 9820 3108 9824
rect 3044 9764 3048 9820
rect 3048 9764 3104 9820
rect 3104 9764 3108 9820
rect 3044 9760 3108 9764
rect 3124 9820 3188 9824
rect 3124 9764 3128 9820
rect 3128 9764 3184 9820
rect 3184 9764 3188 9820
rect 3124 9760 3188 9764
rect 4816 9820 4880 9824
rect 4816 9764 4820 9820
rect 4820 9764 4876 9820
rect 4876 9764 4880 9820
rect 4816 9760 4880 9764
rect 4896 9820 4960 9824
rect 4896 9764 4900 9820
rect 4900 9764 4956 9820
rect 4956 9764 4960 9820
rect 4896 9760 4960 9764
rect 4976 9820 5040 9824
rect 4976 9764 4980 9820
rect 4980 9764 5036 9820
rect 5036 9764 5040 9820
rect 4976 9760 5040 9764
rect 5056 9820 5120 9824
rect 5056 9764 5060 9820
rect 5060 9764 5116 9820
rect 5116 9764 5120 9820
rect 5056 9760 5120 9764
rect 6748 9820 6812 9824
rect 6748 9764 6752 9820
rect 6752 9764 6808 9820
rect 6808 9764 6812 9820
rect 6748 9760 6812 9764
rect 6828 9820 6892 9824
rect 6828 9764 6832 9820
rect 6832 9764 6888 9820
rect 6888 9764 6892 9820
rect 6828 9760 6892 9764
rect 6908 9820 6972 9824
rect 6908 9764 6912 9820
rect 6912 9764 6968 9820
rect 6968 9764 6972 9820
rect 6908 9760 6972 9764
rect 6988 9820 7052 9824
rect 6988 9764 6992 9820
rect 6992 9764 7048 9820
rect 7048 9764 7052 9820
rect 6988 9760 7052 9764
rect 8680 9820 8744 9824
rect 8680 9764 8684 9820
rect 8684 9764 8740 9820
rect 8740 9764 8744 9820
rect 8680 9760 8744 9764
rect 8760 9820 8824 9824
rect 8760 9764 8764 9820
rect 8764 9764 8820 9820
rect 8820 9764 8824 9820
rect 8760 9760 8824 9764
rect 8840 9820 8904 9824
rect 8840 9764 8844 9820
rect 8844 9764 8900 9820
rect 8900 9764 8904 9820
rect 8840 9760 8904 9764
rect 8920 9820 8984 9824
rect 8920 9764 8924 9820
rect 8924 9764 8980 9820
rect 8980 9764 8984 9820
rect 8920 9760 8984 9764
rect 1918 9276 1982 9280
rect 1918 9220 1922 9276
rect 1922 9220 1978 9276
rect 1978 9220 1982 9276
rect 1918 9216 1982 9220
rect 1998 9276 2062 9280
rect 1998 9220 2002 9276
rect 2002 9220 2058 9276
rect 2058 9220 2062 9276
rect 1998 9216 2062 9220
rect 2078 9276 2142 9280
rect 2078 9220 2082 9276
rect 2082 9220 2138 9276
rect 2138 9220 2142 9276
rect 2078 9216 2142 9220
rect 2158 9276 2222 9280
rect 2158 9220 2162 9276
rect 2162 9220 2218 9276
rect 2218 9220 2222 9276
rect 2158 9216 2222 9220
rect 3850 9276 3914 9280
rect 3850 9220 3854 9276
rect 3854 9220 3910 9276
rect 3910 9220 3914 9276
rect 3850 9216 3914 9220
rect 3930 9276 3994 9280
rect 3930 9220 3934 9276
rect 3934 9220 3990 9276
rect 3990 9220 3994 9276
rect 3930 9216 3994 9220
rect 4010 9276 4074 9280
rect 4010 9220 4014 9276
rect 4014 9220 4070 9276
rect 4070 9220 4074 9276
rect 4010 9216 4074 9220
rect 4090 9276 4154 9280
rect 4090 9220 4094 9276
rect 4094 9220 4150 9276
rect 4150 9220 4154 9276
rect 4090 9216 4154 9220
rect 5782 9276 5846 9280
rect 5782 9220 5786 9276
rect 5786 9220 5842 9276
rect 5842 9220 5846 9276
rect 5782 9216 5846 9220
rect 5862 9276 5926 9280
rect 5862 9220 5866 9276
rect 5866 9220 5922 9276
rect 5922 9220 5926 9276
rect 5862 9216 5926 9220
rect 5942 9276 6006 9280
rect 5942 9220 5946 9276
rect 5946 9220 6002 9276
rect 6002 9220 6006 9276
rect 5942 9216 6006 9220
rect 6022 9276 6086 9280
rect 6022 9220 6026 9276
rect 6026 9220 6082 9276
rect 6082 9220 6086 9276
rect 6022 9216 6086 9220
rect 7714 9276 7778 9280
rect 7714 9220 7718 9276
rect 7718 9220 7774 9276
rect 7774 9220 7778 9276
rect 7714 9216 7778 9220
rect 7794 9276 7858 9280
rect 7794 9220 7798 9276
rect 7798 9220 7854 9276
rect 7854 9220 7858 9276
rect 7794 9216 7858 9220
rect 7874 9276 7938 9280
rect 7874 9220 7878 9276
rect 7878 9220 7934 9276
rect 7934 9220 7938 9276
rect 7874 9216 7938 9220
rect 7954 9276 8018 9280
rect 7954 9220 7958 9276
rect 7958 9220 8014 9276
rect 8014 9220 8018 9276
rect 7954 9216 8018 9220
rect 2884 8732 2948 8736
rect 2884 8676 2888 8732
rect 2888 8676 2944 8732
rect 2944 8676 2948 8732
rect 2884 8672 2948 8676
rect 2964 8732 3028 8736
rect 2964 8676 2968 8732
rect 2968 8676 3024 8732
rect 3024 8676 3028 8732
rect 2964 8672 3028 8676
rect 3044 8732 3108 8736
rect 3044 8676 3048 8732
rect 3048 8676 3104 8732
rect 3104 8676 3108 8732
rect 3044 8672 3108 8676
rect 3124 8732 3188 8736
rect 3124 8676 3128 8732
rect 3128 8676 3184 8732
rect 3184 8676 3188 8732
rect 3124 8672 3188 8676
rect 4816 8732 4880 8736
rect 4816 8676 4820 8732
rect 4820 8676 4876 8732
rect 4876 8676 4880 8732
rect 4816 8672 4880 8676
rect 4896 8732 4960 8736
rect 4896 8676 4900 8732
rect 4900 8676 4956 8732
rect 4956 8676 4960 8732
rect 4896 8672 4960 8676
rect 4976 8732 5040 8736
rect 4976 8676 4980 8732
rect 4980 8676 5036 8732
rect 5036 8676 5040 8732
rect 4976 8672 5040 8676
rect 5056 8732 5120 8736
rect 5056 8676 5060 8732
rect 5060 8676 5116 8732
rect 5116 8676 5120 8732
rect 5056 8672 5120 8676
rect 6748 8732 6812 8736
rect 6748 8676 6752 8732
rect 6752 8676 6808 8732
rect 6808 8676 6812 8732
rect 6748 8672 6812 8676
rect 6828 8732 6892 8736
rect 6828 8676 6832 8732
rect 6832 8676 6888 8732
rect 6888 8676 6892 8732
rect 6828 8672 6892 8676
rect 6908 8732 6972 8736
rect 6908 8676 6912 8732
rect 6912 8676 6968 8732
rect 6968 8676 6972 8732
rect 6908 8672 6972 8676
rect 6988 8732 7052 8736
rect 6988 8676 6992 8732
rect 6992 8676 7048 8732
rect 7048 8676 7052 8732
rect 6988 8672 7052 8676
rect 8680 8732 8744 8736
rect 8680 8676 8684 8732
rect 8684 8676 8740 8732
rect 8740 8676 8744 8732
rect 8680 8672 8744 8676
rect 8760 8732 8824 8736
rect 8760 8676 8764 8732
rect 8764 8676 8820 8732
rect 8820 8676 8824 8732
rect 8760 8672 8824 8676
rect 8840 8732 8904 8736
rect 8840 8676 8844 8732
rect 8844 8676 8900 8732
rect 8900 8676 8904 8732
rect 8840 8672 8904 8676
rect 8920 8732 8984 8736
rect 8920 8676 8924 8732
rect 8924 8676 8980 8732
rect 8980 8676 8984 8732
rect 8920 8672 8984 8676
rect 1918 8188 1982 8192
rect 1918 8132 1922 8188
rect 1922 8132 1978 8188
rect 1978 8132 1982 8188
rect 1918 8128 1982 8132
rect 1998 8188 2062 8192
rect 1998 8132 2002 8188
rect 2002 8132 2058 8188
rect 2058 8132 2062 8188
rect 1998 8128 2062 8132
rect 2078 8188 2142 8192
rect 2078 8132 2082 8188
rect 2082 8132 2138 8188
rect 2138 8132 2142 8188
rect 2078 8128 2142 8132
rect 2158 8188 2222 8192
rect 2158 8132 2162 8188
rect 2162 8132 2218 8188
rect 2218 8132 2222 8188
rect 2158 8128 2222 8132
rect 3850 8188 3914 8192
rect 3850 8132 3854 8188
rect 3854 8132 3910 8188
rect 3910 8132 3914 8188
rect 3850 8128 3914 8132
rect 3930 8188 3994 8192
rect 3930 8132 3934 8188
rect 3934 8132 3990 8188
rect 3990 8132 3994 8188
rect 3930 8128 3994 8132
rect 4010 8188 4074 8192
rect 4010 8132 4014 8188
rect 4014 8132 4070 8188
rect 4070 8132 4074 8188
rect 4010 8128 4074 8132
rect 4090 8188 4154 8192
rect 4090 8132 4094 8188
rect 4094 8132 4150 8188
rect 4150 8132 4154 8188
rect 4090 8128 4154 8132
rect 5782 8188 5846 8192
rect 5782 8132 5786 8188
rect 5786 8132 5842 8188
rect 5842 8132 5846 8188
rect 5782 8128 5846 8132
rect 5862 8188 5926 8192
rect 5862 8132 5866 8188
rect 5866 8132 5922 8188
rect 5922 8132 5926 8188
rect 5862 8128 5926 8132
rect 5942 8188 6006 8192
rect 5942 8132 5946 8188
rect 5946 8132 6002 8188
rect 6002 8132 6006 8188
rect 5942 8128 6006 8132
rect 6022 8188 6086 8192
rect 6022 8132 6026 8188
rect 6026 8132 6082 8188
rect 6082 8132 6086 8188
rect 6022 8128 6086 8132
rect 7714 8188 7778 8192
rect 7714 8132 7718 8188
rect 7718 8132 7774 8188
rect 7774 8132 7778 8188
rect 7714 8128 7778 8132
rect 7794 8188 7858 8192
rect 7794 8132 7798 8188
rect 7798 8132 7854 8188
rect 7854 8132 7858 8188
rect 7794 8128 7858 8132
rect 7874 8188 7938 8192
rect 7874 8132 7878 8188
rect 7878 8132 7934 8188
rect 7934 8132 7938 8188
rect 7874 8128 7938 8132
rect 7954 8188 8018 8192
rect 7954 8132 7958 8188
rect 7958 8132 8014 8188
rect 8014 8132 8018 8188
rect 7954 8128 8018 8132
rect 2884 7644 2948 7648
rect 2884 7588 2888 7644
rect 2888 7588 2944 7644
rect 2944 7588 2948 7644
rect 2884 7584 2948 7588
rect 2964 7644 3028 7648
rect 2964 7588 2968 7644
rect 2968 7588 3024 7644
rect 3024 7588 3028 7644
rect 2964 7584 3028 7588
rect 3044 7644 3108 7648
rect 3044 7588 3048 7644
rect 3048 7588 3104 7644
rect 3104 7588 3108 7644
rect 3044 7584 3108 7588
rect 3124 7644 3188 7648
rect 3124 7588 3128 7644
rect 3128 7588 3184 7644
rect 3184 7588 3188 7644
rect 3124 7584 3188 7588
rect 4816 7644 4880 7648
rect 4816 7588 4820 7644
rect 4820 7588 4876 7644
rect 4876 7588 4880 7644
rect 4816 7584 4880 7588
rect 4896 7644 4960 7648
rect 4896 7588 4900 7644
rect 4900 7588 4956 7644
rect 4956 7588 4960 7644
rect 4896 7584 4960 7588
rect 4976 7644 5040 7648
rect 4976 7588 4980 7644
rect 4980 7588 5036 7644
rect 5036 7588 5040 7644
rect 4976 7584 5040 7588
rect 5056 7644 5120 7648
rect 5056 7588 5060 7644
rect 5060 7588 5116 7644
rect 5116 7588 5120 7644
rect 5056 7584 5120 7588
rect 6748 7644 6812 7648
rect 6748 7588 6752 7644
rect 6752 7588 6808 7644
rect 6808 7588 6812 7644
rect 6748 7584 6812 7588
rect 6828 7644 6892 7648
rect 6828 7588 6832 7644
rect 6832 7588 6888 7644
rect 6888 7588 6892 7644
rect 6828 7584 6892 7588
rect 6908 7644 6972 7648
rect 6908 7588 6912 7644
rect 6912 7588 6968 7644
rect 6968 7588 6972 7644
rect 6908 7584 6972 7588
rect 6988 7644 7052 7648
rect 6988 7588 6992 7644
rect 6992 7588 7048 7644
rect 7048 7588 7052 7644
rect 6988 7584 7052 7588
rect 8680 7644 8744 7648
rect 8680 7588 8684 7644
rect 8684 7588 8740 7644
rect 8740 7588 8744 7644
rect 8680 7584 8744 7588
rect 8760 7644 8824 7648
rect 8760 7588 8764 7644
rect 8764 7588 8820 7644
rect 8820 7588 8824 7644
rect 8760 7584 8824 7588
rect 8840 7644 8904 7648
rect 8840 7588 8844 7644
rect 8844 7588 8900 7644
rect 8900 7588 8904 7644
rect 8840 7584 8904 7588
rect 8920 7644 8984 7648
rect 8920 7588 8924 7644
rect 8924 7588 8980 7644
rect 8980 7588 8984 7644
rect 8920 7584 8984 7588
rect 1918 7100 1982 7104
rect 1918 7044 1922 7100
rect 1922 7044 1978 7100
rect 1978 7044 1982 7100
rect 1918 7040 1982 7044
rect 1998 7100 2062 7104
rect 1998 7044 2002 7100
rect 2002 7044 2058 7100
rect 2058 7044 2062 7100
rect 1998 7040 2062 7044
rect 2078 7100 2142 7104
rect 2078 7044 2082 7100
rect 2082 7044 2138 7100
rect 2138 7044 2142 7100
rect 2078 7040 2142 7044
rect 2158 7100 2222 7104
rect 2158 7044 2162 7100
rect 2162 7044 2218 7100
rect 2218 7044 2222 7100
rect 2158 7040 2222 7044
rect 3850 7100 3914 7104
rect 3850 7044 3854 7100
rect 3854 7044 3910 7100
rect 3910 7044 3914 7100
rect 3850 7040 3914 7044
rect 3930 7100 3994 7104
rect 3930 7044 3934 7100
rect 3934 7044 3990 7100
rect 3990 7044 3994 7100
rect 3930 7040 3994 7044
rect 4010 7100 4074 7104
rect 4010 7044 4014 7100
rect 4014 7044 4070 7100
rect 4070 7044 4074 7100
rect 4010 7040 4074 7044
rect 4090 7100 4154 7104
rect 4090 7044 4094 7100
rect 4094 7044 4150 7100
rect 4150 7044 4154 7100
rect 4090 7040 4154 7044
rect 5782 7100 5846 7104
rect 5782 7044 5786 7100
rect 5786 7044 5842 7100
rect 5842 7044 5846 7100
rect 5782 7040 5846 7044
rect 5862 7100 5926 7104
rect 5862 7044 5866 7100
rect 5866 7044 5922 7100
rect 5922 7044 5926 7100
rect 5862 7040 5926 7044
rect 5942 7100 6006 7104
rect 5942 7044 5946 7100
rect 5946 7044 6002 7100
rect 6002 7044 6006 7100
rect 5942 7040 6006 7044
rect 6022 7100 6086 7104
rect 6022 7044 6026 7100
rect 6026 7044 6082 7100
rect 6082 7044 6086 7100
rect 6022 7040 6086 7044
rect 7714 7100 7778 7104
rect 7714 7044 7718 7100
rect 7718 7044 7774 7100
rect 7774 7044 7778 7100
rect 7714 7040 7778 7044
rect 7794 7100 7858 7104
rect 7794 7044 7798 7100
rect 7798 7044 7854 7100
rect 7854 7044 7858 7100
rect 7794 7040 7858 7044
rect 7874 7100 7938 7104
rect 7874 7044 7878 7100
rect 7878 7044 7934 7100
rect 7934 7044 7938 7100
rect 7874 7040 7938 7044
rect 7954 7100 8018 7104
rect 7954 7044 7958 7100
rect 7958 7044 8014 7100
rect 8014 7044 8018 7100
rect 7954 7040 8018 7044
rect 2884 6556 2948 6560
rect 2884 6500 2888 6556
rect 2888 6500 2944 6556
rect 2944 6500 2948 6556
rect 2884 6496 2948 6500
rect 2964 6556 3028 6560
rect 2964 6500 2968 6556
rect 2968 6500 3024 6556
rect 3024 6500 3028 6556
rect 2964 6496 3028 6500
rect 3044 6556 3108 6560
rect 3044 6500 3048 6556
rect 3048 6500 3104 6556
rect 3104 6500 3108 6556
rect 3044 6496 3108 6500
rect 3124 6556 3188 6560
rect 3124 6500 3128 6556
rect 3128 6500 3184 6556
rect 3184 6500 3188 6556
rect 3124 6496 3188 6500
rect 4816 6556 4880 6560
rect 4816 6500 4820 6556
rect 4820 6500 4876 6556
rect 4876 6500 4880 6556
rect 4816 6496 4880 6500
rect 4896 6556 4960 6560
rect 4896 6500 4900 6556
rect 4900 6500 4956 6556
rect 4956 6500 4960 6556
rect 4896 6496 4960 6500
rect 4976 6556 5040 6560
rect 4976 6500 4980 6556
rect 4980 6500 5036 6556
rect 5036 6500 5040 6556
rect 4976 6496 5040 6500
rect 5056 6556 5120 6560
rect 5056 6500 5060 6556
rect 5060 6500 5116 6556
rect 5116 6500 5120 6556
rect 5056 6496 5120 6500
rect 6748 6556 6812 6560
rect 6748 6500 6752 6556
rect 6752 6500 6808 6556
rect 6808 6500 6812 6556
rect 6748 6496 6812 6500
rect 6828 6556 6892 6560
rect 6828 6500 6832 6556
rect 6832 6500 6888 6556
rect 6888 6500 6892 6556
rect 6828 6496 6892 6500
rect 6908 6556 6972 6560
rect 6908 6500 6912 6556
rect 6912 6500 6968 6556
rect 6968 6500 6972 6556
rect 6908 6496 6972 6500
rect 6988 6556 7052 6560
rect 6988 6500 6992 6556
rect 6992 6500 7048 6556
rect 7048 6500 7052 6556
rect 6988 6496 7052 6500
rect 8680 6556 8744 6560
rect 8680 6500 8684 6556
rect 8684 6500 8740 6556
rect 8740 6500 8744 6556
rect 8680 6496 8744 6500
rect 8760 6556 8824 6560
rect 8760 6500 8764 6556
rect 8764 6500 8820 6556
rect 8820 6500 8824 6556
rect 8760 6496 8824 6500
rect 8840 6556 8904 6560
rect 8840 6500 8844 6556
rect 8844 6500 8900 6556
rect 8900 6500 8904 6556
rect 8840 6496 8904 6500
rect 8920 6556 8984 6560
rect 8920 6500 8924 6556
rect 8924 6500 8980 6556
rect 8980 6500 8984 6556
rect 8920 6496 8984 6500
rect 1918 6012 1982 6016
rect 1918 5956 1922 6012
rect 1922 5956 1978 6012
rect 1978 5956 1982 6012
rect 1918 5952 1982 5956
rect 1998 6012 2062 6016
rect 1998 5956 2002 6012
rect 2002 5956 2058 6012
rect 2058 5956 2062 6012
rect 1998 5952 2062 5956
rect 2078 6012 2142 6016
rect 2078 5956 2082 6012
rect 2082 5956 2138 6012
rect 2138 5956 2142 6012
rect 2078 5952 2142 5956
rect 2158 6012 2222 6016
rect 2158 5956 2162 6012
rect 2162 5956 2218 6012
rect 2218 5956 2222 6012
rect 2158 5952 2222 5956
rect 3850 6012 3914 6016
rect 3850 5956 3854 6012
rect 3854 5956 3910 6012
rect 3910 5956 3914 6012
rect 3850 5952 3914 5956
rect 3930 6012 3994 6016
rect 3930 5956 3934 6012
rect 3934 5956 3990 6012
rect 3990 5956 3994 6012
rect 3930 5952 3994 5956
rect 4010 6012 4074 6016
rect 4010 5956 4014 6012
rect 4014 5956 4070 6012
rect 4070 5956 4074 6012
rect 4010 5952 4074 5956
rect 4090 6012 4154 6016
rect 4090 5956 4094 6012
rect 4094 5956 4150 6012
rect 4150 5956 4154 6012
rect 4090 5952 4154 5956
rect 5782 6012 5846 6016
rect 5782 5956 5786 6012
rect 5786 5956 5842 6012
rect 5842 5956 5846 6012
rect 5782 5952 5846 5956
rect 5862 6012 5926 6016
rect 5862 5956 5866 6012
rect 5866 5956 5922 6012
rect 5922 5956 5926 6012
rect 5862 5952 5926 5956
rect 5942 6012 6006 6016
rect 5942 5956 5946 6012
rect 5946 5956 6002 6012
rect 6002 5956 6006 6012
rect 5942 5952 6006 5956
rect 6022 6012 6086 6016
rect 6022 5956 6026 6012
rect 6026 5956 6082 6012
rect 6082 5956 6086 6012
rect 6022 5952 6086 5956
rect 7714 6012 7778 6016
rect 7714 5956 7718 6012
rect 7718 5956 7774 6012
rect 7774 5956 7778 6012
rect 7714 5952 7778 5956
rect 7794 6012 7858 6016
rect 7794 5956 7798 6012
rect 7798 5956 7854 6012
rect 7854 5956 7858 6012
rect 7794 5952 7858 5956
rect 7874 6012 7938 6016
rect 7874 5956 7878 6012
rect 7878 5956 7934 6012
rect 7934 5956 7938 6012
rect 7874 5952 7938 5956
rect 7954 6012 8018 6016
rect 7954 5956 7958 6012
rect 7958 5956 8014 6012
rect 8014 5956 8018 6012
rect 7954 5952 8018 5956
rect 2884 5468 2948 5472
rect 2884 5412 2888 5468
rect 2888 5412 2944 5468
rect 2944 5412 2948 5468
rect 2884 5408 2948 5412
rect 2964 5468 3028 5472
rect 2964 5412 2968 5468
rect 2968 5412 3024 5468
rect 3024 5412 3028 5468
rect 2964 5408 3028 5412
rect 3044 5468 3108 5472
rect 3044 5412 3048 5468
rect 3048 5412 3104 5468
rect 3104 5412 3108 5468
rect 3044 5408 3108 5412
rect 3124 5468 3188 5472
rect 3124 5412 3128 5468
rect 3128 5412 3184 5468
rect 3184 5412 3188 5468
rect 3124 5408 3188 5412
rect 4816 5468 4880 5472
rect 4816 5412 4820 5468
rect 4820 5412 4876 5468
rect 4876 5412 4880 5468
rect 4816 5408 4880 5412
rect 4896 5468 4960 5472
rect 4896 5412 4900 5468
rect 4900 5412 4956 5468
rect 4956 5412 4960 5468
rect 4896 5408 4960 5412
rect 4976 5468 5040 5472
rect 4976 5412 4980 5468
rect 4980 5412 5036 5468
rect 5036 5412 5040 5468
rect 4976 5408 5040 5412
rect 5056 5468 5120 5472
rect 5056 5412 5060 5468
rect 5060 5412 5116 5468
rect 5116 5412 5120 5468
rect 5056 5408 5120 5412
rect 6748 5468 6812 5472
rect 6748 5412 6752 5468
rect 6752 5412 6808 5468
rect 6808 5412 6812 5468
rect 6748 5408 6812 5412
rect 6828 5468 6892 5472
rect 6828 5412 6832 5468
rect 6832 5412 6888 5468
rect 6888 5412 6892 5468
rect 6828 5408 6892 5412
rect 6908 5468 6972 5472
rect 6908 5412 6912 5468
rect 6912 5412 6968 5468
rect 6968 5412 6972 5468
rect 6908 5408 6972 5412
rect 6988 5468 7052 5472
rect 6988 5412 6992 5468
rect 6992 5412 7048 5468
rect 7048 5412 7052 5468
rect 6988 5408 7052 5412
rect 8680 5468 8744 5472
rect 8680 5412 8684 5468
rect 8684 5412 8740 5468
rect 8740 5412 8744 5468
rect 8680 5408 8744 5412
rect 8760 5468 8824 5472
rect 8760 5412 8764 5468
rect 8764 5412 8820 5468
rect 8820 5412 8824 5468
rect 8760 5408 8824 5412
rect 8840 5468 8904 5472
rect 8840 5412 8844 5468
rect 8844 5412 8900 5468
rect 8900 5412 8904 5468
rect 8840 5408 8904 5412
rect 8920 5468 8984 5472
rect 8920 5412 8924 5468
rect 8924 5412 8980 5468
rect 8980 5412 8984 5468
rect 8920 5408 8984 5412
rect 1918 4924 1982 4928
rect 1918 4868 1922 4924
rect 1922 4868 1978 4924
rect 1978 4868 1982 4924
rect 1918 4864 1982 4868
rect 1998 4924 2062 4928
rect 1998 4868 2002 4924
rect 2002 4868 2058 4924
rect 2058 4868 2062 4924
rect 1998 4864 2062 4868
rect 2078 4924 2142 4928
rect 2078 4868 2082 4924
rect 2082 4868 2138 4924
rect 2138 4868 2142 4924
rect 2078 4864 2142 4868
rect 2158 4924 2222 4928
rect 2158 4868 2162 4924
rect 2162 4868 2218 4924
rect 2218 4868 2222 4924
rect 2158 4864 2222 4868
rect 3850 4924 3914 4928
rect 3850 4868 3854 4924
rect 3854 4868 3910 4924
rect 3910 4868 3914 4924
rect 3850 4864 3914 4868
rect 3930 4924 3994 4928
rect 3930 4868 3934 4924
rect 3934 4868 3990 4924
rect 3990 4868 3994 4924
rect 3930 4864 3994 4868
rect 4010 4924 4074 4928
rect 4010 4868 4014 4924
rect 4014 4868 4070 4924
rect 4070 4868 4074 4924
rect 4010 4864 4074 4868
rect 4090 4924 4154 4928
rect 4090 4868 4094 4924
rect 4094 4868 4150 4924
rect 4150 4868 4154 4924
rect 4090 4864 4154 4868
rect 5782 4924 5846 4928
rect 5782 4868 5786 4924
rect 5786 4868 5842 4924
rect 5842 4868 5846 4924
rect 5782 4864 5846 4868
rect 5862 4924 5926 4928
rect 5862 4868 5866 4924
rect 5866 4868 5922 4924
rect 5922 4868 5926 4924
rect 5862 4864 5926 4868
rect 5942 4924 6006 4928
rect 5942 4868 5946 4924
rect 5946 4868 6002 4924
rect 6002 4868 6006 4924
rect 5942 4864 6006 4868
rect 6022 4924 6086 4928
rect 6022 4868 6026 4924
rect 6026 4868 6082 4924
rect 6082 4868 6086 4924
rect 6022 4864 6086 4868
rect 7714 4924 7778 4928
rect 7714 4868 7718 4924
rect 7718 4868 7774 4924
rect 7774 4868 7778 4924
rect 7714 4864 7778 4868
rect 7794 4924 7858 4928
rect 7794 4868 7798 4924
rect 7798 4868 7854 4924
rect 7854 4868 7858 4924
rect 7794 4864 7858 4868
rect 7874 4924 7938 4928
rect 7874 4868 7878 4924
rect 7878 4868 7934 4924
rect 7934 4868 7938 4924
rect 7874 4864 7938 4868
rect 7954 4924 8018 4928
rect 7954 4868 7958 4924
rect 7958 4868 8014 4924
rect 8014 4868 8018 4924
rect 7954 4864 8018 4868
rect 2884 4380 2948 4384
rect 2884 4324 2888 4380
rect 2888 4324 2944 4380
rect 2944 4324 2948 4380
rect 2884 4320 2948 4324
rect 2964 4380 3028 4384
rect 2964 4324 2968 4380
rect 2968 4324 3024 4380
rect 3024 4324 3028 4380
rect 2964 4320 3028 4324
rect 3044 4380 3108 4384
rect 3044 4324 3048 4380
rect 3048 4324 3104 4380
rect 3104 4324 3108 4380
rect 3044 4320 3108 4324
rect 3124 4380 3188 4384
rect 3124 4324 3128 4380
rect 3128 4324 3184 4380
rect 3184 4324 3188 4380
rect 3124 4320 3188 4324
rect 4816 4380 4880 4384
rect 4816 4324 4820 4380
rect 4820 4324 4876 4380
rect 4876 4324 4880 4380
rect 4816 4320 4880 4324
rect 4896 4380 4960 4384
rect 4896 4324 4900 4380
rect 4900 4324 4956 4380
rect 4956 4324 4960 4380
rect 4896 4320 4960 4324
rect 4976 4380 5040 4384
rect 4976 4324 4980 4380
rect 4980 4324 5036 4380
rect 5036 4324 5040 4380
rect 4976 4320 5040 4324
rect 5056 4380 5120 4384
rect 5056 4324 5060 4380
rect 5060 4324 5116 4380
rect 5116 4324 5120 4380
rect 5056 4320 5120 4324
rect 6748 4380 6812 4384
rect 6748 4324 6752 4380
rect 6752 4324 6808 4380
rect 6808 4324 6812 4380
rect 6748 4320 6812 4324
rect 6828 4380 6892 4384
rect 6828 4324 6832 4380
rect 6832 4324 6888 4380
rect 6888 4324 6892 4380
rect 6828 4320 6892 4324
rect 6908 4380 6972 4384
rect 6908 4324 6912 4380
rect 6912 4324 6968 4380
rect 6968 4324 6972 4380
rect 6908 4320 6972 4324
rect 6988 4380 7052 4384
rect 6988 4324 6992 4380
rect 6992 4324 7048 4380
rect 7048 4324 7052 4380
rect 6988 4320 7052 4324
rect 8680 4380 8744 4384
rect 8680 4324 8684 4380
rect 8684 4324 8740 4380
rect 8740 4324 8744 4380
rect 8680 4320 8744 4324
rect 8760 4380 8824 4384
rect 8760 4324 8764 4380
rect 8764 4324 8820 4380
rect 8820 4324 8824 4380
rect 8760 4320 8824 4324
rect 8840 4380 8904 4384
rect 8840 4324 8844 4380
rect 8844 4324 8900 4380
rect 8900 4324 8904 4380
rect 8840 4320 8904 4324
rect 8920 4380 8984 4384
rect 8920 4324 8924 4380
rect 8924 4324 8980 4380
rect 8980 4324 8984 4380
rect 8920 4320 8984 4324
rect 1918 3836 1982 3840
rect 1918 3780 1922 3836
rect 1922 3780 1978 3836
rect 1978 3780 1982 3836
rect 1918 3776 1982 3780
rect 1998 3836 2062 3840
rect 1998 3780 2002 3836
rect 2002 3780 2058 3836
rect 2058 3780 2062 3836
rect 1998 3776 2062 3780
rect 2078 3836 2142 3840
rect 2078 3780 2082 3836
rect 2082 3780 2138 3836
rect 2138 3780 2142 3836
rect 2078 3776 2142 3780
rect 2158 3836 2222 3840
rect 2158 3780 2162 3836
rect 2162 3780 2218 3836
rect 2218 3780 2222 3836
rect 2158 3776 2222 3780
rect 3850 3836 3914 3840
rect 3850 3780 3854 3836
rect 3854 3780 3910 3836
rect 3910 3780 3914 3836
rect 3850 3776 3914 3780
rect 3930 3836 3994 3840
rect 3930 3780 3934 3836
rect 3934 3780 3990 3836
rect 3990 3780 3994 3836
rect 3930 3776 3994 3780
rect 4010 3836 4074 3840
rect 4010 3780 4014 3836
rect 4014 3780 4070 3836
rect 4070 3780 4074 3836
rect 4010 3776 4074 3780
rect 4090 3836 4154 3840
rect 4090 3780 4094 3836
rect 4094 3780 4150 3836
rect 4150 3780 4154 3836
rect 4090 3776 4154 3780
rect 5782 3836 5846 3840
rect 5782 3780 5786 3836
rect 5786 3780 5842 3836
rect 5842 3780 5846 3836
rect 5782 3776 5846 3780
rect 5862 3836 5926 3840
rect 5862 3780 5866 3836
rect 5866 3780 5922 3836
rect 5922 3780 5926 3836
rect 5862 3776 5926 3780
rect 5942 3836 6006 3840
rect 5942 3780 5946 3836
rect 5946 3780 6002 3836
rect 6002 3780 6006 3836
rect 5942 3776 6006 3780
rect 6022 3836 6086 3840
rect 6022 3780 6026 3836
rect 6026 3780 6082 3836
rect 6082 3780 6086 3836
rect 6022 3776 6086 3780
rect 7714 3836 7778 3840
rect 7714 3780 7718 3836
rect 7718 3780 7774 3836
rect 7774 3780 7778 3836
rect 7714 3776 7778 3780
rect 7794 3836 7858 3840
rect 7794 3780 7798 3836
rect 7798 3780 7854 3836
rect 7854 3780 7858 3836
rect 7794 3776 7858 3780
rect 7874 3836 7938 3840
rect 7874 3780 7878 3836
rect 7878 3780 7934 3836
rect 7934 3780 7938 3836
rect 7874 3776 7938 3780
rect 7954 3836 8018 3840
rect 7954 3780 7958 3836
rect 7958 3780 8014 3836
rect 8014 3780 8018 3836
rect 7954 3776 8018 3780
rect 2884 3292 2948 3296
rect 2884 3236 2888 3292
rect 2888 3236 2944 3292
rect 2944 3236 2948 3292
rect 2884 3232 2948 3236
rect 2964 3292 3028 3296
rect 2964 3236 2968 3292
rect 2968 3236 3024 3292
rect 3024 3236 3028 3292
rect 2964 3232 3028 3236
rect 3044 3292 3108 3296
rect 3044 3236 3048 3292
rect 3048 3236 3104 3292
rect 3104 3236 3108 3292
rect 3044 3232 3108 3236
rect 3124 3292 3188 3296
rect 3124 3236 3128 3292
rect 3128 3236 3184 3292
rect 3184 3236 3188 3292
rect 3124 3232 3188 3236
rect 4816 3292 4880 3296
rect 4816 3236 4820 3292
rect 4820 3236 4876 3292
rect 4876 3236 4880 3292
rect 4816 3232 4880 3236
rect 4896 3292 4960 3296
rect 4896 3236 4900 3292
rect 4900 3236 4956 3292
rect 4956 3236 4960 3292
rect 4896 3232 4960 3236
rect 4976 3292 5040 3296
rect 4976 3236 4980 3292
rect 4980 3236 5036 3292
rect 5036 3236 5040 3292
rect 4976 3232 5040 3236
rect 5056 3292 5120 3296
rect 5056 3236 5060 3292
rect 5060 3236 5116 3292
rect 5116 3236 5120 3292
rect 5056 3232 5120 3236
rect 6748 3292 6812 3296
rect 6748 3236 6752 3292
rect 6752 3236 6808 3292
rect 6808 3236 6812 3292
rect 6748 3232 6812 3236
rect 6828 3292 6892 3296
rect 6828 3236 6832 3292
rect 6832 3236 6888 3292
rect 6888 3236 6892 3292
rect 6828 3232 6892 3236
rect 6908 3292 6972 3296
rect 6908 3236 6912 3292
rect 6912 3236 6968 3292
rect 6968 3236 6972 3292
rect 6908 3232 6972 3236
rect 6988 3292 7052 3296
rect 6988 3236 6992 3292
rect 6992 3236 7048 3292
rect 7048 3236 7052 3292
rect 6988 3232 7052 3236
rect 8680 3292 8744 3296
rect 8680 3236 8684 3292
rect 8684 3236 8740 3292
rect 8740 3236 8744 3292
rect 8680 3232 8744 3236
rect 8760 3292 8824 3296
rect 8760 3236 8764 3292
rect 8764 3236 8820 3292
rect 8820 3236 8824 3292
rect 8760 3232 8824 3236
rect 8840 3292 8904 3296
rect 8840 3236 8844 3292
rect 8844 3236 8900 3292
rect 8900 3236 8904 3292
rect 8840 3232 8904 3236
rect 8920 3292 8984 3296
rect 8920 3236 8924 3292
rect 8924 3236 8980 3292
rect 8980 3236 8984 3292
rect 8920 3232 8984 3236
rect 1918 2748 1982 2752
rect 1918 2692 1922 2748
rect 1922 2692 1978 2748
rect 1978 2692 1982 2748
rect 1918 2688 1982 2692
rect 1998 2748 2062 2752
rect 1998 2692 2002 2748
rect 2002 2692 2058 2748
rect 2058 2692 2062 2748
rect 1998 2688 2062 2692
rect 2078 2748 2142 2752
rect 2078 2692 2082 2748
rect 2082 2692 2138 2748
rect 2138 2692 2142 2748
rect 2078 2688 2142 2692
rect 2158 2748 2222 2752
rect 2158 2692 2162 2748
rect 2162 2692 2218 2748
rect 2218 2692 2222 2748
rect 2158 2688 2222 2692
rect 3850 2748 3914 2752
rect 3850 2692 3854 2748
rect 3854 2692 3910 2748
rect 3910 2692 3914 2748
rect 3850 2688 3914 2692
rect 3930 2748 3994 2752
rect 3930 2692 3934 2748
rect 3934 2692 3990 2748
rect 3990 2692 3994 2748
rect 3930 2688 3994 2692
rect 4010 2748 4074 2752
rect 4010 2692 4014 2748
rect 4014 2692 4070 2748
rect 4070 2692 4074 2748
rect 4010 2688 4074 2692
rect 4090 2748 4154 2752
rect 4090 2692 4094 2748
rect 4094 2692 4150 2748
rect 4150 2692 4154 2748
rect 4090 2688 4154 2692
rect 5782 2748 5846 2752
rect 5782 2692 5786 2748
rect 5786 2692 5842 2748
rect 5842 2692 5846 2748
rect 5782 2688 5846 2692
rect 5862 2748 5926 2752
rect 5862 2692 5866 2748
rect 5866 2692 5922 2748
rect 5922 2692 5926 2748
rect 5862 2688 5926 2692
rect 5942 2748 6006 2752
rect 5942 2692 5946 2748
rect 5946 2692 6002 2748
rect 6002 2692 6006 2748
rect 5942 2688 6006 2692
rect 6022 2748 6086 2752
rect 6022 2692 6026 2748
rect 6026 2692 6082 2748
rect 6082 2692 6086 2748
rect 6022 2688 6086 2692
rect 7714 2748 7778 2752
rect 7714 2692 7718 2748
rect 7718 2692 7774 2748
rect 7774 2692 7778 2748
rect 7714 2688 7778 2692
rect 7794 2748 7858 2752
rect 7794 2692 7798 2748
rect 7798 2692 7854 2748
rect 7854 2692 7858 2748
rect 7794 2688 7858 2692
rect 7874 2748 7938 2752
rect 7874 2692 7878 2748
rect 7878 2692 7934 2748
rect 7934 2692 7938 2748
rect 7874 2688 7938 2692
rect 7954 2748 8018 2752
rect 7954 2692 7958 2748
rect 7958 2692 8014 2748
rect 8014 2692 8018 2748
rect 7954 2688 8018 2692
rect 2884 2204 2948 2208
rect 2884 2148 2888 2204
rect 2888 2148 2944 2204
rect 2944 2148 2948 2204
rect 2884 2144 2948 2148
rect 2964 2204 3028 2208
rect 2964 2148 2968 2204
rect 2968 2148 3024 2204
rect 3024 2148 3028 2204
rect 2964 2144 3028 2148
rect 3044 2204 3108 2208
rect 3044 2148 3048 2204
rect 3048 2148 3104 2204
rect 3104 2148 3108 2204
rect 3044 2144 3108 2148
rect 3124 2204 3188 2208
rect 3124 2148 3128 2204
rect 3128 2148 3184 2204
rect 3184 2148 3188 2204
rect 3124 2144 3188 2148
rect 4816 2204 4880 2208
rect 4816 2148 4820 2204
rect 4820 2148 4876 2204
rect 4876 2148 4880 2204
rect 4816 2144 4880 2148
rect 4896 2204 4960 2208
rect 4896 2148 4900 2204
rect 4900 2148 4956 2204
rect 4956 2148 4960 2204
rect 4896 2144 4960 2148
rect 4976 2204 5040 2208
rect 4976 2148 4980 2204
rect 4980 2148 5036 2204
rect 5036 2148 5040 2204
rect 4976 2144 5040 2148
rect 5056 2204 5120 2208
rect 5056 2148 5060 2204
rect 5060 2148 5116 2204
rect 5116 2148 5120 2204
rect 5056 2144 5120 2148
rect 6748 2204 6812 2208
rect 6748 2148 6752 2204
rect 6752 2148 6808 2204
rect 6808 2148 6812 2204
rect 6748 2144 6812 2148
rect 6828 2204 6892 2208
rect 6828 2148 6832 2204
rect 6832 2148 6888 2204
rect 6888 2148 6892 2204
rect 6828 2144 6892 2148
rect 6908 2204 6972 2208
rect 6908 2148 6912 2204
rect 6912 2148 6968 2204
rect 6968 2148 6972 2204
rect 6908 2144 6972 2148
rect 6988 2204 7052 2208
rect 6988 2148 6992 2204
rect 6992 2148 7048 2204
rect 7048 2148 7052 2204
rect 6988 2144 7052 2148
rect 8680 2204 8744 2208
rect 8680 2148 8684 2204
rect 8684 2148 8740 2204
rect 8740 2148 8744 2204
rect 8680 2144 8744 2148
rect 8760 2204 8824 2208
rect 8760 2148 8764 2204
rect 8764 2148 8820 2204
rect 8820 2148 8824 2204
rect 8760 2144 8824 2148
rect 8840 2204 8904 2208
rect 8840 2148 8844 2204
rect 8844 2148 8900 2204
rect 8900 2148 8904 2204
rect 8840 2144 8904 2148
rect 8920 2204 8984 2208
rect 8920 2148 8924 2204
rect 8924 2148 8980 2204
rect 8980 2148 8984 2204
rect 8920 2144 8984 2148
<< metal4 >>
rect 1910 19072 2230 19632
rect 1910 19008 1918 19072
rect 1982 19008 1998 19072
rect 2062 19008 2078 19072
rect 2142 19008 2158 19072
rect 2222 19008 2230 19072
rect 1910 17984 2230 19008
rect 1910 17920 1918 17984
rect 1982 17920 1998 17984
rect 2062 17920 2078 17984
rect 2142 17920 2158 17984
rect 2222 17920 2230 17984
rect 1910 16896 2230 17920
rect 1910 16832 1918 16896
rect 1982 16832 1998 16896
rect 2062 16832 2078 16896
rect 2142 16832 2158 16896
rect 2222 16832 2230 16896
rect 1910 15808 2230 16832
rect 1910 15744 1918 15808
rect 1982 15744 1998 15808
rect 2062 15744 2078 15808
rect 2142 15744 2158 15808
rect 2222 15744 2230 15808
rect 1910 14720 2230 15744
rect 1910 14656 1918 14720
rect 1982 14656 1998 14720
rect 2062 14656 2078 14720
rect 2142 14656 2158 14720
rect 2222 14656 2230 14720
rect 1910 13632 2230 14656
rect 1910 13568 1918 13632
rect 1982 13568 1998 13632
rect 2062 13568 2078 13632
rect 2142 13568 2158 13632
rect 2222 13568 2230 13632
rect 1910 12544 2230 13568
rect 1910 12480 1918 12544
rect 1982 12480 1998 12544
rect 2062 12480 2078 12544
rect 2142 12480 2158 12544
rect 2222 12480 2230 12544
rect 1910 11456 2230 12480
rect 1910 11392 1918 11456
rect 1982 11392 1998 11456
rect 2062 11392 2078 11456
rect 2142 11392 2158 11456
rect 2222 11392 2230 11456
rect 1910 10368 2230 11392
rect 1910 10304 1918 10368
rect 1982 10304 1998 10368
rect 2062 10304 2078 10368
rect 2142 10304 2158 10368
rect 2222 10304 2230 10368
rect 1910 9280 2230 10304
rect 1910 9216 1918 9280
rect 1982 9216 1998 9280
rect 2062 9216 2078 9280
rect 2142 9216 2158 9280
rect 2222 9216 2230 9280
rect 1910 8192 2230 9216
rect 1910 8128 1918 8192
rect 1982 8128 1998 8192
rect 2062 8128 2078 8192
rect 2142 8128 2158 8192
rect 2222 8128 2230 8192
rect 1910 7104 2230 8128
rect 1910 7040 1918 7104
rect 1982 7040 1998 7104
rect 2062 7040 2078 7104
rect 2142 7040 2158 7104
rect 2222 7040 2230 7104
rect 1910 6016 2230 7040
rect 1910 5952 1918 6016
rect 1982 5952 1998 6016
rect 2062 5952 2078 6016
rect 2142 5952 2158 6016
rect 2222 5952 2230 6016
rect 1910 4928 2230 5952
rect 1910 4864 1918 4928
rect 1982 4864 1998 4928
rect 2062 4864 2078 4928
rect 2142 4864 2158 4928
rect 2222 4864 2230 4928
rect 1910 3840 2230 4864
rect 1910 3776 1918 3840
rect 1982 3776 1998 3840
rect 2062 3776 2078 3840
rect 2142 3776 2158 3840
rect 2222 3776 2230 3840
rect 1910 2752 2230 3776
rect 1910 2688 1918 2752
rect 1982 2688 1998 2752
rect 2062 2688 2078 2752
rect 2142 2688 2158 2752
rect 2222 2688 2230 2752
rect 1910 2128 2230 2688
rect 2876 19616 3196 19632
rect 2876 19552 2884 19616
rect 2948 19552 2964 19616
rect 3028 19552 3044 19616
rect 3108 19552 3124 19616
rect 3188 19552 3196 19616
rect 2876 18528 3196 19552
rect 2876 18464 2884 18528
rect 2948 18464 2964 18528
rect 3028 18464 3044 18528
rect 3108 18464 3124 18528
rect 3188 18464 3196 18528
rect 2876 17440 3196 18464
rect 2876 17376 2884 17440
rect 2948 17376 2964 17440
rect 3028 17376 3044 17440
rect 3108 17376 3124 17440
rect 3188 17376 3196 17440
rect 2876 16352 3196 17376
rect 2876 16288 2884 16352
rect 2948 16288 2964 16352
rect 3028 16288 3044 16352
rect 3108 16288 3124 16352
rect 3188 16288 3196 16352
rect 2876 15264 3196 16288
rect 2876 15200 2884 15264
rect 2948 15200 2964 15264
rect 3028 15200 3044 15264
rect 3108 15200 3124 15264
rect 3188 15200 3196 15264
rect 2876 14176 3196 15200
rect 2876 14112 2884 14176
rect 2948 14112 2964 14176
rect 3028 14112 3044 14176
rect 3108 14112 3124 14176
rect 3188 14112 3196 14176
rect 2876 13088 3196 14112
rect 2876 13024 2884 13088
rect 2948 13024 2964 13088
rect 3028 13024 3044 13088
rect 3108 13024 3124 13088
rect 3188 13024 3196 13088
rect 2876 12000 3196 13024
rect 2876 11936 2884 12000
rect 2948 11936 2964 12000
rect 3028 11936 3044 12000
rect 3108 11936 3124 12000
rect 3188 11936 3196 12000
rect 2876 10912 3196 11936
rect 2876 10848 2884 10912
rect 2948 10848 2964 10912
rect 3028 10848 3044 10912
rect 3108 10848 3124 10912
rect 3188 10848 3196 10912
rect 2876 9824 3196 10848
rect 2876 9760 2884 9824
rect 2948 9760 2964 9824
rect 3028 9760 3044 9824
rect 3108 9760 3124 9824
rect 3188 9760 3196 9824
rect 2876 8736 3196 9760
rect 2876 8672 2884 8736
rect 2948 8672 2964 8736
rect 3028 8672 3044 8736
rect 3108 8672 3124 8736
rect 3188 8672 3196 8736
rect 2876 7648 3196 8672
rect 2876 7584 2884 7648
rect 2948 7584 2964 7648
rect 3028 7584 3044 7648
rect 3108 7584 3124 7648
rect 3188 7584 3196 7648
rect 2876 6560 3196 7584
rect 2876 6496 2884 6560
rect 2948 6496 2964 6560
rect 3028 6496 3044 6560
rect 3108 6496 3124 6560
rect 3188 6496 3196 6560
rect 2876 5472 3196 6496
rect 2876 5408 2884 5472
rect 2948 5408 2964 5472
rect 3028 5408 3044 5472
rect 3108 5408 3124 5472
rect 3188 5408 3196 5472
rect 2876 4384 3196 5408
rect 2876 4320 2884 4384
rect 2948 4320 2964 4384
rect 3028 4320 3044 4384
rect 3108 4320 3124 4384
rect 3188 4320 3196 4384
rect 2876 3296 3196 4320
rect 2876 3232 2884 3296
rect 2948 3232 2964 3296
rect 3028 3232 3044 3296
rect 3108 3232 3124 3296
rect 3188 3232 3196 3296
rect 2876 2208 3196 3232
rect 2876 2144 2884 2208
rect 2948 2144 2964 2208
rect 3028 2144 3044 2208
rect 3108 2144 3124 2208
rect 3188 2144 3196 2208
rect 2876 2128 3196 2144
rect 3842 19072 4162 19632
rect 3842 19008 3850 19072
rect 3914 19008 3930 19072
rect 3994 19008 4010 19072
rect 4074 19008 4090 19072
rect 4154 19008 4162 19072
rect 3842 17984 4162 19008
rect 3842 17920 3850 17984
rect 3914 17920 3930 17984
rect 3994 17920 4010 17984
rect 4074 17920 4090 17984
rect 4154 17920 4162 17984
rect 3842 16896 4162 17920
rect 3842 16832 3850 16896
rect 3914 16832 3930 16896
rect 3994 16832 4010 16896
rect 4074 16832 4090 16896
rect 4154 16832 4162 16896
rect 3842 15808 4162 16832
rect 3842 15744 3850 15808
rect 3914 15744 3930 15808
rect 3994 15744 4010 15808
rect 4074 15744 4090 15808
rect 4154 15744 4162 15808
rect 3842 14720 4162 15744
rect 3842 14656 3850 14720
rect 3914 14656 3930 14720
rect 3994 14656 4010 14720
rect 4074 14656 4090 14720
rect 4154 14656 4162 14720
rect 3842 13632 4162 14656
rect 3842 13568 3850 13632
rect 3914 13568 3930 13632
rect 3994 13568 4010 13632
rect 4074 13568 4090 13632
rect 4154 13568 4162 13632
rect 3842 12544 4162 13568
rect 3842 12480 3850 12544
rect 3914 12480 3930 12544
rect 3994 12480 4010 12544
rect 4074 12480 4090 12544
rect 4154 12480 4162 12544
rect 3842 11456 4162 12480
rect 3842 11392 3850 11456
rect 3914 11392 3930 11456
rect 3994 11392 4010 11456
rect 4074 11392 4090 11456
rect 4154 11392 4162 11456
rect 3842 10368 4162 11392
rect 3842 10304 3850 10368
rect 3914 10304 3930 10368
rect 3994 10304 4010 10368
rect 4074 10304 4090 10368
rect 4154 10304 4162 10368
rect 3842 9280 4162 10304
rect 3842 9216 3850 9280
rect 3914 9216 3930 9280
rect 3994 9216 4010 9280
rect 4074 9216 4090 9280
rect 4154 9216 4162 9280
rect 3842 8192 4162 9216
rect 3842 8128 3850 8192
rect 3914 8128 3930 8192
rect 3994 8128 4010 8192
rect 4074 8128 4090 8192
rect 4154 8128 4162 8192
rect 3842 7104 4162 8128
rect 3842 7040 3850 7104
rect 3914 7040 3930 7104
rect 3994 7040 4010 7104
rect 4074 7040 4090 7104
rect 4154 7040 4162 7104
rect 3842 6016 4162 7040
rect 3842 5952 3850 6016
rect 3914 5952 3930 6016
rect 3994 5952 4010 6016
rect 4074 5952 4090 6016
rect 4154 5952 4162 6016
rect 3842 4928 4162 5952
rect 3842 4864 3850 4928
rect 3914 4864 3930 4928
rect 3994 4864 4010 4928
rect 4074 4864 4090 4928
rect 4154 4864 4162 4928
rect 3842 3840 4162 4864
rect 3842 3776 3850 3840
rect 3914 3776 3930 3840
rect 3994 3776 4010 3840
rect 4074 3776 4090 3840
rect 4154 3776 4162 3840
rect 3842 2752 4162 3776
rect 3842 2688 3850 2752
rect 3914 2688 3930 2752
rect 3994 2688 4010 2752
rect 4074 2688 4090 2752
rect 4154 2688 4162 2752
rect 3842 2128 4162 2688
rect 4808 19616 5128 19632
rect 4808 19552 4816 19616
rect 4880 19552 4896 19616
rect 4960 19552 4976 19616
rect 5040 19552 5056 19616
rect 5120 19552 5128 19616
rect 4808 18528 5128 19552
rect 4808 18464 4816 18528
rect 4880 18464 4896 18528
rect 4960 18464 4976 18528
rect 5040 18464 5056 18528
rect 5120 18464 5128 18528
rect 4808 17440 5128 18464
rect 4808 17376 4816 17440
rect 4880 17376 4896 17440
rect 4960 17376 4976 17440
rect 5040 17376 5056 17440
rect 5120 17376 5128 17440
rect 4808 16352 5128 17376
rect 4808 16288 4816 16352
rect 4880 16288 4896 16352
rect 4960 16288 4976 16352
rect 5040 16288 5056 16352
rect 5120 16288 5128 16352
rect 4808 15264 5128 16288
rect 4808 15200 4816 15264
rect 4880 15200 4896 15264
rect 4960 15200 4976 15264
rect 5040 15200 5056 15264
rect 5120 15200 5128 15264
rect 4808 14176 5128 15200
rect 4808 14112 4816 14176
rect 4880 14112 4896 14176
rect 4960 14112 4976 14176
rect 5040 14112 5056 14176
rect 5120 14112 5128 14176
rect 4808 13088 5128 14112
rect 4808 13024 4816 13088
rect 4880 13024 4896 13088
rect 4960 13024 4976 13088
rect 5040 13024 5056 13088
rect 5120 13024 5128 13088
rect 4808 12000 5128 13024
rect 4808 11936 4816 12000
rect 4880 11936 4896 12000
rect 4960 11936 4976 12000
rect 5040 11936 5056 12000
rect 5120 11936 5128 12000
rect 4808 10912 5128 11936
rect 4808 10848 4816 10912
rect 4880 10848 4896 10912
rect 4960 10848 4976 10912
rect 5040 10848 5056 10912
rect 5120 10848 5128 10912
rect 4808 9824 5128 10848
rect 4808 9760 4816 9824
rect 4880 9760 4896 9824
rect 4960 9760 4976 9824
rect 5040 9760 5056 9824
rect 5120 9760 5128 9824
rect 4808 8736 5128 9760
rect 4808 8672 4816 8736
rect 4880 8672 4896 8736
rect 4960 8672 4976 8736
rect 5040 8672 5056 8736
rect 5120 8672 5128 8736
rect 4808 7648 5128 8672
rect 4808 7584 4816 7648
rect 4880 7584 4896 7648
rect 4960 7584 4976 7648
rect 5040 7584 5056 7648
rect 5120 7584 5128 7648
rect 4808 6560 5128 7584
rect 4808 6496 4816 6560
rect 4880 6496 4896 6560
rect 4960 6496 4976 6560
rect 5040 6496 5056 6560
rect 5120 6496 5128 6560
rect 4808 5472 5128 6496
rect 4808 5408 4816 5472
rect 4880 5408 4896 5472
rect 4960 5408 4976 5472
rect 5040 5408 5056 5472
rect 5120 5408 5128 5472
rect 4808 4384 5128 5408
rect 4808 4320 4816 4384
rect 4880 4320 4896 4384
rect 4960 4320 4976 4384
rect 5040 4320 5056 4384
rect 5120 4320 5128 4384
rect 4808 3296 5128 4320
rect 4808 3232 4816 3296
rect 4880 3232 4896 3296
rect 4960 3232 4976 3296
rect 5040 3232 5056 3296
rect 5120 3232 5128 3296
rect 4808 2208 5128 3232
rect 4808 2144 4816 2208
rect 4880 2144 4896 2208
rect 4960 2144 4976 2208
rect 5040 2144 5056 2208
rect 5120 2144 5128 2208
rect 4808 2128 5128 2144
rect 5774 19072 6094 19632
rect 5774 19008 5782 19072
rect 5846 19008 5862 19072
rect 5926 19008 5942 19072
rect 6006 19008 6022 19072
rect 6086 19008 6094 19072
rect 5774 17984 6094 19008
rect 5774 17920 5782 17984
rect 5846 17920 5862 17984
rect 5926 17920 5942 17984
rect 6006 17920 6022 17984
rect 6086 17920 6094 17984
rect 5774 16896 6094 17920
rect 5774 16832 5782 16896
rect 5846 16832 5862 16896
rect 5926 16832 5942 16896
rect 6006 16832 6022 16896
rect 6086 16832 6094 16896
rect 5774 15808 6094 16832
rect 5774 15744 5782 15808
rect 5846 15744 5862 15808
rect 5926 15744 5942 15808
rect 6006 15744 6022 15808
rect 6086 15744 6094 15808
rect 5774 14720 6094 15744
rect 5774 14656 5782 14720
rect 5846 14656 5862 14720
rect 5926 14656 5942 14720
rect 6006 14656 6022 14720
rect 6086 14656 6094 14720
rect 5774 13632 6094 14656
rect 5774 13568 5782 13632
rect 5846 13568 5862 13632
rect 5926 13568 5942 13632
rect 6006 13568 6022 13632
rect 6086 13568 6094 13632
rect 5774 12544 6094 13568
rect 5774 12480 5782 12544
rect 5846 12480 5862 12544
rect 5926 12480 5942 12544
rect 6006 12480 6022 12544
rect 6086 12480 6094 12544
rect 5774 11456 6094 12480
rect 5774 11392 5782 11456
rect 5846 11392 5862 11456
rect 5926 11392 5942 11456
rect 6006 11392 6022 11456
rect 6086 11392 6094 11456
rect 5774 10368 6094 11392
rect 5774 10304 5782 10368
rect 5846 10304 5862 10368
rect 5926 10304 5942 10368
rect 6006 10304 6022 10368
rect 6086 10304 6094 10368
rect 5774 9280 6094 10304
rect 5774 9216 5782 9280
rect 5846 9216 5862 9280
rect 5926 9216 5942 9280
rect 6006 9216 6022 9280
rect 6086 9216 6094 9280
rect 5774 8192 6094 9216
rect 5774 8128 5782 8192
rect 5846 8128 5862 8192
rect 5926 8128 5942 8192
rect 6006 8128 6022 8192
rect 6086 8128 6094 8192
rect 5774 7104 6094 8128
rect 5774 7040 5782 7104
rect 5846 7040 5862 7104
rect 5926 7040 5942 7104
rect 6006 7040 6022 7104
rect 6086 7040 6094 7104
rect 5774 6016 6094 7040
rect 5774 5952 5782 6016
rect 5846 5952 5862 6016
rect 5926 5952 5942 6016
rect 6006 5952 6022 6016
rect 6086 5952 6094 6016
rect 5774 4928 6094 5952
rect 5774 4864 5782 4928
rect 5846 4864 5862 4928
rect 5926 4864 5942 4928
rect 6006 4864 6022 4928
rect 6086 4864 6094 4928
rect 5774 3840 6094 4864
rect 5774 3776 5782 3840
rect 5846 3776 5862 3840
rect 5926 3776 5942 3840
rect 6006 3776 6022 3840
rect 6086 3776 6094 3840
rect 5774 2752 6094 3776
rect 5774 2688 5782 2752
rect 5846 2688 5862 2752
rect 5926 2688 5942 2752
rect 6006 2688 6022 2752
rect 6086 2688 6094 2752
rect 5774 2128 6094 2688
rect 6740 19616 7060 19632
rect 6740 19552 6748 19616
rect 6812 19552 6828 19616
rect 6892 19552 6908 19616
rect 6972 19552 6988 19616
rect 7052 19552 7060 19616
rect 6740 18528 7060 19552
rect 6740 18464 6748 18528
rect 6812 18464 6828 18528
rect 6892 18464 6908 18528
rect 6972 18464 6988 18528
rect 7052 18464 7060 18528
rect 6740 17440 7060 18464
rect 6740 17376 6748 17440
rect 6812 17376 6828 17440
rect 6892 17376 6908 17440
rect 6972 17376 6988 17440
rect 7052 17376 7060 17440
rect 6740 16352 7060 17376
rect 6740 16288 6748 16352
rect 6812 16288 6828 16352
rect 6892 16288 6908 16352
rect 6972 16288 6988 16352
rect 7052 16288 7060 16352
rect 6740 15264 7060 16288
rect 6740 15200 6748 15264
rect 6812 15200 6828 15264
rect 6892 15200 6908 15264
rect 6972 15200 6988 15264
rect 7052 15200 7060 15264
rect 6740 14176 7060 15200
rect 6740 14112 6748 14176
rect 6812 14112 6828 14176
rect 6892 14112 6908 14176
rect 6972 14112 6988 14176
rect 7052 14112 7060 14176
rect 6740 13088 7060 14112
rect 6740 13024 6748 13088
rect 6812 13024 6828 13088
rect 6892 13024 6908 13088
rect 6972 13024 6988 13088
rect 7052 13024 7060 13088
rect 6740 12000 7060 13024
rect 6740 11936 6748 12000
rect 6812 11936 6828 12000
rect 6892 11936 6908 12000
rect 6972 11936 6988 12000
rect 7052 11936 7060 12000
rect 6740 10912 7060 11936
rect 6740 10848 6748 10912
rect 6812 10848 6828 10912
rect 6892 10848 6908 10912
rect 6972 10848 6988 10912
rect 7052 10848 7060 10912
rect 6740 9824 7060 10848
rect 6740 9760 6748 9824
rect 6812 9760 6828 9824
rect 6892 9760 6908 9824
rect 6972 9760 6988 9824
rect 7052 9760 7060 9824
rect 6740 8736 7060 9760
rect 6740 8672 6748 8736
rect 6812 8672 6828 8736
rect 6892 8672 6908 8736
rect 6972 8672 6988 8736
rect 7052 8672 7060 8736
rect 6740 7648 7060 8672
rect 6740 7584 6748 7648
rect 6812 7584 6828 7648
rect 6892 7584 6908 7648
rect 6972 7584 6988 7648
rect 7052 7584 7060 7648
rect 6740 6560 7060 7584
rect 6740 6496 6748 6560
rect 6812 6496 6828 6560
rect 6892 6496 6908 6560
rect 6972 6496 6988 6560
rect 7052 6496 7060 6560
rect 6740 5472 7060 6496
rect 6740 5408 6748 5472
rect 6812 5408 6828 5472
rect 6892 5408 6908 5472
rect 6972 5408 6988 5472
rect 7052 5408 7060 5472
rect 6740 4384 7060 5408
rect 6740 4320 6748 4384
rect 6812 4320 6828 4384
rect 6892 4320 6908 4384
rect 6972 4320 6988 4384
rect 7052 4320 7060 4384
rect 6740 3296 7060 4320
rect 6740 3232 6748 3296
rect 6812 3232 6828 3296
rect 6892 3232 6908 3296
rect 6972 3232 6988 3296
rect 7052 3232 7060 3296
rect 6740 2208 7060 3232
rect 6740 2144 6748 2208
rect 6812 2144 6828 2208
rect 6892 2144 6908 2208
rect 6972 2144 6988 2208
rect 7052 2144 7060 2208
rect 6740 2128 7060 2144
rect 7706 19072 8026 19632
rect 7706 19008 7714 19072
rect 7778 19008 7794 19072
rect 7858 19008 7874 19072
rect 7938 19008 7954 19072
rect 8018 19008 8026 19072
rect 7706 17984 8026 19008
rect 7706 17920 7714 17984
rect 7778 17920 7794 17984
rect 7858 17920 7874 17984
rect 7938 17920 7954 17984
rect 8018 17920 8026 17984
rect 7706 16896 8026 17920
rect 7706 16832 7714 16896
rect 7778 16832 7794 16896
rect 7858 16832 7874 16896
rect 7938 16832 7954 16896
rect 8018 16832 8026 16896
rect 7706 15808 8026 16832
rect 7706 15744 7714 15808
rect 7778 15744 7794 15808
rect 7858 15744 7874 15808
rect 7938 15744 7954 15808
rect 8018 15744 8026 15808
rect 7706 14720 8026 15744
rect 7706 14656 7714 14720
rect 7778 14656 7794 14720
rect 7858 14656 7874 14720
rect 7938 14656 7954 14720
rect 8018 14656 8026 14720
rect 7706 13632 8026 14656
rect 7706 13568 7714 13632
rect 7778 13568 7794 13632
rect 7858 13568 7874 13632
rect 7938 13568 7954 13632
rect 8018 13568 8026 13632
rect 7706 12544 8026 13568
rect 7706 12480 7714 12544
rect 7778 12480 7794 12544
rect 7858 12480 7874 12544
rect 7938 12480 7954 12544
rect 8018 12480 8026 12544
rect 7706 11456 8026 12480
rect 7706 11392 7714 11456
rect 7778 11392 7794 11456
rect 7858 11392 7874 11456
rect 7938 11392 7954 11456
rect 8018 11392 8026 11456
rect 7706 10368 8026 11392
rect 7706 10304 7714 10368
rect 7778 10304 7794 10368
rect 7858 10304 7874 10368
rect 7938 10304 7954 10368
rect 8018 10304 8026 10368
rect 7706 9280 8026 10304
rect 7706 9216 7714 9280
rect 7778 9216 7794 9280
rect 7858 9216 7874 9280
rect 7938 9216 7954 9280
rect 8018 9216 8026 9280
rect 7706 8192 8026 9216
rect 7706 8128 7714 8192
rect 7778 8128 7794 8192
rect 7858 8128 7874 8192
rect 7938 8128 7954 8192
rect 8018 8128 8026 8192
rect 7706 7104 8026 8128
rect 7706 7040 7714 7104
rect 7778 7040 7794 7104
rect 7858 7040 7874 7104
rect 7938 7040 7954 7104
rect 8018 7040 8026 7104
rect 7706 6016 8026 7040
rect 7706 5952 7714 6016
rect 7778 5952 7794 6016
rect 7858 5952 7874 6016
rect 7938 5952 7954 6016
rect 8018 5952 8026 6016
rect 7706 4928 8026 5952
rect 7706 4864 7714 4928
rect 7778 4864 7794 4928
rect 7858 4864 7874 4928
rect 7938 4864 7954 4928
rect 8018 4864 8026 4928
rect 7706 3840 8026 4864
rect 7706 3776 7714 3840
rect 7778 3776 7794 3840
rect 7858 3776 7874 3840
rect 7938 3776 7954 3840
rect 8018 3776 8026 3840
rect 7706 2752 8026 3776
rect 7706 2688 7714 2752
rect 7778 2688 7794 2752
rect 7858 2688 7874 2752
rect 7938 2688 7954 2752
rect 8018 2688 8026 2752
rect 7706 2128 8026 2688
rect 8672 19616 8992 19632
rect 8672 19552 8680 19616
rect 8744 19552 8760 19616
rect 8824 19552 8840 19616
rect 8904 19552 8920 19616
rect 8984 19552 8992 19616
rect 8672 18528 8992 19552
rect 8672 18464 8680 18528
rect 8744 18464 8760 18528
rect 8824 18464 8840 18528
rect 8904 18464 8920 18528
rect 8984 18464 8992 18528
rect 8672 17440 8992 18464
rect 8672 17376 8680 17440
rect 8744 17376 8760 17440
rect 8824 17376 8840 17440
rect 8904 17376 8920 17440
rect 8984 17376 8992 17440
rect 8672 16352 8992 17376
rect 8672 16288 8680 16352
rect 8744 16288 8760 16352
rect 8824 16288 8840 16352
rect 8904 16288 8920 16352
rect 8984 16288 8992 16352
rect 8672 15264 8992 16288
rect 8672 15200 8680 15264
rect 8744 15200 8760 15264
rect 8824 15200 8840 15264
rect 8904 15200 8920 15264
rect 8984 15200 8992 15264
rect 8672 14176 8992 15200
rect 8672 14112 8680 14176
rect 8744 14112 8760 14176
rect 8824 14112 8840 14176
rect 8904 14112 8920 14176
rect 8984 14112 8992 14176
rect 8672 13088 8992 14112
rect 8672 13024 8680 13088
rect 8744 13024 8760 13088
rect 8824 13024 8840 13088
rect 8904 13024 8920 13088
rect 8984 13024 8992 13088
rect 8672 12000 8992 13024
rect 8672 11936 8680 12000
rect 8744 11936 8760 12000
rect 8824 11936 8840 12000
rect 8904 11936 8920 12000
rect 8984 11936 8992 12000
rect 8672 10912 8992 11936
rect 8672 10848 8680 10912
rect 8744 10848 8760 10912
rect 8824 10848 8840 10912
rect 8904 10848 8920 10912
rect 8984 10848 8992 10912
rect 8672 9824 8992 10848
rect 8672 9760 8680 9824
rect 8744 9760 8760 9824
rect 8824 9760 8840 9824
rect 8904 9760 8920 9824
rect 8984 9760 8992 9824
rect 8672 8736 8992 9760
rect 8672 8672 8680 8736
rect 8744 8672 8760 8736
rect 8824 8672 8840 8736
rect 8904 8672 8920 8736
rect 8984 8672 8992 8736
rect 8672 7648 8992 8672
rect 8672 7584 8680 7648
rect 8744 7584 8760 7648
rect 8824 7584 8840 7648
rect 8904 7584 8920 7648
rect 8984 7584 8992 7648
rect 8672 6560 8992 7584
rect 8672 6496 8680 6560
rect 8744 6496 8760 6560
rect 8824 6496 8840 6560
rect 8904 6496 8920 6560
rect 8984 6496 8992 6560
rect 8672 5472 8992 6496
rect 8672 5408 8680 5472
rect 8744 5408 8760 5472
rect 8824 5408 8840 5472
rect 8904 5408 8920 5472
rect 8984 5408 8992 5472
rect 8672 4384 8992 5408
rect 8672 4320 8680 4384
rect 8744 4320 8760 4384
rect 8824 4320 8840 4384
rect 8904 4320 8920 4384
rect 8984 4320 8992 4384
rect 8672 3296 8992 4320
rect 8672 3232 8680 3296
rect 8744 3232 8760 3296
rect 8824 3232 8840 3296
rect 8904 3232 8920 3296
rect 8984 3232 8992 3296
rect 8672 2208 8992 3232
rect 8672 2144 8680 2208
rect 8744 2144 8760 2208
rect 8824 2144 8840 2208
rect 8904 2144 8920 2208
rect 8984 2144 8992 2208
rect 8672 2128 8992 2144
use sky130_fd_sc_hd__mux2_1  _13_ pdk/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1689802698
transform -1 0 2208 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__and3b_1  _14_ pdk/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1689802698
transform 1 0 1380 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nor3b_1  _15_ pdk/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1689802698
transform -1 0 1932 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a2111oi_1  _16_ pdk/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1689802698
transform -1 0 2944 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _17_
timestamp 1689802698
transform -1 0 2208 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _18_ pdk/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1689802698
transform -1 0 2024 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand3b_1  _19_ pdk/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1689802698
transform -1 0 2760 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _20_ pdk/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1689802698
transform 1 0 1564 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_1  _21_ pdk/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1689802698
transform -1 0 2392 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__mux4_1  _22_ pdk/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1689802698
transform 1 0 1380 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _23_
timestamp 1689802698
transform 1 0 1380 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _24_
timestamp 1689802698
transform 1 0 2300 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _25_ pdk/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1689802698
transform 1 0 2300 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_2  _26_ pdk/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1689802698
transform -1 0 3036 0 -1 11968
box -38 -48 682 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_9 pdk/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1689802698
transform 1 0 1932 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_21 pdk/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1689802698
transform 1 0 3036 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 pdk/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1689802698
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1689802698
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1689802698
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53 pdk/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1689802698
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1689802698
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 1689802698
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1689802698
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1689802698
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1689802698
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1689802698
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51 pdk/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1689802698
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1689802698
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1689802698
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1689802698
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_6
timestamp 1689802698
transform 1 0 1656 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_18 pdk/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1689802698
transform 1 0 2760 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_26 pdk/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1689802698
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1689802698
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1689802698
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1689802698
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1689802698
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_77
timestamp 1689802698
transform 1 0 8188 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1689802698
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1689802698
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1689802698
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1689802698
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1689802698
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1689802698
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1689802698
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1689802698
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_6
timestamp 1689802698
transform 1 0 1656 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_18
timestamp 1689802698
transform 1 0 2760 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_26
timestamp 1689802698
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1689802698
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1689802698
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1689802698
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1689802698
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_77
timestamp 1689802698
transform 1 0 8188 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_12
timestamp 1689802698
transform 1 0 2208 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_24
timestamp 1689802698
transform 1 0 3312 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_36
timestamp 1689802698
transform 1 0 4416 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_48
timestamp 1689802698
transform 1 0 5520 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1689802698
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1689802698
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_6
timestamp 1689802698
transform 1 0 1656 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_10
timestamp 1689802698
transform 1 0 2024 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_22
timestamp 1689802698
transform 1 0 3128 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1689802698
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1689802698
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1689802698
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1689802698
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_77
timestamp 1689802698
transform 1 0 8188 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_3
timestamp 1689802698
transform 1 0 1380 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_18
timestamp 1689802698
transform 1 0 2760 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_30
timestamp 1689802698
transform 1 0 3864 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_42
timestamp 1689802698
transform 1 0 4968 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_54
timestamp 1689802698
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1689802698
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1689802698
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_3
timestamp 1689802698
transform 1 0 1380 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_14
timestamp 1689802698
transform 1 0 2392 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_26
timestamp 1689802698
transform 1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1689802698
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1689802698
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1689802698
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 1689802698
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_77
timestamp 1689802698
transform 1 0 8188 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_6
timestamp 1689802698
transform 1 0 1656 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_18
timestamp 1689802698
transform 1 0 2760 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_30
timestamp 1689802698
transform 1 0 3864 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_42
timestamp 1689802698
transform 1 0 4968 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_54
timestamp 1689802698
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1689802698
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 1689802698
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_10
timestamp 1689802698
transform 1 0 2024 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_22
timestamp 1689802698
transform 1 0 3128 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1689802698
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1689802698
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 1689802698
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_65
timestamp 1689802698
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_77
timestamp 1689802698
transform 1 0 8188 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_20
timestamp 1689802698
transform 1 0 2944 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_32
timestamp 1689802698
transform 1 0 4048 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_44
timestamp 1689802698
transform 1 0 5152 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1689802698
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 1689802698
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_6
timestamp 1689802698
transform 1 0 1656 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_18
timestamp 1689802698
transform 1 0 2760 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_26
timestamp 1689802698
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1689802698
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1689802698
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_53
timestamp 1689802698
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_65
timestamp 1689802698
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_77
timestamp 1689802698
transform 1 0 8188 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_9
timestamp 1689802698
transform 1 0 1932 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_21
timestamp 1689802698
transform 1 0 3036 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_33
timestamp 1689802698
transform 1 0 4140 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_45
timestamp 1689802698
transform 1 0 5244 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_53
timestamp 1689802698
transform 1 0 5980 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 1689802698
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_69
timestamp 1689802698
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1689802698
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 1689802698
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1689802698
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1689802698
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_41
timestamp 1689802698
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_53
timestamp 1689802698
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_65
timestamp 1689802698
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_77
timestamp 1689802698
transform 1 0 8188 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_6
timestamp 1689802698
transform 1 0 1656 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_18
timestamp 1689802698
transform 1 0 2760 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_30
timestamp 1689802698
transform 1 0 3864 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_42
timestamp 1689802698
transform 1 0 4968 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_54
timestamp 1689802698
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp 1689802698
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_69
timestamp 1689802698
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1689802698
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp 1689802698
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1689802698
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 1689802698
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_41
timestamp 1689802698
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_53
timestamp 1689802698
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_6
timestamp 1689802698
transform 1 0 1656 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_21
timestamp 1689802698
transform 1 0 3036 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_33
timestamp 1689802698
transform 1 0 4140 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_45
timestamp 1689802698
transform 1 0 5244 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_53
timestamp 1689802698
transform 1 0 5980 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_57
timestamp 1689802698
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_69
timestamp 1689802698
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_3
timestamp 1689802698
transform 1 0 1380 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_11
timestamp 1689802698
transform 1 0 2116 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_16
timestamp 1689802698
transform 1 0 2576 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp 1689802698
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_41
timestamp 1689802698
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_53
timestamp 1689802698
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_65
timestamp 1689802698
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_77
timestamp 1689802698
transform 1 0 8188 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 1689802698
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_15
timestamp 1689802698
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_27
timestamp 1689802698
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_39
timestamp 1689802698
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_51
timestamp 1689802698
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_55
timestamp 1689802698
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_57
timestamp 1689802698
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_69
timestamp 1689802698
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_6
timestamp 1689802698
transform 1 0 1656 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_18
timestamp 1689802698
transform 1 0 2760 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_26
timestamp 1689802698
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_29
timestamp 1689802698
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_41
timestamp 1689802698
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_53
timestamp 1689802698
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_65
timestamp 1689802698
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_77
timestamp 1689802698
transform 1 0 8188 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 1689802698
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_15
timestamp 1689802698
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_27
timestamp 1689802698
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_39
timestamp 1689802698
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_51
timestamp 1689802698
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 1689802698
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_57
timestamp 1689802698
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_69
timestamp 1689802698
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_6
timestamp 1689802698
transform 1 0 1656 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_12
timestamp 1689802698
transform 1 0 2208 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_22
timestamp 1689802698
transform 1 0 3128 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_29
timestamp 1689802698
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_41
timestamp 1689802698
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_53
timestamp 1689802698
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_65
timestamp 1689802698
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_77
timestamp 1689802698
transform 1 0 8188 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_24
timestamp 1689802698
transform 1 0 3312 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_36
timestamp 1689802698
transform 1 0 4416 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_48
timestamp 1689802698
transform 1 0 5520 0 -1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_57
timestamp 1689802698
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_69
timestamp 1689802698
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_6
timestamp 1689802698
transform 1 0 1656 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_18
timestamp 1689802698
transform 1 0 2760 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_26
timestamp 1689802698
transform 1 0 3496 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_29
timestamp 1689802698
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_41
timestamp 1689802698
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_53
timestamp 1689802698
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_65
timestamp 1689802698
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_77
timestamp 1689802698
transform 1 0 8188 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_24
timestamp 1689802698
transform 1 0 3312 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_36
timestamp 1689802698
transform 1 0 4416 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_48
timestamp 1689802698
transform 1 0 5520 0 -1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_57
timestamp 1689802698
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_69
timestamp 1689802698
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_3
timestamp 1689802698
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_15
timestamp 1689802698
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 1689802698
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_29
timestamp 1689802698
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_41
timestamp 1689802698
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_53
timestamp 1689802698
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_65
timestamp 1689802698
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_77
timestamp 1689802698
transform 1 0 8188 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_6
timestamp 1689802698
transform 1 0 1656 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_18
timestamp 1689802698
transform 1 0 2760 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_30
timestamp 1689802698
transform 1 0 3864 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_42
timestamp 1689802698
transform 1 0 4968 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_54
timestamp 1689802698
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_57
timestamp 1689802698
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_69
timestamp 1689802698
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp 1689802698
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_15
timestamp 1689802698
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 1689802698
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_29
timestamp 1689802698
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_41
timestamp 1689802698
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_53
timestamp 1689802698
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_65
timestamp 1689802698
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_77
timestamp 1689802698
transform 1 0 8188 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_3
timestamp 1689802698
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_15
timestamp 1689802698
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_27
timestamp 1689802698
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_39
timestamp 1689802698
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_51
timestamp 1689802698
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_55
timestamp 1689802698
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_57
timestamp 1689802698
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_69
timestamp 1689802698
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_6
timestamp 1689802698
transform 1 0 1656 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_18
timestamp 1689802698
transform 1 0 2760 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_26
timestamp 1689802698
transform 1 0 3496 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_29
timestamp 1689802698
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_41
timestamp 1689802698
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_53
timestamp 1689802698
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_65
timestamp 1689802698
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_77
timestamp 1689802698
transform 1 0 8188 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_13
timestamp 1689802698
transform 1 0 2300 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_25
timestamp 1689802698
transform 1 0 3404 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_33
timestamp 1689802698
transform 1 0 4140 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_45
timestamp 1689802698
transform 1 0 5244 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_53
timestamp 1689802698
transform 1 0 5980 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_61
timestamp 1689802698
transform 1 0 6716 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_73
timestamp 1689802698
transform 1 0 7820 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_77
timestamp 1689802698
transform 1 0 8188 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input1 pdk/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1689802698
transform 1 0 1748 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1689802698
transform -1 0 1656 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1689802698
transform -1 0 1656 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1689802698
transform -1 0 1656 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1689802698
transform -1 0 1656 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1689802698
transform -1 0 1656 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1689802698
transform -1 0 1932 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1689802698
transform 1 0 2024 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1689802698
transform -1 0 1656 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1689802698
transform -1 0 1656 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1689802698
transform -1 0 1656 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1689802698
transform -1 0 1656 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1689802698
transform -1 0 1656 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1689802698
transform -1 0 1656 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1689802698
transform -1 0 1656 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1689802698
transform -1 0 1656 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input17 pdk/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1689802698
transform 1 0 1380 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input18 pdk/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1689802698
transform 1 0 3772 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input19
timestamp 1689802698
transform -1 0 6716 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input20 pdk/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1689802698
transform -1 0 8556 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  output21 pdk/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1689802698
transform 1 0 7084 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1689802698
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1689802698
transform -1 0 8832 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1689802698
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1689802698
transform -1 0 8832 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1689802698
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1689802698
transform -1 0 8832 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1689802698
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1689802698
transform -1 0 8832 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1689802698
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1689802698
transform -1 0 8832 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1689802698
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1689802698
transform -1 0 8832 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1689802698
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1689802698
transform -1 0 8832 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1689802698
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1689802698
transform -1 0 8832 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1689802698
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1689802698
transform -1 0 8832 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1689802698
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1689802698
transform -1 0 8832 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1689802698
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1689802698
transform -1 0 8832 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1689802698
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1689802698
transform -1 0 8832 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1689802698
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1689802698
transform -1 0 8832 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1689802698
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1689802698
transform -1 0 8832 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1689802698
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1689802698
transform -1 0 8832 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1689802698
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1689802698
transform -1 0 8832 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1689802698
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1689802698
transform -1 0 8832 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1689802698
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1689802698
transform -1 0 8832 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1689802698
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1689802698
transform -1 0 8832 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1689802698
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1689802698
transform -1 0 8832 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1689802698
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1689802698
transform -1 0 8832 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1689802698
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1689802698
transform -1 0 8832 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1689802698
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1689802698
transform -1 0 8832 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1689802698
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1689802698
transform -1 0 8832 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1689802698
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1689802698
transform -1 0 8832 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1689802698
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1689802698
transform -1 0 8832 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1689802698
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1689802698
transform -1 0 8832 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1689802698
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1689802698
transform -1 0 8832 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1689802698
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1689802698
transform -1 0 8832 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1689802698
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1689802698
transform -1 0 8832 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1689802698
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1689802698
transform -1 0 8832 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1689802698
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1689802698
transform -1 0 8832 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64 pdk/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1689802698
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1689802698
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1689802698
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1689802698
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1689802698
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1689802698
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1689802698
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1689802698
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1689802698
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1689802698
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1689802698
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1689802698
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1689802698
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1689802698
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1689802698
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1689802698
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1689802698
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1689802698
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1689802698
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1689802698
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1689802698
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1689802698
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1689802698
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1689802698
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1689802698
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1689802698
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1689802698
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1689802698
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1689802698
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1689802698
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1689802698
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1689802698
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1689802698
transform 1 0 3680 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1689802698
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
<< labels >>
flabel metal3 s 0 20952 800 21072 0 FreeSans 480 0 0 0 data_in[0]
port 0 nsew signal input
flabel metal3 s 0 7352 800 7472 0 FreeSans 480 0 0 0 data_in[10]
port 1 nsew signal input
flabel metal3 s 0 5992 800 6112 0 FreeSans 480 0 0 0 data_in[11]
port 2 nsew signal input
flabel metal3 s 0 4632 800 4752 0 FreeSans 480 0 0 0 data_in[12]
port 3 nsew signal input
flabel metal3 s 0 3272 800 3392 0 FreeSans 480 0 0 0 data_in[13]
port 4 nsew signal input
flabel metal3 s 0 1912 800 2032 0 FreeSans 480 0 0 0 data_in[14]
port 5 nsew signal input
flabel metal3 s 0 552 800 672 0 FreeSans 480 0 0 0 data_in[15]
port 6 nsew signal input
flabel metal3 s 0 19592 800 19712 0 FreeSans 480 0 0 0 data_in[1]
port 7 nsew signal input
flabel metal3 s 0 18232 800 18352 0 FreeSans 480 0 0 0 data_in[2]
port 8 nsew signal input
flabel metal3 s 0 16872 800 16992 0 FreeSans 480 0 0 0 data_in[3]
port 9 nsew signal input
flabel metal3 s 0 15512 800 15632 0 FreeSans 480 0 0 0 data_in[4]
port 10 nsew signal input
flabel metal3 s 0 14152 800 14272 0 FreeSans 480 0 0 0 data_in[5]
port 11 nsew signal input
flabel metal3 s 0 12792 800 12912 0 FreeSans 480 0 0 0 data_in[6]
port 12 nsew signal input
flabel metal3 s 0 11432 800 11552 0 FreeSans 480 0 0 0 data_in[7]
port 13 nsew signal input
flabel metal3 s 0 10072 800 10192 0 FreeSans 480 0 0 0 data_in[8]
port 14 nsew signal input
flabel metal3 s 0 8712 800 8832 0 FreeSans 480 0 0 0 data_in[9]
port 15 nsew signal input
flabel metal2 s 1214 21200 1270 22000 0 FreeSans 224 90 0 0 select[0]
port 16 nsew signal input
flabel metal2 s 3698 21200 3754 22000 0 FreeSans 224 90 0 0 select[1]
port 17 nsew signal input
flabel metal2 s 6182 21200 6238 22000 0 FreeSans 224 90 0 0 select[2]
port 18 nsew signal input
flabel metal2 s 8666 21200 8722 22000 0 FreeSans 224 90 0 0 select[3]
port 19 nsew signal input
flabel metal4 s 1910 2128 2230 19632 0 FreeSans 1920 90 0 0 vccd1
port 20 nsew power bidirectional
flabel metal4 s 3842 2128 4162 19632 0 FreeSans 1920 90 0 0 vccd1
port 20 nsew power bidirectional
flabel metal4 s 5774 2128 6094 19632 0 FreeSans 1920 90 0 0 vccd1
port 20 nsew power bidirectional
flabel metal4 s 7706 2128 8026 19632 0 FreeSans 1920 90 0 0 vccd1
port 20 nsew power bidirectional
flabel metal4 s 2876 2128 3196 19632 0 FreeSans 1920 90 0 0 vssd1
port 21 nsew ground bidirectional
flabel metal4 s 4808 2128 5128 19632 0 FreeSans 1920 90 0 0 vssd1
port 21 nsew ground bidirectional
flabel metal4 s 6740 2128 7060 19632 0 FreeSans 1920 90 0 0 vssd1
port 21 nsew ground bidirectional
flabel metal4 s 8672 2128 8992 19632 0 FreeSans 1920 90 0 0 vssd1
port 21 nsew ground bidirectional
flabel metal3 s 9200 10888 10000 11008 0 FreeSans 480 0 0 0 y
port 22 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 10000 22000
<< end >>
