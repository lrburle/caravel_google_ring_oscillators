magic
tech sky130A
magscale 1 2
timestamp 1713454761
<< nwell >>
rect 0 1674 1180 1748
rect 1342 1674 3267 1748
rect 0 1086 3267 1674
rect 0 921 112 1086
rect 0 819 177 921
rect 2077 804 2291 1086
rect 2078 744 2291 804
rect 3073 772 3103 807
rect 3222 744 3267 1086
<< ndiff >>
rect 3159 442 3193 476
<< locali >>
rect 2 2172 3268 2492
rect 1 1086 3267 1406
rect 175 567 250 578
rect 175 550 214 567
rect 627 550 705 578
rect 1060 572 1099 578
rect 1002 550 1041 572
rect 1370 550 1409 578
rect 1740 550 1780 573
rect 2075 572 2113 576
rect 2074 550 2113 572
rect 150 320 2113 550
rect 1 0 3267 320
<< viali >>
rect 3159 1720 3193 1754
rect 3160 1460 3194 1494
rect 3159 998 3193 1032
rect 3159 442 3193 476
<< metal1 >>
rect 2 2172 3268 2492
rect 1317 1755 1352 2172
rect 1463 1933 1537 1942
rect 1463 1877 1472 1933
rect 1528 1877 1537 1933
rect 2636 1908 2920 1915
rect 2648 1902 2920 1908
rect 1463 1872 1537 1877
rect 2602 1881 2920 1902
rect 1463 1868 1514 1872
rect 2602 1868 2648 1881
rect 2681 1846 2746 1853
rect 2681 1828 2688 1846
rect 1565 1794 2688 1828
rect 2740 1794 2746 1846
rect 2681 1788 2746 1794
rect 1317 1754 1381 1755
rect 1317 1741 1392 1754
rect 1317 1720 1409 1741
rect 2521 1708 2527 1766
rect 2579 1708 2585 1766
rect 1189 1635 1195 1693
rect 1247 1680 1253 1693
rect 2311 1689 2379 1695
rect 2311 1680 2317 1689
rect 1247 1646 2317 1680
rect 1247 1635 1253 1646
rect 2311 1631 2317 1646
rect 2375 1631 2379 1689
rect 2886 1645 2920 1881
rect 2995 1722 3119 1754
rect 2995 1721 3027 1722
rect 3085 1686 3119 1722
rect 3087 1646 3119 1686
rect 2311 1625 2379 1631
rect 3142 1448 3148 1506
rect 3206 1448 3212 1506
rect 1 1086 3267 1406
rect 3141 986 3147 1044
rect 3205 986 3211 1044
rect 1920 861 1984 870
rect 1936 848 1984 861
rect 2313 864 2381 870
rect 1936 811 2113 848
rect 1936 806 1984 811
rect 175 550 214 578
rect 627 550 705 578
rect 1060 572 1099 578
rect 1002 550 1041 572
rect 1370 550 1409 578
rect 2076 576 2113 811
rect 2313 806 2319 864
rect 2377 806 2381 864
rect 2887 819 2921 846
rect 2887 812 2922 819
rect 2888 809 2922 812
rect 2313 800 2381 806
rect 2887 806 2922 809
rect 3065 807 3086 852
rect 2521 790 2585 796
rect 2521 772 2527 790
rect 2515 738 2527 772
rect 2579 738 2585 790
rect 2521 732 2585 738
rect 2676 716 2746 722
rect 2676 698 2682 716
rect 2215 664 2682 698
rect 2215 621 2249 664
rect 2676 658 2682 664
rect 2740 658 2746 716
rect 2676 652 2746 658
rect 2887 624 2920 806
rect 3065 772 3103 807
rect 2994 738 3103 772
rect 2602 623 2636 624
rect 2648 623 2920 624
rect 2075 572 2113 576
rect 2074 550 2113 572
rect 2197 615 2265 621
rect 2197 557 2203 615
rect 2261 557 2265 615
rect 2602 590 2920 623
rect 2197 551 2265 557
rect 150 320 2113 550
rect 1 0 3267 320
<< via1 >>
rect 1472 1877 1528 1933
rect 2688 1794 2740 1846
rect 2527 1708 2579 1766
rect 1195 1635 1247 1693
rect 2317 1631 2375 1689
rect 3148 1494 3206 1506
rect 3148 1460 3160 1494
rect 3160 1460 3194 1494
rect 3194 1460 3206 1494
rect 3148 1448 3206 1460
rect 3147 1032 3205 1044
rect 3147 998 3159 1032
rect 3159 998 3193 1032
rect 3193 998 3205 1032
rect 3147 986 3205 998
rect 2319 806 2377 864
rect 2527 738 2579 790
rect 2682 658 2740 716
rect 2203 557 2261 615
<< metal2 >>
rect 1463 1933 1537 1942
rect 1463 1877 1472 1933
rect 1528 1877 1537 1933
rect 1463 1868 1537 1877
rect 2681 1846 2746 1853
rect 2681 1840 2688 1846
rect 2458 1806 2688 1840
rect 1195 1693 1251 1702
rect 1195 1626 1251 1635
rect 2311 1689 2379 1695
rect 2311 1631 2317 1689
rect 2375 1631 2379 1689
rect 2311 1625 2379 1631
rect 2328 870 2362 1625
rect 2313 864 2381 870
rect 2313 806 2319 864
rect 2377 806 2381 864
rect 2313 800 2381 806
rect 2458 772 2490 1806
rect 2681 1794 2688 1806
rect 2740 1794 2746 1846
rect 2681 1788 2746 1794
rect 2521 1708 2527 1766
rect 2579 1708 2585 1766
rect 2521 1701 2585 1708
rect 2527 1666 2561 1701
rect 2527 1631 2562 1666
rect 2527 1596 2722 1631
rect 2521 790 2585 796
rect 2521 772 2527 790
rect 2458 738 2527 772
rect 2579 738 2585 790
rect 2521 732 2585 738
rect 2687 722 2722 1596
rect 3139 1506 3215 1515
rect 3139 1448 3148 1506
rect 3206 1448 3215 1506
rect 3139 1439 3215 1448
rect 3138 1044 3214 1053
rect 3138 986 3147 1044
rect 3205 986 3214 1044
rect 3138 977 3214 986
rect 2676 716 2746 722
rect 2676 658 2682 716
rect 2740 658 2746 716
rect 500 547 534 657
rect 2676 652 2746 658
rect 2215 621 2249 622
rect 2197 615 2265 621
rect 2197 557 2203 615
rect 2261 557 2265 615
rect 2197 551 2265 557
rect 2197 547 2249 551
rect 500 513 2249 547
<< via2 >>
rect 1472 1877 1528 1933
rect 1195 1635 1247 1693
rect 1247 1635 1251 1693
rect 3148 1448 3206 1506
rect 3147 986 3205 1044
<< metal3 >>
rect 1189 1693 1256 2492
rect 1463 1935 1537 1942
rect 1463 1933 1860 1935
rect 1463 1877 1472 1933
rect 1528 1877 1860 1933
rect 1463 1875 1860 1877
rect 1463 1868 1537 1875
rect 1189 1635 1195 1693
rect 1251 1635 1256 1693
rect 1189 1626 1256 1635
rect 1800 775 1860 1875
rect 3139 1506 3215 2492
rect 3139 1448 3148 1506
rect 3206 1448 3215 1506
rect 3139 1439 3215 1448
rect 1032 715 1452 775
rect 1392 713 1452 715
rect 1640 715 1860 775
rect 3138 1044 3214 1053
rect 3138 986 3147 1044
rect 3205 986 3214 1044
rect 1640 713 1701 715
rect 1392 655 1701 713
rect 1392 652 1664 655
rect 3138 0 3214 986
use scs130hd_mpr2ea_8  scs130hd_mpr2ea_8_0
timestamp 1712673195
transform 1 0 150 0 1 559
box -38 -48 1970 592
use sky130_osu_sc_12T_hs__fill_2  sky130_osu_sc_12T_hs__fill_2_0
timestamp 1713287902
transform 1 0 1728 0 -1 2233
box -7 0 161 897
use sky130_osu_sc_12T_hs__fill_8  sky130_osu_sc_12T_hs__fill_8_0
timestamp 1713287902
transform 1 0 1899 0 -1 2233
box -9 0 179 897
use sky130_osu_sc_12T_hs__inv_1  sky130_osu_sc_12T_hs__inv_1_1
timestamp 1713454387
transform 1 0 2840 0 1 259
box -10 0 199 902
use sky130_osu_sc_12T_hs__inv_1  sky130_osu_sc_12T_hs__inv_1_2
timestamp 1713454387
transform 1 0 3038 0 1 260
box -10 0 199 902
use sky130_osu_sc_12T_hs__inv_1  sky130_osu_sc_12T_hs__inv_1_3
timestamp 1713454387
transform 1 0 3039 0 -1 2232
box -10 0 199 902
use sky130_osu_sc_12T_hs__inv_1  sky130_osu_sc_12T_hs__inv_1_4
timestamp 1713454387
transform 1 0 2840 0 -1 2233
box -10 0 199 902
use sky130_osu_sc_12T_hs__mux2_1  sky130_osu_sc_12T_hs__mux2_1_0
timestamp 1713287902
transform 1 0 2291 0 1 259
box -10 0 552 902
use sky130_osu_sc_12T_hs__mux2_1  sky130_osu_sc_12T_hs__mux2_1_1
timestamp 1713287902
transform 1 0 1168 0 -1 2233
box -10 0 552 902
use sky130_osu_sc_12T_hs__mux2_1  sky130_osu_sc_12T_hs__mux2_1_2
timestamp 1713287902
transform 1 0 2291 0 -1 2233
box -10 0 552 902
<< labels >>
rlabel metal1 76 1151 76 1151 1 vccd1
port 6 n
rlabel metal1 53 293 53 293 1 vssd1
port 5 n
rlabel metal2 2347 837 2347 837 1 sel
port 7 n
rlabel viali 3159 1720 3193 1754 1 Y0
port 9 n
rlabel metal1 1565 1794 1594 1828 1 in
port 8 n
rlabel metal1 53 2200 53 2200 1 vssd1
port 5 n
rlabel metal1 3159 442 3193 476 1 Y1
port 10 n
<< end >>
